//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2017 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------

`ifndef HQM_MRA_CONNECT_CHK_SEQ__SV
`define HQM_MRA_CONNECT_CHK_SEQ__SV

//-----------------------------------------------------------------------------------
// File        : hqm_mra_connect_chk_seq.sv
// Author      : Neeraj Shete
//
// Description : This sequence does the connectivity checks of mra pins driven to HQM.
//               Values are checked within RTL at the points where mra pins are used 
//               within HQM.
//               The RTL points where to check are listed within file below:
//               - tools/mbist/hqm_memory_info.sim_rep.txt
//               - tools/mbist/hqm_memory_info.sim_trim.txt
//-----------------------------------------------------------------------------------

import hqm_tb_sequences_pkg::*;

import "DPI-C" context SLA_VPI_put_value =
  function void hqm_mra_seq_put_value(input chandle handle, input logic [0:0] value);

import "DPI-C" context SLA_VPI_get_value =
  function void hqm_mra_seq_get_value(input chandle handle, output logic [0:0] value);

class hqm_mra_connect_chk_seq extends sla_sequence_base;

  `ovm_object_utils(hqm_mra_connect_chk_seq)
  hqm_reset_sequences_pkg::hqm_cold_reset_sequence  cold_reset;
  pcie_seqlib_pkg::hqm_sla_pcie_init_seq            hqm_pcie_init_seq;

  string mra_ip_bit_q[$], mra_op_bit_q[$];
  string unique_mra_ip_bit_q[$];
  string fuse_mode_check = "";
  bit    mra_ip_val_q[$];
  int    checked_no_of_pins = 0;

  string mem_trim_fuse_ip_bit_q[$], mem_trim_fuse_op_bit_q[$];
  string unique_mem_trim_fuse_ip_bit_q[$];
  bit    mem_trim_fuse_ip_val_q[$];
  int    checked_no_of_mem_trim_pins = 0;


  //----------------------------------------------
  //-- new()
  //----------------------------------------------  
  function new(string name = "hqm_mra_connect_chk_seq");
    super.new(name); 
    mra_ip_bit_q.delete();
    mra_op_bit_q.delete();
    reset_mra_drive();
    reset_mem_trim_fuse_drive();
    if(!$value$plusargs("HQM_FUSE_MODE_CHECK=%s",fuse_mode_check)) fuse_mode_check = "hqm_mra_fuses_check";
  endfunction

  //----------------------------------------------
  //-- body()
  //----------------------------------------------  
  virtual task body();

    // ---------------------------------------------------------------------------------
    // -- Inline include of the file generated by script '' 
    // ---------------------------------------------------------------------------------
    `include "hqm_mra_ip_op_populated_array.svh";

    // ---------------------------------------------------------------------------------
    // -- Inline include of the file generated by script '' 
    // ---------------------------------------------------------------------------------
    `include "hqm_mem_trim_fuse_ip_op_populated_array.svh";
    
    unique_mra_ip_bit_q = mra_ip_bit_q.unique;
    unique_mem_trim_fuse_ip_bit_q = mem_trim_fuse_ip_bit_q.unique;

    if(fuse_mode_check == "hqm_mra_fuses_check") begin
       `ovm_info(get_full_name(), $psprintf(" ------------ Starting MRA fuse array connectivity check ------------- "), OVM_LOW)
       `ovm_info(get_full_name(), $psprintf(" With unique_mra_ip_bit_q size(0x%0x) ", unique_mra_ip_bit_q.size()), OVM_LOW)
       `ovm_info(get_full_name(), $psprintf(" --------------------------------------------------------------------- "), OVM_LOW)
       drive_mra_fuse_walking_ones();
       drive_mra_fuse_walking_zeros();
       drive_mra_fuse_all_zeros();
       drive_mra_fuse_all_ones();
    end else begin
       `ovm_info(get_full_name(), $psprintf(" ------------ Starting mem trim fuse array connectivity check ------------- "), OVM_LOW)
       `ovm_info(get_full_name(), $psprintf(" With unique_mem_trim_fuse_ip_bit_q size(0x%0x) ", unique_mem_trim_fuse_ip_bit_q.size()), OVM_LOW)
       `ovm_info(get_full_name(), $psprintf(" --------------------------------------------------------------------- "), OVM_LOW)
       drive_mem_trim_fuse_walking_ones();
       drive_mem_trim_fuse_walking_zeros();
       drive_mem_trim_fuse_all_zeros();
       drive_mem_trim_fuse_all_ones();
    end

  endtask : body

  function mem_trim_fuse_ip_op_chk();
    chandle             mra_bit_handle;
    string debug_msg = "";
    bit    sig_val, exp_val;
    foreach(mem_trim_fuse_ip_bit_q[k]) begin
       mra_bit_handle = SLA_VPI_get_handle_by_name(mem_trim_fuse_ip_bit_q[k],0);
       hqm_mra_seq_get_value(mra_bit_handle, exp_val);
       mra_bit_handle = SLA_VPI_get_handle_by_name(mem_trim_fuse_op_bit_q[k],0);
       hqm_mra_seq_get_value(mra_bit_handle, sig_val);
       debug_msg = $psprintf("obs_val (0x%0x) and exp_val(0x%0x)",sig_val,exp_val);
       if(sig_val==exp_val) `ovm_info(get_full_name(), $sformatf("Mem margin fuse pin %s value check passed for %s", mem_trim_fuse_op_bit_q[k], debug_msg),OVM_LOW) 
       else                 `ovm_error(get_full_name(),$sformatf("Mem margin fuse pin %s value check failed for %s", mem_trim_fuse_op_bit_q[k], debug_msg))
    end
  endfunction : mem_trim_fuse_ip_op_chk

  task drive_mra_fuse_all_zeros();
      `ovm_info(get_full_name(), $psprintf(" ------ drive_mra_fuse_all_zeros ----- "), OVM_LOW);
      reset_mra_drive();
      foreach(mra_ip_bit_q[i])     begin    mra_ip_val_q.push_back(0);   end
      drive_and_chk_mra_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
  endtask : drive_mra_fuse_all_zeros

  task drive_mra_fuse_all_ones();
      `ovm_info(get_full_name(), $psprintf(" ------ drive_mra_fuse_all_ones ----- "), OVM_LOW);
      reset_mra_drive();
      foreach(mra_ip_bit_q[i])     begin    mra_ip_val_q.push_back(1);   end
      drive_and_chk_mra_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
  endtask : drive_mra_fuse_all_ones

  task drive_mra_fuse_walking_zeros();
    foreach(unique_mra_ip_bit_q[i]) begin
      `ovm_info(get_full_name(), $psprintf("drive_mra_fuse_walking_zeros: selected input signal is %s", unique_mra_ip_bit_q[i]), OVM_LOW);
      reset_mra_drive();
      for(int k=0; k<mra_ip_bit_q.size(); k++) begin
         mra_ip_val_q.push_back(mra_ip_bit_q[k] != unique_mra_ip_bit_q[i]);
      end
      drive_and_chk_mra_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
    end
  endtask : drive_mra_fuse_walking_zeros

  task drive_mra_fuse_walking_ones();
    foreach(unique_mra_ip_bit_q[i]) begin
      `ovm_info(get_full_name(), $psprintf("drive_mra_fuse_walking_ones: selected input signal is %s", unique_mra_ip_bit_q[i]), OVM_LOW);
      reset_mra_drive();
      for(int k=0; k<mra_ip_bit_q.size(); k++) begin
         mra_ip_val_q.push_back(mra_ip_bit_q[k] == unique_mra_ip_bit_q[i]);
      end
      drive_and_chk_mra_bits();
      repeat(50) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
    end
  endtask : drive_mra_fuse_walking_ones

  task drive_mem_trim_fuse_all_ones();
      `ovm_info(get_full_name(), $psprintf(" --------- drive_mem_trim_fuse_all_ones --------- "), OVM_LOW);
      reset_mem_trim_fuse_drive();
      foreach(mem_trim_fuse_ip_bit_q[i]) begin mem_trim_fuse_ip_val_q.push_back(1); end
      drive_and_chk_mem_trim_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
  endtask : drive_mem_trim_fuse_all_ones

  task drive_mem_trim_fuse_all_zeros();
      `ovm_info(get_full_name(), $psprintf(" --------- drive_mem_trim_fuse_all_zeros --------- "), OVM_LOW);
      reset_mem_trim_fuse_drive();
      foreach(mem_trim_fuse_ip_bit_q[i]) begin mem_trim_fuse_ip_val_q.push_back(0); end
      drive_and_chk_mem_trim_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
  endtask : drive_mem_trim_fuse_all_zeros

  task drive_mem_trim_fuse_walking_zeros();
    foreach(unique_mem_trim_fuse_ip_bit_q[i]) begin
      `ovm_info(get_full_name(), $psprintf("drive_mem_trim_fuse_walking_zeros: selected input signal is %s", unique_mem_trim_fuse_ip_bit_q[i]), OVM_LOW);
      reset_mem_trim_fuse_drive();
      for(int k=0; k<mem_trim_fuse_ip_bit_q.size(); k++) begin
         mem_trim_fuse_ip_val_q.push_back(mem_trim_fuse_ip_bit_q[k] != unique_mem_trim_fuse_ip_bit_q[i]);
      end
      drive_and_chk_mem_trim_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
    end
  endtask : drive_mem_trim_fuse_walking_zeros

  task drive_mem_trim_fuse_walking_ones();
    foreach(unique_mem_trim_fuse_ip_bit_q[i]) begin
      `ovm_info(get_full_name(), $psprintf("drive_mem_trim_fuse_walking_ones: selected input signal is %s", unique_mem_trim_fuse_ip_bit_q[i]), OVM_LOW);
      reset_mem_trim_fuse_drive();
      for(int k=0; k<mem_trim_fuse_ip_bit_q.size(); k++) begin
         mem_trim_fuse_ip_val_q.push_back(mem_trim_fuse_ip_bit_q[k] == unique_mem_trim_fuse_ip_bit_q[i]);
      end
      drive_and_chk_mem_trim_bits();
      repeat(100) begin @(sla_tb_env::sys_clk_r); end // -- Added some delay before next drive -- //
    end
  endtask : drive_mem_trim_fuse_walking_ones

  task drive_and_chk_mem_trim_bits();

    `ovm_info(get_full_name(), $psprintf(" -------- Starting drive_and_chk_mem_trim_bits ---------"), OVM_LOW)

    foreach(mem_trim_fuse_ip_bit_q[i]) begin
       automatic string pin_name = mem_trim_fuse_ip_bit_q[i];
       automatic bit    val      = mem_trim_fuse_ip_val_q[i];
       fork  begin set_val(pin_name,val, .trim_fuse(1)); end  join_none
    end

    `ovm_info(get_full_name(), $psprintf("Drove all input pins mem_trim_fuse_ip_bit_q.size() (0x%0x)", mem_trim_fuse_ip_bit_q.size()), OVM_LOW)
  
    // -- `ovm_do(cold_reset);
    // -- `ovm_do(hqm_pcie_init_seq);

    foreach(mem_trim_fuse_op_bit_q[i]) begin
       automatic string pin_name = mem_trim_fuse_op_bit_q[i];
       automatic bit    val      = mem_trim_fuse_ip_val_q[i];
       fork  begin chk_val(pin_name,val, .trim_fuse(1)); checked_no_of_mem_trim_pins++; end  join_none
    end

    `ovm_info(get_full_name(), $psprintf("Waiting to check connectivity of all pins checked_no_of_mem_trim_pins (0x%0x), mem_trim_fuse_op_bit_q.size() (0x%0x)", checked_no_of_mem_trim_pins, mem_trim_fuse_op_bit_q.size()), OVM_LOW)

    wait (checked_no_of_mem_trim_pins == mem_trim_fuse_op_bit_q.size());

    `ovm_info(get_full_name(), $psprintf("Done checking connectivity of all pins checked_no_of_mem_trim_pins (0x%0x), mem_trim_fuse_op_bit_q.size() (0x%0x)", checked_no_of_mem_trim_pins, mem_trim_fuse_op_bit_q.size()), OVM_LOW)

    `ovm_info(get_full_name(), $psprintf(" -------- Done drive_and_chk_mem_trim_bits ---------"), OVM_LOW)

  endtask : drive_and_chk_mem_trim_bits


  function reset_mem_trim_fuse_drive();
    mem_trim_fuse_ip_val_q.delete();
    checked_no_of_mem_trim_pins = 0;
    `ovm_info(get_full_name(), $sformatf("Done deleting mem_trim_fuse_ip_val_q -> size(0x%0x) and set checked_no_of_mem_trim_pins to (0x%0x)", mem_trim_fuse_ip_val_q.size(),checked_no_of_mem_trim_pins), OVM_LOW)
  endfunction : reset_mem_trim_fuse_drive

  function reset_mra_drive();
    mra_ip_val_q.delete();
    checked_no_of_pins = 0;
    `ovm_info(get_full_name(), $sformatf("Done deleting mra_ip_val_q -> size(0x%0x) and set checked_no_of_pins to (0x%0x)", mra_ip_val_q.size(),checked_no_of_pins), OVM_LOW)
  endfunction : reset_mra_drive

  task drive_and_chk_mra_bits();

    `ovm_info(get_full_name(), $psprintf(" -------- Starting drive_and_chk_mra_bits ---------"), OVM_LOW)

    foreach(mra_ip_bit_q[i]) begin
       automatic string pin_name = mra_ip_bit_q[i];
       automatic bit    val      = mra_ip_val_q[i];
       fork  begin set_val(pin_name,val); end  join_none
    end

    `ovm_info(get_full_name(), $psprintf("Drove all input pins mra_ip_bit_q.size() (0x%0x)", mra_ip_bit_q.size()), OVM_LOW)
  
    // -- `ovm_do(cold_reset);
    // -- `ovm_do(hqm_pcie_init_seq);

    foreach(mra_op_bit_q[i]) begin
       automatic string pin_name = mra_op_bit_q[i];
       automatic bit    val      = mra_ip_val_q[i];
       fork  begin chk_val(pin_name,val); checked_no_of_pins++; end  join_none
    end

    `ovm_info(get_full_name(), $psprintf("Waiting to check connectivity of all pins checked_no_of_pins (0x%0x), mra_op_bit_q.size() (0x%0x)", checked_no_of_pins, mra_op_bit_q.size()), OVM_LOW)

    wait (checked_no_of_pins == mra_op_bit_q.size());

    `ovm_info(get_full_name(), $psprintf("Done checking connectivity of all pins checked_no_of_pins (0x%0x), mra_op_bit_q.size() (0x%0x)", checked_no_of_pins, mra_op_bit_q.size()), OVM_LOW)

    `ovm_info(get_full_name(), $psprintf(" -------- Done drive_and_chk_mra_bits ---------"), OVM_LOW)

  endtask : drive_and_chk_mra_bits

  task set_val(string pin_name, bit sig_val, bit trim_fuse = 0);
    chandle             mra_bit_handle;
    string              debug_msg="";
    string              hdr_str  ="";

    mra_bit_handle = SLA_VPI_get_handle_by_name(pin_name,0);
    hqm_mra_seq_put_value(mra_bit_handle, sig_val);
    debug_msg = $psprintf("set_val (0x%0x)",sig_val);

    if(trim_fuse)  hdr_str = "MEM trim fuse"; else hdr_str = "MRA pin";
    `ovm_info(get_full_name(), $sformatf("%s %s: %s", hdr_str, pin_name, debug_msg),OVM_LOW) 
  endtask

  task chk_val(string pin_name, bit exp_val, bit trim_fuse = 0, int clk_ticks = 1000);
    chandle             mra_bit_handle;
    string              debug_msg = "", hdr_str = "";
    bit                 sig_val;

    repeat(clk_ticks) begin @(sla_tb_env::sys_clk_r); end

// --    for(int i = 0; i<10; i++) begin
       mra_bit_handle = SLA_VPI_get_handle_by_name(pin_name,0);
       hqm_mra_seq_get_value(mra_bit_handle, sig_val);
       debug_msg = $psprintf("obs_val (0x%0x) and exp_val(0x%0x)",sig_val,exp_val);
  
       if(trim_fuse)  hdr_str = "MEM trim fuse"; else hdr_str = "MRA pin";
       // -- `ovm_info(get_full_name(), $sformatf("%s %s value @clk_tick %0d is, %s", hdr_str, pin_name, i, debug_msg),OVM_DEBUG) 

       // -- if(sig_val != exp_val) break;
   
// --    end

    if(sig_val==exp_val) `ovm_info(get_full_name(), $sformatf("%s %s value check passed for %s", hdr_str, pin_name, debug_msg),OVM_LOW) 
    else                 `ovm_error(get_full_name(),$sformatf("%s %s value check failed for %s", hdr_str, pin_name, debug_msg))

  endtask

endclass : hqm_mra_connect_chk_seq

`endif
