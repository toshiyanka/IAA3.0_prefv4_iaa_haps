
`ifndef HQM_RESET_PKG__SV
`define HQM_RESET_PKG__SV

package hqm_reset_pkg;

   import ovm_pkg::*;
   import sla_pkg::*;

  `include "ovm_macros.svh"
  `include "sla_macros.svh"

  `include "hqm_reset_types.sv"
  `include "hqm_reset_transaction.sv"
  `include "hqm_reset_config.sv"
  `include "hqm_reset_driver.sv"
  `include "hqm_reset_monitor.sv"
  `include "hqm_reset_sequencer.sv"
  `include "hqm_reset_agent.sv"

endpackage

`endif
