module ctech_lib_clk_inv (
   input logic clk,
   output logic clkout
);
   d04gin00ld0c0 ctech_lib_dcszo (.clk(clk), .clkout(clkout));
endmodule
