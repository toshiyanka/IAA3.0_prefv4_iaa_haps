// File output was printed on: Thursday, March 21, 2013 4:21:02 PM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
//              TAP name,      Opcode,   DR_length
//
Create_Reg_Model (IPLEVEL_STAP,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (IPLEVEL_STAP,   8'hC,      'd32     );   // opcode is SLVIDCODE [0xC]
Create_Reg_Model (IPLEVEL_STAP,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
