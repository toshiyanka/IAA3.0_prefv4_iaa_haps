//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2022 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------

module hqm_mem_ctech_doublesync_rstb (
   input  logic clk,
   input  logic rstb,
   input  logic d,
   output logic o
);
ctech_lib_doublesync_rstb ctech_lib_doublesync_rstb (.clk(clk), .d(d), .rstb(rstb), .o(o));
endmodule

module hqm_mem_ctech_buf (
   input logic a,
   output logic o
);
ctech_lib_buf ctech_lib_buf(.a(a), .o(o));
endmodule

