module bogus_verilog;
endmodule //bogus_verilog;