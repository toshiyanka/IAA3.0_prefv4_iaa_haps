//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// AW_lsfr_load
//
// implements a LSFR counter using the following paramters & inputs.
//   WIDTH	(1 to 50) Word length of counter
//   enable     0:stop counting  1:enable counting
//   load_seed  0:do not use input seed (use default seed)  1:use input seed
//   seed       is WIDTH wide and used to seed LSFR when enabled
//   output     LSFR counter output 
//
//-----------------------------------------------------------------------------------------------------

module hqm_AW_lsfr_load
       import hqm_AW_pkg::*; #(

	 parameter WIDTH	= 2
) (
	 input	logic			clk
	,input	logic			rst_n
	,input	logic			enable
	,input	logic			load_seed
	,input	logic	[WIDTH-1:0]	seed
	,output	logic	[WIDTH-1:0]	count
);

DW03_lfsr_load #(WIDTH) i_DW03_lfsr_load ( 

	 .clk	(clk)
	,.reset	(rst_n) 
	,.cen	(enable)
	,.load	(load_seed)
	,.data	(seed)
	,.count	(count) 
);

endmodule 

