VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf156b040e2r2w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf156b040e2r2w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 37.8 BY 46.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 23.64 13.628 24.84 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.444 23.64 17.488 24.84 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 20.76 13.628 21.96 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.612 20.76 17.656 21.96 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 23.64 15.428 24.84 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.644 23.64 15.688 24.84 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 23.64 15.856 24.84 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 23.64 16.116 24.84 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 23.64 16.416 24.84 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 23.64 17.228 24.84 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 23.64 14.316 24.84 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.64 14.616 24.84 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 23.64 19.028 24.84 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 23.64 19.288 24.84 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 23.64 19.716 24.84 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 23.64 20.016 24.84 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 23.64 20.828 24.84 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 23.64 21.088 24.84 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.612 23.64 17.656 24.84 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 23.64 18.216 24.84 ;
    END
  END rdaddrp1_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 23.64 14.872 24.84 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 23.64 18.472 24.84 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 23.64 15.128 24.84 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 23.64 18.728 24.84 ;
    END
  END sdl_initp1
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.644 20.76 15.688 21.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 20.76 15.856 21.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 20.76 16.116 21.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 20.76 16.416 21.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 20.76 17.228 21.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.444 20.76 17.488 21.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 20.76 14.316 21.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 20.76 14.616 21.96 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 20.76 19.716 21.96 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 20.76 20.016 21.96 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 20.76 20.828 21.96 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 20.76 21.088 21.96 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 20.76 21.256 21.96 ;
    END
  END wraddrp1[4]
  PIN wraddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 20.76 21.516 21.96 ;
    END
  END wraddrp1[5]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 20.76 18.216 21.96 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 20.76 18.472 21.96 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 0.36 16.116 1.56 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 30.6 15.772 31.8 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 30.6 15.856 31.8 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 30.6 18.816 31.8 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 30.6 19.028 31.8 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 31.56 16.928 32.76 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 31.56 17.016 32.76 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 31.56 19.628 32.76 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 31.56 17.916 32.76 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 32.52 15.772 33.72 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 32.52 15.856 33.72 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 2.28 18.556 3.48 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 32.52 18.816 33.72 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 32.52 19.028 33.72 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 33.48 16.928 34.68 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 33.48 17.016 34.68 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 33.48 19.628 34.68 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 33.48 17.916 34.68 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 34.44 15.772 35.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 34.44 15.856 35.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 34.44 18.816 35.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 34.44 19.028 35.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 2.28 18.728 3.48 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 35.4 16.928 36.6 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 35.4 17.016 36.6 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 35.4 19.628 36.6 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 35.4 17.916 36.6 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 36.36 15.772 37.56 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 36.36 15.856 37.56 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 36.36 18.816 37.56 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 36.36 19.028 37.56 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 37.32 16.928 38.52 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 37.32 17.016 38.52 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 3.24 16.672 4.44 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 37.32 19.628 38.52 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 37.32 17.916 38.52 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 38.28 15.772 39.48 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 38.28 15.856 39.48 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 38.28 18.816 39.48 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 38.28 19.028 39.48 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 39.24 16.928 40.44 ;
    END
  END wrdatap0[136]
  PIN wrdatap0[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 39.24 17.016 40.44 ;
    END
  END wrdatap0[137]
  PIN wrdatap0[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 39.24 19.628 40.44 ;
    END
  END wrdatap0[138]
  PIN wrdatap0[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 39.24 17.916 40.44 ;
    END
  END wrdatap0[139]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 3.24 16.756 4.44 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 40.2 15.772 41.4 ;
    END
  END wrdatap0[140]
  PIN wrdatap0[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 40.2 15.856 41.4 ;
    END
  END wrdatap0[141]
  PIN wrdatap0[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 40.2 18.816 41.4 ;
    END
  END wrdatap0[142]
  PIN wrdatap0[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 40.2 19.028 41.4 ;
    END
  END wrdatap0[143]
  PIN wrdatap0[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 41.16 16.928 42.36 ;
    END
  END wrdatap0[144]
  PIN wrdatap0[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 41.16 17.016 42.36 ;
    END
  END wrdatap0[145]
  PIN wrdatap0[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 41.16 19.628 42.36 ;
    END
  END wrdatap0[146]
  PIN wrdatap0[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 41.16 17.916 42.36 ;
    END
  END wrdatap0[147]
  PIN wrdatap0[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 42.12 15.772 43.32 ;
    END
  END wrdatap0[148]
  PIN wrdatap0[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 42.12 15.856 43.32 ;
    END
  END wrdatap0[149]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 3.24 19.456 4.44 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 42.12 18.816 43.32 ;
    END
  END wrdatap0[150]
  PIN wrdatap0[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 42.12 19.028 43.32 ;
    END
  END wrdatap0[151]
  PIN wrdatap0[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 43.08 16.928 44.28 ;
    END
  END wrdatap0[152]
  PIN wrdatap0[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 43.08 17.016 44.28 ;
    END
  END wrdatap0[153]
  PIN wrdatap0[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 43.08 19.628 44.28 ;
    END
  END wrdatap0[154]
  PIN wrdatap0[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 43.08 17.916 44.28 ;
    END
  END wrdatap0[155]
  PIN wrdatap0[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 44.04 15.772 45.24 ;
    END
  END wrdatap0[156]
  PIN wrdatap0[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 44.04 15.856 45.24 ;
    END
  END wrdatap0[157]
  PIN wrdatap0[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 44.04 18.816 45.24 ;
    END
  END wrdatap0[158]
  PIN wrdatap0[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 44.04 19.028 45.24 ;
    END
  END wrdatap0[159]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 3.24 19.628 4.44 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 4.2 17.572 5.4 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 4.2 15.772 5.4 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 4.2 18.556 5.4 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 4.2 18.728 5.4 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 0.36 16.328 1.56 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 5.16 16.672 6.36 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 5.16 16.756 6.36 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 5.16 19.456 6.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 5.16 19.628 6.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 6.12 17.572 7.32 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 6.12 15.772 7.32 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 6.12 18.556 7.32 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 6.12 18.728 7.32 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 7.08 16.672 8.28 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 7.08 16.756 8.28 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.36 18.816 1.56 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 7.08 19.456 8.28 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 7.08 19.628 8.28 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 8.04 17.572 9.24 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 8.04 15.772 9.24 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 8.04 18.556 9.24 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 8.04 18.728 9.24 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 9 16.672 10.2 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 9 16.756 10.2 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 9 19.456 10.2 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 9 19.628 10.2 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.36 19.028 1.56 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 9.96 17.572 11.16 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 9.96 15.772 11.16 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 9.96 18.556 11.16 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 9.96 18.728 11.16 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 10.92 16.672 12.12 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 10.92 16.756 12.12 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 10.92 19.456 12.12 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 10.92 19.628 12.12 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 11.88 17.572 13.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 11.88 15.772 13.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 1.32 16.756 2.52 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 11.88 18.556 13.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.88 18.728 13.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 12.84 16.672 14.04 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 12.84 16.756 14.04 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 12.84 19.456 14.04 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 12.84 19.628 14.04 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 13.8 17.572 15 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 13.8 15.772 15 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 13.8 18.556 15 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 13.8 18.728 15 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 1.32 16.928 2.52 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 14.76 16.672 15.96 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 14.76 16.756 15.96 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 14.76 19.456 15.96 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 14.76 19.628 15.96 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 15.72 17.572 16.92 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 15.72 15.772 16.92 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 15.72 18.556 16.92 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 15.72 18.728 16.92 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 16.68 16.672 17.88 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 16.68 16.756 17.88 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 1.32 19.456 2.52 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 16.68 19.456 17.88 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 16.68 19.628 17.88 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 17.64 17.572 18.84 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 17.64 15.772 18.84 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 17.64 18.556 18.84 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 17.64 18.728 18.84 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 18.6 16.672 19.8 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 18.6 16.756 19.8 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 18.6 19.456 19.8 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 18.6 19.628 19.8 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 1.32 19.628 2.52 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 25.8 16.756 27 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 25.8 16.928 27 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 25.8 19.628 27 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 25.8 17.916 27 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 26.76 15.772 27.96 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 26.76 15.856 27.96 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.76 18.816 27.96 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.76 19.028 27.96 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 27.72 16.928 28.92 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 27.72 17.016 28.92 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 2.28 17.572 3.48 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 27.72 19.628 28.92 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 27.72 17.916 28.92 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 28.68 15.772 29.88 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 28.68 15.856 29.88 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 28.68 18.816 29.88 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 28.68 19.028 29.88 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 29.64 16.928 30.84 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 29.64 17.016 30.84 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 29.64 19.628 30.84 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 29.64 17.916 30.84 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 2.28 15.772 3.48 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 20.76 15.128 21.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 20.76 15.428 21.96 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 0.36 16.416 1.56 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 30.6 16.028 31.8 ;
    END
  END wrdatap1[100]
  PIN wrdatap1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 30.6 16.116 31.8 ;
    END
  END wrdatap1[101]
  PIN wrdatap1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 30.6 19.116 31.8 ;
    END
  END wrdatap1[102]
  PIN wrdatap1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 30.6 19.288 31.8 ;
    END
  END wrdatap1[103]
  PIN wrdatap1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 31.56 17.228 32.76 ;
    END
  END wrdatap1[104]
  PIN wrdatap1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 31.56 17.316 32.76 ;
    END
  END wrdatap1[105]
  PIN wrdatap1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 31.56 18.128 32.76 ;
    END
  END wrdatap1[106]
  PIN wrdatap1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 31.56 18.216 32.76 ;
    END
  END wrdatap1[107]
  PIN wrdatap1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 32.52 16.028 33.72 ;
    END
  END wrdatap1[108]
  PIN wrdatap1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 32.52 16.116 33.72 ;
    END
  END wrdatap1[109]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 2.28 18.816 3.48 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 32.52 19.116 33.72 ;
    END
  END wrdatap1[110]
  PIN wrdatap1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 32.52 19.288 33.72 ;
    END
  END wrdatap1[111]
  PIN wrdatap1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 33.48 17.228 34.68 ;
    END
  END wrdatap1[112]
  PIN wrdatap1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 33.48 17.316 34.68 ;
    END
  END wrdatap1[113]
  PIN wrdatap1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 33.48 18.128 34.68 ;
    END
  END wrdatap1[114]
  PIN wrdatap1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 33.48 18.216 34.68 ;
    END
  END wrdatap1[115]
  PIN wrdatap1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 34.44 16.028 35.64 ;
    END
  END wrdatap1[116]
  PIN wrdatap1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 34.44 16.116 35.64 ;
    END
  END wrdatap1[117]
  PIN wrdatap1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 34.44 19.116 35.64 ;
    END
  END wrdatap1[118]
  PIN wrdatap1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 34.44 19.288 35.64 ;
    END
  END wrdatap1[119]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 2.28 19.028 3.48 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 35.4 17.228 36.6 ;
    END
  END wrdatap1[120]
  PIN wrdatap1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 35.4 17.316 36.6 ;
    END
  END wrdatap1[121]
  PIN wrdatap1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 35.4 18.128 36.6 ;
    END
  END wrdatap1[122]
  PIN wrdatap1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 35.4 18.216 36.6 ;
    END
  END wrdatap1[123]
  PIN wrdatap1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 36.36 16.028 37.56 ;
    END
  END wrdatap1[124]
  PIN wrdatap1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 36.36 16.116 37.56 ;
    END
  END wrdatap1[125]
  PIN wrdatap1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 36.36 19.116 37.56 ;
    END
  END wrdatap1[126]
  PIN wrdatap1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 36.36 19.288 37.56 ;
    END
  END wrdatap1[127]
  PIN wrdatap1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 37.32 17.228 38.52 ;
    END
  END wrdatap1[128]
  PIN wrdatap1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 37.32 17.316 38.52 ;
    END
  END wrdatap1[129]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 3.24 16.928 4.44 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 37.32 18.128 38.52 ;
    END
  END wrdatap1[130]
  PIN wrdatap1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 37.32 18.216 38.52 ;
    END
  END wrdatap1[131]
  PIN wrdatap1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 38.28 16.028 39.48 ;
    END
  END wrdatap1[132]
  PIN wrdatap1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 38.28 16.116 39.48 ;
    END
  END wrdatap1[133]
  PIN wrdatap1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 38.28 19.116 39.48 ;
    END
  END wrdatap1[134]
  PIN wrdatap1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 38.28 19.288 39.48 ;
    END
  END wrdatap1[135]
  PIN wrdatap1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 39.24 17.228 40.44 ;
    END
  END wrdatap1[136]
  PIN wrdatap1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 39.24 17.316 40.44 ;
    END
  END wrdatap1[137]
  PIN wrdatap1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 39.24 18.128 40.44 ;
    END
  END wrdatap1[138]
  PIN wrdatap1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 39.24 18.216 40.44 ;
    END
  END wrdatap1[139]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 3.24 17.016 4.44 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 40.2 16.028 41.4 ;
    END
  END wrdatap1[140]
  PIN wrdatap1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 40.2 16.116 41.4 ;
    END
  END wrdatap1[141]
  PIN wrdatap1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 40.2 19.116 41.4 ;
    END
  END wrdatap1[142]
  PIN wrdatap1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 40.2 19.288 41.4 ;
    END
  END wrdatap1[143]
  PIN wrdatap1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 41.16 17.228 42.36 ;
    END
  END wrdatap1[144]
  PIN wrdatap1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 41.16 17.316 42.36 ;
    END
  END wrdatap1[145]
  PIN wrdatap1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 41.16 18.128 42.36 ;
    END
  END wrdatap1[146]
  PIN wrdatap1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 41.16 18.216 42.36 ;
    END
  END wrdatap1[147]
  PIN wrdatap1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 42.12 16.028 43.32 ;
    END
  END wrdatap1[148]
  PIN wrdatap1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 42.12 16.116 43.32 ;
    END
  END wrdatap1[149]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 3.24 17.916 4.44 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 42.12 19.116 43.32 ;
    END
  END wrdatap1[150]
  PIN wrdatap1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 42.12 19.288 43.32 ;
    END
  END wrdatap1[151]
  PIN wrdatap1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 43.08 17.228 44.28 ;
    END
  END wrdatap1[152]
  PIN wrdatap1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 43.08 17.316 44.28 ;
    END
  END wrdatap1[153]
  PIN wrdatap1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 43.08 18.128 44.28 ;
    END
  END wrdatap1[154]
  PIN wrdatap1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 43.08 18.216 44.28 ;
    END
  END wrdatap1[155]
  PIN wrdatap1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 44.04 16.028 45.24 ;
    END
  END wrdatap1[156]
  PIN wrdatap1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 44.04 16.116 45.24 ;
    END
  END wrdatap1[157]
  PIN wrdatap1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 44.04 19.116 45.24 ;
    END
  END wrdatap1[158]
  PIN wrdatap1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 44.04 19.288 45.24 ;
    END
  END wrdatap1[159]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 3.24 18.128 4.44 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 4.2 15.856 5.4 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 4.2 16.028 5.4 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 4.2 18.816 5.4 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 4.2 19.028 5.4 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.544 0.36 16.588 1.56 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 5.16 16.928 6.36 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 5.16 17.016 6.36 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 5.16 17.916 6.36 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 5.16 18.128 6.36 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 6.12 15.856 7.32 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 6.12 16.028 7.32 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 6.12 18.816 7.32 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 6.12 19.028 7.32 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 7.08 16.928 8.28 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 7.08 17.016 8.28 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 0.36 19.116 1.56 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 7.08 17.916 8.28 ;
    END
  END wrdatap1[30]
  PIN wrdatap1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 7.08 18.128 8.28 ;
    END
  END wrdatap1[31]
  PIN wrdatap1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 8.04 15.856 9.24 ;
    END
  END wrdatap1[32]
  PIN wrdatap1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 8.04 16.028 9.24 ;
    END
  END wrdatap1[33]
  PIN wrdatap1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.04 18.816 9.24 ;
    END
  END wrdatap1[34]
  PIN wrdatap1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.04 19.028 9.24 ;
    END
  END wrdatap1[35]
  PIN wrdatap1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 9 16.928 10.2 ;
    END
  END wrdatap1[36]
  PIN wrdatap1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 9 17.016 10.2 ;
    END
  END wrdatap1[37]
  PIN wrdatap1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 9 17.916 10.2 ;
    END
  END wrdatap1[38]
  PIN wrdatap1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 9 18.128 10.2 ;
    END
  END wrdatap1[39]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 0.36 19.288 1.56 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 9.96 15.856 11.16 ;
    END
  END wrdatap1[40]
  PIN wrdatap1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 9.96 16.028 11.16 ;
    END
  END wrdatap1[41]
  PIN wrdatap1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 9.96 18.816 11.16 ;
    END
  END wrdatap1[42]
  PIN wrdatap1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 9.96 19.028 11.16 ;
    END
  END wrdatap1[43]
  PIN wrdatap1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 10.92 16.928 12.12 ;
    END
  END wrdatap1[44]
  PIN wrdatap1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 10.92 17.016 12.12 ;
    END
  END wrdatap1[45]
  PIN wrdatap1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 10.92 17.916 12.12 ;
    END
  END wrdatap1[46]
  PIN wrdatap1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 10.92 18.128 12.12 ;
    END
  END wrdatap1[47]
  PIN wrdatap1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 11.88 15.856 13.08 ;
    END
  END wrdatap1[48]
  PIN wrdatap1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 11.88 16.028 13.08 ;
    END
  END wrdatap1[49]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 1.32 17.016 2.52 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 11.88 18.816 13.08 ;
    END
  END wrdatap1[50]
  PIN wrdatap1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 11.88 19.028 13.08 ;
    END
  END wrdatap1[51]
  PIN wrdatap1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 12.84 16.928 14.04 ;
    END
  END wrdatap1[52]
  PIN wrdatap1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 12.84 17.016 14.04 ;
    END
  END wrdatap1[53]
  PIN wrdatap1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 12.84 17.916 14.04 ;
    END
  END wrdatap1[54]
  PIN wrdatap1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 12.84 18.128 14.04 ;
    END
  END wrdatap1[55]
  PIN wrdatap1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 13.8 15.856 15 ;
    END
  END wrdatap1[56]
  PIN wrdatap1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 13.8 16.028 15 ;
    END
  END wrdatap1[57]
  PIN wrdatap1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 13.8 18.816 15 ;
    END
  END wrdatap1[58]
  PIN wrdatap1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 13.8 19.028 15 ;
    END
  END wrdatap1[59]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 1.32 17.228 2.52 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 14.76 16.928 15.96 ;
    END
  END wrdatap1[60]
  PIN wrdatap1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 14.76 17.016 15.96 ;
    END
  END wrdatap1[61]
  PIN wrdatap1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 14.76 17.916 15.96 ;
    END
  END wrdatap1[62]
  PIN wrdatap1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 14.76 18.128 15.96 ;
    END
  END wrdatap1[63]
  PIN wrdatap1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 15.72 15.856 16.92 ;
    END
  END wrdatap1[64]
  PIN wrdatap1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 15.72 16.028 16.92 ;
    END
  END wrdatap1[65]
  PIN wrdatap1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 15.72 18.816 16.92 ;
    END
  END wrdatap1[66]
  PIN wrdatap1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 15.72 19.028 16.92 ;
    END
  END wrdatap1[67]
  PIN wrdatap1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 16.68 16.928 17.88 ;
    END
  END wrdatap1[68]
  PIN wrdatap1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 16.68 17.016 17.88 ;
    END
  END wrdatap1[69]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 1.32 17.916 2.52 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 16.68 17.916 17.88 ;
    END
  END wrdatap1[70]
  PIN wrdatap1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 16.68 18.128 17.88 ;
    END
  END wrdatap1[71]
  PIN wrdatap1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 17.64 15.856 18.84 ;
    END
  END wrdatap1[72]
  PIN wrdatap1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 17.64 16.028 18.84 ;
    END
  END wrdatap1[73]
  PIN wrdatap1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 17.64 18.816 18.84 ;
    END
  END wrdatap1[74]
  PIN wrdatap1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 17.64 19.028 18.84 ;
    END
  END wrdatap1[75]
  PIN wrdatap1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 18.6 16.928 19.8 ;
    END
  END wrdatap1[76]
  PIN wrdatap1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 18.6 17.016 19.8 ;
    END
  END wrdatap1[77]
  PIN wrdatap1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 18.6 17.916 19.8 ;
    END
  END wrdatap1[78]
  PIN wrdatap1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 18.6 18.128 19.8 ;
    END
  END wrdatap1[79]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 1.32 18.128 2.52 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 25.8 17.016 27 ;
    END
  END wrdatap1[80]
  PIN wrdatap1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 25.8 17.316 27 ;
    END
  END wrdatap1[81]
  PIN wrdatap1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 25.8 18.128 27 ;
    END
  END wrdatap1[82]
  PIN wrdatap1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.344 25.8 18.388 27 ;
    END
  END wrdatap1[83]
  PIN wrdatap1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 26.76 16.028 27.96 ;
    END
  END wrdatap1[84]
  PIN wrdatap1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 26.76 16.116 27.96 ;
    END
  END wrdatap1[85]
  PIN wrdatap1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 26.76 19.116 27.96 ;
    END
  END wrdatap1[86]
  PIN wrdatap1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 26.76 19.288 27.96 ;
    END
  END wrdatap1[87]
  PIN wrdatap1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 27.72 17.228 28.92 ;
    END
  END wrdatap1[88]
  PIN wrdatap1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 27.72 17.316 28.92 ;
    END
  END wrdatap1[89]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 2.28 15.856 3.48 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 27.72 18.128 28.92 ;
    END
  END wrdatap1[90]
  PIN wrdatap1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 27.72 18.216 28.92 ;
    END
  END wrdatap1[91]
  PIN wrdatap1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 28.68 16.028 29.88 ;
    END
  END wrdatap1[92]
  PIN wrdatap1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 28.68 16.116 29.88 ;
    END
  END wrdatap1[93]
  PIN wrdatap1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 28.68 19.116 29.88 ;
    END
  END wrdatap1[94]
  PIN wrdatap1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 28.68 19.288 29.88 ;
    END
  END wrdatap1[95]
  PIN wrdatap1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 29.64 17.228 30.84 ;
    END
  END wrdatap1[96]
  PIN wrdatap1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 29.64 17.316 30.84 ;
    END
  END wrdatap1[97]
  PIN wrdatap1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 29.64 18.128 30.84 ;
    END
  END wrdatap1[98]
  PIN wrdatap1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 29.64 18.216 30.84 ;
    END
  END wrdatap1[99]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 2.28 16.028 3.48 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 20.76 19.028 21.96 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 20.76 19.288 21.96 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 20.76 14.872 21.96 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 20.76 18.728 21.96 ;
    END
  END wrenp1
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 0.36 13.628 1.56 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 30.6 15.128 31.8 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 30.6 15.216 31.8 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 30.6 21.516 31.8 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 30.6 21.728 31.8 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 31.56 13.888 32.76 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 31.56 13.972 32.76 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 31.56 20.528 32.76 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 31.56 20.616 32.76 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 32.52 15.128 33.72 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 32.52 15.216 33.72 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 2.28 21.428 3.48 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 32.52 21.516 33.72 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 32.52 21.728 33.72 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 33.48 13.888 34.68 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 33.48 13.972 34.68 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 33.48 20.528 34.68 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 33.48 20.616 34.68 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 34.44 15.128 35.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 34.44 15.216 35.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 34.44 21.516 35.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 34.44 21.728 35.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 2.28 21.516 3.48 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 35.4 13.888 36.6 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 35.4 13.972 36.6 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 35.4 20.528 36.6 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 35.4 20.616 36.6 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 36.36 15.128 37.56 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 36.36 15.216 37.56 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 36.36 21.516 37.56 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 36.36 21.728 37.56 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 37.32 13.888 38.52 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 37.32 13.972 38.52 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.24 13.716 4.44 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 37.32 20.528 38.52 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 37.32 20.616 38.52 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 38.28 15.128 39.48 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 38.28 15.216 39.48 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 38.28 21.516 39.48 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 38.28 21.728 39.48 ;
    END
  END rddatap0[135]
  PIN rddatap0[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 39.24 13.888 40.44 ;
    END
  END rddatap0[136]
  PIN rddatap0[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 39.24 13.972 40.44 ;
    END
  END rddatap0[137]
  PIN rddatap0[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 39.24 20.528 40.44 ;
    END
  END rddatap0[138]
  PIN rddatap0[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 39.24 20.616 40.44 ;
    END
  END rddatap0[139]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 3.24 13.888 4.44 ;
    END
  END rddatap0[13]
  PIN rddatap0[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 40.2 15.128 41.4 ;
    END
  END rddatap0[140]
  PIN rddatap0[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 40.2 15.216 41.4 ;
    END
  END rddatap0[141]
  PIN rddatap0[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 40.2 21.516 41.4 ;
    END
  END rddatap0[142]
  PIN rddatap0[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 40.2 21.728 41.4 ;
    END
  END rddatap0[143]
  PIN rddatap0[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 41.16 13.888 42.36 ;
    END
  END rddatap0[144]
  PIN rddatap0[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 41.16 13.972 42.36 ;
    END
  END rddatap0[145]
  PIN rddatap0[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 41.16 20.528 42.36 ;
    END
  END rddatap0[146]
  PIN rddatap0[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 41.16 20.616 42.36 ;
    END
  END rddatap0[147]
  PIN rddatap0[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 42.12 15.128 43.32 ;
    END
  END rddatap0[148]
  PIN rddatap0[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 42.12 15.216 43.32 ;
    END
  END rddatap0[149]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 3.24 20.272 4.44 ;
    END
  END rddatap0[14]
  PIN rddatap0[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 42.12 21.516 43.32 ;
    END
  END rddatap0[150]
  PIN rddatap0[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 42.12 21.728 43.32 ;
    END
  END rddatap0[151]
  PIN rddatap0[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 43.08 13.888 44.28 ;
    END
  END rddatap0[152]
  PIN rddatap0[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 43.08 13.972 44.28 ;
    END
  END rddatap0[153]
  PIN rddatap0[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 43.08 20.528 44.28 ;
    END
  END rddatap0[154]
  PIN rddatap0[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 43.08 20.616 44.28 ;
    END
  END rddatap0[155]
  PIN rddatap0[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 44.04 15.128 45.24 ;
    END
  END rddatap0[156]
  PIN rddatap0[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 44.04 15.216 45.24 ;
    END
  END rddatap0[157]
  PIN rddatap0[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 44.04 21.516 45.24 ;
    END
  END rddatap0[158]
  PIN rddatap0[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 44.04 21.728 45.24 ;
    END
  END rddatap0[159]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 3.24 20.356 4.44 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 4.2 14.956 5.4 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 4.2 15.128 5.4 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 4.2 21.428 5.4 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 4.2 21.516 5.4 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.36 13.716 1.56 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 5.16 13.716 6.36 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 5.16 13.888 6.36 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 5.16 20.272 6.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 5.16 20.356 6.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 6.12 14.956 7.32 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 6.12 15.128 7.32 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 6.12 21.428 7.32 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 6.12 21.516 7.32 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 7.08 13.716 8.28 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 7.08 13.888 8.28 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 0.36 21.428 1.56 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 7.08 20.272 8.28 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 7.08 20.356 8.28 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 8.04 14.956 9.24 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 8.04 15.128 9.24 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 8.04 21.428 9.24 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 8.04 21.516 9.24 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 9 13.716 10.2 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 9 13.888 10.2 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 9 20.272 10.2 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 9 20.356 10.2 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 0.36 21.516 1.56 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 9.96 14.956 11.16 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 9.96 15.128 11.16 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 9.96 21.428 11.16 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 9.96 21.516 11.16 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 10.92 13.716 12.12 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 10.92 13.888 12.12 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 10.92 20.272 12.12 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 10.92 20.356 12.12 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 11.88 14.956 13.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 11.88 15.128 13.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 1.32 14.228 2.52 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 11.88 21.428 13.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 11.88 21.516 13.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 12.84 13.716 14.04 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 12.84 13.888 14.04 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 12.84 20.272 14.04 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 12.84 20.356 14.04 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 13.8 14.956 15 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 13.8 15.128 15 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 13.8 21.428 15 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 13.8 21.516 15 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 1.32 14.316 2.52 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 14.76 13.716 15.96 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 14.76 13.888 15.96 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 14.76 20.272 15.96 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 14.76 20.356 15.96 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 15.72 14.956 16.92 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 15.72 15.128 16.92 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 15.72 21.428 16.92 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 15.72 21.516 16.92 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 16.68 13.716 17.88 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 16.68 13.888 17.88 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 1.32 20.272 2.52 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 16.68 20.272 17.88 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 16.68 20.356 17.88 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 17.64 14.956 18.84 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 17.64 15.128 18.84 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 17.64 21.428 18.84 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 17.64 21.516 18.84 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 18.6 13.716 19.8 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 18.6 13.888 19.8 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 18.6 20.272 19.8 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 18.6 20.356 19.8 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 1.32 20.356 2.52 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 25.8 13.888 27 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 25.8 13.972 27 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 25.8 20.528 27 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 25.8 20.616 27 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 26.76 15.128 27.96 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 26.76 15.216 27.96 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 26.76 21.516 27.96 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 26.76 21.728 27.96 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 27.72 13.888 28.92 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 27.72 13.972 28.92 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 2.28 14.956 3.48 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 27.72 20.528 28.92 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 27.72 20.616 28.92 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 28.68 15.128 29.88 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 28.68 15.216 29.88 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 28.68 21.516 29.88 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 28.68 21.728 29.88 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 29.64 13.888 30.84 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 29.64 13.972 30.84 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 29.64 20.528 30.84 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 29.64 20.616 30.84 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 2.28 15.128 3.48 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 0.36 13.888 1.56 ;
    END
  END rddatap1[0]
  PIN rddatap1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 30.6 15.428 31.8 ;
    END
  END rddatap1[100]
  PIN rddatap1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 30.6 15.516 31.8 ;
    END
  END rddatap1[101]
  PIN rddatap1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 30.6 21.816 31.8 ;
    END
  END rddatap1[102]
  PIN rddatap1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 30.6 20.016 31.8 ;
    END
  END rddatap1[103]
  PIN rddatap1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 31.56 14.056 32.76 ;
    END
  END rddatap1[104]
  PIN rddatap1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 31.56 14.228 32.76 ;
    END
  END rddatap1[105]
  PIN rddatap1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 31.56 20.828 32.76 ;
    END
  END rddatap1[106]
  PIN rddatap1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 31.56 20.916 32.76 ;
    END
  END rddatap1[107]
  PIN rddatap1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 32.52 15.428 33.72 ;
    END
  END rddatap1[108]
  PIN rddatap1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 32.52 15.516 33.72 ;
    END
  END rddatap1[109]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 2.28 21.728 3.48 ;
    END
  END rddatap1[10]
  PIN rddatap1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 32.52 21.816 33.72 ;
    END
  END rddatap1[110]
  PIN rddatap1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 32.52 20.016 33.72 ;
    END
  END rddatap1[111]
  PIN rddatap1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 33.48 14.056 34.68 ;
    END
  END rddatap1[112]
  PIN rddatap1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 33.48 14.228 34.68 ;
    END
  END rddatap1[113]
  PIN rddatap1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 33.48 20.828 34.68 ;
    END
  END rddatap1[114]
  PIN rddatap1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 33.48 20.916 34.68 ;
    END
  END rddatap1[115]
  PIN rddatap1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 34.44 15.428 35.64 ;
    END
  END rddatap1[116]
  PIN rddatap1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 34.44 15.516 35.64 ;
    END
  END rddatap1[117]
  PIN rddatap1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 34.44 21.816 35.64 ;
    END
  END rddatap1[118]
  PIN rddatap1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 34.44 20.016 35.64 ;
    END
  END rddatap1[119]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.28 21.816 3.48 ;
    END
  END rddatap1[11]
  PIN rddatap1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 35.4 14.056 36.6 ;
    END
  END rddatap1[120]
  PIN rddatap1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 35.4 14.228 36.6 ;
    END
  END rddatap1[121]
  PIN rddatap1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 35.4 20.828 36.6 ;
    END
  END rddatap1[122]
  PIN rddatap1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 35.4 20.916 36.6 ;
    END
  END rddatap1[123]
  PIN rddatap1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 36.36 15.428 37.56 ;
    END
  END rddatap1[124]
  PIN rddatap1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 36.36 15.516 37.56 ;
    END
  END rddatap1[125]
  PIN rddatap1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 36.36 21.816 37.56 ;
    END
  END rddatap1[126]
  PIN rddatap1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 36.36 20.016 37.56 ;
    END
  END rddatap1[127]
  PIN rddatap1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 37.32 14.056 38.52 ;
    END
  END rddatap1[128]
  PIN rddatap1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 37.32 14.228 38.52 ;
    END
  END rddatap1[129]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.24 13.972 4.44 ;
    END
  END rddatap1[12]
  PIN rddatap1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 37.32 20.828 38.52 ;
    END
  END rddatap1[130]
  PIN rddatap1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 37.32 20.916 38.52 ;
    END
  END rddatap1[131]
  PIN rddatap1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 38.28 15.428 39.48 ;
    END
  END rddatap1[132]
  PIN rddatap1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 38.28 15.516 39.48 ;
    END
  END rddatap1[133]
  PIN rddatap1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 38.28 21.816 39.48 ;
    END
  END rddatap1[134]
  PIN rddatap1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 38.28 20.016 39.48 ;
    END
  END rddatap1[135]
  PIN rddatap1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 39.24 14.056 40.44 ;
    END
  END rddatap1[136]
  PIN rddatap1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 39.24 14.228 40.44 ;
    END
  END rddatap1[137]
  PIN rddatap1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 39.24 20.828 40.44 ;
    END
  END rddatap1[138]
  PIN rddatap1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 39.24 20.916 40.44 ;
    END
  END rddatap1[139]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 3.24 14.056 4.44 ;
    END
  END rddatap1[13]
  PIN rddatap1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 40.2 15.428 41.4 ;
    END
  END rddatap1[140]
  PIN rddatap1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 40.2 15.516 41.4 ;
    END
  END rddatap1[141]
  PIN rddatap1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 40.2 21.816 41.4 ;
    END
  END rddatap1[142]
  PIN rddatap1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 40.2 20.016 41.4 ;
    END
  END rddatap1[143]
  PIN rddatap1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 41.16 14.056 42.36 ;
    END
  END rddatap1[144]
  PIN rddatap1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 41.16 14.228 42.36 ;
    END
  END rddatap1[145]
  PIN rddatap1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 41.16 20.828 42.36 ;
    END
  END rddatap1[146]
  PIN rddatap1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 41.16 20.916 42.36 ;
    END
  END rddatap1[147]
  PIN rddatap1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 42.12 15.428 43.32 ;
    END
  END rddatap1[148]
  PIN rddatap1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 42.12 15.516 43.32 ;
    END
  END rddatap1[149]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 3.24 20.528 4.44 ;
    END
  END rddatap1[14]
  PIN rddatap1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 42.12 21.816 43.32 ;
    END
  END rddatap1[150]
  PIN rddatap1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 42.12 20.016 43.32 ;
    END
  END rddatap1[151]
  PIN rddatap1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 43.08 14.056 44.28 ;
    END
  END rddatap1[152]
  PIN rddatap1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 43.08 14.228 44.28 ;
    END
  END rddatap1[153]
  PIN rddatap1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 43.08 20.828 44.28 ;
    END
  END rddatap1[154]
  PIN rddatap1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 43.08 20.916 44.28 ;
    END
  END rddatap1[155]
  PIN rddatap1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 44.04 15.428 45.24 ;
    END
  END rddatap1[156]
  PIN rddatap1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 44.04 15.516 45.24 ;
    END
  END rddatap1[157]
  PIN rddatap1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 44.04 21.816 45.24 ;
    END
  END rddatap1[158]
  PIN rddatap1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 44.04 20.016 45.24 ;
    END
  END rddatap1[159]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 3.24 20.616 4.44 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 4.2 15.216 5.4 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.2 15.428 5.4 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 4.2 21.728 5.4 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 4.2 21.816 5.4 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.36 13.972 1.56 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 5.16 13.972 6.36 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 5.16 14.056 6.36 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 5.16 20.528 6.36 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 5.16 20.616 6.36 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 6.12 15.216 7.32 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6.12 15.428 7.32 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 6.12 21.728 7.32 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 6.12 21.816 7.32 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 7.08 13.972 8.28 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 7.08 14.056 8.28 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 0.36 21.728 1.56 ;
    END
  END rddatap1[2]
  PIN rddatap1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 7.08 20.528 8.28 ;
    END
  END rddatap1[30]
  PIN rddatap1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 7.08 20.616 8.28 ;
    END
  END rddatap1[31]
  PIN rddatap1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 8.04 15.216 9.24 ;
    END
  END rddatap1[32]
  PIN rddatap1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.04 15.428 9.24 ;
    END
  END rddatap1[33]
  PIN rddatap1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 8.04 21.728 9.24 ;
    END
  END rddatap1[34]
  PIN rddatap1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 8.04 21.816 9.24 ;
    END
  END rddatap1[35]
  PIN rddatap1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 9 13.972 10.2 ;
    END
  END rddatap1[36]
  PIN rddatap1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 9 14.056 10.2 ;
    END
  END rddatap1[37]
  PIN rddatap1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 9 20.528 10.2 ;
    END
  END rddatap1[38]
  PIN rddatap1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 9 20.616 10.2 ;
    END
  END rddatap1[39]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 0.36 21.816 1.56 ;
    END
  END rddatap1[3]
  PIN rddatap1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 9.96 15.216 11.16 ;
    END
  END rddatap1[40]
  PIN rddatap1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 9.96 15.428 11.16 ;
    END
  END rddatap1[41]
  PIN rddatap1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 9.96 21.728 11.16 ;
    END
  END rddatap1[42]
  PIN rddatap1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 9.96 21.816 11.16 ;
    END
  END rddatap1[43]
  PIN rddatap1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 10.92 13.972 12.12 ;
    END
  END rddatap1[44]
  PIN rddatap1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 10.92 14.056 12.12 ;
    END
  END rddatap1[45]
  PIN rddatap1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 10.92 20.528 12.12 ;
    END
  END rddatap1[46]
  PIN rddatap1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 10.92 20.616 12.12 ;
    END
  END rddatap1[47]
  PIN rddatap1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 11.88 15.216 13.08 ;
    END
  END rddatap1[48]
  PIN rddatap1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 11.88 15.428 13.08 ;
    END
  END rddatap1[49]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 1.32 14.528 2.52 ;
    END
  END rddatap1[4]
  PIN rddatap1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 11.88 21.728 13.08 ;
    END
  END rddatap1[50]
  PIN rddatap1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 11.88 21.816 13.08 ;
    END
  END rddatap1[51]
  PIN rddatap1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 12.84 13.972 14.04 ;
    END
  END rddatap1[52]
  PIN rddatap1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 12.84 14.056 14.04 ;
    END
  END rddatap1[53]
  PIN rddatap1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 12.84 20.528 14.04 ;
    END
  END rddatap1[54]
  PIN rddatap1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 12.84 20.616 14.04 ;
    END
  END rddatap1[55]
  PIN rddatap1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 13.8 15.216 15 ;
    END
  END rddatap1[56]
  PIN rddatap1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 13.8 15.428 15 ;
    END
  END rddatap1[57]
  PIN rddatap1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 13.8 21.728 15 ;
    END
  END rddatap1[58]
  PIN rddatap1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 13.8 21.816 15 ;
    END
  END rddatap1[59]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 1.32 14.616 2.52 ;
    END
  END rddatap1[5]
  PIN rddatap1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 14.76 13.972 15.96 ;
    END
  END rddatap1[60]
  PIN rddatap1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 14.76 14.056 15.96 ;
    END
  END rddatap1[61]
  PIN rddatap1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 14.76 20.528 15.96 ;
    END
  END rddatap1[62]
  PIN rddatap1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 14.76 20.616 15.96 ;
    END
  END rddatap1[63]
  PIN rddatap1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 15.72 15.216 16.92 ;
    END
  END rddatap1[64]
  PIN rddatap1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 15.72 15.428 16.92 ;
    END
  END rddatap1[65]
  PIN rddatap1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 15.72 21.728 16.92 ;
    END
  END rddatap1[66]
  PIN rddatap1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 15.72 21.816 16.92 ;
    END
  END rddatap1[67]
  PIN rddatap1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 16.68 13.972 17.88 ;
    END
  END rddatap1[68]
  PIN rddatap1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 16.68 14.056 17.88 ;
    END
  END rddatap1[69]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 1.32 20.528 2.52 ;
    END
  END rddatap1[6]
  PIN rddatap1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 16.68 20.528 17.88 ;
    END
  END rddatap1[70]
  PIN rddatap1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 16.68 20.616 17.88 ;
    END
  END rddatap1[71]
  PIN rddatap1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 17.64 15.216 18.84 ;
    END
  END rddatap1[72]
  PIN rddatap1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 17.64 15.428 18.84 ;
    END
  END rddatap1[73]
  PIN rddatap1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 17.64 21.728 18.84 ;
    END
  END rddatap1[74]
  PIN rddatap1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 17.64 21.816 18.84 ;
    END
  END rddatap1[75]
  PIN rddatap1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 18.6 13.972 19.8 ;
    END
  END rddatap1[76]
  PIN rddatap1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 18.6 14.056 19.8 ;
    END
  END rddatap1[77]
  PIN rddatap1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 18.6 20.528 19.8 ;
    END
  END rddatap1[78]
  PIN rddatap1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 18.6 20.616 19.8 ;
    END
  END rddatap1[79]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.32 20.616 2.52 ;
    END
  END rddatap1[7]
  PIN rddatap1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 25.8 14.056 27 ;
    END
  END rddatap1[80]
  PIN rddatap1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 25.8 14.228 27 ;
    END
  END rddatap1[81]
  PIN rddatap1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 25.8 20.916 27 ;
    END
  END rddatap1[82]
  PIN rddatap1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 25.8 21.172 27 ;
    END
  END rddatap1[83]
  PIN rddatap1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 26.76 15.428 27.96 ;
    END
  END rddatap1[84]
  PIN rddatap1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 26.76 15.516 27.96 ;
    END
  END rddatap1[85]
  PIN rddatap1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 26.76 21.816 27.96 ;
    END
  END rddatap1[86]
  PIN rddatap1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 26.76 20.016 27.96 ;
    END
  END rddatap1[87]
  PIN rddatap1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 27.72 14.056 28.92 ;
    END
  END rddatap1[88]
  PIN rddatap1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 27.72 14.228 28.92 ;
    END
  END rddatap1[89]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 2.28 15.216 3.48 ;
    END
  END rddatap1[8]
  PIN rddatap1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 27.72 20.828 28.92 ;
    END
  END rddatap1[90]
  PIN rddatap1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 27.72 20.916 28.92 ;
    END
  END rddatap1[91]
  PIN rddatap1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 28.68 15.428 29.88 ;
    END
  END rddatap1[92]
  PIN rddatap1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 28.68 15.516 29.88 ;
    END
  END rddatap1[93]
  PIN rddatap1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 28.68 21.816 29.88 ;
    END
  END rddatap1[94]
  PIN rddatap1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 28.68 20.016 29.88 ;
    END
  END rddatap1[95]
  PIN rddatap1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 29.64 14.056 30.84 ;
    END
  END rddatap1[96]
  PIN rddatap1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 29.64 14.228 30.84 ;
    END
  END rddatap1[97]
  PIN rddatap1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 29.64 20.828 30.84 ;
    END
  END rddatap1[98]
  PIN rddatap1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 29.64 20.916 30.84 ;
    END
  END rddatap1[99]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 2.28 15.428 3.48 ;
    END
  END rddatap1[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 46.02 ;
        RECT 2.662 0.06 2.738 46.02 ;
        RECT 4.462 0.06 4.538 46.02 ;
        RECT 6.262 0.06 6.338 46.02 ;
        RECT 8.062 0.06 8.138 46.02 ;
        RECT 9.862 0.06 9.938 46.02 ;
        RECT 11.662 0.06 11.738 46.02 ;
        RECT 13.462 0.06 13.538 46.02 ;
        RECT 15.262 0.06 15.338 46.02 ;
        RECT 17.062 0.06 17.138 46.02 ;
        RECT 18.862 0.06 18.938 46.02 ;
        RECT 20.662 0.06 20.738 46.02 ;
        RECT 22.462 0.06 22.538 46.02 ;
        RECT 24.262 0.06 24.338 46.02 ;
        RECT 26.062 0.06 26.138 46.02 ;
        RECT 27.862 0.06 27.938 46.02 ;
        RECT 29.662 0.06 29.738 46.02 ;
        RECT 31.462 0.06 31.538 46.02 ;
        RECT 33.262 0.06 33.338 46.02 ;
        RECT 35.062 0.06 35.138 46.02 ;
        RECT 36.862 0.06 36.938 46.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 46.02 ;
        RECT 3.562 0.06 3.638 46.02 ;
        RECT 5.362 0.06 5.438 46.02 ;
        RECT 7.162 0.06 7.238 46.02 ;
        RECT 8.962 0.06 9.038 46.02 ;
        RECT 10.762 0.06 10.838 46.02 ;
        RECT 12.562 0.06 12.638 46.02 ;
        RECT 14.362 0.06 14.438 46.02 ;
        RECT 16.162 0.06 16.238 46.02 ;
        RECT 17.962 0.06 18.038 46.02 ;
        RECT 19.762 0.06 19.838 46.02 ;
        RECT 21.562 0.06 21.638 46.02 ;
        RECT 23.362 0.06 23.438 46.02 ;
        RECT 25.162 0.06 25.238 46.02 ;
        RECT 26.962 0.06 27.038 46.02 ;
        RECT 28.762 0.06 28.838 46.02 ;
        RECT 30.562 0.06 30.638 46.02 ;
        RECT 32.362 0.06 32.438 46.02 ;
        RECT 34.162 0.06 34.238 46.02 ;
        RECT 35.962 0.06 36.038 46.02 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 37.816 46.094 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 37.82 46.1 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 37.8705 46.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 37.835 46.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 37.87 46.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 37.859 46.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 37.89 46.142 ;
    LAYER m7 SPACING 0 ;
      RECT 36.938 46.14 37.84 46.2 ;
      RECT 36.938 -0.06 37.892 46.14 ;
      RECT 36.938 -0.12 37.84 -0.06 ;
      RECT 36.038 -0.12 36.862 46.2 ;
      RECT 35.138 -0.12 35.962 46.2 ;
      RECT 34.238 -0.12 35.062 46.2 ;
      RECT 33.338 -0.12 34.162 46.2 ;
      RECT 32.438 -0.12 33.262 46.2 ;
      RECT 31.538 -0.12 32.362 46.2 ;
      RECT 30.638 -0.12 31.462 46.2 ;
      RECT 29.738 -0.12 30.562 46.2 ;
      RECT 28.838 -0.12 29.662 46.2 ;
      RECT 27.938 -0.12 28.762 46.2 ;
      RECT 27.038 -0.12 27.862 46.2 ;
      RECT 26.138 -0.12 26.962 46.2 ;
      RECT 25.238 -0.12 26.062 46.2 ;
      RECT 24.338 -0.12 25.162 46.2 ;
      RECT 23.438 -0.12 24.262 46.2 ;
      RECT 22.538 -0.12 23.362 46.2 ;
      RECT 21.638 45.24 22.462 46.2 ;
      RECT 21.638 44.04 21.684 45.24 ;
      RECT 21.728 44.04 21.772 45.24 ;
      RECT 21.816 44.04 22.462 45.24 ;
      RECT 21.638 43.32 22.462 44.04 ;
      RECT 21.638 42.12 21.684 43.32 ;
      RECT 21.728 42.12 21.772 43.32 ;
      RECT 21.816 42.12 22.462 43.32 ;
      RECT 21.638 41.4 22.462 42.12 ;
      RECT 21.638 40.2 21.684 41.4 ;
      RECT 21.728 40.2 21.772 41.4 ;
      RECT 21.816 40.2 22.462 41.4 ;
      RECT 21.638 39.48 22.462 40.2 ;
      RECT 21.638 38.28 21.684 39.48 ;
      RECT 21.728 38.28 21.772 39.48 ;
      RECT 21.816 38.28 22.462 39.48 ;
      RECT 21.638 37.56 22.462 38.28 ;
      RECT 21.638 36.36 21.684 37.56 ;
      RECT 21.728 36.36 21.772 37.56 ;
      RECT 21.816 36.36 22.462 37.56 ;
      RECT 21.638 35.64 22.462 36.36 ;
      RECT 21.638 34.44 21.684 35.64 ;
      RECT 21.728 34.44 21.772 35.64 ;
      RECT 21.816 34.44 22.462 35.64 ;
      RECT 21.638 33.72 22.462 34.44 ;
      RECT 21.638 32.52 21.684 33.72 ;
      RECT 21.728 32.52 21.772 33.72 ;
      RECT 21.816 32.52 22.462 33.72 ;
      RECT 21.638 31.8 22.462 32.52 ;
      RECT 21.638 30.6 21.684 31.8 ;
      RECT 21.728 30.6 21.772 31.8 ;
      RECT 21.816 30.6 22.462 31.8 ;
      RECT 21.638 29.88 22.462 30.6 ;
      RECT 21.638 28.68 21.684 29.88 ;
      RECT 21.728 28.68 21.772 29.88 ;
      RECT 21.816 28.68 22.462 29.88 ;
      RECT 21.638 27.96 22.462 28.68 ;
      RECT 21.638 26.76 21.684 27.96 ;
      RECT 21.728 26.76 21.772 27.96 ;
      RECT 21.816 26.76 22.462 27.96 ;
      RECT 21.638 18.84 22.462 26.76 ;
      RECT 21.638 17.64 21.684 18.84 ;
      RECT 21.728 17.64 21.772 18.84 ;
      RECT 21.816 17.64 22.462 18.84 ;
      RECT 21.638 16.92 22.462 17.64 ;
      RECT 21.638 15.72 21.684 16.92 ;
      RECT 21.728 15.72 21.772 16.92 ;
      RECT 21.816 15.72 22.462 16.92 ;
      RECT 21.638 15 22.462 15.72 ;
      RECT 21.638 13.8 21.684 15 ;
      RECT 21.728 13.8 21.772 15 ;
      RECT 21.816 13.8 22.462 15 ;
      RECT 21.638 13.08 22.462 13.8 ;
      RECT 21.638 11.88 21.684 13.08 ;
      RECT 21.728 11.88 21.772 13.08 ;
      RECT 21.816 11.88 22.462 13.08 ;
      RECT 21.638 11.16 22.462 11.88 ;
      RECT 21.638 9.96 21.684 11.16 ;
      RECT 21.728 9.96 21.772 11.16 ;
      RECT 21.816 9.96 22.462 11.16 ;
      RECT 21.638 9.24 22.462 9.96 ;
      RECT 21.638 8.04 21.684 9.24 ;
      RECT 21.728 8.04 21.772 9.24 ;
      RECT 21.816 8.04 22.462 9.24 ;
      RECT 21.638 7.32 22.462 8.04 ;
      RECT 21.638 6.12 21.684 7.32 ;
      RECT 21.728 6.12 21.772 7.32 ;
      RECT 21.816 6.12 22.462 7.32 ;
      RECT 21.638 5.4 22.462 6.12 ;
      RECT 21.638 4.2 21.684 5.4 ;
      RECT 21.728 4.2 21.772 5.4 ;
      RECT 21.816 4.2 22.462 5.4 ;
      RECT 21.638 3.48 22.462 4.2 ;
      RECT 21.638 2.28 21.684 3.48 ;
      RECT 21.728 2.28 21.772 3.48 ;
      RECT 21.816 2.28 22.462 3.48 ;
      RECT 21.638 1.56 22.462 2.28 ;
      RECT 21.638 0.36 21.684 1.56 ;
      RECT 21.728 0.36 21.772 1.56 ;
      RECT 21.816 0.36 22.462 1.56 ;
      RECT 21.638 -0.12 22.462 0.36 ;
      RECT 20.738 45.24 21.562 46.2 ;
      RECT 20.738 44.28 21.472 45.24 ;
      RECT 21.516 44.04 21.562 45.24 ;
      RECT 20.916 44.04 21.472 44.28 ;
      RECT 20.916 43.32 21.562 44.04 ;
      RECT 20.738 43.08 20.784 44.28 ;
      RECT 20.828 43.08 20.872 44.28 ;
      RECT 20.916 43.08 21.472 43.32 ;
      RECT 20.738 42.36 21.472 43.08 ;
      RECT 21.516 42.12 21.562 43.32 ;
      RECT 20.916 42.12 21.472 42.36 ;
      RECT 20.916 41.4 21.562 42.12 ;
      RECT 20.738 41.16 20.784 42.36 ;
      RECT 20.828 41.16 20.872 42.36 ;
      RECT 20.916 41.16 21.472 41.4 ;
      RECT 20.738 40.44 21.472 41.16 ;
      RECT 21.516 40.2 21.562 41.4 ;
      RECT 20.916 40.2 21.472 40.44 ;
      RECT 20.916 39.48 21.562 40.2 ;
      RECT 20.738 39.24 20.784 40.44 ;
      RECT 20.828 39.24 20.872 40.44 ;
      RECT 20.916 39.24 21.472 39.48 ;
      RECT 20.738 38.52 21.472 39.24 ;
      RECT 21.516 38.28 21.562 39.48 ;
      RECT 20.916 38.28 21.472 38.52 ;
      RECT 20.916 37.56 21.562 38.28 ;
      RECT 20.738 37.32 20.784 38.52 ;
      RECT 20.828 37.32 20.872 38.52 ;
      RECT 20.916 37.32 21.472 37.56 ;
      RECT 20.738 36.6 21.472 37.32 ;
      RECT 21.516 36.36 21.562 37.56 ;
      RECT 20.916 36.36 21.472 36.6 ;
      RECT 20.916 35.64 21.562 36.36 ;
      RECT 20.738 35.4 20.784 36.6 ;
      RECT 20.828 35.4 20.872 36.6 ;
      RECT 20.916 35.4 21.472 35.64 ;
      RECT 20.738 34.68 21.472 35.4 ;
      RECT 21.516 34.44 21.562 35.64 ;
      RECT 20.916 34.44 21.472 34.68 ;
      RECT 20.916 33.72 21.562 34.44 ;
      RECT 20.738 33.48 20.784 34.68 ;
      RECT 20.828 33.48 20.872 34.68 ;
      RECT 20.916 33.48 21.472 33.72 ;
      RECT 20.738 32.76 21.472 33.48 ;
      RECT 21.516 32.52 21.562 33.72 ;
      RECT 20.916 32.52 21.472 32.76 ;
      RECT 20.916 31.8 21.562 32.52 ;
      RECT 20.738 31.56 20.784 32.76 ;
      RECT 20.828 31.56 20.872 32.76 ;
      RECT 20.916 31.56 21.472 31.8 ;
      RECT 20.738 30.84 21.472 31.56 ;
      RECT 21.516 30.6 21.562 31.8 ;
      RECT 20.916 30.6 21.472 30.84 ;
      RECT 20.916 29.88 21.562 30.6 ;
      RECT 20.738 29.64 20.784 30.84 ;
      RECT 20.828 29.64 20.872 30.84 ;
      RECT 20.916 29.64 21.472 29.88 ;
      RECT 20.738 28.92 21.472 29.64 ;
      RECT 21.516 28.68 21.562 29.88 ;
      RECT 20.916 28.68 21.472 28.92 ;
      RECT 20.916 27.96 21.562 28.68 ;
      RECT 20.738 27.72 20.784 28.92 ;
      RECT 20.828 27.72 20.872 28.92 ;
      RECT 20.916 27.72 21.472 27.96 ;
      RECT 20.738 27 21.472 27.72 ;
      RECT 21.516 26.76 21.562 27.96 ;
      RECT 21.172 26.76 21.472 27 ;
      RECT 20.738 25.8 20.872 27 ;
      RECT 20.916 25.8 21.128 27 ;
      RECT 21.172 25.8 21.562 26.76 ;
      RECT 20.738 24.84 21.562 25.8 ;
      RECT 20.738 23.64 20.784 24.84 ;
      RECT 20.828 23.64 21.044 24.84 ;
      RECT 21.088 23.64 21.562 24.84 ;
      RECT 20.738 21.96 21.562 23.64 ;
      RECT 20.738 20.76 20.784 21.96 ;
      RECT 20.828 20.76 21.044 21.96 ;
      RECT 21.088 20.76 21.212 21.96 ;
      RECT 21.256 20.76 21.472 21.96 ;
      RECT 21.516 20.76 21.562 21.96 ;
      RECT 20.738 18.84 21.562 20.76 ;
      RECT 20.738 17.64 21.384 18.84 ;
      RECT 21.428 17.64 21.472 18.84 ;
      RECT 21.516 17.64 21.562 18.84 ;
      RECT 20.738 16.92 21.562 17.64 ;
      RECT 20.738 15.72 21.384 16.92 ;
      RECT 21.428 15.72 21.472 16.92 ;
      RECT 21.516 15.72 21.562 16.92 ;
      RECT 20.738 15 21.562 15.72 ;
      RECT 20.738 13.8 21.384 15 ;
      RECT 21.428 13.8 21.472 15 ;
      RECT 21.516 13.8 21.562 15 ;
      RECT 20.738 13.08 21.562 13.8 ;
      RECT 20.738 11.88 21.384 13.08 ;
      RECT 21.428 11.88 21.472 13.08 ;
      RECT 21.516 11.88 21.562 13.08 ;
      RECT 20.738 11.16 21.562 11.88 ;
      RECT 20.738 9.96 21.384 11.16 ;
      RECT 21.428 9.96 21.472 11.16 ;
      RECT 21.516 9.96 21.562 11.16 ;
      RECT 20.738 9.24 21.562 9.96 ;
      RECT 20.738 8.04 21.384 9.24 ;
      RECT 21.428 8.04 21.472 9.24 ;
      RECT 21.516 8.04 21.562 9.24 ;
      RECT 20.738 7.32 21.562 8.04 ;
      RECT 20.738 6.12 21.384 7.32 ;
      RECT 21.428 6.12 21.472 7.32 ;
      RECT 21.516 6.12 21.562 7.32 ;
      RECT 20.738 5.4 21.562 6.12 ;
      RECT 20.738 4.2 21.384 5.4 ;
      RECT 21.428 4.2 21.472 5.4 ;
      RECT 21.516 4.2 21.562 5.4 ;
      RECT 20.738 3.48 21.562 4.2 ;
      RECT 20.738 2.28 21.384 3.48 ;
      RECT 21.428 2.28 21.472 3.48 ;
      RECT 21.516 2.28 21.562 3.48 ;
      RECT 20.738 1.56 21.562 2.28 ;
      RECT 20.738 0.36 21.384 1.56 ;
      RECT 21.428 0.36 21.472 1.56 ;
      RECT 21.516 0.36 21.562 1.56 ;
      RECT 20.738 -0.12 21.562 0.36 ;
      RECT 19.838 45.24 20.662 46.2 ;
      RECT 20.016 44.28 20.662 45.24 ;
      RECT 19.838 44.04 19.972 45.24 ;
      RECT 20.016 44.04 20.484 44.28 ;
      RECT 19.838 43.32 20.484 44.04 ;
      RECT 20.528 43.08 20.572 44.28 ;
      RECT 20.616 43.08 20.662 44.28 ;
      RECT 20.016 43.08 20.484 43.32 ;
      RECT 20.016 42.36 20.662 43.08 ;
      RECT 19.838 42.12 19.972 43.32 ;
      RECT 20.016 42.12 20.484 42.36 ;
      RECT 19.838 41.4 20.484 42.12 ;
      RECT 20.528 41.16 20.572 42.36 ;
      RECT 20.616 41.16 20.662 42.36 ;
      RECT 20.016 41.16 20.484 41.4 ;
      RECT 20.016 40.44 20.662 41.16 ;
      RECT 19.838 40.2 19.972 41.4 ;
      RECT 20.016 40.2 20.484 40.44 ;
      RECT 19.838 39.48 20.484 40.2 ;
      RECT 20.528 39.24 20.572 40.44 ;
      RECT 20.616 39.24 20.662 40.44 ;
      RECT 20.016 39.24 20.484 39.48 ;
      RECT 20.016 38.52 20.662 39.24 ;
      RECT 19.838 38.28 19.972 39.48 ;
      RECT 20.016 38.28 20.484 38.52 ;
      RECT 19.838 37.56 20.484 38.28 ;
      RECT 20.528 37.32 20.572 38.52 ;
      RECT 20.616 37.32 20.662 38.52 ;
      RECT 20.016 37.32 20.484 37.56 ;
      RECT 20.016 36.6 20.662 37.32 ;
      RECT 19.838 36.36 19.972 37.56 ;
      RECT 20.016 36.36 20.484 36.6 ;
      RECT 19.838 35.64 20.484 36.36 ;
      RECT 20.528 35.4 20.572 36.6 ;
      RECT 20.616 35.4 20.662 36.6 ;
      RECT 20.016 35.4 20.484 35.64 ;
      RECT 20.016 34.68 20.662 35.4 ;
      RECT 19.838 34.44 19.972 35.64 ;
      RECT 20.016 34.44 20.484 34.68 ;
      RECT 19.838 33.72 20.484 34.44 ;
      RECT 20.528 33.48 20.572 34.68 ;
      RECT 20.616 33.48 20.662 34.68 ;
      RECT 20.016 33.48 20.484 33.72 ;
      RECT 20.016 32.76 20.662 33.48 ;
      RECT 19.838 32.52 19.972 33.72 ;
      RECT 20.016 32.52 20.484 32.76 ;
      RECT 19.838 31.8 20.484 32.52 ;
      RECT 20.528 31.56 20.572 32.76 ;
      RECT 20.616 31.56 20.662 32.76 ;
      RECT 20.016 31.56 20.484 31.8 ;
      RECT 20.016 30.84 20.662 31.56 ;
      RECT 19.838 30.6 19.972 31.8 ;
      RECT 20.016 30.6 20.484 30.84 ;
      RECT 19.838 29.88 20.484 30.6 ;
      RECT 20.528 29.64 20.572 30.84 ;
      RECT 20.616 29.64 20.662 30.84 ;
      RECT 20.016 29.64 20.484 29.88 ;
      RECT 20.016 28.92 20.662 29.64 ;
      RECT 19.838 28.68 19.972 29.88 ;
      RECT 20.016 28.68 20.484 28.92 ;
      RECT 19.838 27.96 20.484 28.68 ;
      RECT 20.528 27.72 20.572 28.92 ;
      RECT 20.616 27.72 20.662 28.92 ;
      RECT 20.016 27.72 20.484 27.96 ;
      RECT 20.016 27 20.662 27.72 ;
      RECT 19.838 26.76 19.972 27.96 ;
      RECT 20.016 26.76 20.484 27 ;
      RECT 20.528 25.8 20.572 27 ;
      RECT 20.616 25.8 20.662 27 ;
      RECT 19.838 25.8 20.484 26.76 ;
      RECT 19.838 24.84 20.662 25.8 ;
      RECT 19.838 23.64 19.972 24.84 ;
      RECT 20.016 23.64 20.662 24.84 ;
      RECT 19.838 21.96 20.662 23.64 ;
      RECT 19.838 20.76 19.972 21.96 ;
      RECT 20.016 20.76 20.662 21.96 ;
      RECT 19.838 19.8 20.662 20.76 ;
      RECT 19.838 18.6 20.228 19.8 ;
      RECT 20.272 18.6 20.312 19.8 ;
      RECT 20.356 18.6 20.484 19.8 ;
      RECT 20.528 18.6 20.572 19.8 ;
      RECT 20.616 18.6 20.662 19.8 ;
      RECT 19.838 17.88 20.662 18.6 ;
      RECT 19.838 16.68 20.228 17.88 ;
      RECT 20.272 16.68 20.312 17.88 ;
      RECT 20.356 16.68 20.484 17.88 ;
      RECT 20.528 16.68 20.572 17.88 ;
      RECT 20.616 16.68 20.662 17.88 ;
      RECT 19.838 15.96 20.662 16.68 ;
      RECT 19.838 14.76 20.228 15.96 ;
      RECT 20.272 14.76 20.312 15.96 ;
      RECT 20.356 14.76 20.484 15.96 ;
      RECT 20.528 14.76 20.572 15.96 ;
      RECT 20.616 14.76 20.662 15.96 ;
      RECT 19.838 14.04 20.662 14.76 ;
      RECT 19.838 12.84 20.228 14.04 ;
      RECT 20.272 12.84 20.312 14.04 ;
      RECT 20.356 12.84 20.484 14.04 ;
      RECT 20.528 12.84 20.572 14.04 ;
      RECT 20.616 12.84 20.662 14.04 ;
      RECT 19.838 12.12 20.662 12.84 ;
      RECT 19.838 10.92 20.228 12.12 ;
      RECT 20.272 10.92 20.312 12.12 ;
      RECT 20.356 10.92 20.484 12.12 ;
      RECT 20.528 10.92 20.572 12.12 ;
      RECT 20.616 10.92 20.662 12.12 ;
      RECT 19.838 10.2 20.662 10.92 ;
      RECT 19.838 9 20.228 10.2 ;
      RECT 20.272 9 20.312 10.2 ;
      RECT 20.356 9 20.484 10.2 ;
      RECT 20.528 9 20.572 10.2 ;
      RECT 20.616 9 20.662 10.2 ;
      RECT 19.838 8.28 20.662 9 ;
      RECT 19.838 7.08 20.228 8.28 ;
      RECT 20.272 7.08 20.312 8.28 ;
      RECT 20.356 7.08 20.484 8.28 ;
      RECT 20.528 7.08 20.572 8.28 ;
      RECT 20.616 7.08 20.662 8.28 ;
      RECT 19.838 6.36 20.662 7.08 ;
      RECT 19.838 5.16 20.228 6.36 ;
      RECT 20.272 5.16 20.312 6.36 ;
      RECT 20.356 5.16 20.484 6.36 ;
      RECT 20.528 5.16 20.572 6.36 ;
      RECT 20.616 5.16 20.662 6.36 ;
      RECT 19.838 4.44 20.662 5.16 ;
      RECT 19.838 3.24 20.228 4.44 ;
      RECT 20.272 3.24 20.312 4.44 ;
      RECT 20.356 3.24 20.484 4.44 ;
      RECT 20.528 3.24 20.572 4.44 ;
      RECT 20.616 3.24 20.662 4.44 ;
      RECT 19.838 2.52 20.662 3.24 ;
      RECT 19.838 1.32 20.228 2.52 ;
      RECT 20.272 1.32 20.312 2.52 ;
      RECT 20.356 1.32 20.484 2.52 ;
      RECT 20.528 1.32 20.572 2.52 ;
      RECT 20.616 1.32 20.662 2.52 ;
      RECT 19.838 -0.12 20.662 1.32 ;
      RECT 18.938 45.24 19.762 46.2 ;
      RECT 19.288 44.28 19.762 45.24 ;
      RECT 18.938 44.04 18.984 45.24 ;
      RECT 19.028 44.04 19.072 45.24 ;
      RECT 19.116 44.04 19.244 45.24 ;
      RECT 19.288 44.04 19.584 44.28 ;
      RECT 18.938 43.32 19.584 44.04 ;
      RECT 19.628 43.08 19.762 44.28 ;
      RECT 19.288 43.08 19.584 43.32 ;
      RECT 19.288 42.36 19.762 43.08 ;
      RECT 18.938 42.12 18.984 43.32 ;
      RECT 19.028 42.12 19.072 43.32 ;
      RECT 19.116 42.12 19.244 43.32 ;
      RECT 19.288 42.12 19.584 42.36 ;
      RECT 18.938 41.4 19.584 42.12 ;
      RECT 19.628 41.16 19.762 42.36 ;
      RECT 19.288 41.16 19.584 41.4 ;
      RECT 19.288 40.44 19.762 41.16 ;
      RECT 18.938 40.2 18.984 41.4 ;
      RECT 19.028 40.2 19.072 41.4 ;
      RECT 19.116 40.2 19.244 41.4 ;
      RECT 19.288 40.2 19.584 40.44 ;
      RECT 18.938 39.48 19.584 40.2 ;
      RECT 19.628 39.24 19.762 40.44 ;
      RECT 19.288 39.24 19.584 39.48 ;
      RECT 19.288 38.52 19.762 39.24 ;
      RECT 18.938 38.28 18.984 39.48 ;
      RECT 19.028 38.28 19.072 39.48 ;
      RECT 19.116 38.28 19.244 39.48 ;
      RECT 19.288 38.28 19.584 38.52 ;
      RECT 18.938 37.56 19.584 38.28 ;
      RECT 19.628 37.32 19.762 38.52 ;
      RECT 19.288 37.32 19.584 37.56 ;
      RECT 19.288 36.6 19.762 37.32 ;
      RECT 18.938 36.36 18.984 37.56 ;
      RECT 19.028 36.36 19.072 37.56 ;
      RECT 19.116 36.36 19.244 37.56 ;
      RECT 19.288 36.36 19.584 36.6 ;
      RECT 18.938 35.64 19.584 36.36 ;
      RECT 19.628 35.4 19.762 36.6 ;
      RECT 19.288 35.4 19.584 35.64 ;
      RECT 19.288 34.68 19.762 35.4 ;
      RECT 18.938 34.44 18.984 35.64 ;
      RECT 19.028 34.44 19.072 35.64 ;
      RECT 19.116 34.44 19.244 35.64 ;
      RECT 19.288 34.44 19.584 34.68 ;
      RECT 18.938 33.72 19.584 34.44 ;
      RECT 19.628 33.48 19.762 34.68 ;
      RECT 19.288 33.48 19.584 33.72 ;
      RECT 19.288 32.76 19.762 33.48 ;
      RECT 18.938 32.52 18.984 33.72 ;
      RECT 19.028 32.52 19.072 33.72 ;
      RECT 19.116 32.52 19.244 33.72 ;
      RECT 19.288 32.52 19.584 32.76 ;
      RECT 18.938 31.8 19.584 32.52 ;
      RECT 19.628 31.56 19.762 32.76 ;
      RECT 19.288 31.56 19.584 31.8 ;
      RECT 19.288 30.84 19.762 31.56 ;
      RECT 18.938 30.6 18.984 31.8 ;
      RECT 19.028 30.6 19.072 31.8 ;
      RECT 19.116 30.6 19.244 31.8 ;
      RECT 19.288 30.6 19.584 30.84 ;
      RECT 18.938 29.88 19.584 30.6 ;
      RECT 19.628 29.64 19.762 30.84 ;
      RECT 19.288 29.64 19.584 29.88 ;
      RECT 19.288 28.92 19.762 29.64 ;
      RECT 18.938 28.68 18.984 29.88 ;
      RECT 19.028 28.68 19.072 29.88 ;
      RECT 19.116 28.68 19.244 29.88 ;
      RECT 19.288 28.68 19.584 28.92 ;
      RECT 18.938 27.96 19.584 28.68 ;
      RECT 19.628 27.72 19.762 28.92 ;
      RECT 19.288 27.72 19.584 27.96 ;
      RECT 19.288 27 19.762 27.72 ;
      RECT 18.938 26.76 18.984 27.96 ;
      RECT 19.028 26.76 19.072 27.96 ;
      RECT 19.116 26.76 19.244 27.96 ;
      RECT 19.288 26.76 19.584 27 ;
      RECT 19.628 25.8 19.762 27 ;
      RECT 18.938 25.8 19.584 26.76 ;
      RECT 18.938 24.84 19.762 25.8 ;
      RECT 18.938 23.64 18.984 24.84 ;
      RECT 19.028 23.64 19.244 24.84 ;
      RECT 19.288 23.64 19.672 24.84 ;
      RECT 19.716 23.64 19.762 24.84 ;
      RECT 18.938 21.96 19.762 23.64 ;
      RECT 18.938 20.76 18.984 21.96 ;
      RECT 19.028 20.76 19.244 21.96 ;
      RECT 19.288 20.76 19.672 21.96 ;
      RECT 19.716 20.76 19.762 21.96 ;
      RECT 18.938 19.8 19.762 20.76 ;
      RECT 18.938 18.84 19.412 19.8 ;
      RECT 19.456 18.6 19.584 19.8 ;
      RECT 19.628 18.6 19.762 19.8 ;
      RECT 19.028 18.6 19.412 18.84 ;
      RECT 19.028 17.88 19.762 18.6 ;
      RECT 18.938 17.64 18.984 18.84 ;
      RECT 19.028 17.64 19.412 17.88 ;
      RECT 18.938 16.92 19.412 17.64 ;
      RECT 19.456 16.68 19.584 17.88 ;
      RECT 19.628 16.68 19.762 17.88 ;
      RECT 19.028 16.68 19.412 16.92 ;
      RECT 19.028 15.96 19.762 16.68 ;
      RECT 18.938 15.72 18.984 16.92 ;
      RECT 19.028 15.72 19.412 15.96 ;
      RECT 18.938 15 19.412 15.72 ;
      RECT 19.456 14.76 19.584 15.96 ;
      RECT 19.628 14.76 19.762 15.96 ;
      RECT 19.028 14.76 19.412 15 ;
      RECT 19.028 14.04 19.762 14.76 ;
      RECT 18.938 13.8 18.984 15 ;
      RECT 19.028 13.8 19.412 14.04 ;
      RECT 18.938 13.08 19.412 13.8 ;
      RECT 19.456 12.84 19.584 14.04 ;
      RECT 19.628 12.84 19.762 14.04 ;
      RECT 19.028 12.84 19.412 13.08 ;
      RECT 19.028 12.12 19.762 12.84 ;
      RECT 18.938 11.88 18.984 13.08 ;
      RECT 19.028 11.88 19.412 12.12 ;
      RECT 18.938 11.16 19.412 11.88 ;
      RECT 19.456 10.92 19.584 12.12 ;
      RECT 19.628 10.92 19.762 12.12 ;
      RECT 19.028 10.92 19.412 11.16 ;
      RECT 19.028 10.2 19.762 10.92 ;
      RECT 18.938 9.96 18.984 11.16 ;
      RECT 19.028 9.96 19.412 10.2 ;
      RECT 18.938 9.24 19.412 9.96 ;
      RECT 19.456 9 19.584 10.2 ;
      RECT 19.628 9 19.762 10.2 ;
      RECT 19.028 9 19.412 9.24 ;
      RECT 19.028 8.28 19.762 9 ;
      RECT 18.938 8.04 18.984 9.24 ;
      RECT 19.028 8.04 19.412 8.28 ;
      RECT 18.938 7.32 19.412 8.04 ;
      RECT 19.456 7.08 19.584 8.28 ;
      RECT 19.628 7.08 19.762 8.28 ;
      RECT 19.028 7.08 19.412 7.32 ;
      RECT 19.028 6.36 19.762 7.08 ;
      RECT 18.938 6.12 18.984 7.32 ;
      RECT 19.028 6.12 19.412 6.36 ;
      RECT 18.938 5.4 19.412 6.12 ;
      RECT 19.456 5.16 19.584 6.36 ;
      RECT 19.628 5.16 19.762 6.36 ;
      RECT 19.028 5.16 19.412 5.4 ;
      RECT 19.028 4.44 19.762 5.16 ;
      RECT 18.938 4.2 18.984 5.4 ;
      RECT 19.028 4.2 19.412 4.44 ;
      RECT 18.938 3.48 19.412 4.2 ;
      RECT 19.456 3.24 19.584 4.44 ;
      RECT 19.628 3.24 19.762 4.44 ;
      RECT 19.028 3.24 19.412 3.48 ;
      RECT 19.028 2.52 19.762 3.24 ;
      RECT 18.938 2.28 18.984 3.48 ;
      RECT 19.028 2.28 19.412 2.52 ;
      RECT 18.938 1.56 19.412 2.28 ;
      RECT 19.456 1.32 19.584 2.52 ;
      RECT 19.628 1.32 19.762 2.52 ;
      RECT 19.288 1.32 19.412 1.56 ;
      RECT 18.938 0.36 18.984 1.56 ;
      RECT 19.028 0.36 19.072 1.56 ;
      RECT 19.116 0.36 19.244 1.56 ;
      RECT 19.288 0.36 19.762 1.32 ;
      RECT 18.938 -0.12 19.762 0.36 ;
      RECT 18.038 45.24 18.862 46.2 ;
      RECT 18.038 44.28 18.772 45.24 ;
      RECT 18.816 44.04 18.862 45.24 ;
      RECT 18.216 44.04 18.772 44.28 ;
      RECT 18.216 43.32 18.862 44.04 ;
      RECT 18.038 43.08 18.084 44.28 ;
      RECT 18.128 43.08 18.172 44.28 ;
      RECT 18.216 43.08 18.772 43.32 ;
      RECT 18.038 42.36 18.772 43.08 ;
      RECT 18.816 42.12 18.862 43.32 ;
      RECT 18.216 42.12 18.772 42.36 ;
      RECT 18.216 41.4 18.862 42.12 ;
      RECT 18.038 41.16 18.084 42.36 ;
      RECT 18.128 41.16 18.172 42.36 ;
      RECT 18.216 41.16 18.772 41.4 ;
      RECT 18.038 40.44 18.772 41.16 ;
      RECT 18.816 40.2 18.862 41.4 ;
      RECT 18.216 40.2 18.772 40.44 ;
      RECT 18.216 39.48 18.862 40.2 ;
      RECT 18.038 39.24 18.084 40.44 ;
      RECT 18.128 39.24 18.172 40.44 ;
      RECT 18.216 39.24 18.772 39.48 ;
      RECT 18.038 38.52 18.772 39.24 ;
      RECT 18.816 38.28 18.862 39.48 ;
      RECT 18.216 38.28 18.772 38.52 ;
      RECT 18.216 37.56 18.862 38.28 ;
      RECT 18.038 37.32 18.084 38.52 ;
      RECT 18.128 37.32 18.172 38.52 ;
      RECT 18.216 37.32 18.772 37.56 ;
      RECT 18.038 36.6 18.772 37.32 ;
      RECT 18.816 36.36 18.862 37.56 ;
      RECT 18.216 36.36 18.772 36.6 ;
      RECT 18.216 35.64 18.862 36.36 ;
      RECT 18.038 35.4 18.084 36.6 ;
      RECT 18.128 35.4 18.172 36.6 ;
      RECT 18.216 35.4 18.772 35.64 ;
      RECT 18.038 34.68 18.772 35.4 ;
      RECT 18.816 34.44 18.862 35.64 ;
      RECT 18.216 34.44 18.772 34.68 ;
      RECT 18.216 33.72 18.862 34.44 ;
      RECT 18.038 33.48 18.084 34.68 ;
      RECT 18.128 33.48 18.172 34.68 ;
      RECT 18.216 33.48 18.772 33.72 ;
      RECT 18.038 32.76 18.772 33.48 ;
      RECT 18.816 32.52 18.862 33.72 ;
      RECT 18.216 32.52 18.772 32.76 ;
      RECT 18.216 31.8 18.862 32.52 ;
      RECT 18.038 31.56 18.084 32.76 ;
      RECT 18.128 31.56 18.172 32.76 ;
      RECT 18.216 31.56 18.772 31.8 ;
      RECT 18.038 30.84 18.772 31.56 ;
      RECT 18.816 30.6 18.862 31.8 ;
      RECT 18.216 30.6 18.772 30.84 ;
      RECT 18.216 29.88 18.862 30.6 ;
      RECT 18.038 29.64 18.084 30.84 ;
      RECT 18.128 29.64 18.172 30.84 ;
      RECT 18.216 29.64 18.772 29.88 ;
      RECT 18.038 28.92 18.772 29.64 ;
      RECT 18.816 28.68 18.862 29.88 ;
      RECT 18.216 28.68 18.772 28.92 ;
      RECT 18.216 27.96 18.862 28.68 ;
      RECT 18.038 27.72 18.084 28.92 ;
      RECT 18.128 27.72 18.172 28.92 ;
      RECT 18.216 27.72 18.772 27.96 ;
      RECT 18.038 27 18.772 27.72 ;
      RECT 18.816 26.76 18.862 27.96 ;
      RECT 18.388 26.76 18.772 27 ;
      RECT 18.038 25.8 18.084 27 ;
      RECT 18.128 25.8 18.344 27 ;
      RECT 18.388 25.8 18.862 26.76 ;
      RECT 18.038 24.84 18.862 25.8 ;
      RECT 18.038 23.64 18.172 24.84 ;
      RECT 18.216 23.64 18.428 24.84 ;
      RECT 18.472 23.64 18.684 24.84 ;
      RECT 18.728 23.64 18.862 24.84 ;
      RECT 18.038 21.96 18.862 23.64 ;
      RECT 18.038 20.76 18.172 21.96 ;
      RECT 18.216 20.76 18.428 21.96 ;
      RECT 18.472 20.76 18.684 21.96 ;
      RECT 18.728 20.76 18.862 21.96 ;
      RECT 18.038 19.8 18.862 20.76 ;
      RECT 18.128 18.84 18.862 19.8 ;
      RECT 18.038 18.6 18.084 19.8 ;
      RECT 18.128 18.6 18.512 18.84 ;
      RECT 18.038 17.88 18.512 18.6 ;
      RECT 18.556 17.64 18.684 18.84 ;
      RECT 18.728 17.64 18.772 18.84 ;
      RECT 18.816 17.64 18.862 18.84 ;
      RECT 18.128 17.64 18.512 17.88 ;
      RECT 18.128 16.92 18.862 17.64 ;
      RECT 18.038 16.68 18.084 17.88 ;
      RECT 18.128 16.68 18.512 16.92 ;
      RECT 18.038 15.96 18.512 16.68 ;
      RECT 18.556 15.72 18.684 16.92 ;
      RECT 18.728 15.72 18.772 16.92 ;
      RECT 18.816 15.72 18.862 16.92 ;
      RECT 18.128 15.72 18.512 15.96 ;
      RECT 18.128 15 18.862 15.72 ;
      RECT 18.038 14.76 18.084 15.96 ;
      RECT 18.128 14.76 18.512 15 ;
      RECT 18.038 14.04 18.512 14.76 ;
      RECT 18.556 13.8 18.684 15 ;
      RECT 18.728 13.8 18.772 15 ;
      RECT 18.816 13.8 18.862 15 ;
      RECT 18.128 13.8 18.512 14.04 ;
      RECT 18.128 13.08 18.862 13.8 ;
      RECT 18.038 12.84 18.084 14.04 ;
      RECT 18.128 12.84 18.512 13.08 ;
      RECT 18.038 12.12 18.512 12.84 ;
      RECT 18.556 11.88 18.684 13.08 ;
      RECT 18.728 11.88 18.772 13.08 ;
      RECT 18.816 11.88 18.862 13.08 ;
      RECT 18.128 11.88 18.512 12.12 ;
      RECT 18.128 11.16 18.862 11.88 ;
      RECT 18.038 10.92 18.084 12.12 ;
      RECT 18.128 10.92 18.512 11.16 ;
      RECT 18.038 10.2 18.512 10.92 ;
      RECT 18.556 9.96 18.684 11.16 ;
      RECT 18.728 9.96 18.772 11.16 ;
      RECT 18.816 9.96 18.862 11.16 ;
      RECT 18.128 9.96 18.512 10.2 ;
      RECT 18.128 9.24 18.862 9.96 ;
      RECT 18.038 9 18.084 10.2 ;
      RECT 18.128 9 18.512 9.24 ;
      RECT 18.038 8.28 18.512 9 ;
      RECT 18.556 8.04 18.684 9.24 ;
      RECT 18.728 8.04 18.772 9.24 ;
      RECT 18.816 8.04 18.862 9.24 ;
      RECT 18.128 8.04 18.512 8.28 ;
      RECT 18.128 7.32 18.862 8.04 ;
      RECT 18.038 7.08 18.084 8.28 ;
      RECT 18.128 7.08 18.512 7.32 ;
      RECT 18.038 6.36 18.512 7.08 ;
      RECT 18.556 6.12 18.684 7.32 ;
      RECT 18.728 6.12 18.772 7.32 ;
      RECT 18.816 6.12 18.862 7.32 ;
      RECT 18.128 6.12 18.512 6.36 ;
      RECT 18.128 5.4 18.862 6.12 ;
      RECT 18.038 5.16 18.084 6.36 ;
      RECT 18.128 5.16 18.512 5.4 ;
      RECT 18.038 4.44 18.512 5.16 ;
      RECT 18.556 4.2 18.684 5.4 ;
      RECT 18.728 4.2 18.772 5.4 ;
      RECT 18.816 4.2 18.862 5.4 ;
      RECT 18.128 4.2 18.512 4.44 ;
      RECT 18.128 3.48 18.862 4.2 ;
      RECT 18.038 3.24 18.084 4.44 ;
      RECT 18.128 3.24 18.512 3.48 ;
      RECT 18.038 2.52 18.512 3.24 ;
      RECT 18.556 2.28 18.684 3.48 ;
      RECT 18.728 2.28 18.772 3.48 ;
      RECT 18.816 2.28 18.862 3.48 ;
      RECT 18.128 2.28 18.512 2.52 ;
      RECT 18.128 1.56 18.862 2.28 ;
      RECT 18.038 1.32 18.084 2.52 ;
      RECT 18.128 1.32 18.772 1.56 ;
      RECT 18.816 0.36 18.862 1.56 ;
      RECT 18.038 0.36 18.772 1.32 ;
      RECT 18.038 -0.12 18.862 0.36 ;
      RECT 17.138 44.28 17.962 46.2 ;
      RECT 17.138 43.08 17.184 44.28 ;
      RECT 17.228 43.08 17.272 44.28 ;
      RECT 17.316 43.08 17.872 44.28 ;
      RECT 17.916 43.08 17.962 44.28 ;
      RECT 17.138 42.36 17.962 43.08 ;
      RECT 17.138 41.16 17.184 42.36 ;
      RECT 17.228 41.16 17.272 42.36 ;
      RECT 17.316 41.16 17.872 42.36 ;
      RECT 17.916 41.16 17.962 42.36 ;
      RECT 17.138 40.44 17.962 41.16 ;
      RECT 17.138 39.24 17.184 40.44 ;
      RECT 17.228 39.24 17.272 40.44 ;
      RECT 17.316 39.24 17.872 40.44 ;
      RECT 17.916 39.24 17.962 40.44 ;
      RECT 17.138 38.52 17.962 39.24 ;
      RECT 17.138 37.32 17.184 38.52 ;
      RECT 17.228 37.32 17.272 38.52 ;
      RECT 17.316 37.32 17.872 38.52 ;
      RECT 17.916 37.32 17.962 38.52 ;
      RECT 17.138 36.6 17.962 37.32 ;
      RECT 17.138 35.4 17.184 36.6 ;
      RECT 17.228 35.4 17.272 36.6 ;
      RECT 17.316 35.4 17.872 36.6 ;
      RECT 17.916 35.4 17.962 36.6 ;
      RECT 17.138 34.68 17.962 35.4 ;
      RECT 17.138 33.48 17.184 34.68 ;
      RECT 17.228 33.48 17.272 34.68 ;
      RECT 17.316 33.48 17.872 34.68 ;
      RECT 17.916 33.48 17.962 34.68 ;
      RECT 17.138 32.76 17.962 33.48 ;
      RECT 17.138 31.56 17.184 32.76 ;
      RECT 17.228 31.56 17.272 32.76 ;
      RECT 17.316 31.56 17.872 32.76 ;
      RECT 17.916 31.56 17.962 32.76 ;
      RECT 17.138 30.84 17.962 31.56 ;
      RECT 17.138 29.64 17.184 30.84 ;
      RECT 17.228 29.64 17.272 30.84 ;
      RECT 17.316 29.64 17.872 30.84 ;
      RECT 17.916 29.64 17.962 30.84 ;
      RECT 17.138 28.92 17.962 29.64 ;
      RECT 17.138 27.72 17.184 28.92 ;
      RECT 17.228 27.72 17.272 28.92 ;
      RECT 17.316 27.72 17.872 28.92 ;
      RECT 17.916 27.72 17.962 28.92 ;
      RECT 17.138 27 17.962 27.72 ;
      RECT 17.138 25.8 17.272 27 ;
      RECT 17.316 25.8 17.872 27 ;
      RECT 17.916 25.8 17.962 27 ;
      RECT 17.138 24.84 17.962 25.8 ;
      RECT 17.138 23.64 17.184 24.84 ;
      RECT 17.228 23.64 17.444 24.84 ;
      RECT 17.488 23.64 17.612 24.84 ;
      RECT 17.656 23.64 17.962 24.84 ;
      RECT 17.138 21.96 17.962 23.64 ;
      RECT 17.138 20.76 17.184 21.96 ;
      RECT 17.228 20.76 17.444 21.96 ;
      RECT 17.488 20.76 17.612 21.96 ;
      RECT 17.656 20.76 17.962 21.96 ;
      RECT 17.138 19.8 17.962 20.76 ;
      RECT 17.138 18.84 17.872 19.8 ;
      RECT 17.916 18.6 17.962 19.8 ;
      RECT 17.572 18.6 17.872 18.84 ;
      RECT 17.572 17.88 17.962 18.6 ;
      RECT 17.138 17.64 17.528 18.84 ;
      RECT 17.572 17.64 17.872 17.88 ;
      RECT 17.138 16.92 17.872 17.64 ;
      RECT 17.916 16.68 17.962 17.88 ;
      RECT 17.572 16.68 17.872 16.92 ;
      RECT 17.572 15.96 17.962 16.68 ;
      RECT 17.138 15.72 17.528 16.92 ;
      RECT 17.572 15.72 17.872 15.96 ;
      RECT 17.138 15 17.872 15.72 ;
      RECT 17.916 14.76 17.962 15.96 ;
      RECT 17.572 14.76 17.872 15 ;
      RECT 17.572 14.04 17.962 14.76 ;
      RECT 17.138 13.8 17.528 15 ;
      RECT 17.572 13.8 17.872 14.04 ;
      RECT 17.138 13.08 17.872 13.8 ;
      RECT 17.916 12.84 17.962 14.04 ;
      RECT 17.572 12.84 17.872 13.08 ;
      RECT 17.572 12.12 17.962 12.84 ;
      RECT 17.138 11.88 17.528 13.08 ;
      RECT 17.572 11.88 17.872 12.12 ;
      RECT 17.138 11.16 17.872 11.88 ;
      RECT 17.916 10.92 17.962 12.12 ;
      RECT 17.572 10.92 17.872 11.16 ;
      RECT 17.572 10.2 17.962 10.92 ;
      RECT 17.138 9.96 17.528 11.16 ;
      RECT 17.572 9.96 17.872 10.2 ;
      RECT 17.138 9.24 17.872 9.96 ;
      RECT 17.916 9 17.962 10.2 ;
      RECT 17.572 9 17.872 9.24 ;
      RECT 17.572 8.28 17.962 9 ;
      RECT 17.138 8.04 17.528 9.24 ;
      RECT 17.572 8.04 17.872 8.28 ;
      RECT 17.138 7.32 17.872 8.04 ;
      RECT 17.916 7.08 17.962 8.28 ;
      RECT 17.572 7.08 17.872 7.32 ;
      RECT 17.572 6.36 17.962 7.08 ;
      RECT 17.138 6.12 17.528 7.32 ;
      RECT 17.572 6.12 17.872 6.36 ;
      RECT 17.138 5.4 17.872 6.12 ;
      RECT 17.916 5.16 17.962 6.36 ;
      RECT 17.572 5.16 17.872 5.4 ;
      RECT 17.572 4.44 17.962 5.16 ;
      RECT 17.138 4.2 17.528 5.4 ;
      RECT 17.572 4.2 17.872 4.44 ;
      RECT 17.138 3.48 17.872 4.2 ;
      RECT 17.916 3.24 17.962 4.44 ;
      RECT 17.572 3.24 17.872 3.48 ;
      RECT 17.138 2.52 17.528 3.48 ;
      RECT 17.572 2.52 17.962 3.24 ;
      RECT 17.228 2.28 17.528 2.52 ;
      RECT 17.572 2.28 17.872 2.52 ;
      RECT 17.138 1.32 17.184 2.52 ;
      RECT 17.916 1.32 17.962 2.52 ;
      RECT 17.228 1.32 17.872 2.28 ;
      RECT 17.138 -0.12 17.962 1.32 ;
      RECT 16.238 44.28 17.062 46.2 ;
      RECT 16.238 43.08 16.884 44.28 ;
      RECT 16.928 43.08 16.972 44.28 ;
      RECT 17.016 43.08 17.062 44.28 ;
      RECT 16.238 42.36 17.062 43.08 ;
      RECT 16.238 41.16 16.884 42.36 ;
      RECT 16.928 41.16 16.972 42.36 ;
      RECT 17.016 41.16 17.062 42.36 ;
      RECT 16.238 40.44 17.062 41.16 ;
      RECT 16.238 39.24 16.884 40.44 ;
      RECT 16.928 39.24 16.972 40.44 ;
      RECT 17.016 39.24 17.062 40.44 ;
      RECT 16.238 38.52 17.062 39.24 ;
      RECT 16.238 37.32 16.884 38.52 ;
      RECT 16.928 37.32 16.972 38.52 ;
      RECT 17.016 37.32 17.062 38.52 ;
      RECT 16.238 36.6 17.062 37.32 ;
      RECT 16.238 35.4 16.884 36.6 ;
      RECT 16.928 35.4 16.972 36.6 ;
      RECT 17.016 35.4 17.062 36.6 ;
      RECT 16.238 34.68 17.062 35.4 ;
      RECT 16.238 33.48 16.884 34.68 ;
      RECT 16.928 33.48 16.972 34.68 ;
      RECT 17.016 33.48 17.062 34.68 ;
      RECT 16.238 32.76 17.062 33.48 ;
      RECT 16.238 31.56 16.884 32.76 ;
      RECT 16.928 31.56 16.972 32.76 ;
      RECT 17.016 31.56 17.062 32.76 ;
      RECT 16.238 30.84 17.062 31.56 ;
      RECT 16.238 29.64 16.884 30.84 ;
      RECT 16.928 29.64 16.972 30.84 ;
      RECT 17.016 29.64 17.062 30.84 ;
      RECT 16.238 28.92 17.062 29.64 ;
      RECT 16.238 27.72 16.884 28.92 ;
      RECT 16.928 27.72 16.972 28.92 ;
      RECT 17.016 27.72 17.062 28.92 ;
      RECT 16.238 27 17.062 27.72 ;
      RECT 16.238 25.8 16.712 27 ;
      RECT 16.756 25.8 16.884 27 ;
      RECT 16.928 25.8 16.972 27 ;
      RECT 17.016 25.8 17.062 27 ;
      RECT 16.238 24.84 17.062 25.8 ;
      RECT 16.238 23.64 16.372 24.84 ;
      RECT 16.416 23.64 17.062 24.84 ;
      RECT 16.238 21.96 17.062 23.64 ;
      RECT 16.238 20.76 16.372 21.96 ;
      RECT 16.416 20.76 17.062 21.96 ;
      RECT 16.238 19.8 17.062 20.76 ;
      RECT 16.238 18.6 16.628 19.8 ;
      RECT 16.672 18.6 16.712 19.8 ;
      RECT 16.756 18.6 16.884 19.8 ;
      RECT 16.928 18.6 16.972 19.8 ;
      RECT 17.016 18.6 17.062 19.8 ;
      RECT 16.238 17.88 17.062 18.6 ;
      RECT 16.238 16.68 16.628 17.88 ;
      RECT 16.672 16.68 16.712 17.88 ;
      RECT 16.756 16.68 16.884 17.88 ;
      RECT 16.928 16.68 16.972 17.88 ;
      RECT 17.016 16.68 17.062 17.88 ;
      RECT 16.238 15.96 17.062 16.68 ;
      RECT 16.238 14.76 16.628 15.96 ;
      RECT 16.672 14.76 16.712 15.96 ;
      RECT 16.756 14.76 16.884 15.96 ;
      RECT 16.928 14.76 16.972 15.96 ;
      RECT 17.016 14.76 17.062 15.96 ;
      RECT 16.238 14.04 17.062 14.76 ;
      RECT 16.238 12.84 16.628 14.04 ;
      RECT 16.672 12.84 16.712 14.04 ;
      RECT 16.756 12.84 16.884 14.04 ;
      RECT 16.928 12.84 16.972 14.04 ;
      RECT 17.016 12.84 17.062 14.04 ;
      RECT 16.238 12.12 17.062 12.84 ;
      RECT 16.238 10.92 16.628 12.12 ;
      RECT 16.672 10.92 16.712 12.12 ;
      RECT 16.756 10.92 16.884 12.12 ;
      RECT 16.928 10.92 16.972 12.12 ;
      RECT 17.016 10.92 17.062 12.12 ;
      RECT 16.238 10.2 17.062 10.92 ;
      RECT 16.238 9 16.628 10.2 ;
      RECT 16.672 9 16.712 10.2 ;
      RECT 16.756 9 16.884 10.2 ;
      RECT 16.928 9 16.972 10.2 ;
      RECT 17.016 9 17.062 10.2 ;
      RECT 16.238 8.28 17.062 9 ;
      RECT 16.238 7.08 16.628 8.28 ;
      RECT 16.672 7.08 16.712 8.28 ;
      RECT 16.756 7.08 16.884 8.28 ;
      RECT 16.928 7.08 16.972 8.28 ;
      RECT 17.016 7.08 17.062 8.28 ;
      RECT 16.238 6.36 17.062 7.08 ;
      RECT 16.238 5.16 16.628 6.36 ;
      RECT 16.672 5.16 16.712 6.36 ;
      RECT 16.756 5.16 16.884 6.36 ;
      RECT 16.928 5.16 16.972 6.36 ;
      RECT 17.016 5.16 17.062 6.36 ;
      RECT 16.238 4.44 17.062 5.16 ;
      RECT 16.238 3.24 16.628 4.44 ;
      RECT 16.672 3.24 16.712 4.44 ;
      RECT 16.756 3.24 16.884 4.44 ;
      RECT 16.928 3.24 16.972 4.44 ;
      RECT 17.016 3.24 17.062 4.44 ;
      RECT 16.238 2.52 17.062 3.24 ;
      RECT 16.238 1.56 16.712 2.52 ;
      RECT 16.756 1.32 16.884 2.52 ;
      RECT 16.928 1.32 16.972 2.52 ;
      RECT 17.016 1.32 17.062 2.52 ;
      RECT 16.588 1.32 16.712 1.56 ;
      RECT 16.238 0.36 16.284 1.56 ;
      RECT 16.328 0.36 16.372 1.56 ;
      RECT 16.416 0.36 16.544 1.56 ;
      RECT 16.588 0.36 17.062 1.32 ;
      RECT 16.238 -0.12 17.062 0.36 ;
      RECT 15.338 45.24 16.162 46.2 ;
      RECT 15.338 44.04 15.384 45.24 ;
      RECT 15.428 44.04 15.472 45.24 ;
      RECT 15.516 44.04 15.728 45.24 ;
      RECT 15.772 44.04 15.812 45.24 ;
      RECT 15.856 44.04 15.984 45.24 ;
      RECT 16.028 44.04 16.072 45.24 ;
      RECT 16.116 44.04 16.162 45.24 ;
      RECT 15.338 43.32 16.162 44.04 ;
      RECT 15.338 42.12 15.384 43.32 ;
      RECT 15.428 42.12 15.472 43.32 ;
      RECT 15.516 42.12 15.728 43.32 ;
      RECT 15.772 42.12 15.812 43.32 ;
      RECT 15.856 42.12 15.984 43.32 ;
      RECT 16.028 42.12 16.072 43.32 ;
      RECT 16.116 42.12 16.162 43.32 ;
      RECT 15.338 41.4 16.162 42.12 ;
      RECT 15.338 40.2 15.384 41.4 ;
      RECT 15.428 40.2 15.472 41.4 ;
      RECT 15.516 40.2 15.728 41.4 ;
      RECT 15.772 40.2 15.812 41.4 ;
      RECT 15.856 40.2 15.984 41.4 ;
      RECT 16.028 40.2 16.072 41.4 ;
      RECT 16.116 40.2 16.162 41.4 ;
      RECT 15.338 39.48 16.162 40.2 ;
      RECT 15.338 38.28 15.384 39.48 ;
      RECT 15.428 38.28 15.472 39.48 ;
      RECT 15.516 38.28 15.728 39.48 ;
      RECT 15.772 38.28 15.812 39.48 ;
      RECT 15.856 38.28 15.984 39.48 ;
      RECT 16.028 38.28 16.072 39.48 ;
      RECT 16.116 38.28 16.162 39.48 ;
      RECT 15.338 37.56 16.162 38.28 ;
      RECT 15.338 36.36 15.384 37.56 ;
      RECT 15.428 36.36 15.472 37.56 ;
      RECT 15.516 36.36 15.728 37.56 ;
      RECT 15.772 36.36 15.812 37.56 ;
      RECT 15.856 36.36 15.984 37.56 ;
      RECT 16.028 36.36 16.072 37.56 ;
      RECT 16.116 36.36 16.162 37.56 ;
      RECT 15.338 35.64 16.162 36.36 ;
      RECT 15.338 34.44 15.384 35.64 ;
      RECT 15.428 34.44 15.472 35.64 ;
      RECT 15.516 34.44 15.728 35.64 ;
      RECT 15.772 34.44 15.812 35.64 ;
      RECT 15.856 34.44 15.984 35.64 ;
      RECT 16.028 34.44 16.072 35.64 ;
      RECT 16.116 34.44 16.162 35.64 ;
      RECT 15.338 33.72 16.162 34.44 ;
      RECT 15.338 32.52 15.384 33.72 ;
      RECT 15.428 32.52 15.472 33.72 ;
      RECT 15.516 32.52 15.728 33.72 ;
      RECT 15.772 32.52 15.812 33.72 ;
      RECT 15.856 32.52 15.984 33.72 ;
      RECT 16.028 32.52 16.072 33.72 ;
      RECT 16.116 32.52 16.162 33.72 ;
      RECT 15.338 31.8 16.162 32.52 ;
      RECT 15.338 30.6 15.384 31.8 ;
      RECT 15.428 30.6 15.472 31.8 ;
      RECT 15.516 30.6 15.728 31.8 ;
      RECT 15.772 30.6 15.812 31.8 ;
      RECT 15.856 30.6 15.984 31.8 ;
      RECT 16.028 30.6 16.072 31.8 ;
      RECT 16.116 30.6 16.162 31.8 ;
      RECT 15.338 29.88 16.162 30.6 ;
      RECT 15.338 28.68 15.384 29.88 ;
      RECT 15.428 28.68 15.472 29.88 ;
      RECT 15.516 28.68 15.728 29.88 ;
      RECT 15.772 28.68 15.812 29.88 ;
      RECT 15.856 28.68 15.984 29.88 ;
      RECT 16.028 28.68 16.072 29.88 ;
      RECT 16.116 28.68 16.162 29.88 ;
      RECT 15.338 27.96 16.162 28.68 ;
      RECT 15.338 26.76 15.384 27.96 ;
      RECT 15.428 26.76 15.472 27.96 ;
      RECT 15.516 26.76 15.728 27.96 ;
      RECT 15.772 26.76 15.812 27.96 ;
      RECT 15.856 26.76 15.984 27.96 ;
      RECT 16.028 26.76 16.072 27.96 ;
      RECT 16.116 26.76 16.162 27.96 ;
      RECT 15.338 24.84 16.162 26.76 ;
      RECT 15.338 23.64 15.384 24.84 ;
      RECT 15.428 23.64 15.644 24.84 ;
      RECT 15.688 23.64 15.812 24.84 ;
      RECT 15.856 23.64 16.072 24.84 ;
      RECT 16.116 23.64 16.162 24.84 ;
      RECT 15.338 21.96 16.162 23.64 ;
      RECT 15.338 20.76 15.384 21.96 ;
      RECT 15.428 20.76 15.644 21.96 ;
      RECT 15.688 20.76 15.812 21.96 ;
      RECT 15.856 20.76 16.072 21.96 ;
      RECT 16.116 20.76 16.162 21.96 ;
      RECT 15.338 18.84 16.162 20.76 ;
      RECT 15.338 17.64 15.384 18.84 ;
      RECT 15.428 17.64 15.728 18.84 ;
      RECT 15.772 17.64 15.812 18.84 ;
      RECT 15.856 17.64 15.984 18.84 ;
      RECT 16.028 17.64 16.162 18.84 ;
      RECT 15.338 16.92 16.162 17.64 ;
      RECT 15.338 15.72 15.384 16.92 ;
      RECT 15.428 15.72 15.728 16.92 ;
      RECT 15.772 15.72 15.812 16.92 ;
      RECT 15.856 15.72 15.984 16.92 ;
      RECT 16.028 15.72 16.162 16.92 ;
      RECT 15.338 15 16.162 15.72 ;
      RECT 15.338 13.8 15.384 15 ;
      RECT 15.428 13.8 15.728 15 ;
      RECT 15.772 13.8 15.812 15 ;
      RECT 15.856 13.8 15.984 15 ;
      RECT 16.028 13.8 16.162 15 ;
      RECT 15.338 13.08 16.162 13.8 ;
      RECT 15.338 11.88 15.384 13.08 ;
      RECT 15.428 11.88 15.728 13.08 ;
      RECT 15.772 11.88 15.812 13.08 ;
      RECT 15.856 11.88 15.984 13.08 ;
      RECT 16.028 11.88 16.162 13.08 ;
      RECT 15.338 11.16 16.162 11.88 ;
      RECT 15.338 9.96 15.384 11.16 ;
      RECT 15.428 9.96 15.728 11.16 ;
      RECT 15.772 9.96 15.812 11.16 ;
      RECT 15.856 9.96 15.984 11.16 ;
      RECT 16.028 9.96 16.162 11.16 ;
      RECT 15.338 9.24 16.162 9.96 ;
      RECT 15.338 8.04 15.384 9.24 ;
      RECT 15.428 8.04 15.728 9.24 ;
      RECT 15.772 8.04 15.812 9.24 ;
      RECT 15.856 8.04 15.984 9.24 ;
      RECT 16.028 8.04 16.162 9.24 ;
      RECT 15.338 7.32 16.162 8.04 ;
      RECT 15.338 6.12 15.384 7.32 ;
      RECT 15.428 6.12 15.728 7.32 ;
      RECT 15.772 6.12 15.812 7.32 ;
      RECT 15.856 6.12 15.984 7.32 ;
      RECT 16.028 6.12 16.162 7.32 ;
      RECT 15.338 5.4 16.162 6.12 ;
      RECT 15.338 4.2 15.384 5.4 ;
      RECT 15.428 4.2 15.728 5.4 ;
      RECT 15.772 4.2 15.812 5.4 ;
      RECT 15.856 4.2 15.984 5.4 ;
      RECT 16.028 4.2 16.162 5.4 ;
      RECT 15.338 3.48 16.162 4.2 ;
      RECT 15.338 2.28 15.384 3.48 ;
      RECT 15.428 2.28 15.728 3.48 ;
      RECT 15.772 2.28 15.812 3.48 ;
      RECT 15.856 2.28 15.984 3.48 ;
      RECT 16.028 2.28 16.162 3.48 ;
      RECT 15.338 1.56 16.162 2.28 ;
      RECT 15.338 0.36 16.072 1.56 ;
      RECT 16.116 0.36 16.162 1.56 ;
      RECT 15.338 -0.12 16.162 0.36 ;
      RECT 14.438 45.24 15.262 46.2 ;
      RECT 14.438 44.04 15.084 45.24 ;
      RECT 15.128 44.04 15.172 45.24 ;
      RECT 15.216 44.04 15.262 45.24 ;
      RECT 14.438 43.32 15.262 44.04 ;
      RECT 14.438 42.12 15.084 43.32 ;
      RECT 15.128 42.12 15.172 43.32 ;
      RECT 15.216 42.12 15.262 43.32 ;
      RECT 14.438 41.4 15.262 42.12 ;
      RECT 14.438 40.2 15.084 41.4 ;
      RECT 15.128 40.2 15.172 41.4 ;
      RECT 15.216 40.2 15.262 41.4 ;
      RECT 14.438 39.48 15.262 40.2 ;
      RECT 14.438 38.28 15.084 39.48 ;
      RECT 15.128 38.28 15.172 39.48 ;
      RECT 15.216 38.28 15.262 39.48 ;
      RECT 14.438 37.56 15.262 38.28 ;
      RECT 14.438 36.36 15.084 37.56 ;
      RECT 15.128 36.36 15.172 37.56 ;
      RECT 15.216 36.36 15.262 37.56 ;
      RECT 14.438 35.64 15.262 36.36 ;
      RECT 14.438 34.44 15.084 35.64 ;
      RECT 15.128 34.44 15.172 35.64 ;
      RECT 15.216 34.44 15.262 35.64 ;
      RECT 14.438 33.72 15.262 34.44 ;
      RECT 14.438 32.52 15.084 33.72 ;
      RECT 15.128 32.52 15.172 33.72 ;
      RECT 15.216 32.52 15.262 33.72 ;
      RECT 14.438 31.8 15.262 32.52 ;
      RECT 14.438 30.6 15.084 31.8 ;
      RECT 15.128 30.6 15.172 31.8 ;
      RECT 15.216 30.6 15.262 31.8 ;
      RECT 14.438 29.88 15.262 30.6 ;
      RECT 14.438 28.68 15.084 29.88 ;
      RECT 15.128 28.68 15.172 29.88 ;
      RECT 15.216 28.68 15.262 29.88 ;
      RECT 14.438 27.96 15.262 28.68 ;
      RECT 14.438 26.76 15.084 27.96 ;
      RECT 15.128 26.76 15.172 27.96 ;
      RECT 15.216 26.76 15.262 27.96 ;
      RECT 14.438 24.84 15.262 26.76 ;
      RECT 14.438 23.64 14.572 24.84 ;
      RECT 14.616 23.64 14.828 24.84 ;
      RECT 14.872 23.64 15.084 24.84 ;
      RECT 15.128 23.64 15.262 24.84 ;
      RECT 14.438 21.96 15.262 23.64 ;
      RECT 14.438 20.76 14.572 21.96 ;
      RECT 14.616 20.76 14.828 21.96 ;
      RECT 14.872 20.76 15.084 21.96 ;
      RECT 15.128 20.76 15.262 21.96 ;
      RECT 14.438 18.84 15.262 20.76 ;
      RECT 14.438 17.64 14.912 18.84 ;
      RECT 14.956 17.64 15.084 18.84 ;
      RECT 15.128 17.64 15.172 18.84 ;
      RECT 15.216 17.64 15.262 18.84 ;
      RECT 14.438 16.92 15.262 17.64 ;
      RECT 14.438 15.72 14.912 16.92 ;
      RECT 14.956 15.72 15.084 16.92 ;
      RECT 15.128 15.72 15.172 16.92 ;
      RECT 15.216 15.72 15.262 16.92 ;
      RECT 14.438 15 15.262 15.72 ;
      RECT 14.438 13.8 14.912 15 ;
      RECT 14.956 13.8 15.084 15 ;
      RECT 15.128 13.8 15.172 15 ;
      RECT 15.216 13.8 15.262 15 ;
      RECT 14.438 13.08 15.262 13.8 ;
      RECT 14.438 11.88 14.912 13.08 ;
      RECT 14.956 11.88 15.084 13.08 ;
      RECT 15.128 11.88 15.172 13.08 ;
      RECT 15.216 11.88 15.262 13.08 ;
      RECT 14.438 11.16 15.262 11.88 ;
      RECT 14.438 9.96 14.912 11.16 ;
      RECT 14.956 9.96 15.084 11.16 ;
      RECT 15.128 9.96 15.172 11.16 ;
      RECT 15.216 9.96 15.262 11.16 ;
      RECT 14.438 9.24 15.262 9.96 ;
      RECT 14.438 8.04 14.912 9.24 ;
      RECT 14.956 8.04 15.084 9.24 ;
      RECT 15.128 8.04 15.172 9.24 ;
      RECT 15.216 8.04 15.262 9.24 ;
      RECT 14.438 7.32 15.262 8.04 ;
      RECT 14.438 6.12 14.912 7.32 ;
      RECT 14.956 6.12 15.084 7.32 ;
      RECT 15.128 6.12 15.172 7.32 ;
      RECT 15.216 6.12 15.262 7.32 ;
      RECT 14.438 5.4 15.262 6.12 ;
      RECT 14.438 4.2 14.912 5.4 ;
      RECT 14.956 4.2 15.084 5.4 ;
      RECT 15.128 4.2 15.172 5.4 ;
      RECT 15.216 4.2 15.262 5.4 ;
      RECT 14.438 3.48 15.262 4.2 ;
      RECT 14.438 2.52 14.912 3.48 ;
      RECT 14.956 2.28 15.084 3.48 ;
      RECT 15.128 2.28 15.172 3.48 ;
      RECT 15.216 2.28 15.262 3.48 ;
      RECT 14.616 2.28 14.912 2.52 ;
      RECT 14.438 1.32 14.484 2.52 ;
      RECT 14.528 1.32 14.572 2.52 ;
      RECT 14.616 1.32 15.262 2.28 ;
      RECT 14.438 -0.12 15.262 1.32 ;
      RECT 13.538 44.28 14.362 46.2 ;
      RECT 13.538 43.08 13.844 44.28 ;
      RECT 13.888 43.08 13.928 44.28 ;
      RECT 13.972 43.08 14.012 44.28 ;
      RECT 14.056 43.08 14.184 44.28 ;
      RECT 14.228 43.08 14.362 44.28 ;
      RECT 13.538 42.36 14.362 43.08 ;
      RECT 13.538 41.16 13.844 42.36 ;
      RECT 13.888 41.16 13.928 42.36 ;
      RECT 13.972 41.16 14.012 42.36 ;
      RECT 14.056 41.16 14.184 42.36 ;
      RECT 14.228 41.16 14.362 42.36 ;
      RECT 13.538 40.44 14.362 41.16 ;
      RECT 13.538 39.24 13.844 40.44 ;
      RECT 13.888 39.24 13.928 40.44 ;
      RECT 13.972 39.24 14.012 40.44 ;
      RECT 14.056 39.24 14.184 40.44 ;
      RECT 14.228 39.24 14.362 40.44 ;
      RECT 13.538 38.52 14.362 39.24 ;
      RECT 13.538 37.32 13.844 38.52 ;
      RECT 13.888 37.32 13.928 38.52 ;
      RECT 13.972 37.32 14.012 38.52 ;
      RECT 14.056 37.32 14.184 38.52 ;
      RECT 14.228 37.32 14.362 38.52 ;
      RECT 13.538 36.6 14.362 37.32 ;
      RECT 13.538 35.4 13.844 36.6 ;
      RECT 13.888 35.4 13.928 36.6 ;
      RECT 13.972 35.4 14.012 36.6 ;
      RECT 14.056 35.4 14.184 36.6 ;
      RECT 14.228 35.4 14.362 36.6 ;
      RECT 13.538 34.68 14.362 35.4 ;
      RECT 13.538 33.48 13.844 34.68 ;
      RECT 13.888 33.48 13.928 34.68 ;
      RECT 13.972 33.48 14.012 34.68 ;
      RECT 14.056 33.48 14.184 34.68 ;
      RECT 14.228 33.48 14.362 34.68 ;
      RECT 13.538 32.76 14.362 33.48 ;
      RECT 13.538 31.56 13.844 32.76 ;
      RECT 13.888 31.56 13.928 32.76 ;
      RECT 13.972 31.56 14.012 32.76 ;
      RECT 14.056 31.56 14.184 32.76 ;
      RECT 14.228 31.56 14.362 32.76 ;
      RECT 13.538 30.84 14.362 31.56 ;
      RECT 13.538 29.64 13.844 30.84 ;
      RECT 13.888 29.64 13.928 30.84 ;
      RECT 13.972 29.64 14.012 30.84 ;
      RECT 14.056 29.64 14.184 30.84 ;
      RECT 14.228 29.64 14.362 30.84 ;
      RECT 13.538 28.92 14.362 29.64 ;
      RECT 13.538 27.72 13.844 28.92 ;
      RECT 13.888 27.72 13.928 28.92 ;
      RECT 13.972 27.72 14.012 28.92 ;
      RECT 14.056 27.72 14.184 28.92 ;
      RECT 14.228 27.72 14.362 28.92 ;
      RECT 13.538 27 14.362 27.72 ;
      RECT 13.538 25.8 13.844 27 ;
      RECT 13.888 25.8 13.928 27 ;
      RECT 13.972 25.8 14.012 27 ;
      RECT 14.056 25.8 14.184 27 ;
      RECT 14.228 25.8 14.362 27 ;
      RECT 13.538 24.84 14.362 25.8 ;
      RECT 13.538 23.64 13.584 24.84 ;
      RECT 13.628 23.64 14.272 24.84 ;
      RECT 14.316 23.64 14.362 24.84 ;
      RECT 13.538 21.96 14.362 23.64 ;
      RECT 13.538 20.76 13.584 21.96 ;
      RECT 13.628 20.76 14.272 21.96 ;
      RECT 14.316 20.76 14.362 21.96 ;
      RECT 13.538 19.8 14.362 20.76 ;
      RECT 13.538 18.6 13.672 19.8 ;
      RECT 13.716 18.6 13.844 19.8 ;
      RECT 13.888 18.6 13.928 19.8 ;
      RECT 13.972 18.6 14.012 19.8 ;
      RECT 14.056 18.6 14.362 19.8 ;
      RECT 13.538 17.88 14.362 18.6 ;
      RECT 13.538 16.68 13.672 17.88 ;
      RECT 13.716 16.68 13.844 17.88 ;
      RECT 13.888 16.68 13.928 17.88 ;
      RECT 13.972 16.68 14.012 17.88 ;
      RECT 14.056 16.68 14.362 17.88 ;
      RECT 13.538 15.96 14.362 16.68 ;
      RECT 13.538 14.76 13.672 15.96 ;
      RECT 13.716 14.76 13.844 15.96 ;
      RECT 13.888 14.76 13.928 15.96 ;
      RECT 13.972 14.76 14.012 15.96 ;
      RECT 14.056 14.76 14.362 15.96 ;
      RECT 13.538 14.04 14.362 14.76 ;
      RECT 13.538 12.84 13.672 14.04 ;
      RECT 13.716 12.84 13.844 14.04 ;
      RECT 13.888 12.84 13.928 14.04 ;
      RECT 13.972 12.84 14.012 14.04 ;
      RECT 14.056 12.84 14.362 14.04 ;
      RECT 13.538 12.12 14.362 12.84 ;
      RECT 13.538 10.92 13.672 12.12 ;
      RECT 13.716 10.92 13.844 12.12 ;
      RECT 13.888 10.92 13.928 12.12 ;
      RECT 13.972 10.92 14.012 12.12 ;
      RECT 14.056 10.92 14.362 12.12 ;
      RECT 13.538 10.2 14.362 10.92 ;
      RECT 13.538 9 13.672 10.2 ;
      RECT 13.716 9 13.844 10.2 ;
      RECT 13.888 9 13.928 10.2 ;
      RECT 13.972 9 14.012 10.2 ;
      RECT 14.056 9 14.362 10.2 ;
      RECT 13.538 8.28 14.362 9 ;
      RECT 13.538 7.08 13.672 8.28 ;
      RECT 13.716 7.08 13.844 8.28 ;
      RECT 13.888 7.08 13.928 8.28 ;
      RECT 13.972 7.08 14.012 8.28 ;
      RECT 14.056 7.08 14.362 8.28 ;
      RECT 13.538 6.36 14.362 7.08 ;
      RECT 13.538 5.16 13.672 6.36 ;
      RECT 13.716 5.16 13.844 6.36 ;
      RECT 13.888 5.16 13.928 6.36 ;
      RECT 13.972 5.16 14.012 6.36 ;
      RECT 14.056 5.16 14.362 6.36 ;
      RECT 13.538 4.44 14.362 5.16 ;
      RECT 13.538 3.24 13.672 4.44 ;
      RECT 13.716 3.24 13.844 4.44 ;
      RECT 13.888 3.24 13.928 4.44 ;
      RECT 13.972 3.24 14.012 4.44 ;
      RECT 14.056 3.24 14.362 4.44 ;
      RECT 13.538 2.52 14.362 3.24 ;
      RECT 13.538 1.56 14.184 2.52 ;
      RECT 14.228 1.32 14.272 2.52 ;
      RECT 14.316 1.32 14.362 2.52 ;
      RECT 13.972 1.32 14.184 1.56 ;
      RECT 13.538 0.36 13.584 1.56 ;
      RECT 13.628 0.36 13.672 1.56 ;
      RECT 13.716 0.36 13.844 1.56 ;
      RECT 13.888 0.36 13.928 1.56 ;
      RECT 13.972 0.36 14.362 1.32 ;
      RECT 13.538 -0.12 14.362 0.36 ;
      RECT 12.638 -0.12 13.462 46.2 ;
      RECT 11.738 -0.12 12.562 46.2 ;
      RECT 10.838 -0.12 11.662 46.2 ;
      RECT 9.938 -0.12 10.762 46.2 ;
      RECT 9.038 -0.12 9.862 46.2 ;
      RECT 8.138 -0.12 8.962 46.2 ;
      RECT 7.238 -0.12 8.062 46.2 ;
      RECT 6.338 -0.12 7.162 46.2 ;
      RECT 5.438 -0.12 6.262 46.2 ;
      RECT 4.538 -0.12 5.362 46.2 ;
      RECT 3.638 -0.12 4.462 46.2 ;
      RECT 2.738 -0.12 3.562 46.2 ;
      RECT 1.838 -0.12 2.662 46.2 ;
      RECT 0.938 -0.12 1.762 46.2 ;
      RECT -0.04 46.14 0.862 46.2 ;
      RECT -0.092 -0.06 0.862 46.14 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 37.058 0 37.72 46.08 ;
      RECT 36.158 0 36.742 46.08 ;
      RECT 35.258 0 35.842 46.08 ;
      RECT 34.358 0 34.942 46.08 ;
      RECT 33.458 0 34.042 46.08 ;
      RECT 32.558 0 33.142 46.08 ;
      RECT 31.658 0 32.242 46.08 ;
      RECT 30.758 0 31.342 46.08 ;
      RECT 29.858 0 30.442 46.08 ;
      RECT 28.958 0 29.542 46.08 ;
      RECT 28.058 0 28.642 46.08 ;
      RECT 27.158 0 27.742 46.08 ;
      RECT 26.258 0 26.842 46.08 ;
      RECT 25.358 0 25.942 46.08 ;
      RECT 24.458 0 25.042 46.08 ;
      RECT 23.558 0 24.142 46.08 ;
      RECT 22.658 0 23.242 46.08 ;
      RECT 21.758 45.36 22.342 46.08 ;
      RECT 21.936 43.92 22.342 45.36 ;
      RECT 21.758 43.44 22.342 43.92 ;
      RECT 21.936 42 22.342 43.44 ;
      RECT 21.758 41.52 22.342 42 ;
      RECT 21.936 40.08 22.342 41.52 ;
      RECT 21.758 39.6 22.342 40.08 ;
      RECT 21.936 38.16 22.342 39.6 ;
      RECT 21.758 37.68 22.342 38.16 ;
      RECT 21.936 36.24 22.342 37.68 ;
      RECT 21.758 35.76 22.342 36.24 ;
      RECT 21.936 34.32 22.342 35.76 ;
      RECT 21.758 33.84 22.342 34.32 ;
      RECT 21.936 32.4 22.342 33.84 ;
      RECT 21.758 31.92 22.342 32.4 ;
      RECT 21.936 30.48 22.342 31.92 ;
      RECT 21.758 30 22.342 30.48 ;
      RECT 21.936 28.56 22.342 30 ;
      RECT 21.758 28.08 22.342 28.56 ;
      RECT 21.936 26.64 22.342 28.08 ;
      RECT 21.758 18.96 22.342 26.64 ;
      RECT 21.936 17.52 22.342 18.96 ;
      RECT 21.758 17.04 22.342 17.52 ;
      RECT 21.936 15.6 22.342 17.04 ;
      RECT 21.758 15.12 22.342 15.6 ;
      RECT 21.936 13.68 22.342 15.12 ;
      RECT 21.758 13.2 22.342 13.68 ;
      RECT 21.936 11.76 22.342 13.2 ;
      RECT 21.758 11.28 22.342 11.76 ;
      RECT 21.936 9.84 22.342 11.28 ;
      RECT 21.758 9.36 22.342 9.84 ;
      RECT 21.936 7.92 22.342 9.36 ;
      RECT 21.758 7.44 22.342 7.92 ;
      RECT 21.936 6 22.342 7.44 ;
      RECT 21.758 5.52 22.342 6 ;
      RECT 21.936 4.08 22.342 5.52 ;
      RECT 21.758 3.6 22.342 4.08 ;
      RECT 21.936 2.16 22.342 3.6 ;
      RECT 21.758 1.68 22.342 2.16 ;
      RECT 21.936 0.24 22.342 1.68 ;
      RECT 21.758 0 22.342 0.24 ;
      RECT 20.858 45.36 21.442 46.08 ;
      RECT 20.858 44.4 21.352 45.36 ;
      RECT 21.036 43.92 21.352 44.4 ;
      RECT 21.036 43.44 21.442 43.92 ;
      RECT 21.036 42.96 21.352 43.44 ;
      RECT 20.858 42.48 21.352 42.96 ;
      RECT 21.036 42 21.352 42.48 ;
      RECT 21.036 41.52 21.442 42 ;
      RECT 21.036 41.04 21.352 41.52 ;
      RECT 20.858 40.56 21.352 41.04 ;
      RECT 21.036 40.08 21.352 40.56 ;
      RECT 21.036 39.6 21.442 40.08 ;
      RECT 21.036 39.12 21.352 39.6 ;
      RECT 20.858 38.64 21.352 39.12 ;
      RECT 21.036 38.16 21.352 38.64 ;
      RECT 21.036 37.68 21.442 38.16 ;
      RECT 21.036 37.2 21.352 37.68 ;
      RECT 20.858 36.72 21.352 37.2 ;
      RECT 21.036 36.24 21.352 36.72 ;
      RECT 21.036 35.76 21.442 36.24 ;
      RECT 21.036 35.28 21.352 35.76 ;
      RECT 20.858 34.8 21.352 35.28 ;
      RECT 21.036 34.32 21.352 34.8 ;
      RECT 21.036 33.84 21.442 34.32 ;
      RECT 21.036 33.36 21.352 33.84 ;
      RECT 20.858 32.88 21.352 33.36 ;
      RECT 21.036 32.4 21.352 32.88 ;
      RECT 21.036 31.92 21.442 32.4 ;
      RECT 21.036 31.44 21.352 31.92 ;
      RECT 20.858 30.96 21.352 31.44 ;
      RECT 21.036 30.48 21.352 30.96 ;
      RECT 21.036 30 21.442 30.48 ;
      RECT 21.036 29.52 21.352 30 ;
      RECT 20.858 29.04 21.352 29.52 ;
      RECT 21.036 28.56 21.352 29.04 ;
      RECT 21.036 28.08 21.442 28.56 ;
      RECT 21.036 27.6 21.352 28.08 ;
      RECT 20.858 27.12 21.352 27.6 ;
      RECT 21.292 26.64 21.352 27.12 ;
      RECT 21.292 25.68 21.442 26.64 ;
      RECT 20.858 24.96 21.442 25.68 ;
      RECT 21.208 23.52 21.442 24.96 ;
      RECT 20.858 22.08 21.442 23.52 ;
      RECT 19.958 45.36 20.542 46.08 ;
      RECT 20.136 44.4 20.542 45.36 ;
      RECT 20.136 43.92 20.364 44.4 ;
      RECT 19.958 43.44 20.364 43.92 ;
      RECT 20.136 42.96 20.364 43.44 ;
      RECT 20.136 42.48 20.542 42.96 ;
      RECT 20.136 42 20.364 42.48 ;
      RECT 19.958 41.52 20.364 42 ;
      RECT 20.136 41.04 20.364 41.52 ;
      RECT 20.136 40.56 20.542 41.04 ;
      RECT 20.136 40.08 20.364 40.56 ;
      RECT 19.958 39.6 20.364 40.08 ;
      RECT 20.136 39.12 20.364 39.6 ;
      RECT 20.136 38.64 20.542 39.12 ;
      RECT 20.136 38.16 20.364 38.64 ;
      RECT 19.958 37.68 20.364 38.16 ;
      RECT 20.136 37.2 20.364 37.68 ;
      RECT 20.136 36.72 20.542 37.2 ;
      RECT 20.136 36.24 20.364 36.72 ;
      RECT 19.958 35.76 20.364 36.24 ;
      RECT 20.136 35.28 20.364 35.76 ;
      RECT 20.136 34.8 20.542 35.28 ;
      RECT 20.136 34.32 20.364 34.8 ;
      RECT 19.958 33.84 20.364 34.32 ;
      RECT 20.136 33.36 20.364 33.84 ;
      RECT 20.136 32.88 20.542 33.36 ;
      RECT 20.136 32.4 20.364 32.88 ;
      RECT 19.958 31.92 20.364 32.4 ;
      RECT 20.136 31.44 20.364 31.92 ;
      RECT 20.136 30.96 20.542 31.44 ;
      RECT 20.136 30.48 20.364 30.96 ;
      RECT 19.958 30 20.364 30.48 ;
      RECT 20.136 29.52 20.364 30 ;
      RECT 20.136 29.04 20.542 29.52 ;
      RECT 20.136 28.56 20.364 29.04 ;
      RECT 19.958 28.08 20.364 28.56 ;
      RECT 20.136 27.6 20.364 28.08 ;
      RECT 20.136 27.12 20.542 27.6 ;
      RECT 20.136 26.64 20.364 27.12 ;
      RECT 19.958 25.68 20.364 26.64 ;
      RECT 19.958 24.96 20.542 25.68 ;
      RECT 20.136 23.52 20.542 24.96 ;
      RECT 19.958 22.08 20.542 23.52 ;
      RECT 20.136 20.64 20.542 22.08 ;
      RECT 19.958 19.92 20.542 20.64 ;
      RECT 19.958 18.48 20.108 19.92 ;
      RECT 19.958 18 20.542 18.48 ;
      RECT 19.958 16.56 20.108 18 ;
      RECT 19.958 16.08 20.542 16.56 ;
      RECT 19.958 14.64 20.108 16.08 ;
      RECT 19.958 14.16 20.542 14.64 ;
      RECT 19.958 12.72 20.108 14.16 ;
      RECT 19.958 12.24 20.542 12.72 ;
      RECT 19.958 10.8 20.108 12.24 ;
      RECT 19.958 10.32 20.542 10.8 ;
      RECT 19.958 8.88 20.108 10.32 ;
      RECT 19.958 8.4 20.542 8.88 ;
      RECT 19.958 6.96 20.108 8.4 ;
      RECT 19.958 6.48 20.542 6.96 ;
      RECT 19.958 5.04 20.108 6.48 ;
      RECT 19.958 4.56 20.542 5.04 ;
      RECT 19.958 3.12 20.108 4.56 ;
      RECT 19.958 2.64 20.542 3.12 ;
      RECT 19.958 1.2 20.108 2.64 ;
      RECT 19.958 0 20.542 1.2 ;
      RECT 19.058 45.36 19.642 46.08 ;
      RECT 19.408 44.4 19.642 45.36 ;
      RECT 19.408 43.92 19.464 44.4 ;
      RECT 19.058 43.44 19.464 43.92 ;
      RECT 19.408 42.96 19.464 43.44 ;
      RECT 19.408 42.48 19.642 42.96 ;
      RECT 19.408 42 19.464 42.48 ;
      RECT 19.058 41.52 19.464 42 ;
      RECT 19.408 41.04 19.464 41.52 ;
      RECT 19.408 40.56 19.642 41.04 ;
      RECT 19.408 40.08 19.464 40.56 ;
      RECT 19.058 39.6 19.464 40.08 ;
      RECT 19.408 39.12 19.464 39.6 ;
      RECT 19.408 38.64 19.642 39.12 ;
      RECT 19.408 38.16 19.464 38.64 ;
      RECT 19.058 37.68 19.464 38.16 ;
      RECT 19.408 37.2 19.464 37.68 ;
      RECT 19.408 36.72 19.642 37.2 ;
      RECT 19.408 36.24 19.464 36.72 ;
      RECT 19.058 35.76 19.464 36.24 ;
      RECT 19.408 35.28 19.464 35.76 ;
      RECT 19.408 34.8 19.642 35.28 ;
      RECT 19.408 34.32 19.464 34.8 ;
      RECT 19.058 33.84 19.464 34.32 ;
      RECT 19.408 33.36 19.464 33.84 ;
      RECT 19.408 32.88 19.642 33.36 ;
      RECT 19.408 32.4 19.464 32.88 ;
      RECT 19.058 31.92 19.464 32.4 ;
      RECT 19.408 31.44 19.464 31.92 ;
      RECT 19.408 30.96 19.642 31.44 ;
      RECT 19.408 30.48 19.464 30.96 ;
      RECT 19.058 30 19.464 30.48 ;
      RECT 19.408 29.52 19.464 30 ;
      RECT 19.408 29.04 19.642 29.52 ;
      RECT 19.408 28.56 19.464 29.04 ;
      RECT 19.058 28.08 19.464 28.56 ;
      RECT 19.408 27.6 19.464 28.08 ;
      RECT 19.408 27.12 19.642 27.6 ;
      RECT 19.408 26.64 19.464 27.12 ;
      RECT 19.058 25.68 19.464 26.64 ;
      RECT 19.058 24.96 19.642 25.68 ;
      RECT 19.408 23.52 19.552 24.96 ;
      RECT 19.058 22.08 19.642 23.52 ;
      RECT 19.408 20.64 19.552 22.08 ;
      RECT 19.058 19.92 19.642 20.64 ;
      RECT 19.058 18.96 19.292 19.92 ;
      RECT 19.148 18.48 19.292 18.96 ;
      RECT 19.148 18 19.642 18.48 ;
      RECT 19.148 17.52 19.292 18 ;
      RECT 19.058 17.04 19.292 17.52 ;
      RECT 19.148 16.56 19.292 17.04 ;
      RECT 19.148 16.08 19.642 16.56 ;
      RECT 19.148 15.6 19.292 16.08 ;
      RECT 19.058 15.12 19.292 15.6 ;
      RECT 19.148 14.64 19.292 15.12 ;
      RECT 19.148 14.16 19.642 14.64 ;
      RECT 19.148 13.68 19.292 14.16 ;
      RECT 19.058 13.2 19.292 13.68 ;
      RECT 19.148 12.72 19.292 13.2 ;
      RECT 19.148 12.24 19.642 12.72 ;
      RECT 19.148 11.76 19.292 12.24 ;
      RECT 19.058 11.28 19.292 11.76 ;
      RECT 19.148 10.8 19.292 11.28 ;
      RECT 19.148 10.32 19.642 10.8 ;
      RECT 19.148 9.84 19.292 10.32 ;
      RECT 19.058 9.36 19.292 9.84 ;
      RECT 19.148 8.88 19.292 9.36 ;
      RECT 19.148 8.4 19.642 8.88 ;
      RECT 19.148 7.92 19.292 8.4 ;
      RECT 19.058 7.44 19.292 7.92 ;
      RECT 19.148 6.96 19.292 7.44 ;
      RECT 19.148 6.48 19.642 6.96 ;
      RECT 19.148 6 19.292 6.48 ;
      RECT 19.058 5.52 19.292 6 ;
      RECT 19.148 5.04 19.292 5.52 ;
      RECT 19.148 4.56 19.642 5.04 ;
      RECT 19.148 4.08 19.292 4.56 ;
      RECT 19.058 3.6 19.292 4.08 ;
      RECT 19.148 3.12 19.292 3.6 ;
      RECT 19.148 2.64 19.642 3.12 ;
      RECT 19.148 2.16 19.292 2.64 ;
      RECT 19.058 1.68 19.292 2.16 ;
      RECT 18.158 45.36 18.742 46.08 ;
      RECT 18.158 44.4 18.652 45.36 ;
      RECT 18.336 43.92 18.652 44.4 ;
      RECT 18.336 43.44 18.742 43.92 ;
      RECT 18.336 42.96 18.652 43.44 ;
      RECT 18.158 42.48 18.652 42.96 ;
      RECT 18.336 42 18.652 42.48 ;
      RECT 18.336 41.52 18.742 42 ;
      RECT 18.336 41.04 18.652 41.52 ;
      RECT 18.158 40.56 18.652 41.04 ;
      RECT 18.336 40.08 18.652 40.56 ;
      RECT 18.336 39.6 18.742 40.08 ;
      RECT 18.336 39.12 18.652 39.6 ;
      RECT 18.158 38.64 18.652 39.12 ;
      RECT 18.336 38.16 18.652 38.64 ;
      RECT 18.336 37.68 18.742 38.16 ;
      RECT 18.336 37.2 18.652 37.68 ;
      RECT 18.158 36.72 18.652 37.2 ;
      RECT 18.336 36.24 18.652 36.72 ;
      RECT 18.336 35.76 18.742 36.24 ;
      RECT 18.336 35.28 18.652 35.76 ;
      RECT 18.158 34.8 18.652 35.28 ;
      RECT 18.336 34.32 18.652 34.8 ;
      RECT 18.336 33.84 18.742 34.32 ;
      RECT 18.336 33.36 18.652 33.84 ;
      RECT 18.158 32.88 18.652 33.36 ;
      RECT 18.336 32.4 18.652 32.88 ;
      RECT 18.336 31.92 18.742 32.4 ;
      RECT 18.336 31.44 18.652 31.92 ;
      RECT 18.158 30.96 18.652 31.44 ;
      RECT 18.336 30.48 18.652 30.96 ;
      RECT 18.336 30 18.742 30.48 ;
      RECT 18.336 29.52 18.652 30 ;
      RECT 18.158 29.04 18.652 29.52 ;
      RECT 18.336 28.56 18.652 29.04 ;
      RECT 18.336 28.08 18.742 28.56 ;
      RECT 18.336 27.6 18.652 28.08 ;
      RECT 18.158 27.12 18.652 27.6 ;
      RECT 18.508 26.64 18.652 27.12 ;
      RECT 18.508 25.68 18.742 26.64 ;
      RECT 18.158 24.96 18.742 25.68 ;
      RECT 17.258 44.4 17.842 46.08 ;
      RECT 17.436 42.96 17.752 44.4 ;
      RECT 17.258 42.48 17.842 42.96 ;
      RECT 17.436 41.04 17.752 42.48 ;
      RECT 17.258 40.56 17.842 41.04 ;
      RECT 17.436 39.12 17.752 40.56 ;
      RECT 17.258 38.64 17.842 39.12 ;
      RECT 17.436 37.2 17.752 38.64 ;
      RECT 17.258 36.72 17.842 37.2 ;
      RECT 17.436 35.28 17.752 36.72 ;
      RECT 17.258 34.8 17.842 35.28 ;
      RECT 17.436 33.36 17.752 34.8 ;
      RECT 17.258 32.88 17.842 33.36 ;
      RECT 17.436 31.44 17.752 32.88 ;
      RECT 17.258 30.96 17.842 31.44 ;
      RECT 17.436 29.52 17.752 30.96 ;
      RECT 17.258 29.04 17.842 29.52 ;
      RECT 17.436 27.6 17.752 29.04 ;
      RECT 17.258 27.12 17.842 27.6 ;
      RECT 17.436 25.68 17.752 27.12 ;
      RECT 17.258 24.96 17.842 25.68 ;
      RECT 17.776 23.52 17.842 24.96 ;
      RECT 17.258 22.08 17.842 23.52 ;
      RECT 17.776 20.64 17.842 22.08 ;
      RECT 17.258 19.92 17.842 20.64 ;
      RECT 17.258 18.96 17.752 19.92 ;
      RECT 17.692 18.48 17.752 18.96 ;
      RECT 17.692 18 17.842 18.48 ;
      RECT 17.258 17.52 17.408 18.96 ;
      RECT 17.692 17.52 17.752 18 ;
      RECT 17.258 17.04 17.752 17.52 ;
      RECT 17.692 16.56 17.752 17.04 ;
      RECT 17.692 16.08 17.842 16.56 ;
      RECT 17.258 15.6 17.408 17.04 ;
      RECT 17.692 15.6 17.752 16.08 ;
      RECT 17.258 15.12 17.752 15.6 ;
      RECT 17.692 14.64 17.752 15.12 ;
      RECT 17.692 14.16 17.842 14.64 ;
      RECT 17.258 13.68 17.408 15.12 ;
      RECT 17.692 13.68 17.752 14.16 ;
      RECT 17.258 13.2 17.752 13.68 ;
      RECT 17.692 12.72 17.752 13.2 ;
      RECT 17.692 12.24 17.842 12.72 ;
      RECT 17.258 11.76 17.408 13.2 ;
      RECT 17.692 11.76 17.752 12.24 ;
      RECT 17.258 11.28 17.752 11.76 ;
      RECT 17.692 10.8 17.752 11.28 ;
      RECT 17.692 10.32 17.842 10.8 ;
      RECT 17.258 9.84 17.408 11.28 ;
      RECT 17.692 9.84 17.752 10.32 ;
      RECT 17.258 9.36 17.752 9.84 ;
      RECT 17.692 8.88 17.752 9.36 ;
      RECT 17.692 8.4 17.842 8.88 ;
      RECT 17.258 7.92 17.408 9.36 ;
      RECT 17.692 7.92 17.752 8.4 ;
      RECT 17.258 7.44 17.752 7.92 ;
      RECT 17.692 6.96 17.752 7.44 ;
      RECT 17.692 6.48 17.842 6.96 ;
      RECT 17.258 6 17.408 7.44 ;
      RECT 17.692 6 17.752 6.48 ;
      RECT 17.258 5.52 17.752 6 ;
      RECT 17.692 5.04 17.752 5.52 ;
      RECT 17.692 4.56 17.842 5.04 ;
      RECT 17.258 4.08 17.408 5.52 ;
      RECT 17.692 4.08 17.752 4.56 ;
      RECT 17.258 3.6 17.752 4.08 ;
      RECT 17.692 3.12 17.752 3.6 ;
      RECT 17.258 2.64 17.408 3.6 ;
      RECT 17.692 2.64 17.842 3.12 ;
      RECT 17.348 2.16 17.408 2.64 ;
      RECT 17.692 2.16 17.752 2.64 ;
      RECT 17.348 1.2 17.752 2.16 ;
      RECT 17.258 0 17.842 1.2 ;
      RECT 16.358 44.4 16.942 46.08 ;
      RECT 16.358 42.96 16.764 44.4 ;
      RECT 16.358 42.48 16.942 42.96 ;
      RECT 16.358 41.04 16.764 42.48 ;
      RECT 16.358 40.56 16.942 41.04 ;
      RECT 16.358 39.12 16.764 40.56 ;
      RECT 16.358 38.64 16.942 39.12 ;
      RECT 16.358 37.2 16.764 38.64 ;
      RECT 16.358 36.72 16.942 37.2 ;
      RECT 16.358 35.28 16.764 36.72 ;
      RECT 16.358 34.8 16.942 35.28 ;
      RECT 16.358 33.36 16.764 34.8 ;
      RECT 16.358 32.88 16.942 33.36 ;
      RECT 16.358 31.44 16.764 32.88 ;
      RECT 16.358 30.96 16.942 31.44 ;
      RECT 16.358 29.52 16.764 30.96 ;
      RECT 16.358 29.04 16.942 29.52 ;
      RECT 16.358 27.6 16.764 29.04 ;
      RECT 16.358 27.12 16.942 27.6 ;
      RECT 16.358 25.68 16.592 27.12 ;
      RECT 16.358 24.96 16.942 25.68 ;
      RECT 16.536 23.52 16.942 24.96 ;
      RECT 16.358 22.08 16.942 23.52 ;
      RECT 16.536 20.64 16.942 22.08 ;
      RECT 16.358 19.92 16.942 20.64 ;
      RECT 16.358 18.48 16.508 19.92 ;
      RECT 16.358 18 16.942 18.48 ;
      RECT 16.358 16.56 16.508 18 ;
      RECT 16.358 16.08 16.942 16.56 ;
      RECT 16.358 14.64 16.508 16.08 ;
      RECT 16.358 14.16 16.942 14.64 ;
      RECT 16.358 12.72 16.508 14.16 ;
      RECT 16.358 12.24 16.942 12.72 ;
      RECT 16.358 10.8 16.508 12.24 ;
      RECT 16.358 10.32 16.942 10.8 ;
      RECT 16.358 8.88 16.508 10.32 ;
      RECT 16.358 8.4 16.942 8.88 ;
      RECT 16.358 6.96 16.508 8.4 ;
      RECT 16.358 6.48 16.942 6.96 ;
      RECT 16.358 5.04 16.508 6.48 ;
      RECT 16.358 4.56 16.942 5.04 ;
      RECT 16.358 3.12 16.508 4.56 ;
      RECT 16.358 2.64 16.942 3.12 ;
      RECT 16.358 1.68 16.592 2.64 ;
      RECT 15.458 45.36 16.042 46.08 ;
      RECT 14.558 45.36 15.142 46.08 ;
      RECT 14.558 43.92 14.964 45.36 ;
      RECT 14.558 43.44 15.142 43.92 ;
      RECT 14.558 42 14.964 43.44 ;
      RECT 14.558 41.52 15.142 42 ;
      RECT 14.558 40.08 14.964 41.52 ;
      RECT 14.558 39.6 15.142 40.08 ;
      RECT 14.558 38.16 14.964 39.6 ;
      RECT 14.558 37.68 15.142 38.16 ;
      RECT 14.558 36.24 14.964 37.68 ;
      RECT 14.558 35.76 15.142 36.24 ;
      RECT 14.558 34.32 14.964 35.76 ;
      RECT 14.558 33.84 15.142 34.32 ;
      RECT 14.558 32.4 14.964 33.84 ;
      RECT 14.558 31.92 15.142 32.4 ;
      RECT 14.558 30.48 14.964 31.92 ;
      RECT 14.558 30 15.142 30.48 ;
      RECT 14.558 28.56 14.964 30 ;
      RECT 14.558 28.08 15.142 28.56 ;
      RECT 14.558 26.64 14.964 28.08 ;
      RECT 14.558 24.96 15.142 26.64 ;
      RECT 13.658 44.4 14.242 46.08 ;
      RECT 13.658 42.96 13.724 44.4 ;
      RECT 13.658 42.48 14.242 42.96 ;
      RECT 13.658 41.04 13.724 42.48 ;
      RECT 13.658 40.56 14.242 41.04 ;
      RECT 13.658 39.12 13.724 40.56 ;
      RECT 13.658 38.64 14.242 39.12 ;
      RECT 13.658 37.2 13.724 38.64 ;
      RECT 13.658 36.72 14.242 37.2 ;
      RECT 13.658 35.28 13.724 36.72 ;
      RECT 13.658 34.8 14.242 35.28 ;
      RECT 13.658 33.36 13.724 34.8 ;
      RECT 13.658 32.88 14.242 33.36 ;
      RECT 13.658 31.44 13.724 32.88 ;
      RECT 13.658 30.96 14.242 31.44 ;
      RECT 13.658 29.52 13.724 30.96 ;
      RECT 13.658 29.04 14.242 29.52 ;
      RECT 13.658 27.6 13.724 29.04 ;
      RECT 13.658 27.12 14.242 27.6 ;
      RECT 13.658 25.68 13.724 27.12 ;
      RECT 13.658 24.96 14.242 25.68 ;
      RECT 13.748 23.52 14.152 24.96 ;
      RECT 13.658 22.08 14.242 23.52 ;
      RECT 13.748 20.64 14.152 22.08 ;
      RECT 13.658 19.92 14.242 20.64 ;
      RECT 14.176 18.48 14.242 19.92 ;
      RECT 13.658 18 14.242 18.48 ;
      RECT 14.176 16.56 14.242 18 ;
      RECT 13.658 16.08 14.242 16.56 ;
      RECT 14.176 14.64 14.242 16.08 ;
      RECT 13.658 14.16 14.242 14.64 ;
      RECT 14.176 12.72 14.242 14.16 ;
      RECT 13.658 12.24 14.242 12.72 ;
      RECT 14.176 10.8 14.242 12.24 ;
      RECT 13.658 10.32 14.242 10.8 ;
      RECT 14.176 8.88 14.242 10.32 ;
      RECT 13.658 8.4 14.242 8.88 ;
      RECT 14.176 6.96 14.242 8.4 ;
      RECT 13.658 6.48 14.242 6.96 ;
      RECT 14.176 5.04 14.242 6.48 ;
      RECT 13.658 4.56 14.242 5.04 ;
      RECT 14.176 3.12 14.242 4.56 ;
      RECT 13.658 2.64 14.242 3.12 ;
      RECT 13.658 1.68 14.064 2.64 ;
      RECT 12.758 0 13.342 46.08 ;
      RECT 11.858 0 12.442 46.08 ;
      RECT 10.958 0 11.542 46.08 ;
      RECT 10.058 0 10.642 46.08 ;
      RECT 9.158 0 9.742 46.08 ;
      RECT 8.258 0 8.842 46.08 ;
      RECT 7.358 0 7.942 46.08 ;
      RECT 6.458 0 7.042 46.08 ;
      RECT 5.558 0 6.142 46.08 ;
      RECT 4.658 0 5.242 46.08 ;
      RECT 3.758 0 4.342 46.08 ;
      RECT 2.858 0 3.442 46.08 ;
      RECT 1.958 0 2.542 46.08 ;
      RECT 1.058 0 1.642 46.08 ;
      RECT 0.08 0 0.742 46.08 ;
      RECT 15.458 43.44 16.042 43.92 ;
      RECT 15.458 41.52 16.042 42 ;
      RECT 15.458 39.6 16.042 40.08 ;
      RECT 15.458 37.68 16.042 38.16 ;
      RECT 15.458 35.76 16.042 36.24 ;
      RECT 15.458 33.84 16.042 34.32 ;
      RECT 15.458 31.92 16.042 32.4 ;
      RECT 15.458 30 16.042 30.48 ;
      RECT 15.458 28.08 16.042 28.56 ;
      RECT 15.458 24.96 16.042 26.64 ;
      RECT 18.158 22.08 18.742 23.52 ;
      RECT 15.458 22.08 16.042 23.52 ;
      RECT 14.558 22.08 15.142 23.52 ;
      RECT 20.858 18.96 21.442 20.64 ;
      RECT 20.858 17.52 21.264 18.96 ;
      RECT 20.858 17.04 21.442 17.52 ;
      RECT 20.858 15.6 21.264 17.04 ;
      RECT 20.858 15.12 21.442 15.6 ;
      RECT 20.858 13.68 21.264 15.12 ;
      RECT 20.858 13.2 21.442 13.68 ;
      RECT 20.858 11.76 21.264 13.2 ;
      RECT 20.858 11.28 21.442 11.76 ;
      RECT 20.858 9.84 21.264 11.28 ;
      RECT 20.858 9.36 21.442 9.84 ;
      RECT 20.858 7.92 21.264 9.36 ;
      RECT 20.858 7.44 21.442 7.92 ;
      RECT 20.858 6 21.264 7.44 ;
      RECT 20.858 5.52 21.442 6 ;
      RECT 20.858 4.08 21.264 5.52 ;
      RECT 20.858 3.6 21.442 4.08 ;
      RECT 20.858 2.16 21.264 3.6 ;
      RECT 20.858 1.68 21.442 2.16 ;
      RECT 20.858 0.24 21.264 1.68 ;
      RECT 20.858 0 21.442 0.24 ;
      RECT 18.158 19.92 18.742 20.64 ;
      RECT 18.248 18.96 18.742 19.92 ;
      RECT 18.248 18.48 18.392 18.96 ;
      RECT 18.158 18 18.392 18.48 ;
      RECT 18.248 17.52 18.392 18 ;
      RECT 18.248 17.04 18.742 17.52 ;
      RECT 18.248 16.56 18.392 17.04 ;
      RECT 18.158 16.08 18.392 16.56 ;
      RECT 18.248 15.6 18.392 16.08 ;
      RECT 18.248 15.12 18.742 15.6 ;
      RECT 18.248 14.64 18.392 15.12 ;
      RECT 18.158 14.16 18.392 14.64 ;
      RECT 18.248 13.68 18.392 14.16 ;
      RECT 18.248 13.2 18.742 13.68 ;
      RECT 18.248 12.72 18.392 13.2 ;
      RECT 18.158 12.24 18.392 12.72 ;
      RECT 18.248 11.76 18.392 12.24 ;
      RECT 18.248 11.28 18.742 11.76 ;
      RECT 18.248 10.8 18.392 11.28 ;
      RECT 18.158 10.32 18.392 10.8 ;
      RECT 18.248 9.84 18.392 10.32 ;
      RECT 18.248 9.36 18.742 9.84 ;
      RECT 18.248 8.88 18.392 9.36 ;
      RECT 18.158 8.4 18.392 8.88 ;
      RECT 18.248 7.92 18.392 8.4 ;
      RECT 18.248 7.44 18.742 7.92 ;
      RECT 18.248 6.96 18.392 7.44 ;
      RECT 18.158 6.48 18.392 6.96 ;
      RECT 18.248 6 18.392 6.48 ;
      RECT 18.248 5.52 18.742 6 ;
      RECT 18.248 5.04 18.392 5.52 ;
      RECT 18.158 4.56 18.392 5.04 ;
      RECT 18.248 4.08 18.392 4.56 ;
      RECT 18.248 3.6 18.742 4.08 ;
      RECT 18.248 3.12 18.392 3.6 ;
      RECT 18.158 2.64 18.392 3.12 ;
      RECT 18.248 2.16 18.392 2.64 ;
      RECT 18.248 1.68 18.742 2.16 ;
      RECT 18.248 1.2 18.652 1.68 ;
      RECT 18.158 0.24 18.652 1.2 ;
      RECT 18.158 0 18.742 0.24 ;
      RECT 15.458 18.96 16.042 20.64 ;
      RECT 15.548 17.52 15.608 18.96 ;
      RECT 15.458 17.04 16.042 17.52 ;
      RECT 15.548 15.6 15.608 17.04 ;
      RECT 15.458 15.12 16.042 15.6 ;
      RECT 15.548 13.68 15.608 15.12 ;
      RECT 15.458 13.2 16.042 13.68 ;
      RECT 15.548 11.76 15.608 13.2 ;
      RECT 15.458 11.28 16.042 11.76 ;
      RECT 15.548 9.84 15.608 11.28 ;
      RECT 15.458 9.36 16.042 9.84 ;
      RECT 15.548 7.92 15.608 9.36 ;
      RECT 15.458 7.44 16.042 7.92 ;
      RECT 15.548 6 15.608 7.44 ;
      RECT 15.458 5.52 16.042 6 ;
      RECT 15.548 4.08 15.608 5.52 ;
      RECT 15.458 3.6 16.042 4.08 ;
      RECT 15.548 2.16 15.608 3.6 ;
      RECT 15.458 1.68 16.042 2.16 ;
      RECT 15.458 0.24 15.952 1.68 ;
      RECT 15.458 0 16.042 0.24 ;
      RECT 14.558 18.96 15.142 20.64 ;
      RECT 14.558 17.52 14.792 18.96 ;
      RECT 14.558 17.04 15.142 17.52 ;
      RECT 14.558 15.6 14.792 17.04 ;
      RECT 14.558 15.12 15.142 15.6 ;
      RECT 14.558 13.68 14.792 15.12 ;
      RECT 14.558 13.2 15.142 13.68 ;
      RECT 14.558 11.76 14.792 13.2 ;
      RECT 14.558 11.28 15.142 11.76 ;
      RECT 14.558 9.84 14.792 11.28 ;
      RECT 14.558 9.36 15.142 9.84 ;
      RECT 14.558 7.92 14.792 9.36 ;
      RECT 14.558 7.44 15.142 7.92 ;
      RECT 14.558 6 14.792 7.44 ;
      RECT 14.558 5.52 15.142 6 ;
      RECT 14.558 4.08 14.792 5.52 ;
      RECT 14.558 3.6 15.142 4.08 ;
      RECT 14.558 2.64 14.792 3.6 ;
      RECT 14.736 2.16 14.792 2.64 ;
      RECT 14.736 1.2 15.142 2.16 ;
      RECT 14.558 0 15.142 1.2 ;
      RECT 19.408 0.24 19.642 1.2 ;
      RECT 19.058 0 19.642 0.24 ;
      RECT 16.708 0.24 16.942 1.2 ;
      RECT 16.358 0 16.942 0.24 ;
      RECT 14.092 0.24 14.242 1.2 ;
      RECT 13.658 0 14.242 0.24 ;
    LAYER m0 ;
      RECT 0 0.002 37.8 46.078 ;
    LAYER m1 ;
      RECT 0 0 37.8 46.08 ;
    LAYER m2 ;
      RECT 0 0.015 37.8 46.065 ;
    LAYER m3 ;
      RECT 0.015 0 37.785 46.08 ;
    LAYER m4 ;
      RECT 0 0.02 37.8 46.06 ;
    LAYER m5 ;
      RECT 0.012 0 37.788 46.08 ;
    LAYER m6 ;
      RECT 0 0.012 37.8 46.068 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf156b040e2r2w0cbbehbaa4acw

END LIBRARY
