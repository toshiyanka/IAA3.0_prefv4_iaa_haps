// Create a constraint class
// Arg 1: Unique class name
// Arg 2: Name of picker to apply constraints to
// Arg 3: Instance name of picker - can be anything you choose to reference the picker instance
`constraint_wrapper_class_begin(test_constraints)
`constraint_wrapper_class_end






