VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf066b128e2r1w0cbbehsaa4acw
  CLASS BLOCK ;
  FOREIGN arf066b128e2r1w0cbbehsaa4acw ;
  ORIGIN 0 0 ;
  SIZE 45 BY 22.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 11.16 0.388 12.36 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 11.16 4.156 12.36 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 9 0.388 10.2 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 11.16 1.928 12.36 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 11.16 2.188 12.36 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 11.16 2.356 12.36 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 11.16 2.616 12.36 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 11.16 2.916 12.36 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 11.16 3.172 12.36 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 11.16 3.988 12.36 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 11.16 0.556 12.36 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 11.16 0.816 12.36 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 11.16 5.528 12.36 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 11.16 5.788 12.36 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 11.16 5.956 12.36 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 11.16 6.216 12.36 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 11.16 6.516 12.36 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 11.16 0.472 12.36 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 11.16 0.728 12.36 ;
    END
  END rdaddrp1[6]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 11.16 4.416 12.36 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 11.16 4.716 12.36 ;
    END
  END rdaddrp1_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 11.16 1.116 12.36 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 11.16 4.972 12.36 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 11.16 1.628 12.36 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 11.16 5.228 12.36 ;
    END
  END sdl_initp1
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 9 2.188 10.2 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 9 2.356 10.2 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 9 2.916 10.2 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 9 3.172 10.2 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 9 3.988 10.2 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 9 4.156 10.2 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 9 4.416 10.2 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 9 0.556 10.2 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 9 0.816 10.2 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.244 0.12 1.288 1.32 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 2.52 2.356 3.72 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.52 2.528 3.72 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 3 1.628 4.2 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 3 1.716 4.2 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.48 2.616 4.68 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 3.48 2.828 4.68 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 3.96 1.372 5.16 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 3.96 1.456 5.16 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 4.44 2.356 5.64 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 4.44 2.528 5.64 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 0.12 1.372 1.32 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 4.92 1.628 6.12 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 4.92 1.716 6.12 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.4 2.616 6.6 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.4 2.828 6.6 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 5.88 1.372 7.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 5.88 1.456 7.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 6.36 2.356 7.56 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6.36 2.528 7.56 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 6.84 1.628 8.04 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 6.84 1.716 8.04 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.6 2.272 1.8 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 7.32 2.616 8.52 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 7.32 2.828 8.52 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 7.8 1.372 9 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 7.8 1.456 9 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 13.08 2.828 14.28 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 13.08 1.716 14.28 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 13.56 1.372 14.76 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 13.56 1.456 14.76 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 14.04 2.528 15.24 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.04 2.616 15.24 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 0.6 2.356 1.8 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 14.52 1.628 15.72 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 14.52 1.716 15.72 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 15 2.356 16.2 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 15 2.828 16.2 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 15.48 1.372 16.68 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 15.48 1.456 16.68 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 15.96 2.528 17.16 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 15.96 2.616 17.16 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 16.44 1.628 17.64 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 16.44 1.716 17.64 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 1.08 1.628 2.28 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 16.92 2.356 18.12 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 16.92 2.828 18.12 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 17.4 1.372 18.6 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 17.4 1.456 18.6 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 17.88 2.528 19.08 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 17.88 2.616 19.08 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 18.36 1.628 19.56 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 18.36 1.716 19.56 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 18.84 2.356 20.04 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 18.84 2.828 20.04 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 1.08 1.716 2.28 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 19.32 1.372 20.52 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 19.32 1.456 20.52 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 19.8 2.528 21 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.8 2.616 21 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 20.28 1.628 21.48 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 20.28 1.716 21.48 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 20.76 2.356 21.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 20.76 2.828 21.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 1.56 2.616 2.76 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 1.56 2.828 2.76 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 2.04 1.372 3.24 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 2.04 1.456 3.24 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 9 1.628 10.2 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 9 1.928 10.2 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 9 1.116 10.2 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 0.12 3.256 1.32 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 2.52 4.716 3.72 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 2.52 4.888 3.72 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 3 3.988 4.2 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 3 4.072 4.2 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 3.48 5.228 4.68 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 3.48 5.316 4.68 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 3.96 3.428 5.16 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.96 3.516 5.16 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 4.44 4.716 5.64 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 4.44 4.888 5.64 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.12 3.428 1.32 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 4.92 3.988 6.12 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 4.92 4.072 6.12 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 5.4 5.228 6.6 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 5.4 5.316 6.6 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 5.88 3.428 7.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.88 3.516 7.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 6.36 4.716 7.56 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 6.36 4.888 7.56 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 6.84 3.988 8.04 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.84 4.072 8.04 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 0.6 4.628 1.8 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 7.32 5.228 8.52 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 7.32 5.316 8.52 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 7.8 3.428 9 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.8 3.516 9 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 13.08 4.072 14.28 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 13.08 4.328 14.28 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 13.56 3.516 14.76 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 13.56 3.728 14.76 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 14.04 5.228 15.24 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 14.04 5.316 15.24 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 0.6 4.716 1.8 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 14.52 3.428 15.72 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 14.52 3.988 15.72 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 15 4.716 16.2 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 15 4.888 16.2 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 15.48 3.516 16.68 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 15.48 3.728 16.68 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 15.96 5.228 17.16 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 15.96 5.316 17.16 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.44 3.428 17.64 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 16.44 3.988 17.64 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 1.08 3.988 2.28 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 16.92 4.716 18.12 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 16.92 4.888 18.12 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 17.4 3.516 18.6 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 17.4 3.728 18.6 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 17.88 5.228 19.08 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 17.88 5.316 19.08 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 18.36 3.428 19.56 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 18.36 3.988 19.56 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 18.84 4.716 20.04 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 18.84 4.888 20.04 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 1.08 4.072 2.28 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.32 3.516 20.52 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 19.32 3.728 20.52 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 19.8 5.228 21 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 19.8 5.316 21 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.28 3.428 21.48 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 20.28 3.988 21.48 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 20.76 4.716 21.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 20.76 4.888 21.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 1.56 5.228 2.76 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 1.56 5.316 2.76 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.04 3.428 3.24 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 2.04 3.516 3.24 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 0.12 3.516 1.32 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 2.52 4.972 3.72 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 2.52 5.056 3.72 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 3 4.156 4.2 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 3 4.328 4.2 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 3.48 5.528 4.68 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 3.48 5.616 4.68 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.96 3.728 5.16 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 3.96 3.816 5.16 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 4.44 4.972 5.64 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 4.44 5.056 5.64 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.12 3.728 1.32 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 4.92 4.156 6.12 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 4.92 4.328 6.12 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 5.4 5.528 6.6 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 5.4 5.616 6.6 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 5.88 3.728 7.08 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 5.88 3.816 7.08 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 6.36 4.972 7.56 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 6.36 5.056 7.56 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 6.84 4.156 8.04 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6.84 4.328 8.04 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 0.6 4.888 1.8 ;
    END
  END rddatap1[2]
  PIN rddatap1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 7.32 5.528 8.52 ;
    END
  END rddatap1[30]
  PIN rddatap1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 7.32 5.616 8.52 ;
    END
  END rddatap1[31]
  PIN rddatap1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 7.8 3.728 9 ;
    END
  END rddatap1[32]
  PIN rddatap1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 7.8 3.816 9 ;
    END
  END rddatap1[33]
  PIN rddatap1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 13.08 4.628 14.28 ;
    END
  END rddatap1[34]
  PIN rddatap1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 13.08 4.888 14.28 ;
    END
  END rddatap1[35]
  PIN rddatap1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 13.56 3.816 14.76 ;
    END
  END rddatap1[36]
  PIN rddatap1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 13.56 5.056 14.76 ;
    END
  END rddatap1[37]
  PIN rddatap1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 14.04 5.528 15.24 ;
    END
  END rddatap1[38]
  PIN rddatap1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 14.04 5.616 15.24 ;
    END
  END rddatap1[39]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 0.6 4.972 1.8 ;
    END
  END rddatap1[3]
  PIN rddatap1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 14.52 4.072 15.72 ;
    END
  END rddatap1[40]
  PIN rddatap1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 14.52 4.156 15.72 ;
    END
  END rddatap1[41]
  PIN rddatap1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 15 4.972 16.2 ;
    END
  END rddatap1[42]
  PIN rddatap1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 15 5.056 16.2 ;
    END
  END rddatap1[43]
  PIN rddatap1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 15.48 3.816 16.68 ;
    END
  END rddatap1[44]
  PIN rddatap1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 15.48 4.328 16.68 ;
    END
  END rddatap1[45]
  PIN rddatap1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 15.96 5.528 17.16 ;
    END
  END rddatap1[46]
  PIN rddatap1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 15.96 5.616 17.16 ;
    END
  END rddatap1[47]
  PIN rddatap1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.44 4.072 17.64 ;
    END
  END rddatap1[48]
  PIN rddatap1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 16.44 4.156 17.64 ;
    END
  END rddatap1[49]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 1.08 4.156 2.28 ;
    END
  END rddatap1[4]
  PIN rddatap1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 16.92 4.972 18.12 ;
    END
  END rddatap1[50]
  PIN rddatap1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 16.92 5.056 18.12 ;
    END
  END rddatap1[51]
  PIN rddatap1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 17.4 3.816 18.6 ;
    END
  END rddatap1[52]
  PIN rddatap1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 17.4 4.328 18.6 ;
    END
  END rddatap1[53]
  PIN rddatap1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 17.88 5.528 19.08 ;
    END
  END rddatap1[54]
  PIN rddatap1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 17.88 5.616 19.08 ;
    END
  END rddatap1[55]
  PIN rddatap1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 18.36 4.072 19.56 ;
    END
  END rddatap1[56]
  PIN rddatap1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 18.36 4.156 19.56 ;
    END
  END rddatap1[57]
  PIN rddatap1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 18.84 4.972 20.04 ;
    END
  END rddatap1[58]
  PIN rddatap1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 18.84 5.056 20.04 ;
    END
  END rddatap1[59]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 1.08 4.328 2.28 ;
    END
  END rddatap1[5]
  PIN rddatap1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 19.32 3.816 20.52 ;
    END
  END rddatap1[60]
  PIN rddatap1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 19.32 4.328 20.52 ;
    END
  END rddatap1[61]
  PIN rddatap1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 19.8 5.528 21 ;
    END
  END rddatap1[62]
  PIN rddatap1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 19.8 5.616 21 ;
    END
  END rddatap1[63]
  PIN rddatap1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 20.28 4.072 21.48 ;
    END
  END rddatap1[64]
  PIN rddatap1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 20.28 4.156 21.48 ;
    END
  END rddatap1[65]
  PIN rddatap1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 20.76 4.972 21.96 ;
    END
  END rddatap1[66]
  PIN rddatap1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 20.76 5.056 21.96 ;
    END
  END rddatap1[67]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 1.56 5.528 2.76 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 1.56 5.616 2.76 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 2.04 3.728 3.24 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 2.04 3.816 3.24 ;
    END
  END rddatap1[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 22.02 ;
        RECT 2.662 0.06 2.738 22.02 ;
        RECT 4.462 0.06 4.538 22.02 ;
        RECT 6.262 0.06 6.338 22.02 ;
        RECT 8.062 0.06 8.138 22.02 ;
        RECT 9.862 0.06 9.938 22.02 ;
        RECT 11.662 0.06 11.738 22.02 ;
        RECT 13.462 0.06 13.538 22.02 ;
        RECT 15.262 0.06 15.338 22.02 ;
        RECT 17.062 0.06 17.138 22.02 ;
        RECT 18.862 0.06 18.938 22.02 ;
        RECT 20.662 0.06 20.738 22.02 ;
        RECT 22.462 0.06 22.538 22.02 ;
        RECT 24.262 0.06 24.338 22.02 ;
        RECT 26.062 0.06 26.138 22.02 ;
        RECT 27.862 0.06 27.938 22.02 ;
        RECT 29.662 0.06 29.738 22.02 ;
        RECT 31.462 0.06 31.538 22.02 ;
        RECT 33.262 0.06 33.338 22.02 ;
        RECT 35.062 0.06 35.138 22.02 ;
        RECT 36.862 0.06 36.938 22.02 ;
        RECT 38.662 0.06 38.738 22.02 ;
        RECT 40.462 0.06 40.538 22.02 ;
        RECT 42.262 0.06 42.338 22.02 ;
        RECT 44.062 0.06 44.138 22.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 22.02 ;
        RECT 3.562 0.06 3.638 22.02 ;
        RECT 5.362 0.06 5.438 22.02 ;
        RECT 7.162 0.06 7.238 22.02 ;
        RECT 8.962 0.06 9.038 22.02 ;
        RECT 10.762 0.06 10.838 22.02 ;
        RECT 12.562 0.06 12.638 22.02 ;
        RECT 14.362 0.06 14.438 22.02 ;
        RECT 16.162 0.06 16.238 22.02 ;
        RECT 17.962 0.06 18.038 22.02 ;
        RECT 19.762 0.06 19.838 22.02 ;
        RECT 21.562 0.06 21.638 22.02 ;
        RECT 23.362 0.06 23.438 22.02 ;
        RECT 25.162 0.06 25.238 22.02 ;
        RECT 26.962 0.06 27.038 22.02 ;
        RECT 28.762 0.06 28.838 22.02 ;
        RECT 30.562 0.06 30.638 22.02 ;
        RECT 32.362 0.06 32.438 22.02 ;
        RECT 34.162 0.06 34.238 22.02 ;
        RECT 35.962 0.06 36.038 22.02 ;
        RECT 37.762 0.06 37.838 22.02 ;
        RECT 39.562 0.06 39.638 22.02 ;
        RECT 41.362 0.06 41.438 22.02 ;
        RECT 43.162 0.06 43.238 22.02 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 45.016 22.094 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 45.02 22.1 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 45.0705 22.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 45.035 22.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 45.07 22.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 45.059 22.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 45.09 22.142 ;
    LAYER m7 SPACING 0 ;
      RECT 44.138 22.14 45.04 22.2 ;
      RECT 44.138 -0.06 45.092 22.14 ;
      RECT 44.138 -0.12 45.04 -0.06 ;
      RECT 43.238 -0.12 44.062 22.2 ;
      RECT 42.338 -0.12 43.162 22.2 ;
      RECT 41.438 -0.12 42.262 22.2 ;
      RECT 40.538 -0.12 41.362 22.2 ;
      RECT 39.638 -0.12 40.462 22.2 ;
      RECT 38.738 -0.12 39.562 22.2 ;
      RECT 37.838 -0.12 38.662 22.2 ;
      RECT 36.938 -0.12 37.762 22.2 ;
      RECT 36.038 -0.12 36.862 22.2 ;
      RECT 35.138 -0.12 35.962 22.2 ;
      RECT 34.238 -0.12 35.062 22.2 ;
      RECT 33.338 -0.12 34.162 22.2 ;
      RECT 32.438 -0.12 33.262 22.2 ;
      RECT 31.538 -0.12 32.362 22.2 ;
      RECT 30.638 -0.12 31.462 22.2 ;
      RECT 29.738 -0.12 30.562 22.2 ;
      RECT 28.838 -0.12 29.662 22.2 ;
      RECT 27.938 -0.12 28.762 22.2 ;
      RECT 27.038 -0.12 27.862 22.2 ;
      RECT 26.138 -0.12 26.962 22.2 ;
      RECT 25.238 -0.12 26.062 22.2 ;
      RECT 24.338 -0.12 25.162 22.2 ;
      RECT 23.438 -0.12 24.262 22.2 ;
      RECT 22.538 -0.12 23.362 22.2 ;
      RECT 21.638 -0.12 22.462 22.2 ;
      RECT 20.738 -0.12 21.562 22.2 ;
      RECT 19.838 -0.12 20.662 22.2 ;
      RECT 18.938 -0.12 19.762 22.2 ;
      RECT 18.038 -0.12 18.862 22.2 ;
      RECT 17.138 -0.12 17.962 22.2 ;
      RECT 16.238 -0.12 17.062 22.2 ;
      RECT 15.338 -0.12 16.162 22.2 ;
      RECT 14.438 -0.12 15.262 22.2 ;
      RECT 13.538 -0.12 14.362 22.2 ;
      RECT 12.638 -0.12 13.462 22.2 ;
      RECT 11.738 -0.12 12.562 22.2 ;
      RECT 10.838 -0.12 11.662 22.2 ;
      RECT 9.938 -0.12 10.762 22.2 ;
      RECT 9.038 -0.12 9.862 22.2 ;
      RECT 8.138 -0.12 8.962 22.2 ;
      RECT 7.238 -0.12 8.062 22.2 ;
      RECT 6.338 12.36 7.162 22.2 ;
      RECT 6.338 11.16 6.472 12.36 ;
      RECT 6.516 11.16 7.162 12.36 ;
      RECT 6.338 -0.12 7.162 11.16 ;
      RECT 5.438 21 6.262 22.2 ;
      RECT 5.438 19.8 5.484 21 ;
      RECT 5.528 19.8 5.572 21 ;
      RECT 5.616 19.8 6.262 21 ;
      RECT 5.438 19.08 6.262 19.8 ;
      RECT 5.438 17.88 5.484 19.08 ;
      RECT 5.528 17.88 5.572 19.08 ;
      RECT 5.616 17.88 6.262 19.08 ;
      RECT 5.438 17.16 6.262 17.88 ;
      RECT 5.438 15.96 5.484 17.16 ;
      RECT 5.528 15.96 5.572 17.16 ;
      RECT 5.616 15.96 6.262 17.16 ;
      RECT 5.438 15.24 6.262 15.96 ;
      RECT 5.438 14.04 5.484 15.24 ;
      RECT 5.528 14.04 5.572 15.24 ;
      RECT 5.616 14.04 6.262 15.24 ;
      RECT 5.438 12.36 6.262 14.04 ;
      RECT 5.438 11.16 5.484 12.36 ;
      RECT 5.528 11.16 5.744 12.36 ;
      RECT 5.788 11.16 5.912 12.36 ;
      RECT 5.956 11.16 6.172 12.36 ;
      RECT 6.216 11.16 6.262 12.36 ;
      RECT 5.438 8.52 6.262 11.16 ;
      RECT 5.438 7.32 5.484 8.52 ;
      RECT 5.528 7.32 5.572 8.52 ;
      RECT 5.616 7.32 6.262 8.52 ;
      RECT 5.438 6.6 6.262 7.32 ;
      RECT 5.438 5.4 5.484 6.6 ;
      RECT 5.528 5.4 5.572 6.6 ;
      RECT 5.616 5.4 6.262 6.6 ;
      RECT 5.438 4.68 6.262 5.4 ;
      RECT 5.438 3.48 5.484 4.68 ;
      RECT 5.528 3.48 5.572 4.68 ;
      RECT 5.616 3.48 6.262 4.68 ;
      RECT 5.438 2.76 6.262 3.48 ;
      RECT 5.438 1.56 5.484 2.76 ;
      RECT 5.528 1.56 5.572 2.76 ;
      RECT 5.616 1.56 6.262 2.76 ;
      RECT 5.438 -0.12 6.262 1.56 ;
      RECT 4.538 21.96 5.362 22.2 ;
      RECT 5.056 21 5.362 21.96 ;
      RECT 4.538 20.76 4.672 21.96 ;
      RECT 4.716 20.76 4.844 21.96 ;
      RECT 4.888 20.76 4.928 21.96 ;
      RECT 4.972 20.76 5.012 21.96 ;
      RECT 5.056 20.76 5.184 21 ;
      RECT 4.538 20.04 5.184 20.76 ;
      RECT 5.228 19.8 5.272 21 ;
      RECT 5.316 19.8 5.362 21 ;
      RECT 5.056 19.8 5.184 20.04 ;
      RECT 5.056 19.08 5.362 19.8 ;
      RECT 4.538 18.84 4.672 20.04 ;
      RECT 4.716 18.84 4.844 20.04 ;
      RECT 4.888 18.84 4.928 20.04 ;
      RECT 4.972 18.84 5.012 20.04 ;
      RECT 5.056 18.84 5.184 19.08 ;
      RECT 4.538 18.12 5.184 18.84 ;
      RECT 5.228 17.88 5.272 19.08 ;
      RECT 5.316 17.88 5.362 19.08 ;
      RECT 5.056 17.88 5.184 18.12 ;
      RECT 5.056 17.16 5.362 17.88 ;
      RECT 4.538 16.92 4.672 18.12 ;
      RECT 4.716 16.92 4.844 18.12 ;
      RECT 4.888 16.92 4.928 18.12 ;
      RECT 4.972 16.92 5.012 18.12 ;
      RECT 5.056 16.92 5.184 17.16 ;
      RECT 4.538 16.2 5.184 16.92 ;
      RECT 5.228 15.96 5.272 17.16 ;
      RECT 5.316 15.96 5.362 17.16 ;
      RECT 5.056 15.96 5.184 16.2 ;
      RECT 5.056 15.24 5.362 15.96 ;
      RECT 4.538 15 4.672 16.2 ;
      RECT 4.716 15 4.844 16.2 ;
      RECT 4.888 15 4.928 16.2 ;
      RECT 4.972 15 5.012 16.2 ;
      RECT 5.056 15 5.184 15.24 ;
      RECT 4.538 14.76 5.184 15 ;
      RECT 4.538 14.28 5.012 14.76 ;
      RECT 5.228 14.04 5.272 15.24 ;
      RECT 5.316 14.04 5.362 15.24 ;
      RECT 5.056 14.04 5.184 14.76 ;
      RECT 4.888 13.56 5.012 14.28 ;
      RECT 5.056 13.56 5.362 14.04 ;
      RECT 4.538 13.08 4.584 14.28 ;
      RECT 4.628 13.08 4.844 14.28 ;
      RECT 4.888 13.08 5.362 13.56 ;
      RECT 4.538 12.36 5.362 13.08 ;
      RECT 4.538 11.16 4.672 12.36 ;
      RECT 4.716 11.16 4.928 12.36 ;
      RECT 4.972 11.16 5.184 12.36 ;
      RECT 5.228 11.16 5.362 12.36 ;
      RECT 4.538 8.52 5.362 11.16 ;
      RECT 4.538 7.56 5.184 8.52 ;
      RECT 5.228 7.32 5.272 8.52 ;
      RECT 5.316 7.32 5.362 8.52 ;
      RECT 5.056 7.32 5.184 7.56 ;
      RECT 5.056 6.6 5.362 7.32 ;
      RECT 4.538 6.36 4.672 7.56 ;
      RECT 4.716 6.36 4.844 7.56 ;
      RECT 4.888 6.36 4.928 7.56 ;
      RECT 4.972 6.36 5.012 7.56 ;
      RECT 5.056 6.36 5.184 6.6 ;
      RECT 4.538 5.64 5.184 6.36 ;
      RECT 5.228 5.4 5.272 6.6 ;
      RECT 5.316 5.4 5.362 6.6 ;
      RECT 5.056 5.4 5.184 5.64 ;
      RECT 5.056 4.68 5.362 5.4 ;
      RECT 4.538 4.44 4.672 5.64 ;
      RECT 4.716 4.44 4.844 5.64 ;
      RECT 4.888 4.44 4.928 5.64 ;
      RECT 4.972 4.44 5.012 5.64 ;
      RECT 5.056 4.44 5.184 4.68 ;
      RECT 4.538 3.72 5.184 4.44 ;
      RECT 5.228 3.48 5.272 4.68 ;
      RECT 5.316 3.48 5.362 4.68 ;
      RECT 5.056 3.48 5.184 3.72 ;
      RECT 5.056 2.76 5.362 3.48 ;
      RECT 4.538 2.52 4.672 3.72 ;
      RECT 4.716 2.52 4.844 3.72 ;
      RECT 4.888 2.52 4.928 3.72 ;
      RECT 4.972 2.52 5.012 3.72 ;
      RECT 5.056 2.52 5.184 2.76 ;
      RECT 4.538 1.8 5.184 2.52 ;
      RECT 5.228 1.56 5.272 2.76 ;
      RECT 5.316 1.56 5.362 2.76 ;
      RECT 4.972 1.56 5.184 1.8 ;
      RECT 4.538 0.6 4.584 1.8 ;
      RECT 4.628 0.6 4.672 1.8 ;
      RECT 4.716 0.6 4.844 1.8 ;
      RECT 4.888 0.6 4.928 1.8 ;
      RECT 4.972 0.6 5.362 1.56 ;
      RECT 4.538 -0.12 5.362 0.6 ;
      RECT 3.638 21.48 4.462 22.2 ;
      RECT 3.638 20.52 3.944 21.48 ;
      RECT 4.156 20.52 4.462 21.48 ;
      RECT 3.988 20.28 4.028 21.48 ;
      RECT 4.072 20.28 4.112 21.48 ;
      RECT 3.816 20.28 3.944 20.52 ;
      RECT 4.156 20.28 4.284 20.52 ;
      RECT 3.816 19.56 4.284 20.28 ;
      RECT 3.638 19.32 3.684 20.52 ;
      RECT 3.728 19.32 3.772 20.52 ;
      RECT 4.328 19.32 4.462 20.52 ;
      RECT 3.816 19.32 3.944 19.56 ;
      RECT 4.156 19.32 4.284 19.56 ;
      RECT 3.638 18.6 3.944 19.32 ;
      RECT 4.156 18.6 4.462 19.32 ;
      RECT 3.988 18.36 4.028 19.56 ;
      RECT 4.072 18.36 4.112 19.56 ;
      RECT 3.816 18.36 3.944 18.6 ;
      RECT 4.156 18.36 4.284 18.6 ;
      RECT 3.816 17.64 4.284 18.36 ;
      RECT 3.638 17.4 3.684 18.6 ;
      RECT 3.728 17.4 3.772 18.6 ;
      RECT 4.328 17.4 4.462 18.6 ;
      RECT 3.816 17.4 3.944 17.64 ;
      RECT 4.156 17.4 4.284 17.64 ;
      RECT 3.638 16.68 3.944 17.4 ;
      RECT 4.156 16.68 4.462 17.4 ;
      RECT 3.988 16.44 4.028 17.64 ;
      RECT 4.072 16.44 4.112 17.64 ;
      RECT 3.816 16.44 3.944 16.68 ;
      RECT 4.156 16.44 4.284 16.68 ;
      RECT 3.816 15.72 4.284 16.44 ;
      RECT 3.638 15.48 3.684 16.68 ;
      RECT 3.728 15.48 3.772 16.68 ;
      RECT 4.328 15.48 4.462 16.68 ;
      RECT 3.816 15.48 3.944 15.72 ;
      RECT 4.156 15.48 4.284 15.72 ;
      RECT 3.638 14.76 3.944 15.48 ;
      RECT 3.988 14.52 4.028 15.72 ;
      RECT 4.072 14.52 4.112 15.72 ;
      RECT 4.156 14.52 4.462 15.48 ;
      RECT 3.816 14.52 3.944 14.76 ;
      RECT 3.816 14.28 4.462 14.52 ;
      RECT 3.638 13.56 3.684 14.76 ;
      RECT 3.728 13.56 3.772 14.76 ;
      RECT 3.816 13.56 4.028 14.28 ;
      RECT 4.072 13.08 4.284 14.28 ;
      RECT 4.328 13.08 4.462 14.28 ;
      RECT 3.638 13.08 4.028 13.56 ;
      RECT 3.638 12.36 4.462 13.08 ;
      RECT 3.638 11.16 3.944 12.36 ;
      RECT 3.988 11.16 4.112 12.36 ;
      RECT 4.156 11.16 4.372 12.36 ;
      RECT 4.416 11.16 4.462 12.36 ;
      RECT 3.638 10.2 4.462 11.16 ;
      RECT 3.638 9 3.944 10.2 ;
      RECT 3.988 9 4.112 10.2 ;
      RECT 4.156 9 4.372 10.2 ;
      RECT 4.416 9 4.462 10.2 ;
      RECT 3.816 8.04 4.462 9 ;
      RECT 3.638 7.8 3.684 9 ;
      RECT 3.728 7.8 3.772 9 ;
      RECT 3.816 7.8 3.944 8.04 ;
      RECT 3.638 7.08 3.944 7.8 ;
      RECT 3.988 6.84 4.028 8.04 ;
      RECT 4.072 6.84 4.112 8.04 ;
      RECT 4.156 6.84 4.284 8.04 ;
      RECT 4.328 6.84 4.462 8.04 ;
      RECT 3.816 6.84 3.944 7.08 ;
      RECT 3.816 6.12 4.462 6.84 ;
      RECT 3.638 5.88 3.684 7.08 ;
      RECT 3.728 5.88 3.772 7.08 ;
      RECT 3.816 5.88 3.944 6.12 ;
      RECT 3.638 5.16 3.944 5.88 ;
      RECT 3.988 4.92 4.028 6.12 ;
      RECT 4.072 4.92 4.112 6.12 ;
      RECT 4.156 4.92 4.284 6.12 ;
      RECT 4.328 4.92 4.462 6.12 ;
      RECT 3.816 4.92 3.944 5.16 ;
      RECT 3.816 4.2 4.462 4.92 ;
      RECT 3.638 3.96 3.684 5.16 ;
      RECT 3.728 3.96 3.772 5.16 ;
      RECT 3.816 3.96 3.944 4.2 ;
      RECT 3.638 3.24 3.944 3.96 ;
      RECT 3.988 3 4.028 4.2 ;
      RECT 4.072 3 4.112 4.2 ;
      RECT 4.156 3 4.284 4.2 ;
      RECT 4.328 3 4.462 4.2 ;
      RECT 3.816 3 3.944 3.24 ;
      RECT 3.816 2.28 4.462 3 ;
      RECT 3.638 2.04 3.684 3.24 ;
      RECT 3.728 2.04 3.772 3.24 ;
      RECT 3.816 2.04 3.944 2.28 ;
      RECT 3.638 1.32 3.944 2.04 ;
      RECT 3.988 1.08 4.028 2.28 ;
      RECT 4.072 1.08 4.112 2.28 ;
      RECT 4.156 1.08 4.284 2.28 ;
      RECT 4.328 1.08 4.462 2.28 ;
      RECT 3.728 1.08 3.944 1.32 ;
      RECT 3.638 0.12 3.684 1.32 ;
      RECT 3.728 0.12 4.462 1.08 ;
      RECT 3.638 -0.12 4.462 0.12 ;
      RECT 2.738 21.96 3.562 22.2 ;
      RECT 2.828 21.48 3.562 21.96 ;
      RECT 2.738 20.76 2.784 21.96 ;
      RECT 2.828 20.76 3.384 21.48 ;
      RECT 3.428 20.52 3.562 21.48 ;
      RECT 2.738 20.28 3.384 20.76 ;
      RECT 3.428 20.28 3.472 20.52 ;
      RECT 2.738 20.04 3.472 20.28 ;
      RECT 2.828 19.56 3.472 20.04 ;
      RECT 3.516 19.32 3.562 20.52 ;
      RECT 3.428 19.32 3.472 19.56 ;
      RECT 2.738 18.84 2.784 20.04 ;
      RECT 2.828 18.84 3.384 19.56 ;
      RECT 3.428 18.6 3.562 19.32 ;
      RECT 2.738 18.36 3.384 18.84 ;
      RECT 3.428 18.36 3.472 18.6 ;
      RECT 2.738 18.12 3.472 18.36 ;
      RECT 2.828 17.64 3.472 18.12 ;
      RECT 3.516 17.4 3.562 18.6 ;
      RECT 3.428 17.4 3.472 17.64 ;
      RECT 2.738 16.92 2.784 18.12 ;
      RECT 2.828 16.92 3.384 17.64 ;
      RECT 3.428 16.68 3.562 17.4 ;
      RECT 2.738 16.44 3.384 16.92 ;
      RECT 3.428 16.44 3.472 16.68 ;
      RECT 2.738 16.2 3.472 16.44 ;
      RECT 2.828 15.72 3.472 16.2 ;
      RECT 3.516 15.48 3.562 16.68 ;
      RECT 3.428 15.48 3.472 15.72 ;
      RECT 2.738 15 2.784 16.2 ;
      RECT 2.828 15 3.384 15.72 ;
      RECT 3.428 14.76 3.562 15.48 ;
      RECT 2.738 14.52 3.384 15 ;
      RECT 3.428 14.52 3.472 14.76 ;
      RECT 2.738 14.28 3.472 14.52 ;
      RECT 3.516 13.56 3.562 14.76 ;
      RECT 2.828 13.56 3.472 14.28 ;
      RECT 2.738 13.08 2.784 14.28 ;
      RECT 2.828 13.08 3.562 13.56 ;
      RECT 2.738 12.36 3.562 13.08 ;
      RECT 2.738 11.16 2.872 12.36 ;
      RECT 2.916 11.16 3.128 12.36 ;
      RECT 3.172 11.16 3.562 12.36 ;
      RECT 2.738 10.2 3.562 11.16 ;
      RECT 2.738 9 2.872 10.2 ;
      RECT 2.916 9 3.128 10.2 ;
      RECT 3.172 9 3.562 10.2 ;
      RECT 2.738 8.52 3.384 9 ;
      RECT 3.428 7.8 3.472 9 ;
      RECT 3.516 7.8 3.562 9 ;
      RECT 2.828 7.8 3.384 8.52 ;
      RECT 2.738 7.32 2.784 8.52 ;
      RECT 2.828 7.32 3.562 7.8 ;
      RECT 2.738 7.08 3.562 7.32 ;
      RECT 2.738 6.6 3.384 7.08 ;
      RECT 3.428 5.88 3.472 7.08 ;
      RECT 3.516 5.88 3.562 7.08 ;
      RECT 2.828 5.88 3.384 6.6 ;
      RECT 2.738 5.4 2.784 6.6 ;
      RECT 2.828 5.4 3.562 5.88 ;
      RECT 2.738 5.16 3.562 5.4 ;
      RECT 2.738 4.68 3.384 5.16 ;
      RECT 3.428 3.96 3.472 5.16 ;
      RECT 3.516 3.96 3.562 5.16 ;
      RECT 2.828 3.96 3.384 4.68 ;
      RECT 2.738 3.48 2.784 4.68 ;
      RECT 2.828 3.48 3.562 3.96 ;
      RECT 2.738 3.24 3.562 3.48 ;
      RECT 2.738 2.76 3.384 3.24 ;
      RECT 3.428 2.04 3.472 3.24 ;
      RECT 3.516 2.04 3.562 3.24 ;
      RECT 2.828 2.04 3.384 2.76 ;
      RECT 2.738 1.56 2.784 2.76 ;
      RECT 2.828 1.56 3.562 2.04 ;
      RECT 2.738 1.32 3.562 1.56 ;
      RECT 2.738 0.12 3.212 1.32 ;
      RECT 3.256 0.12 3.384 1.32 ;
      RECT 3.428 0.12 3.472 1.32 ;
      RECT 3.516 0.12 3.562 1.32 ;
      RECT 2.738 -0.12 3.562 0.12 ;
      RECT 1.838 21.96 2.662 22.2 ;
      RECT 2.356 21 2.662 21.96 ;
      RECT 1.838 20.76 2.312 21.96 ;
      RECT 2.356 20.76 2.484 21 ;
      RECT 1.838 20.04 2.484 20.76 ;
      RECT 2.528 19.8 2.572 21 ;
      RECT 2.616 19.8 2.662 21 ;
      RECT 2.356 19.8 2.484 20.04 ;
      RECT 2.356 19.08 2.662 19.8 ;
      RECT 1.838 18.84 2.312 20.04 ;
      RECT 2.356 18.84 2.484 19.08 ;
      RECT 1.838 18.12 2.484 18.84 ;
      RECT 2.528 17.88 2.572 19.08 ;
      RECT 2.616 17.88 2.662 19.08 ;
      RECT 2.356 17.88 2.484 18.12 ;
      RECT 2.356 17.16 2.662 17.88 ;
      RECT 1.838 16.92 2.312 18.12 ;
      RECT 2.356 16.92 2.484 17.16 ;
      RECT 1.838 16.2 2.484 16.92 ;
      RECT 2.528 15.96 2.572 17.16 ;
      RECT 2.616 15.96 2.662 17.16 ;
      RECT 2.356 15.96 2.484 16.2 ;
      RECT 2.356 15.24 2.662 15.96 ;
      RECT 1.838 15 2.312 16.2 ;
      RECT 2.356 15 2.484 15.24 ;
      RECT 2.528 14.04 2.572 15.24 ;
      RECT 2.616 14.04 2.662 15.24 ;
      RECT 1.838 14.04 2.484 15 ;
      RECT 1.838 12.36 2.662 14.04 ;
      RECT 1.838 11.16 1.884 12.36 ;
      RECT 1.928 11.16 2.144 12.36 ;
      RECT 2.188 11.16 2.312 12.36 ;
      RECT 2.356 11.16 2.572 12.36 ;
      RECT 2.616 11.16 2.662 12.36 ;
      RECT 1.838 10.2 2.662 11.16 ;
      RECT 1.838 9 1.884 10.2 ;
      RECT 1.928 9 2.144 10.2 ;
      RECT 2.188 9 2.312 10.2 ;
      RECT 2.356 9 2.662 10.2 ;
      RECT 1.838 8.52 2.662 9 ;
      RECT 1.838 7.56 2.572 8.52 ;
      RECT 2.616 7.32 2.662 8.52 ;
      RECT 2.528 7.32 2.572 7.56 ;
      RECT 2.528 6.6 2.662 7.32 ;
      RECT 1.838 6.36 2.312 7.56 ;
      RECT 2.356 6.36 2.484 7.56 ;
      RECT 2.528 6.36 2.572 6.6 ;
      RECT 1.838 5.64 2.572 6.36 ;
      RECT 2.616 5.4 2.662 6.6 ;
      RECT 2.528 5.4 2.572 5.64 ;
      RECT 2.528 4.68 2.662 5.4 ;
      RECT 1.838 4.44 2.312 5.64 ;
      RECT 2.356 4.44 2.484 5.64 ;
      RECT 2.528 4.44 2.572 4.68 ;
      RECT 1.838 3.72 2.572 4.44 ;
      RECT 2.616 3.48 2.662 4.68 ;
      RECT 2.528 3.48 2.572 3.72 ;
      RECT 2.528 2.76 2.662 3.48 ;
      RECT 1.838 2.52 2.312 3.72 ;
      RECT 2.356 2.52 2.484 3.72 ;
      RECT 2.528 2.52 2.572 2.76 ;
      RECT 1.838 1.8 2.572 2.52 ;
      RECT 2.616 1.56 2.662 2.76 ;
      RECT 2.356 1.56 2.572 1.8 ;
      RECT 1.838 0.6 2.228 1.8 ;
      RECT 2.272 0.6 2.312 1.8 ;
      RECT 2.356 0.6 2.662 1.56 ;
      RECT 1.838 -0.12 2.662 0.6 ;
      RECT 0.938 21.48 1.762 22.2 ;
      RECT 0.938 20.52 1.584 21.48 ;
      RECT 1.628 20.28 1.672 21.48 ;
      RECT 1.716 20.28 1.762 21.48 ;
      RECT 1.456 20.28 1.584 20.52 ;
      RECT 1.456 19.56 1.762 20.28 ;
      RECT 0.938 19.32 1.328 20.52 ;
      RECT 1.372 19.32 1.412 20.52 ;
      RECT 1.456 19.32 1.584 19.56 ;
      RECT 0.938 18.6 1.584 19.32 ;
      RECT 1.628 18.36 1.672 19.56 ;
      RECT 1.716 18.36 1.762 19.56 ;
      RECT 1.456 18.36 1.584 18.6 ;
      RECT 1.456 17.64 1.762 18.36 ;
      RECT 0.938 17.4 1.328 18.6 ;
      RECT 1.372 17.4 1.412 18.6 ;
      RECT 1.456 17.4 1.584 17.64 ;
      RECT 0.938 16.68 1.584 17.4 ;
      RECT 1.628 16.44 1.672 17.64 ;
      RECT 1.716 16.44 1.762 17.64 ;
      RECT 1.456 16.44 1.584 16.68 ;
      RECT 1.456 15.72 1.762 16.44 ;
      RECT 0.938 15.48 1.328 16.68 ;
      RECT 1.372 15.48 1.412 16.68 ;
      RECT 1.456 15.48 1.584 15.72 ;
      RECT 0.938 14.76 1.584 15.48 ;
      RECT 1.628 14.52 1.672 15.72 ;
      RECT 1.716 14.52 1.762 15.72 ;
      RECT 1.456 14.52 1.584 14.76 ;
      RECT 1.456 14.28 1.762 14.52 ;
      RECT 0.938 13.56 1.328 14.76 ;
      RECT 1.372 13.56 1.412 14.76 ;
      RECT 1.456 13.56 1.672 14.28 ;
      RECT 1.716 13.08 1.762 14.28 ;
      RECT 0.938 13.08 1.672 13.56 ;
      RECT 0.938 12.36 1.762 13.08 ;
      RECT 0.938 11.16 1.072 12.36 ;
      RECT 1.116 11.16 1.584 12.36 ;
      RECT 1.628 11.16 1.762 12.36 ;
      RECT 0.938 10.2 1.762 11.16 ;
      RECT 0.938 9 1.072 10.2 ;
      RECT 1.116 9 1.584 10.2 ;
      RECT 1.628 9 1.762 10.2 ;
      RECT 1.456 8.04 1.762 9 ;
      RECT 0.938 7.8 1.328 9 ;
      RECT 1.372 7.8 1.412 9 ;
      RECT 1.456 7.8 1.584 8.04 ;
      RECT 0.938 7.08 1.584 7.8 ;
      RECT 1.628 6.84 1.672 8.04 ;
      RECT 1.716 6.84 1.762 8.04 ;
      RECT 1.456 6.84 1.584 7.08 ;
      RECT 1.456 6.12 1.762 6.84 ;
      RECT 0.938 5.88 1.328 7.08 ;
      RECT 1.372 5.88 1.412 7.08 ;
      RECT 1.456 5.88 1.584 6.12 ;
      RECT 0.938 5.16 1.584 5.88 ;
      RECT 1.628 4.92 1.672 6.12 ;
      RECT 1.716 4.92 1.762 6.12 ;
      RECT 1.456 4.92 1.584 5.16 ;
      RECT 1.456 4.2 1.762 4.92 ;
      RECT 0.938 3.96 1.328 5.16 ;
      RECT 1.372 3.96 1.412 5.16 ;
      RECT 1.456 3.96 1.584 4.2 ;
      RECT 0.938 3.24 1.584 3.96 ;
      RECT 1.628 3 1.672 4.2 ;
      RECT 1.716 3 1.762 4.2 ;
      RECT 1.456 3 1.584 3.24 ;
      RECT 1.456 2.28 1.762 3 ;
      RECT 0.938 2.04 1.328 3.24 ;
      RECT 1.372 2.04 1.412 3.24 ;
      RECT 1.456 2.04 1.584 2.28 ;
      RECT 0.938 1.32 1.584 2.04 ;
      RECT 1.628 1.08 1.672 2.28 ;
      RECT 1.716 1.08 1.762 2.28 ;
      RECT 1.372 1.08 1.584 1.32 ;
      RECT 0.938 0.12 1.244 1.32 ;
      RECT 1.288 0.12 1.328 1.32 ;
      RECT 1.372 0.12 1.762 1.08 ;
      RECT 0.938 -0.12 1.762 0.12 ;
      RECT -0.04 22.14 0.862 22.2 ;
      RECT -0.092 12.36 0.862 22.14 ;
      RECT -0.092 11.16 0.344 12.36 ;
      RECT 0.388 11.16 0.428 12.36 ;
      RECT 0.472 11.16 0.512 12.36 ;
      RECT 0.556 11.16 0.684 12.36 ;
      RECT 0.728 11.16 0.772 12.36 ;
      RECT 0.816 11.16 0.862 12.36 ;
      RECT -0.092 10.2 0.862 11.16 ;
      RECT -0.092 9 0.344 10.2 ;
      RECT 0.388 9 0.512 10.2 ;
      RECT 0.556 9 0.772 10.2 ;
      RECT 0.816 9 0.862 10.2 ;
      RECT -0.092 -0.06 0.862 9 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 44.258 0 44.92 22.08 ;
      RECT 43.358 0 43.942 22.08 ;
      RECT 42.458 0 43.042 22.08 ;
      RECT 41.558 0 42.142 22.08 ;
      RECT 40.658 0 41.242 22.08 ;
      RECT 39.758 0 40.342 22.08 ;
      RECT 38.858 0 39.442 22.08 ;
      RECT 37.958 0 38.542 22.08 ;
      RECT 37.058 0 37.642 22.08 ;
      RECT 36.158 0 36.742 22.08 ;
      RECT 35.258 0 35.842 22.08 ;
      RECT 34.358 0 34.942 22.08 ;
      RECT 33.458 0 34.042 22.08 ;
      RECT 32.558 0 33.142 22.08 ;
      RECT 31.658 0 32.242 22.08 ;
      RECT 30.758 0 31.342 22.08 ;
      RECT 29.858 0 30.442 22.08 ;
      RECT 28.958 0 29.542 22.08 ;
      RECT 28.058 0 28.642 22.08 ;
      RECT 27.158 0 27.742 22.08 ;
      RECT 26.258 0 26.842 22.08 ;
      RECT 25.358 0 25.942 22.08 ;
      RECT 24.458 0 25.042 22.08 ;
      RECT 23.558 0 24.142 22.08 ;
      RECT 22.658 0 23.242 22.08 ;
      RECT 21.758 0 22.342 22.08 ;
      RECT 20.858 0 21.442 22.08 ;
      RECT 19.958 0 20.542 22.08 ;
      RECT 19.058 0 19.642 22.08 ;
      RECT 18.158 0 18.742 22.08 ;
      RECT 17.258 0 17.842 22.08 ;
      RECT 16.358 0 16.942 22.08 ;
      RECT 15.458 0 16.042 22.08 ;
      RECT 14.558 0 15.142 22.08 ;
      RECT 13.658 0 14.242 22.08 ;
      RECT 12.758 0 13.342 22.08 ;
      RECT 11.858 0 12.442 22.08 ;
      RECT 10.958 0 11.542 22.08 ;
      RECT 10.058 0 10.642 22.08 ;
      RECT 9.158 0 9.742 22.08 ;
      RECT 8.258 0 8.842 22.08 ;
      RECT 7.358 0 7.942 22.08 ;
      RECT 6.458 12.48 7.042 22.08 ;
      RECT 6.636 11.04 7.042 12.48 ;
      RECT 6.458 0 7.042 11.04 ;
      RECT 5.558 21.12 6.142 22.08 ;
      RECT 5.736 19.68 6.142 21.12 ;
      RECT 5.558 19.2 6.142 19.68 ;
      RECT 5.736 17.76 6.142 19.2 ;
      RECT 5.558 17.28 6.142 17.76 ;
      RECT 5.736 15.84 6.142 17.28 ;
      RECT 5.558 15.36 6.142 15.84 ;
      RECT 5.736 13.92 6.142 15.36 ;
      RECT 5.558 12.48 6.142 13.92 ;
      RECT 5.176 21.12 5.242 22.08 ;
      RECT 3.758 21.6 4.342 22.08 ;
      RECT 3.758 20.64 3.824 21.6 ;
      RECT 4.276 20.64 4.342 21.6 ;
      RECT 2.948 21.6 3.442 22.08 ;
      RECT 2.948 20.64 3.264 21.6 ;
      RECT 2.858 20.16 3.264 20.64 ;
      RECT 2.948 19.68 3.352 20.16 ;
      RECT 2.948 18.72 3.264 19.68 ;
      RECT 2.858 18.24 3.264 18.72 ;
      RECT 2.948 17.76 3.352 18.24 ;
      RECT 2.948 16.8 3.264 17.76 ;
      RECT 2.858 16.32 3.264 16.8 ;
      RECT 2.948 15.84 3.352 16.32 ;
      RECT 2.948 14.88 3.264 15.84 ;
      RECT 2.858 14.4 3.264 14.88 ;
      RECT 2.948 13.44 3.352 14.4 ;
      RECT 2.948 12.96 3.442 13.44 ;
      RECT 2.858 12.48 3.442 12.96 ;
      RECT 3.292 11.04 3.442 12.48 ;
      RECT 2.858 10.32 3.442 11.04 ;
      RECT 3.292 9.12 3.442 10.32 ;
      RECT 2.476 21.12 2.542 22.08 ;
      RECT 1.958 20.64 2.192 22.08 ;
      RECT 1.958 20.16 2.364 20.64 ;
      RECT 1.958 18.72 2.192 20.16 ;
      RECT 1.958 18.24 2.364 18.72 ;
      RECT 1.958 16.8 2.192 18.24 ;
      RECT 1.958 16.32 2.364 16.8 ;
      RECT 1.958 14.88 2.192 16.32 ;
      RECT 1.958 13.92 2.364 14.88 ;
      RECT 1.958 12.48 2.542 13.92 ;
      RECT 1.058 21.6 1.642 22.08 ;
      RECT 1.058 20.64 1.464 21.6 ;
      RECT 1.058 19.2 1.208 20.64 ;
      RECT 1.058 18.72 1.464 19.2 ;
      RECT 1.058 17.28 1.208 18.72 ;
      RECT 1.058 16.8 1.464 17.28 ;
      RECT 1.058 15.36 1.208 16.8 ;
      RECT 1.058 14.88 1.464 15.36 ;
      RECT 1.058 13.44 1.208 14.88 ;
      RECT 1.058 12.96 1.552 13.44 ;
      RECT 1.058 12.48 1.642 12.96 ;
      RECT 1.236 11.04 1.464 12.48 ;
      RECT 1.058 10.32 1.642 11.04 ;
      RECT 1.236 9.12 1.464 10.32 ;
      RECT 0.08 12.48 0.742 22.08 ;
      RECT 0.08 11.04 0.224 12.48 ;
      RECT 0.08 10.32 0.742 11.04 ;
      RECT 0.08 8.88 0.224 10.32 ;
      RECT 0.08 0 0.742 8.88 ;
      RECT 4.658 20.16 5.064 20.64 ;
      RECT 3.936 19.68 4.164 20.16 ;
      RECT 1.576 19.68 1.642 20.16 ;
      RECT 5.176 19.2 5.242 19.68 ;
      RECT 2.476 19.2 2.542 19.68 ;
      RECT 4.276 18.72 4.342 19.2 ;
      RECT 3.758 18.72 3.824 19.2 ;
      RECT 4.658 18.24 5.064 18.72 ;
      RECT 3.936 17.76 4.164 18.24 ;
      RECT 1.576 17.76 1.642 18.24 ;
      RECT 5.176 17.28 5.242 17.76 ;
      RECT 2.476 17.28 2.542 17.76 ;
      RECT 4.276 16.8 4.342 17.28 ;
      RECT 3.758 16.8 3.824 17.28 ;
      RECT 4.658 16.32 5.064 16.8 ;
      RECT 3.936 15.84 4.164 16.32 ;
      RECT 1.576 15.84 1.642 16.32 ;
      RECT 5.176 15.36 5.242 15.84 ;
      RECT 2.476 15.36 2.542 15.84 ;
      RECT 4.276 14.4 4.342 15.36 ;
      RECT 3.758 14.88 3.824 15.36 ;
      RECT 4.658 14.4 4.892 14.88 ;
      RECT 5.176 13.44 5.242 13.92 ;
      RECT 5.008 12.96 5.242 13.44 ;
      RECT 4.658 12.48 5.242 12.96 ;
      RECT 3.758 12.96 3.908 13.44 ;
      RECT 3.758 12.48 4.342 12.96 ;
      RECT 3.758 11.04 3.824 12.48 ;
      RECT 3.758 10.32 4.342 11.04 ;
      RECT 3.758 9.12 3.824 10.32 ;
      RECT 5.558 8.64 6.142 11.04 ;
      RECT 5.736 7.2 6.142 8.64 ;
      RECT 5.558 6.72 6.142 7.2 ;
      RECT 5.736 5.28 6.142 6.72 ;
      RECT 5.558 4.8 6.142 5.28 ;
      RECT 5.736 3.36 6.142 4.8 ;
      RECT 5.558 2.88 6.142 3.36 ;
      RECT 5.736 1.44 6.142 2.88 ;
      RECT 5.558 0 6.142 1.44 ;
      RECT 4.658 8.64 5.242 11.04 ;
      RECT 4.658 7.68 5.064 8.64 ;
      RECT 1.958 10.32 2.542 11.04 ;
      RECT 2.476 8.88 2.542 10.32 ;
      RECT 1.958 8.64 2.542 8.88 ;
      RECT 1.958 7.68 2.452 8.64 ;
      RECT 1.958 6.24 2.192 7.68 ;
      RECT 1.958 5.76 2.452 6.24 ;
      RECT 1.958 4.32 2.192 5.76 ;
      RECT 1.958 3.84 2.452 4.32 ;
      RECT 1.958 2.4 2.192 3.84 ;
      RECT 1.958 1.92 2.452 2.4 ;
      RECT 1.958 0.48 2.108 1.92 ;
      RECT 2.476 0.48 2.542 1.44 ;
      RECT 1.958 0 2.542 0.48 ;
      RECT 3.936 8.16 4.342 8.88 ;
      RECT 2.858 8.64 3.264 8.88 ;
      RECT 2.948 7.68 3.264 8.64 ;
      RECT 2.948 7.2 3.442 7.68 ;
      RECT 2.858 6.72 3.264 7.2 ;
      RECT 2.948 5.76 3.264 6.72 ;
      RECT 2.948 5.28 3.442 5.76 ;
      RECT 2.858 4.8 3.264 5.28 ;
      RECT 2.948 3.84 3.264 4.8 ;
      RECT 2.948 3.36 3.442 3.84 ;
      RECT 2.858 2.88 3.264 3.36 ;
      RECT 2.948 1.92 3.264 2.88 ;
      RECT 2.948 1.44 3.442 1.92 ;
      RECT 2.858 0 3.092 1.44 ;
      RECT 1.576 8.16 1.642 8.88 ;
      RECT 1.058 7.68 1.208 8.88 ;
      RECT 1.058 7.2 1.464 7.68 ;
      RECT 1.058 5.76 1.208 7.2 ;
      RECT 1.058 5.28 1.464 5.76 ;
      RECT 1.058 3.84 1.208 5.28 ;
      RECT 1.058 3.36 1.464 3.84 ;
      RECT 1.058 1.92 1.208 3.36 ;
      RECT 1.058 1.44 1.464 1.92 ;
      RECT 1.058 0 1.124 1.44 ;
      RECT 3.758 7.2 3.824 7.68 ;
      RECT 5.176 6.72 5.242 7.2 ;
      RECT 3.936 6.24 4.342 6.72 ;
      RECT 1.576 6.24 1.642 6.72 ;
      RECT 4.658 5.76 5.064 6.24 ;
      RECT 3.758 5.28 3.824 5.76 ;
      RECT 5.176 4.8 5.242 5.28 ;
      RECT 3.936 4.32 4.342 4.8 ;
      RECT 1.576 4.32 1.642 4.8 ;
      RECT 4.658 3.84 5.064 4.32 ;
      RECT 3.758 3.36 3.824 3.84 ;
      RECT 5.176 2.88 5.242 3.36 ;
      RECT 3.936 2.4 4.342 2.88 ;
      RECT 1.576 2.4 1.642 2.88 ;
      RECT 4.658 1.92 5.064 2.4 ;
      RECT 3.758 1.44 3.824 1.92 ;
      RECT 5.092 0.48 5.242 1.44 ;
      RECT 4.658 0 5.242 0.48 ;
      RECT 3.848 0 4.342 0.96 ;
      RECT 1.492 0 1.642 0.96 ;
    LAYER m0 ;
      RECT 0 0.002 45 22.078 ;
    LAYER m1 ;
      RECT 0 0 45 22.08 ;
    LAYER m2 ;
      RECT 0 0.015 45 22.065 ;
    LAYER m3 ;
      RECT 0.015 0 44.985 22.08 ;
    LAYER m4 ;
      RECT 0 0.02 45 22.06 ;
    LAYER m5 ;
      RECT 0.012 0 44.988 22.08 ;
    LAYER m6 ;
      RECT 0 0.012 45 22.068 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf066b128e2r1w0cbbehsaa4acw

END LIBRARY
