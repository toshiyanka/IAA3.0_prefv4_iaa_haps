module ctech_lib_power_switch (a, o);
     input a;
     output o;
   d04pws00ld0b0 ctech_lib_dcszo (.a(a),.o(o));
endmodule
