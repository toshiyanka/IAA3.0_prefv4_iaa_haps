`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

(* inserted_by="VISA IT" *) .visaRt_probe_from_i_hqm_master_visa_block(visaPrbsTo_i_hqm_visa_mux_top_vcfn),


`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
