//              TAP name,       Opcode,   DR_length
//
Create_Reg_Model (IPLEVEL_STAP,  8'hFF,      'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (IPLEVEL_STAP,  8'hC,       'd32     );   // opcode is SLVIDCODE [0xC]
//
