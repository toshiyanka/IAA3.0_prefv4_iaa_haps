package PowerGatingParamsPkg;	

	parameter int MAX_SIP = 128;
	parameter int MAX_FAB = 128;
	parameter int MAX_FET = 128;
endpackage: PowerGatingParamsPkg
