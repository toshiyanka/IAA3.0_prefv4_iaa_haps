//=====================================================================================================================
//
// iommu_cust_params.vh
//
// Contacts            : Chintan Panirwala & Camron Rust
// Original Author(s)  : Chintan Panirwala & Camron Rust
// Original Date       : 3/2014
//
// -- Intel Proprietary
// -- Copyright (C) 2016 Intel Corporation
// -- All Rights Reserved
//
// This file contains all customer defined parameters.
//
//=====================================================================================================================

//=====================================================================================================================
// All additional parameters added to this file need to also be added to the bind statement at the bottom of iommu.sv.
// The FPV reference model needs to have these parameters passed in for proper functionality at integration.
//=====================================================================================================================



//=====================================================================================================================
// All additional parameters added to this file need to also be added to the bind statement at the bottom of iommu.sv.
// The FPV reference model needs to have these parameters passed in for proper functionality at integration.
//=====================================================================================================================

