module dump_hier_test();
endmodule
