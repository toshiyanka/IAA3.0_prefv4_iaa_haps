/*
================================================================================
  Copyright (c) 2011 Intel Corporation, all rights reserved.

  THIS PROGRAM IS AN UNPUBLISHED WORK FULLY PROTECTED BY COPYRIGHT LAWS AND IS 
  CONSIDERED A TRADE SECRET BELONGING TO THE INTEL CORPORATION.
================================================================================

  Author          : 
  Email           : 
  Phone           : 
  Date            : 

================================================================================
  Description     : One line description of this class
  
Write your wordy description here.
================================================================================
*/

//Minimum Subset an Agent should contain
`include "PGCBAgentTypes.svh"
`include "PGCBAgentDriver.svh"
//col change
`include "PGCBAgentDriver_Col.svh"
//END col change
`include "PGCBAgentSeqItem.svh"
`include "PGCBAgentSequencer.svh"
`include "PGCBAgentFabricResponder.svh"
`include "PGCBAgentSIPResponder.svh"
`include "PGCBAgentSeqLib.svh"
`include "PGCBAgent.svh"
`include "PGCBAgentResponseSeqItem.svh"
`include "PGCBAgentSIPFSM.svh"
`include "PGCBAgentFabricFSM.svh"
//col change
`include "PGCBAgentSIPFSM_Col.svh"
`include "PGCBAgentFabricFSM_Col.svh"
//END col change


