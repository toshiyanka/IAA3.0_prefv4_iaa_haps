# Text_Tag % Vendor Intel % Product c73p4rfshdxrom % Techno P1273.1 % Tag_Spec 1.0 % ECCN US_3E002 % Signature debc08ffedd3027797a0273bd28a69585f4c0a48 % Version r1.0.0_m1.18 % _View_Id lef % Date_Time 20160216_100949 
################################################################################
# Intel Confidential                                                           #
################################################################################
# Copyright 2014 Intel Corporation.                                            #
# The information contained herein is the proprietary and confidential         #
# information of Intel or its licensors, and is supplied subject to, and       #
# may be used only in accordance with, previously executed agreements          #
# with Intel ,                                                                 #
# EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING:                                #
# (1) ALL MATERIALS FURNISHED BY INTEL HEREUNDER ARE PROVIDED "AS IS"          #
#      WITHOUT WARRANTY OF ANY KIND;                                           #
# (2) INTEL SPECIFICALLY DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS    #
#      FOR A PARTICULAR PURPOSE OR MERCHANTABILITY; AND                        #
# (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF SUBSTITUTES,    #
#      LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR                           #
#      FOR ANY OTHER SPECIAL, CONSEQUENTIAL OR INCIDENTAL DAMAGES,             #
#      HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY, CONTRACT,               #
#      TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                        #
################################################################################
################################################################################
#                                                                              #
# Vendor: Intel                                                                #
# Product: c73p4rfshdxrom                                                      #
# Version: r1.0.0_m1.18                                                        #
# Technology: p1273.1                                                          #
# Celltype: IP                                                                 #
# IP_Owner: Intel DTS CMO                                                      #
# Date_Time: YYYYMMDD_HHMMSS                                                   #
#                                                                              #
################################################################################
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

SITE c73p1rfshdxrom2048x32hb4img108
  SIZE 75.432 by 49.476 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END c73p1rfshdxrom2048x32hb4img108


MACRO c73p1rfshdxrom2048x32hb4img108
     FOREIGN c73p1rfshdxrom2048x32hb4img108 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 75.432 by 49.476 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE c73p1rfshdxrom2048x32hb4img108 ;
     PIN iar[10]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 21.068 0.308 21.1 ;
          END
     END iar[10]
     PIN iar[0]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 21.754 0.308 21.786 ;
          END
     END iar[0]
     PIN iar[1]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 22.496 0.308 22.528 ;
          END
     END iar[1]
     PIN iar[2]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 23.126 0.308 23.158 ;
          END
     END iar[2]
     PIN iar[4]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 23.812 0.308 23.844 ;
          END
     END iar[4]
     PIN iar[3]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 24.442 0.308 24.474 ;
          END
     END iar[3]
     PIN iar[7]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 25.744 0.308 25.776 ;
          END
     END iar[7]
     PIN iar[6]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 26.43 0.308 26.462 ;
          END
     END iar[6]
     PIN iar[5]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 27.004 0.308 27.036 ;
          END
     END iar[5]
     PIN iar[9]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 27.802 0.308 27.834 ;
          END
     END iar[9]
     PIN iar[8]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 28.432 0.308 28.464 ;
          END
     END iar[8]
     PIN iren
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 25.184 0.308 25.216 ;
          END
     END iren
     PIN ickr
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 24.946 0.308 24.978 ;
          END
     END ickr
     PIN ipwreninb
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 48.718 0.308 48.75 ;
          END
     END ipwreninb
     PIN opwrenoutb
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 0.95 0.308 0.982 ;
          END
     END opwrenoutb
     PIN odout[0]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 1.062 0.308 1.094 ;
          END
     END odout[0]
     PIN odout[1]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 2.434 0.308 2.466 ;
          END
     END odout[1]
     PIN odout[2]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 3.694 0.308 3.726 ;
          END
     END odout[2]
     PIN odout[3]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 4.94 0.308 4.972 ;
          END
     END odout[3]
     PIN odout[4]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 6.088 0.308 6.12 ;
          END
     END odout[4]
     PIN odout[5]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 7.334 0.308 7.366 ;
          END
     END odout[5]
     PIN odout[6]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 8.594 0.308 8.626 ;
          END
     END odout[6]
     PIN odout[7]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 9.84 0.308 9.872 ;
          END
     END odout[7]
     PIN odout[8]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 11.212 0.308 11.244 ;
          END
     END odout[8]
     PIN odout[9]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 12.234 0.308 12.266 ;
          END
     END odout[9]
     PIN odout[10]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 13.494 0.308 13.526 ;
          END
     END odout[10]
     PIN odout[11]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 14.866 0.308 14.898 ;
          END
     END odout[11]
     PIN odout[12]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 16.224 0.308 16.256 ;
          END
     END odout[12]
     PIN odout[13]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 17.372 0.308 17.404 ;
          END
     END odout[13]
     PIN odout[14]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 18.618 0.308 18.65 ;
          END
     END odout[14]
     PIN odout[15]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 19.99 0.308 20.022 ;
          END
     END odout[15]
     PIN odout[16]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 29.342 0.308 29.374 ;
          END
     END odout[16]
     PIN odout[17]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 30.588 0.308 30.62 ;
          END
     END odout[17]
     PIN odout[18]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 31.624 0.308 31.656 ;
          END
     END odout[18]
     PIN odout[19]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 32.982 0.308 33.014 ;
          END
     END odout[19]
     PIN odout[20]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 34.354 0.308 34.386 ;
          END
     END odout[20]
     PIN odout[21]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 35.614 0.308 35.646 ;
          END
     END odout[21]
     PIN odout[22]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 36.748 0.308 36.78 ;
          END
     END odout[22]
     PIN odout[23]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 38.008 0.308 38.04 ;
          END
     END odout[23]
     PIN odout[24]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 39.254 0.308 39.286 ;
          END
     END odout[24]
     PIN odout[25]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 40.514 0.308 40.546 ;
          END
     END odout[25]
     PIN odout[26]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 41.76 0.308 41.792 ;
          END
     END odout[26]
     PIN odout[27]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 43.02 0.308 43.052 ;
          END
     END odout[27]
     PIN odout[28]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 44.154 0.308 44.186 ;
          END
     END odout[28]
     PIN odout[29]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 45.526 0.308 45.558 ;
          END
     END odout[29]
     PIN odout[30]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 46.898 0.308 46.93 ;
          END
     END odout[30]
     PIN odout[31]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 48.144 0.308 48.176 ;
          END
     END odout[31]
     PIN vccd_1p0
     SHAPE ABUTMENT ;
     USE   POWER ;
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0.42 0.654 74.894 0.7 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.852 14.274 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.064 2.832 1.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.34 13.678 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.474 13.354 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.722 14 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.914 74.894 1.96 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.16 13.678 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.294 13.354 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.542 14 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.734 74.894 10.78 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.932 14.274 10.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.144 2.832 11.228 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.42 13.678 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.554 13.354 11.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.802 14 11.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.994 74.894 12.04 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.192 14.274 12.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.404 2.832 12.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.68 13.678 12.726 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.814 13.354 12.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.062 14 13.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.254 74.894 13.3 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.452 14.274 13.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.664 2.832 13.748 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.94 13.678 13.986 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.074 13.354 14.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.322 14 14.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.514 74.894 14.56 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.712 14.274 14.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.924 2.832 15.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.2 13.678 15.246 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.334 13.354 15.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.582 14 15.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.774 74.894 15.82 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.972 14.274 16.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.184 2.832 16.268 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.46 13.678 16.506 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.594 13.354 16.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.842 14 16.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.034 74.894 17.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.232 14.274 17.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.444 2.832 17.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.72 13.678 17.766 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.854 13.354 17.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.102 14 18.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.294 74.894 18.34 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.492 14.274 18.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.704 2.832 18.788 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.98 13.678 19.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.114 13.354 19.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.362 14 19.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.554 74.894 19.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.752 14.274 19.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.964 2.832 20.048 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.112 14.274 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.324 2.832 2.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.6 13.678 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.734 13.354 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.982 14 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.24 13.678 20.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.374 13.354 20.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.622 14 20.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.744 74.894 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.964 74.894 21.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.168 74.894 21.214 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.372 74.894 21.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.57 6.19 21.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.64 74.894 21.68 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.768 74.894 21.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.402 74.894 22.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.67 74.894 22.724 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.086 74.894 23.126 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.83 74.894 23.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.326 74.894 24.366 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.194 74.894 25.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.566 74.894 25.606 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.062 74.894 26.102 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.558 74.894 26.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.93 74.894 26.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.178 74.894 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.542 74.894 27.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.686 74.894 27.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.826 74.894 27.872 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.976 74.894 28.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.116 74.894 28.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.276 74.894 28.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.41 74.894 28.464 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.558 74.894 28.604 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.692 74.894 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.878 74.894 28.924 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.076 14.274 29.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.288 2.832 29.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.564 13.678 29.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.698 13.354 29.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.946 14 29.992 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.174 74.894 3.22 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.372 14.274 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.584 2.832 3.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.86 13.678 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.994 13.354 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.138 74.894 30.184 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.336 14.274 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.548 2.832 30.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.824 13.678 30.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.958 13.354 30.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.206 14 31.252 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.398 74.894 31.444 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.596 14.274 31.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.808 2.832 31.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.084 13.678 32.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.218 13.354 32.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.466 14 32.512 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.658 74.894 32.704 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.856 14.274 32.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.068 2.832 33.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.344 13.678 33.39 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.478 13.354 33.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.726 14 33.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.918 74.894 33.964 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.116 14.274 34.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.328 2.832 34.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.604 13.678 34.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.738 13.354 34.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.986 14 35.032 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.178 74.894 35.224 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.376 14.274 35.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.588 2.832 35.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.864 13.678 35.91 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.998 13.354 36.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.246 14 36.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.438 74.894 36.484 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.636 14.274 36.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.848 2.832 36.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.124 13.678 37.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.258 13.354 37.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.506 14 37.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.698 74.894 37.744 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.896 14.274 37.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.108 2.832 38.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.384 13.678 38.43 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.518 13.354 38.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.766 14 38.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.958 74.894 39.004 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.156 14.274 39.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.368 2.832 39.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.644 13.678 39.69 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.778 13.354 39.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.242 14 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.434 74.894 4.48 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.632 14.274 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.844 2.832 4.928 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.026 14 40.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.218 74.894 40.264 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.416 14.274 40.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.628 2.832 40.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.904 13.678 40.95 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.038 13.354 41.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.286 14 41.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.478 74.894 41.524 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.676 14.274 41.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.888 2.832 41.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.164 13.678 42.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.298 13.354 42.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.546 14 42.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.738 74.894 42.784 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.936 14.274 42.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.148 2.832 43.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.424 13.678 43.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.558 13.354 43.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.806 14 43.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.998 74.894 44.044 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.196 14.274 44.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.408 2.832 44.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.684 13.678 44.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.818 13.354 44.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.066 14 45.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.258 74.894 45.304 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.456 14.274 45.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.668 2.832 45.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.944 13.678 45.99 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.078 13.354 46.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.326 14 46.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.518 74.894 46.564 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.716 14.274 46.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.928 2.832 47.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.204 13.678 47.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.338 13.354 47.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.586 14 47.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.778 74.894 47.824 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.976 14.274 48.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.188 2.832 48.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.464 13.678 48.51 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.598 13.354 48.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.846 14 48.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.12 13.678 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.254 13.354 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.502 14 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.694 74.894 5.74 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.892 14.274 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.104 2.832 6.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.38 13.678 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.514 13.354 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.762 14 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.954 74.894 7 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.152 14.274 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.364 2.832 7.448 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.64 13.678 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.774 13.354 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.022 14 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.214 74.894 8.26 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.412 14.274 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.624 2.832 8.708 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.9 13.678 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.034 13.354 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.282 14 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.474 74.894 9.52 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.672 14.274 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.884 2.832 9.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 1.722 31.052 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 10.542 31.052 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 11.802 31.052 11.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 13.062 31.052 13.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 14.322 31.052 14.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 15.582 31.052 15.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 16.842 31.052 16.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 18.102 31.052 18.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 19.362 31.052 19.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 2.982 31.052 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 20.622 31.052 20.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 29.946 31.052 29.992 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 31.206 31.052 31.252 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 32.466 31.052 32.512 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 33.726 31.052 33.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 34.986 31.052 35.032 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 36.246 31.052 36.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 37.506 31.052 37.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 38.766 31.052 38.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 4.242 31.052 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 40.026 31.052 40.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 41.286 31.052 41.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 42.546 31.052 42.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 43.806 31.052 43.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 45.066 31.052 45.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 46.326 31.052 46.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 47.586 31.052 47.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 48.846 31.052 48.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 5.502 31.052 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 6.762 31.052 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 8.022 31.052 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 9.282 31.052 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 0.852 31.326 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 10.932 31.326 10.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 12.192 31.326 12.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 13.452 31.326 13.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 14.712 31.326 14.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 15.972 31.326 16.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 17.232 31.326 17.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 18.492 31.326 18.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 19.752 31.326 19.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 2.112 31.326 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 29.076 31.326 29.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 3.372 31.326 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 30.336 31.326 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 31.596 31.326 31.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 32.856 31.326 32.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 34.116 31.326 34.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 35.376 31.326 35.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 36.636 31.326 36.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 37.896 31.326 37.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 39.156 31.326 39.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 4.632 31.326 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 40.416 31.326 40.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 41.676 31.326 41.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 42.936 31.326 42.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 44.196 31.326 44.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 45.456 31.326 45.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 46.716 31.326 46.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 47.976 31.326 48.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 5.892 31.326 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 7.152 31.326 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 8.412 31.326 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 9.672 31.326 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 1.474 30.406 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 10.294 30.406 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 11.554 30.406 11.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 12.814 30.406 12.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 14.074 30.406 14.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 15.334 30.406 15.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 16.594 30.406 16.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 17.854 30.406 17.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 19.114 30.406 19.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 2.734 30.406 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 20.374 30.406 20.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 29.698 30.406 29.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 3.994 30.406 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 30.958 30.406 30.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 32.218 30.406 32.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 33.478 30.406 33.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 34.738 30.406 34.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 35.998 30.406 36.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 37.258 30.406 37.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 38.518 30.406 38.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 39.778 30.406 39.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 41.038 30.406 41.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 42.298 30.406 42.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 43.558 30.406 43.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 44.818 30.406 44.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 46.078 30.406 46.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 47.338 30.406 47.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 48.598 30.406 48.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 5.254 30.406 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 6.514 30.406 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 7.774 30.406 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 9.034 30.406 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 1.34 30.73 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 10.16 30.73 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 11.42 30.73 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 12.68 30.73 12.726 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 13.94 30.73 13.986 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 15.2 30.73 15.246 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 16.46 30.73 16.506 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 17.72 30.73 17.766 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 18.98 30.73 19.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 2.6 30.73 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 20.24 30.73 20.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 29.564 30.73 29.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 3.86 30.73 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 30.824 30.73 30.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 32.084 30.73 32.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 33.344 30.73 33.39 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 34.604 30.73 34.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 35.864 30.73 35.91 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 37.124 30.73 37.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 38.384 30.73 38.43 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 39.644 30.73 39.69 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 40.904 30.73 40.95 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 42.164 30.73 42.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 43.424 30.73 43.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 44.684 30.73 44.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 45.944 30.73 45.99 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 47.204 30.73 47.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 48.464 30.73 48.51 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 5.12 30.73 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 6.38 30.73 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 7.64 30.73 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 8.9 30.73 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 1.722 48.104 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 10.542 48.104 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 11.802 48.104 11.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 13.062 48.104 13.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 14.322 48.104 14.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 15.582 48.104 15.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 16.842 48.104 16.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 18.102 48.104 18.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 19.362 48.104 19.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 2.982 48.104 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 20.622 48.104 20.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 29.946 48.104 29.992 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 31.206 48.104 31.252 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 32.466 48.104 32.512 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 33.726 48.104 33.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 34.986 48.104 35.032 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 36.246 48.104 36.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 37.506 48.104 37.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 38.766 48.104 38.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 4.242 48.104 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 40.026 48.104 40.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 41.286 48.104 41.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 42.546 48.104 42.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 43.806 48.104 43.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 45.066 48.104 45.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 46.326 48.104 46.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 47.586 48.104 47.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 48.846 48.104 48.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 5.502 48.104 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 6.762 48.104 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 8.022 48.104 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 9.282 48.104 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 0.852 48.378 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 10.932 48.378 10.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 12.192 48.378 12.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 13.452 48.378 13.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 14.712 48.378 14.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 15.972 48.378 16.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 17.232 48.378 17.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 18.492 48.378 18.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 19.752 48.378 19.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 2.112 48.378 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 29.076 48.378 29.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 3.372 48.378 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 30.336 48.378 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 31.596 48.378 31.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 32.856 48.378 32.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 34.116 48.378 34.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 35.376 48.378 35.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 36.636 48.378 36.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 37.896 48.378 37.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 39.156 48.378 39.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 4.632 48.378 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 40.416 48.378 40.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 41.676 48.378 41.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 42.936 48.378 42.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 44.196 48.378 44.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 45.456 48.378 45.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 46.716 48.378 46.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 47.976 48.378 48.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 5.892 48.378 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 7.152 48.378 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 8.412 48.378 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 9.672 48.378 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 1.474 47.458 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 10.294 47.458 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 11.554 47.458 11.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 12.814 47.458 12.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 14.074 47.458 14.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 15.334 47.458 15.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 16.594 47.458 16.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 17.854 47.458 17.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 19.114 47.458 19.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 2.734 47.458 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 20.374 47.458 20.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 29.698 47.458 29.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 3.994 47.458 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 30.958 47.458 30.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 32.218 47.458 32.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 33.478 47.458 33.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 34.738 47.458 34.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 35.998 47.458 36.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 37.258 47.458 37.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 38.518 47.458 38.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 39.778 47.458 39.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 41.038 47.458 41.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 42.298 47.458 42.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 43.558 47.458 43.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 44.818 47.458 44.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 46.078 47.458 46.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 47.338 47.458 47.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 48.598 47.458 48.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 5.254 47.458 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 6.514 47.458 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 7.774 47.458 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 9.034 47.458 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 1.34 47.782 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 10.16 47.782 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 11.42 47.782 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 12.68 47.782 12.726 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 13.94 47.782 13.986 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 15.2 47.782 15.246 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 16.46 47.782 16.506 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 17.72 47.782 17.766 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 18.98 47.782 19.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 2.6 47.782 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 20.24 47.782 20.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 29.564 47.782 29.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 3.86 47.782 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 30.824 47.782 30.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 32.084 47.782 32.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 33.344 47.782 33.39 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 34.604 47.782 34.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 35.864 47.782 35.91 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 37.124 47.782 37.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 38.384 47.782 38.43 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 39.644 47.782 39.69 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 40.904 47.782 40.95 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 42.164 47.782 42.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 43.424 47.782 43.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 44.684 47.782 44.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 45.944 47.782 45.99 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 47.204 47.782 47.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 48.464 47.782 48.51 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 5.12 47.782 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 6.38 47.782 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 7.64 47.782 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 8.9 47.782 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 1.722 65.156 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 10.542 65.156 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 11.802 65.156 11.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 13.062 65.156 13.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 14.322 65.156 14.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 15.582 65.156 15.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 16.842 65.156 16.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 18.102 65.156 18.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 19.362 65.156 19.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 2.982 65.156 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 20.622 65.156 20.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 29.946 65.156 29.992 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 31.206 65.156 31.252 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 32.466 65.156 32.512 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 33.726 65.156 33.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 34.986 65.156 35.032 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 36.246 65.156 36.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 37.506 65.156 37.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 38.766 65.156 38.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 4.242 65.156 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 40.026 65.156 40.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 41.286 65.156 41.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 42.546 65.156 42.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 43.806 65.156 43.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 45.066 65.156 45.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 46.326 65.156 46.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 47.586 65.156 47.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 48.846 65.156 48.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 5.502 65.156 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 6.762 65.156 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 8.022 65.156 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 9.282 65.156 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 0.852 65.43 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 10.932 65.43 10.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 12.192 65.43 12.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 13.452 65.43 13.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 14.712 65.43 14.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 15.972 65.43 16.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 17.232 65.43 17.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 18.492 65.43 18.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 19.752 65.43 19.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 2.112 65.43 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 29.076 65.43 29.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 3.372 65.43 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 30.336 65.43 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 31.596 65.43 31.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 32.856 65.43 32.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 34.116 65.43 34.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 35.376 65.43 35.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 36.636 65.43 36.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 37.896 65.43 37.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 39.156 65.43 39.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 4.632 65.43 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 40.416 65.43 40.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 41.676 65.43 41.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 42.936 65.43 42.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 44.196 65.43 44.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 45.456 65.43 45.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 46.716 65.43 46.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 47.976 65.43 48.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 5.892 65.43 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 7.152 65.43 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 8.412 65.43 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 9.672 65.43 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 1.474 64.51 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 10.294 64.51 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 11.554 64.51 11.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 12.814 64.51 12.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 14.074 64.51 14.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 15.334 64.51 15.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 16.594 64.51 16.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 17.854 64.51 17.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 19.114 64.51 19.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 2.734 64.51 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 20.374 64.51 20.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 29.698 64.51 29.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 3.994 64.51 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 30.958 64.51 30.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 32.218 64.51 32.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 33.478 64.51 33.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 34.738 64.51 34.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 35.998 64.51 36.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 37.258 64.51 37.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 38.518 64.51 38.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 39.778 64.51 39.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 41.038 64.51 41.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 42.298 64.51 42.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 43.558 64.51 43.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 44.818 64.51 44.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 46.078 64.51 46.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 47.338 64.51 47.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 48.598 64.51 48.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 5.254 64.51 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 6.514 64.51 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 7.774 64.51 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 9.034 64.51 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 1.34 64.834 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 10.16 64.834 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 11.42 64.834 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 12.68 64.834 12.726 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 13.94 64.834 13.986 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 15.2 64.834 15.246 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 16.46 64.834 16.506 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 17.72 64.834 17.766 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 18.98 64.834 19.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 2.6 64.834 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 20.24 64.834 20.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 29.564 64.834 29.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 3.86 64.834 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 30.824 64.834 30.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 32.084 64.834 32.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 33.344 64.834 33.39 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 34.604 64.834 34.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 35.864 64.834 35.91 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 37.124 64.834 37.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 38.384 64.834 38.43 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 39.644 64.834 39.69 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 40.904 64.834 40.95 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 42.164 64.834 42.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 43.424 64.834 43.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 44.684 64.834 44.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 45.944 64.834 45.99 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 47.204 64.834 47.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 48.464 64.834 48.51 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 5.12 64.834 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 6.38 64.834 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 7.64 64.834 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 8.9 64.834 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 1.722 74.894 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 10.542 74.894 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 11.802 74.894 11.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 13.062 74.894 13.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 14.322 74.894 14.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 15.582 74.894 15.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 16.842 74.894 16.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 18.102 74.894 18.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 19.362 74.894 19.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 2.982 74.894 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 20.622 74.894 20.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 29.946 74.894 29.992 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 31.206 74.894 31.252 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 32.466 74.894 32.512 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 33.726 74.894 33.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 34.986 74.894 35.032 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 36.246 74.894 36.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 37.506 74.894 37.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 38.766 74.894 38.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 4.242 74.894 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 40.026 74.894 40.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 41.286 74.894 41.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 42.546 74.894 42.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 43.806 74.894 43.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 45.066 74.894 45.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 46.326 74.894 46.372 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 47.586 74.894 47.632 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 48.846 74.894 48.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 5.502 74.894 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 6.762 74.894 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 8.022 74.894 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 9.282 74.894 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 0.852 74.894 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 10.932 74.894 10.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 12.192 74.894 12.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 13.452 74.894 13.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 14.712 74.894 14.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 15.972 74.894 16.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 17.232 74.894 17.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 18.492 74.894 18.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 19.752 74.894 19.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 2.112 74.894 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 29.076 74.894 29.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 3.372 74.894 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 30.336 74.894 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 31.596 74.894 31.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 32.856 74.894 32.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 34.116 74.894 34.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 35.376 74.894 35.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 36.636 74.894 36.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 37.896 74.894 37.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 39.156 74.894 39.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 4.632 74.894 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 40.416 74.894 40.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 41.676 74.894 41.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 42.936 74.894 42.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 44.196 74.894 44.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 45.456 74.894 45.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 46.716 74.894 46.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 47.976 74.894 48.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 5.892 74.894 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 7.152 74.894 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 8.412 74.894 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 9.672 74.894 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 1.474 74.894 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 10.294 74.894 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 11.554 74.894 11.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 12.814 74.894 12.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 14.074 74.894 14.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 15.334 74.894 15.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 16.594 74.894 16.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 17.854 74.894 17.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 19.114 74.894 19.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 2.734 74.894 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 20.374 74.894 20.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 29.698 74.894 29.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 3.994 74.894 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 30.958 74.894 30.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 32.218 74.894 32.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 33.478 74.894 33.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 34.738 74.894 34.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 35.998 74.894 36.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 37.258 74.894 37.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 38.518 74.894 38.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 39.778 74.894 39.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 41.038 74.894 41.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 42.298 74.894 42.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 43.558 74.894 43.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 44.818 74.894 44.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 46.078 74.894 46.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 47.338 74.894 47.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 48.598 74.894 48.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 5.254 74.894 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 6.514 74.894 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 7.774 74.894 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 9.034 74.894 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 1.34 74.894 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 10.16 74.894 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 11.42 74.894 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 12.68 74.894 12.726 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 13.94 74.894 13.986 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 15.2 74.894 15.246 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 16.46 74.894 16.506 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 17.72 74.894 17.766 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 18.98 74.894 19.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 2.6 74.894 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 20.24 74.894 20.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 29.564 74.894 29.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 3.86 74.894 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 30.824 74.894 30.87 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 32.084 74.894 32.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 33.344 74.894 33.39 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 34.604 74.894 34.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 35.864 74.894 35.91 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 37.124 74.894 37.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 38.384 74.894 38.43 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 39.644 74.894 39.69 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 40.904 74.894 40.95 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 42.164 74.894 42.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 43.424 74.894 43.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 44.684 74.894 44.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 45.944 74.894 45.99 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 47.204 74.894 47.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 48.464 74.894 48.51 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 5.12 74.894 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 6.38 74.894 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 7.64 74.894 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 8.9 74.894 8.946 ;
          END
     END vccd_1p0
     PIN vss
     SHAPE ABUTMENT ;
     USE   GROUND ;
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 0.894 0.308 0.926 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 1.006 0.308 1.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 11.156 0.308 11.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 12.178 0.308 12.21 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 13.438 0.308 13.47 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 14.81 0.308 14.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 16.168 0.308 16.2 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 17.316 0.308 17.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 18.674 0.308 18.706 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 19.934 0.308 19.966 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 2.378 0.308 2.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 21.012 0.308 21.044 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 21.698 0.308 21.73 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 22.44 0.308 22.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 23.182 0.308 23.214 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 23.756 0.308 23.788 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 24.386 0.308 24.418 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 24.89 0.308 24.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 25.24 0.308 25.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 25.688 0.308 25.72 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 26.374 0.308 26.406 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 26.948 0.308 26.98 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 27.858 0.308 27.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 28.376 0.308 28.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 29.286 0.308 29.318 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 3.638 0.308 3.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 30.532 0.308 30.564 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 31.68 0.308 31.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 32.926 0.308 32.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 34.298 0.308 34.33 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 35.558 0.308 35.59 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 36.692 0.308 36.724 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 37.952 0.308 37.984 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 39.198 0.308 39.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 4.884 0.308 4.916 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 40.458 0.308 40.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 41.704 0.308 41.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 42.964 0.308 42.996 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 44.098 0.308 44.13 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 45.47 0.308 45.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 46.842 0.308 46.874 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 48.088 0.308 48.12 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 48.662 0.308 48.694 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 6.032 0.308 6.064 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 7.278 0.308 7.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 8.538 0.308 8.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 9.784 0.308 9.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.584 14.184 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.788 74.894 0.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.986 74.894 1.04 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.262 74.894 1.316 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.538 74.894 1.578 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.844 14.184 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.082 74.894 10.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.358 74.894 10.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.664 14.184 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.868 74.894 10.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.066 74.894 11.12 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.342 74.894 11.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.618 74.894 11.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.924 14.184 11.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.128 74.894 12.168 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.326 74.894 12.38 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.602 74.894 12.656 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.878 74.894 12.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.184 14.184 13.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.388 74.894 13.428 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.586 74.894 13.64 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.862 74.894 13.916 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.138 74.894 14.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.444 14.184 14.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.648 74.894 14.688 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.846 74.894 14.9 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.122 74.894 15.176 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.398 74.894 15.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.704 14.184 15.75 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.908 74.894 15.948 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.106 74.894 16.16 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.382 74.894 16.436 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.658 74.894 16.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.964 14.184 17.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.168 74.894 17.208 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.366 74.894 17.42 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.642 74.894 17.696 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.918 74.894 17.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.224 14.184 18.27 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.428 74.894 18.468 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.626 74.894 18.68 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.902 74.894 18.956 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.178 74.894 19.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.484 14.184 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.688 74.894 19.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.886 74.894 19.94 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.048 74.894 2.088 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.246 74.894 2.3 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.522 74.894 2.576 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.798 74.894 2.838 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.162 74.894 20.216 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.438 74.894 20.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.894 74.894 20.94 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.034 74.894 21.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.506 74.894 21.546 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.898 74.894 21.944 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.148 74.894 22.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.526 74.894 22.566 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.748 74.894 22.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.21 74.894 23.25 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.458 74.894 23.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.706 74.894 23.746 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.078 74.894 24.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.574 74.894 24.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.822 74.894 24.862 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.07 74.894 25.11 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.442 74.894 25.482 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.938 74.894 25.978 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.186 74.894 26.226 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.434 74.894 26.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.682 74.894 26.722 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.452 74.894 27.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.756 74.894 27.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.488 74.894 28.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.808 14.184 28.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.012 74.894 29.052 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.21 74.894 29.264 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.486 74.894 29.54 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 29.762 74.894 29.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.104 14.184 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.308 74.894 3.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.506 74.894 3.56 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.782 74.894 3.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.068 14.184 30.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.272 74.894 30.312 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.47 74.894 30.524 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 30.746 74.894 30.8 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.022 74.894 31.062 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.328 14.184 31.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.532 74.894 31.572 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 31.73 74.894 31.784 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.006 74.894 32.06 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.282 74.894 32.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.588 14.184 32.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.792 74.894 32.832 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 32.99 74.894 33.044 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.266 74.894 33.32 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.542 74.894 33.582 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 33.848 14.184 33.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.052 74.894 34.092 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.25 74.894 34.304 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.526 74.894 34.58 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 34.802 74.894 34.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.108 14.184 35.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.312 74.894 35.352 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.51 74.894 35.564 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 35.786 74.894 35.84 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.062 74.894 36.102 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.368 14.184 36.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.572 74.894 36.612 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 36.77 74.894 36.824 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.046 74.894 37.1 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.322 74.894 37.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.628 14.184 37.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 37.832 74.894 37.872 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.03 74.894 38.084 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.306 74.894 38.36 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.582 74.894 38.622 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 38.888 14.184 38.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.092 74.894 39.132 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.29 74.894 39.344 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.566 74.894 39.62 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 39.842 74.894 39.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.058 74.894 4.098 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.364 14.184 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.568 74.894 4.608 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.766 74.894 4.82 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.148 14.184 40.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.352 74.894 40.392 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.55 74.894 40.604 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 40.826 74.894 40.88 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.102 74.894 41.142 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.408 14.184 41.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.612 74.894 41.652 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 41.81 74.894 41.864 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.086 74.894 42.14 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.362 74.894 42.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.668 14.184 42.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 42.872 74.894 42.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.07 74.894 43.124 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.346 74.894 43.4 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.622 74.894 43.662 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 43.928 14.184 43.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.132 74.894 44.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.33 74.894 44.384 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.606 74.894 44.66 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 44.882 74.894 44.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.188 14.184 45.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.392 74.894 45.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.59 74.894 45.644 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 45.866 74.894 45.92 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.142 74.894 46.182 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.448 14.184 46.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.652 74.894 46.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 46.85 74.894 46.904 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.126 74.894 47.18 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.402 74.894 47.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.708 14.184 47.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 47.912 74.894 47.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.11 74.894 48.164 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.386 74.894 48.44 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 48.662 74.894 48.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.042 74.894 5.096 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.318 74.894 5.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.624 14.184 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.828 74.894 5.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.026 74.894 6.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.302 74.894 6.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.578 74.894 6.618 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.884 14.184 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.088 74.894 7.128 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.286 74.894 7.34 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.562 74.894 7.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.838 74.894 7.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.144 14.184 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.348 74.894 8.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.546 74.894 8.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.822 74.894 8.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.098 74.894 9.138 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.404 14.184 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.608 74.894 9.648 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.806 74.894 9.86 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 0.584 31.236 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 1.844 31.236 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 10.664 31.236 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 11.924 31.236 11.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 13.184 31.236 13.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 14.444 31.236 14.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 15.704 31.236 15.75 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 16.964 31.236 17.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 18.224 31.236 18.27 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 19.484 31.236 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 28.808 31.236 28.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 3.104 31.236 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 30.068 31.236 30.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 31.328 31.236 31.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 32.588 31.236 32.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 33.848 31.236 33.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 35.108 31.236 35.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 36.368 31.236 36.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 37.628 31.236 37.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 38.888 31.236 38.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 4.364 31.236 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 40.148 31.236 40.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 41.408 31.236 41.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 42.668 31.236 42.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 43.928 31.236 43.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 45.188 31.236 45.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 46.448 31.236 46.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 47.708 31.236 47.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 5.624 31.236 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 6.884 31.236 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 8.144 31.236 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 9.404 31.236 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 0.584 48.288 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 1.844 48.288 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 10.664 48.288 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 11.924 48.288 11.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 13.184 48.288 13.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 14.444 48.288 14.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 15.704 48.288 15.75 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 16.964 48.288 17.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 18.224 48.288 18.27 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 19.484 48.288 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 28.808 48.288 28.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 3.104 48.288 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 30.068 48.288 30.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 31.328 48.288 31.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 32.588 48.288 32.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 33.848 48.288 33.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 35.108 48.288 35.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 36.368 48.288 36.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 37.628 48.288 37.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 38.888 48.288 38.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 4.364 48.288 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 40.148 48.288 40.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 41.408 48.288 41.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 42.668 48.288 42.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 43.928 48.288 43.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 45.188 48.288 45.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 46.448 48.288 46.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 47.708 48.288 47.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 5.624 48.288 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 6.884 48.288 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 8.144 48.288 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 9.404 48.288 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 0.584 65.34 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 1.844 65.34 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 10.664 65.34 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 11.924 65.34 11.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 13.184 65.34 13.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 14.444 65.34 14.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 15.704 65.34 15.75 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 16.964 65.34 17.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 18.224 65.34 18.27 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 19.484 65.34 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 28.808 65.34 28.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 3.104 65.34 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 30.068 65.34 30.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 31.328 65.34 31.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 32.588 65.34 32.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 33.848 65.34 33.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 35.108 65.34 35.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 36.368 65.34 36.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 37.628 65.34 37.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 38.888 65.34 38.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 4.364 65.34 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 40.148 65.34 40.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 41.408 65.34 41.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 42.668 65.34 42.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 43.928 65.34 43.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 45.188 65.34 45.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 46.448 65.34 46.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 47.708 65.34 47.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 5.624 65.34 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 6.884 65.34 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 8.144 65.34 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 9.404 65.34 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 0.584 74.894 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 1.844 74.894 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 10.664 74.894 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 11.924 74.894 11.97 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 13.184 74.894 13.23 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 14.444 74.894 14.49 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 15.704 74.894 15.75 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 16.964 74.894 17.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 18.224 74.894 18.27 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 19.484 74.894 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 28.808 74.894 28.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 3.104 74.894 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 30.068 74.894 30.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 31.328 74.894 31.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 32.588 74.894 32.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 33.848 74.894 33.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 35.108 74.894 35.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 36.368 74.894 36.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 37.628 74.894 37.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 38.888 74.894 38.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 4.364 74.894 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 40.148 74.894 40.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 41.408 74.894 41.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 42.668 74.894 42.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 43.928 74.894 43.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 45.188 74.894 45.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 46.448 74.894 46.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 47.708 74.894 47.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 5.624 74.894 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 6.884 74.894 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 8.144 74.894 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 9.404 74.894 9.45 ;
          END
     END vss
     OBS
          LAYER m0 ;
               POLYGON
                    75.432 49.476 0 49.476 0 0 75.432 0 75.432 49.476 ;
          LAYER m1 ;
               POLYGON
                    75.432 49.476 0 49.476 0 0 75.432 0 75.432 49.476 ;
          LAYER m2 ;
               POLYGON
                    75.432 49.476 0 49.476 0 0 75.432 0 75.432 49.476 ;
          LAYER m3 ;
               POLYGON
                    75.432 49.476 0 49.476 0 0 75.432 0 75.432 49.476 ;
          LAYER m4 ;
               POLYGON
                    75.432 49.476 0 49.476 0 0 75.432 0 75.432 49.476 ;
     END
END c73p1rfshdxrom2048x32hb4img108
END LIBRARY
