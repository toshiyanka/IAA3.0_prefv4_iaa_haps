// This file is `included outside of the tb module in the tb.sv file.
// You can place any definition code here. Macro definitions, typedefs, class/interface definitions, etc are good examples 
`define UTB_DUT_PARAM_PORTMAP
