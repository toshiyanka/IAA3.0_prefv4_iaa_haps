// File output was printed on: Wednesday, March 20, 2013 9:00:22 AM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
// ENUM DECLARATIONS
//------------------------------------------------------------------------
typedef enum int {
   CLTAP    =  'd0,
   STAP0    =  'd1,
   STAP1    =  'd2,
   STAP2    =  'd3,
   STAP3    =  'd4,
   STAP4    =  'd5,
   STAP5    =  'd6,
   STAP6    =  'd7,
   STAP7    =  'd8,
   STAP8    =  'd9,
   STAP9    =  'd10,
   STAP10   =  'd11,
   STAP11   =  'd12,
   STAP12   =  'd13,
   STAP13   =  'd14,
   STAP14   =  'd15,
   STAP15   =  'd16,
   STAP16   =  'd17,
   STAP17   =  'd18,
   STAP18   =  'd19,
   STAP19   =  'd20,
   STAP20   =  'd21,
   STAP21   =  'd22,
   STAP22   =  'd23,
   STAP23   =  'd24,
   STAP24   =  'd25,
   STAP25   =  'd26,
   STAP26   =  'd27,
   STAP27   =  'd28,
   STAP28   =  'd29,
   STAP29   =  'd30,
   NOTAP    =  'hFFFF_FFFF
} Tap_t;


