VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf070b144e1r1w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf070b144e1r1w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 30.6 BY 31.68 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 16.68 14.528 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 14.76 11.916 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 16.68 15.428 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 16.68 15.516 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 16.68 10.028 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 16.68 10.116 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 16.68 10.372 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 16.68 10.628 17.88 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 16.68 10.716 17.88 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 16.68 10.928 17.88 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 16.68 14.616 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 16.68 14.872 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 16.68 15.128 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 16.68 15.216 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 14.76 13.072 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 14.76 13.328 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 14.76 13.416 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 14.76 13.628 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 14.76 13.716 15.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 14.76 13.972 15.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 14.76 14.228 15.96 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 14.76 14.316 15.96 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 14.76 12.172 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 14.76 12.428 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 3.84 14.316 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 3.84 14.528 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 4.56 10.372 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 4.56 10.628 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 5.28 11.616 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 5.28 11.828 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 6 12.428 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 6 12.516 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 6.72 13.072 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 6.72 13.328 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 7.44 13.716 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 7.44 13.972 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 8.16 14.528 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.16 14.616 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 8.88 10.716 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 8.88 10.928 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 9.6 11.828 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 9.6 11.916 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 10.32 12.516 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 10.32 12.728 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 0.96 11.528 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 11.04 13.328 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 11.04 13.416 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 11.76 13.972 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 11.76 14.228 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 12.48 14.616 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 12.48 10.028 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 13.2 11.016 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 13.2 11.272 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 18.72 12.172 19.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 18.72 12.428 19.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 0.96 11.616 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 19.44 11.828 20.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 19.44 11.916 20.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 20.16 13.328 21.36 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 20.16 13.416 21.36 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 20.88 13.972 22.08 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 20.88 14.228 22.08 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 21.6 14.616 22.8 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 21.6 10.028 22.8 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 22.32 11.016 23.52 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 22.32 11.272 23.52 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 1.68 12.172 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 23.04 11.916 24.24 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 23.04 12.172 24.24 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 23.76 12.728 24.96 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 23.76 12.816 24.96 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 24.48 13.416 25.68 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 24.48 13.628 25.68 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 25.2 14.228 26.4 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 25.2 14.316 26.4 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 25.92 10.028 27.12 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 25.92 10.116 27.12 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 1.68 12.428 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 26.64 11.528 27.84 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 26.64 11.616 27.84 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 27.36 12.172 28.56 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 27.36 12.428 28.56 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 28.08 12.816 29.28 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 28.08 13.072 29.28 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 28.8 13.628 30 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 28.8 13.716 30 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 29.52 14.316 30.72 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 29.52 14.528 30.72 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 2.4 12.816 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 30.24 10.372 31.44 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 30.24 10.628 31.44 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 2.4 13.072 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 3.12 13.628 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.12 13.716 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 14.76 12.728 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 14.76 12.816 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 14.76 12.516 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.24 10.372 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.84 14.616 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 3.84 10.028 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 4.56 10.716 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 4.56 10.928 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 5.28 11.916 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 5.28 12.172 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 6 12.728 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 6 12.816 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 6.72 13.416 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 6.72 13.628 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 0.24 10.628 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 7.44 14.228 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 7.44 14.316 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 8.16 10.028 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.16 10.116 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 8.88 11.016 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 8.88 11.272 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 9.6 12.172 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 9.6 12.428 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 10.32 12.816 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 10.32 13.072 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 0.96 11.828 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.04 13.628 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 11.04 13.716 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 11.76 14.316 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 11.76 14.528 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 12.48 10.116 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 12.48 10.372 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 13.2 11.528 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 13.2 11.616 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 18.72 12.516 19.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 18.72 12.728 19.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 0.96 11.916 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 19.44 12.816 20.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 19.44 13.072 20.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 20.16 13.628 21.36 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 20.16 13.716 21.36 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 20.88 14.316 22.08 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 20.88 14.528 22.08 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 21.6 10.116 22.8 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 21.6 10.372 22.8 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 22.32 11.528 23.52 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 22.32 11.616 23.52 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 1.68 12.516 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 23.04 12.428 24.24 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 23.04 12.516 24.24 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 23.76 13.072 24.96 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 23.76 13.328 24.96 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 24.48 13.716 25.68 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 24.48 13.972 25.68 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 25.2 14.528 26.4 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 25.2 14.616 26.4 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 25.92 10.372 27.12 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 25.92 10.628 27.12 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 1.68 12.728 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 26.64 11.828 27.84 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 26.64 11.916 27.84 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 27.36 12.516 28.56 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 27.36 12.728 28.56 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 28.08 13.328 29.28 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 28.08 13.416 29.28 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 28.8 13.972 30 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 28.8 14.228 30 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 29.52 14.616 30.72 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 29.52 10.028 30.72 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 2.4 13.328 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 30.24 10.716 31.44 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 30.24 10.928 31.44 ;
    END
  END rddatap0[71]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 2.4 13.416 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.12 13.972 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 3.12 14.228 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 31.62 ;
        RECT 2.662 0.06 2.738 31.62 ;
        RECT 4.462 0.06 4.538 31.62 ;
        RECT 6.262 0.06 6.338 31.62 ;
        RECT 8.062 0.06 8.138 31.62 ;
        RECT 9.862 0.06 9.938 31.62 ;
        RECT 11.662 0.06 11.738 31.62 ;
        RECT 13.462 0.06 13.538 31.62 ;
        RECT 15.262 0.06 15.338 31.62 ;
        RECT 17.062 0.06 17.138 31.62 ;
        RECT 18.862 0.06 18.938 31.62 ;
        RECT 20.662 0.06 20.738 31.62 ;
        RECT 22.462 0.06 22.538 31.62 ;
        RECT 24.262 0.06 24.338 31.62 ;
        RECT 26.062 0.06 26.138 31.62 ;
        RECT 27.862 0.06 27.938 31.62 ;
        RECT 29.662 0.06 29.738 31.62 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 31.62 ;
        RECT 3.562 0.06 3.638 31.62 ;
        RECT 5.362 0.06 5.438 31.62 ;
        RECT 7.162 0.06 7.238 31.62 ;
        RECT 8.962 0.06 9.038 31.62 ;
        RECT 10.762 0.06 10.838 31.62 ;
        RECT 12.562 0.06 12.638 31.62 ;
        RECT 14.362 0.06 14.438 31.62 ;
        RECT 16.162 0.06 16.238 31.62 ;
        RECT 17.962 0.06 18.038 31.62 ;
        RECT 19.762 0.06 19.838 31.62 ;
        RECT 21.562 0.06 21.638 31.62 ;
        RECT 23.362 0.06 23.438 31.62 ;
        RECT 25.162 0.06 25.238 31.62 ;
        RECT 26.962 0.06 27.038 31.62 ;
        RECT 28.762 0.06 28.838 31.62 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 30.616 31.694 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 30.62 31.7 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 30.6705 31.718 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 30.635 31.75 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 30.67 31.718 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 30.659 31.77 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 30.69 31.742 ;
    LAYER m7 SPACING 0 ;
      RECT 29.738 31.74 30.64 31.8 ;
      RECT 29.738 -0.06 30.692 31.74 ;
      RECT 29.738 -0.12 30.64 -0.06 ;
      RECT 28.838 -0.12 29.662 31.8 ;
      RECT 27.938 -0.12 28.762 31.8 ;
      RECT 27.038 -0.12 27.862 31.8 ;
      RECT 26.138 -0.12 26.962 31.8 ;
      RECT 25.238 -0.12 26.062 31.8 ;
      RECT 24.338 -0.12 25.162 31.8 ;
      RECT 23.438 -0.12 24.262 31.8 ;
      RECT 22.538 -0.12 23.362 31.8 ;
      RECT 21.638 -0.12 22.462 31.8 ;
      RECT 20.738 -0.12 21.562 31.8 ;
      RECT 19.838 -0.12 20.662 31.8 ;
      RECT 18.938 -0.12 19.762 31.8 ;
      RECT 18.038 -0.12 18.862 31.8 ;
      RECT 17.138 -0.12 17.962 31.8 ;
      RECT 16.238 -0.12 17.062 31.8 ;
      RECT 15.338 17.88 16.162 31.8 ;
      RECT 15.338 16.68 15.384 17.88 ;
      RECT 15.428 16.68 15.472 17.88 ;
      RECT 15.516 16.68 16.162 17.88 ;
      RECT 15.338 -0.12 16.162 16.68 ;
      RECT 14.438 30.72 15.262 31.8 ;
      RECT 14.438 29.52 14.484 30.72 ;
      RECT 14.528 29.52 14.572 30.72 ;
      RECT 14.616 29.52 15.262 30.72 ;
      RECT 14.438 26.4 15.262 29.52 ;
      RECT 14.438 25.2 14.484 26.4 ;
      RECT 14.528 25.2 14.572 26.4 ;
      RECT 14.616 25.2 15.262 26.4 ;
      RECT 14.438 22.8 15.262 25.2 ;
      RECT 14.438 22.08 14.572 22.8 ;
      RECT 14.616 21.6 15.262 22.8 ;
      RECT 14.528 21.6 14.572 22.08 ;
      RECT 14.438 20.88 14.484 22.08 ;
      RECT 14.528 20.88 15.262 21.6 ;
      RECT 14.438 17.88 15.262 20.88 ;
      RECT 14.438 16.68 14.484 17.88 ;
      RECT 14.528 16.68 14.572 17.88 ;
      RECT 14.616 16.68 14.828 17.88 ;
      RECT 14.872 16.68 15.084 17.88 ;
      RECT 15.128 16.68 15.172 17.88 ;
      RECT 15.216 16.68 15.262 17.88 ;
      RECT 14.438 13.68 15.262 16.68 ;
      RECT 14.438 12.96 14.572 13.68 ;
      RECT 14.616 12.48 15.262 13.68 ;
      RECT 14.528 12.48 14.572 12.96 ;
      RECT 14.438 11.76 14.484 12.96 ;
      RECT 14.528 11.76 15.262 12.48 ;
      RECT 14.438 9.36 15.262 11.76 ;
      RECT 14.438 8.16 14.484 9.36 ;
      RECT 14.528 8.16 14.572 9.36 ;
      RECT 14.616 8.16 15.262 9.36 ;
      RECT 14.438 5.04 15.262 8.16 ;
      RECT 14.438 3.84 14.484 5.04 ;
      RECT 14.528 3.84 14.572 5.04 ;
      RECT 14.616 3.84 15.262 5.04 ;
      RECT 14.438 -0.12 15.262 3.84 ;
      RECT 13.538 30.72 14.362 31.8 ;
      RECT 13.538 30 14.272 30.72 ;
      RECT 14.316 29.52 14.362 30.72 ;
      RECT 14.228 29.52 14.272 30 ;
      RECT 13.538 28.8 13.584 30 ;
      RECT 13.628 28.8 13.672 30 ;
      RECT 13.716 28.8 13.928 30 ;
      RECT 13.972 28.8 14.184 30 ;
      RECT 14.228 28.8 14.362 29.52 ;
      RECT 13.538 26.4 14.362 28.8 ;
      RECT 13.538 25.68 14.184 26.4 ;
      RECT 14.228 25.2 14.272 26.4 ;
      RECT 14.316 25.2 14.362 26.4 ;
      RECT 13.972 25.2 14.184 25.68 ;
      RECT 13.538 24.48 13.584 25.68 ;
      RECT 13.628 24.48 13.672 25.68 ;
      RECT 13.716 24.48 13.928 25.68 ;
      RECT 13.972 24.48 14.362 25.2 ;
      RECT 13.538 22.08 14.362 24.48 ;
      RECT 13.538 21.36 13.928 22.08 ;
      RECT 13.972 20.88 14.184 22.08 ;
      RECT 14.228 20.88 14.272 22.08 ;
      RECT 14.316 20.88 14.362 22.08 ;
      RECT 13.716 20.88 13.928 21.36 ;
      RECT 13.538 20.16 13.584 21.36 ;
      RECT 13.628 20.16 13.672 21.36 ;
      RECT 13.716 20.16 14.362 20.88 ;
      RECT 13.538 15.96 14.362 20.16 ;
      RECT 13.538 14.76 13.584 15.96 ;
      RECT 13.628 14.76 13.672 15.96 ;
      RECT 13.716 14.76 13.928 15.96 ;
      RECT 13.972 14.76 14.184 15.96 ;
      RECT 14.228 14.76 14.272 15.96 ;
      RECT 14.316 14.76 14.362 15.96 ;
      RECT 13.538 12.96 14.362 14.76 ;
      RECT 13.538 12.24 13.928 12.96 ;
      RECT 13.972 11.76 14.184 12.96 ;
      RECT 14.228 11.76 14.272 12.96 ;
      RECT 14.316 11.76 14.362 12.96 ;
      RECT 13.716 11.76 13.928 12.24 ;
      RECT 13.538 11.04 13.584 12.24 ;
      RECT 13.628 11.04 13.672 12.24 ;
      RECT 13.716 11.04 14.362 11.76 ;
      RECT 13.538 8.64 14.362 11.04 ;
      RECT 13.538 7.92 13.672 8.64 ;
      RECT 13.716 7.44 13.928 8.64 ;
      RECT 13.972 7.44 14.184 8.64 ;
      RECT 14.228 7.44 14.272 8.64 ;
      RECT 14.316 7.44 14.362 8.64 ;
      RECT 13.628 7.44 13.672 7.92 ;
      RECT 13.538 6.72 13.584 7.92 ;
      RECT 13.628 6.72 14.362 7.44 ;
      RECT 13.538 5.04 14.362 6.72 ;
      RECT 13.538 4.32 14.272 5.04 ;
      RECT 14.316 3.84 14.362 5.04 ;
      RECT 14.228 3.84 14.272 4.32 ;
      RECT 13.538 3.12 13.584 4.32 ;
      RECT 13.628 3.12 13.672 4.32 ;
      RECT 13.716 3.12 13.928 4.32 ;
      RECT 13.972 3.12 14.184 4.32 ;
      RECT 14.228 3.12 14.362 3.84 ;
      RECT 13.538 -0.12 14.362 3.12 ;
      RECT 12.638 29.28 13.462 31.8 ;
      RECT 12.638 28.56 12.772 29.28 ;
      RECT 12.816 28.08 13.028 29.28 ;
      RECT 13.072 28.08 13.284 29.28 ;
      RECT 13.328 28.08 13.372 29.28 ;
      RECT 13.416 28.08 13.462 29.28 ;
      RECT 12.728 28.08 12.772 28.56 ;
      RECT 12.638 27.36 12.684 28.56 ;
      RECT 12.728 27.36 13.462 28.08 ;
      RECT 12.638 25.68 13.462 27.36 ;
      RECT 12.638 24.96 13.372 25.68 ;
      RECT 13.416 24.48 13.462 25.68 ;
      RECT 13.328 24.48 13.372 24.96 ;
      RECT 12.638 23.76 12.684 24.96 ;
      RECT 12.728 23.76 12.772 24.96 ;
      RECT 12.816 23.76 13.028 24.96 ;
      RECT 13.072 23.76 13.284 24.96 ;
      RECT 13.328 23.76 13.462 24.48 ;
      RECT 12.638 21.36 13.462 23.76 ;
      RECT 12.638 20.64 13.284 21.36 ;
      RECT 13.328 20.16 13.372 21.36 ;
      RECT 13.416 20.16 13.462 21.36 ;
      RECT 13.072 20.16 13.284 20.64 ;
      RECT 12.638 19.92 12.772 20.64 ;
      RECT 12.816 19.44 13.028 20.64 ;
      RECT 13.072 19.44 13.462 20.16 ;
      RECT 12.728 19.44 12.772 19.92 ;
      RECT 12.638 18.72 12.684 19.92 ;
      RECT 12.728 18.72 13.462 19.44 ;
      RECT 12.638 15.96 13.462 18.72 ;
      RECT 12.638 14.76 12.684 15.96 ;
      RECT 12.728 14.76 12.772 15.96 ;
      RECT 12.816 14.76 13.028 15.96 ;
      RECT 13.072 14.76 13.284 15.96 ;
      RECT 13.328 14.76 13.372 15.96 ;
      RECT 13.416 14.76 13.462 15.96 ;
      RECT 12.638 12.24 13.462 14.76 ;
      RECT 12.638 11.52 13.284 12.24 ;
      RECT 13.328 11.04 13.372 12.24 ;
      RECT 13.416 11.04 13.462 12.24 ;
      RECT 13.072 11.04 13.284 11.52 ;
      RECT 12.638 10.32 12.684 11.52 ;
      RECT 12.728 10.32 12.772 11.52 ;
      RECT 12.816 10.32 13.028 11.52 ;
      RECT 13.072 10.32 13.462 11.04 ;
      RECT 12.638 7.92 13.462 10.32 ;
      RECT 12.638 7.2 13.028 7.92 ;
      RECT 13.072 6.72 13.284 7.92 ;
      RECT 13.328 6.72 13.372 7.92 ;
      RECT 13.416 6.72 13.462 7.92 ;
      RECT 12.816 6.72 13.028 7.2 ;
      RECT 12.638 6 12.684 7.2 ;
      RECT 12.728 6 12.772 7.2 ;
      RECT 12.816 6 13.462 6.72 ;
      RECT 12.638 3.6 13.462 6 ;
      RECT 12.638 2.88 12.772 3.6 ;
      RECT 12.816 2.4 13.028 3.6 ;
      RECT 13.072 2.4 13.284 3.6 ;
      RECT 13.328 2.4 13.372 3.6 ;
      RECT 13.416 2.4 13.462 3.6 ;
      RECT 12.728 2.4 12.772 2.88 ;
      RECT 12.638 1.68 12.684 2.88 ;
      RECT 12.728 1.68 13.462 2.4 ;
      RECT 12.638 -0.12 13.462 1.68 ;
      RECT 11.738 28.56 12.562 31.8 ;
      RECT 11.738 27.84 12.128 28.56 ;
      RECT 12.172 27.36 12.384 28.56 ;
      RECT 12.428 27.36 12.472 28.56 ;
      RECT 12.516 27.36 12.562 28.56 ;
      RECT 11.916 27.36 12.128 27.84 ;
      RECT 11.738 26.64 11.784 27.84 ;
      RECT 11.828 26.64 11.872 27.84 ;
      RECT 11.916 26.64 12.562 27.36 ;
      RECT 11.738 24.24 12.562 26.64 ;
      RECT 11.738 23.04 11.872 24.24 ;
      RECT 11.916 23.04 12.128 24.24 ;
      RECT 12.172 23.04 12.384 24.24 ;
      RECT 12.428 23.04 12.472 24.24 ;
      RECT 12.516 23.04 12.562 24.24 ;
      RECT 11.738 20.64 12.562 23.04 ;
      RECT 11.916 19.92 12.562 20.64 ;
      RECT 11.738 19.44 11.784 20.64 ;
      RECT 11.828 19.44 11.872 20.64 ;
      RECT 11.916 19.44 12.128 19.92 ;
      RECT 12.172 18.72 12.384 19.92 ;
      RECT 12.428 18.72 12.472 19.92 ;
      RECT 12.516 18.72 12.562 19.92 ;
      RECT 11.738 18.72 12.128 19.44 ;
      RECT 11.738 15.96 12.562 18.72 ;
      RECT 11.738 14.76 11.872 15.96 ;
      RECT 11.916 14.76 12.128 15.96 ;
      RECT 12.172 14.76 12.384 15.96 ;
      RECT 12.428 14.76 12.472 15.96 ;
      RECT 12.516 14.76 12.562 15.96 ;
      RECT 11.738 11.52 12.562 14.76 ;
      RECT 11.738 10.8 12.472 11.52 ;
      RECT 12.516 10.32 12.562 11.52 ;
      RECT 12.428 10.32 12.472 10.8 ;
      RECT 11.738 9.6 11.784 10.8 ;
      RECT 11.828 9.6 11.872 10.8 ;
      RECT 11.916 9.6 12.128 10.8 ;
      RECT 12.172 9.6 12.384 10.8 ;
      RECT 12.428 9.6 12.562 10.32 ;
      RECT 11.738 7.2 12.562 9.6 ;
      RECT 11.738 6.48 12.384 7.2 ;
      RECT 12.428 6 12.472 7.2 ;
      RECT 12.516 6 12.562 7.2 ;
      RECT 12.172 6 12.384 6.48 ;
      RECT 11.738 5.28 11.784 6.48 ;
      RECT 11.828 5.28 11.872 6.48 ;
      RECT 11.916 5.28 12.128 6.48 ;
      RECT 12.172 5.28 12.562 6 ;
      RECT 11.738 2.88 12.562 5.28 ;
      RECT 11.738 2.16 12.128 2.88 ;
      RECT 12.172 1.68 12.384 2.88 ;
      RECT 12.428 1.68 12.472 2.88 ;
      RECT 12.516 1.68 12.562 2.88 ;
      RECT 11.916 1.68 12.128 2.16 ;
      RECT 11.738 0.96 11.784 2.16 ;
      RECT 11.828 0.96 11.872 2.16 ;
      RECT 11.916 0.96 12.562 1.68 ;
      RECT 11.738 -0.12 12.562 0.96 ;
      RECT 10.838 31.44 11.662 31.8 ;
      RECT 10.838 30.24 10.884 31.44 ;
      RECT 10.928 30.24 11.662 31.44 ;
      RECT 10.838 27.84 11.662 30.24 ;
      RECT 10.838 26.64 11.484 27.84 ;
      RECT 11.528 26.64 11.572 27.84 ;
      RECT 11.616 26.64 11.662 27.84 ;
      RECT 10.838 23.52 11.662 26.64 ;
      RECT 10.838 22.32 10.972 23.52 ;
      RECT 11.016 22.32 11.228 23.52 ;
      RECT 11.272 22.32 11.484 23.52 ;
      RECT 11.528 22.32 11.572 23.52 ;
      RECT 11.616 22.32 11.662 23.52 ;
      RECT 10.838 17.88 11.662 22.32 ;
      RECT 10.838 16.68 10.884 17.88 ;
      RECT 10.928 16.68 11.662 17.88 ;
      RECT 10.838 14.4 11.662 16.68 ;
      RECT 10.838 13.2 10.972 14.4 ;
      RECT 11.016 13.2 11.228 14.4 ;
      RECT 11.272 13.2 11.484 14.4 ;
      RECT 11.528 13.2 11.572 14.4 ;
      RECT 11.616 13.2 11.662 14.4 ;
      RECT 10.838 10.08 11.662 13.2 ;
      RECT 10.838 8.88 10.884 10.08 ;
      RECT 10.928 8.88 10.972 10.08 ;
      RECT 11.016 8.88 11.228 10.08 ;
      RECT 11.272 8.88 11.662 10.08 ;
      RECT 10.838 6.48 11.662 8.88 ;
      RECT 10.838 5.76 11.572 6.48 ;
      RECT 11.616 5.28 11.662 6.48 ;
      RECT 10.928 5.28 11.572 5.76 ;
      RECT 10.838 4.56 10.884 5.76 ;
      RECT 10.928 4.56 11.662 5.28 ;
      RECT 10.838 2.16 11.662 4.56 ;
      RECT 10.838 0.96 11.484 2.16 ;
      RECT 11.528 0.96 11.572 2.16 ;
      RECT 11.616 0.96 11.662 2.16 ;
      RECT 10.838 -0.12 11.662 0.96 ;
      RECT 9.938 31.44 10.762 31.8 ;
      RECT 9.938 30.72 10.328 31.44 ;
      RECT 10.372 30.24 10.584 31.44 ;
      RECT 10.628 30.24 10.672 31.44 ;
      RECT 10.716 30.24 10.762 31.44 ;
      RECT 10.028 30.24 10.328 30.72 ;
      RECT 9.938 29.52 9.984 30.72 ;
      RECT 10.028 29.52 10.762 30.24 ;
      RECT 9.938 27.12 10.762 29.52 ;
      RECT 9.938 25.92 9.984 27.12 ;
      RECT 10.028 25.92 10.072 27.12 ;
      RECT 10.116 25.92 10.328 27.12 ;
      RECT 10.372 25.92 10.584 27.12 ;
      RECT 10.628 25.92 10.762 27.12 ;
      RECT 9.938 22.8 10.762 25.92 ;
      RECT 9.938 21.6 9.984 22.8 ;
      RECT 10.028 21.6 10.072 22.8 ;
      RECT 10.116 21.6 10.328 22.8 ;
      RECT 10.372 21.6 10.762 22.8 ;
      RECT 9.938 17.88 10.762 21.6 ;
      RECT 9.938 16.68 9.984 17.88 ;
      RECT 10.028 16.68 10.072 17.88 ;
      RECT 10.116 16.68 10.328 17.88 ;
      RECT 10.372 16.68 10.584 17.88 ;
      RECT 10.628 16.68 10.672 17.88 ;
      RECT 10.716 16.68 10.762 17.88 ;
      RECT 9.938 13.68 10.762 16.68 ;
      RECT 9.938 12.48 9.984 13.68 ;
      RECT 10.028 12.48 10.072 13.68 ;
      RECT 10.116 12.48 10.328 13.68 ;
      RECT 10.372 12.48 10.762 13.68 ;
      RECT 9.938 10.08 10.762 12.48 ;
      RECT 9.938 9.36 10.672 10.08 ;
      RECT 10.716 8.88 10.762 10.08 ;
      RECT 10.116 8.88 10.672 9.36 ;
      RECT 9.938 8.16 9.984 9.36 ;
      RECT 10.028 8.16 10.072 9.36 ;
      RECT 10.116 8.16 10.762 8.88 ;
      RECT 9.938 5.76 10.762 8.16 ;
      RECT 9.938 5.04 10.328 5.76 ;
      RECT 10.372 4.56 10.584 5.76 ;
      RECT 10.628 4.56 10.672 5.76 ;
      RECT 10.716 4.56 10.762 5.76 ;
      RECT 10.028 4.56 10.328 5.04 ;
      RECT 9.938 3.84 9.984 5.04 ;
      RECT 10.028 3.84 10.762 4.56 ;
      RECT 9.938 1.44 10.762 3.84 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.328 1.44 ;
      RECT 10.372 0.24 10.584 1.44 ;
      RECT 10.628 0.24 10.762 1.44 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 31.8 ;
      RECT 8.138 -0.12 8.962 31.8 ;
      RECT 7.238 -0.12 8.062 31.8 ;
      RECT 6.338 -0.12 7.162 31.8 ;
      RECT 5.438 -0.12 6.262 31.8 ;
      RECT 4.538 -0.12 5.362 31.8 ;
      RECT 3.638 -0.12 4.462 31.8 ;
      RECT 2.738 -0.12 3.562 31.8 ;
      RECT 1.838 -0.12 2.662 31.8 ;
      RECT 0.938 -0.12 1.762 31.8 ;
      RECT -0.04 31.74 0.862 31.8 ;
      RECT -0.092 -0.06 0.862 31.74 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 29.858 0 30.52 31.68 ;
      RECT 28.958 0 29.542 31.68 ;
      RECT 28.058 0 28.642 31.68 ;
      RECT 27.158 0 27.742 31.68 ;
      RECT 26.258 0 26.842 31.68 ;
      RECT 25.358 0 25.942 31.68 ;
      RECT 24.458 0 25.042 31.68 ;
      RECT 23.558 0 24.142 31.68 ;
      RECT 22.658 0 23.242 31.68 ;
      RECT 21.758 0 22.342 31.68 ;
      RECT 20.858 0 21.442 31.68 ;
      RECT 19.958 0 20.542 31.68 ;
      RECT 19.058 0 19.642 31.68 ;
      RECT 18.158 0 18.742 31.68 ;
      RECT 17.258 0 17.842 31.68 ;
      RECT 16.358 0 16.942 31.68 ;
      RECT 15.458 18 16.042 31.68 ;
      RECT 15.636 16.56 16.042 18 ;
      RECT 15.458 0 16.042 16.56 ;
      RECT 14.558 30.84 15.142 31.68 ;
      RECT 14.736 29.4 15.142 30.84 ;
      RECT 14.558 26.52 15.142 29.4 ;
      RECT 14.736 25.08 15.142 26.52 ;
      RECT 14.558 22.92 15.142 25.08 ;
      RECT 14.736 21.48 15.142 22.92 ;
      RECT 14.648 20.76 15.142 21.48 ;
      RECT 14.558 18 15.142 20.76 ;
      RECT 13.658 30.84 14.242 31.68 ;
      RECT 13.658 30.12 14.152 30.84 ;
      RECT 12.758 29.4 13.342 31.68 ;
      RECT 11.858 28.68 12.442 31.68 ;
      RECT 11.858 27.96 12.008 28.68 ;
      RECT 10.958 31.56 11.542 31.68 ;
      RECT 11.048 30.12 11.542 31.56 ;
      RECT 10.958 27.96 11.542 30.12 ;
      RECT 10.958 26.52 11.364 27.96 ;
      RECT 10.958 23.64 11.542 26.52 ;
      RECT 10.058 31.56 10.642 31.68 ;
      RECT 10.058 30.84 10.208 31.56 ;
      RECT 10.148 30.12 10.208 30.84 ;
      RECT 10.148 29.4 10.642 30.12 ;
      RECT 10.058 27.24 10.642 29.4 ;
      RECT 9.158 0 9.742 31.68 ;
      RECT 8.258 0 8.842 31.68 ;
      RECT 7.358 0 7.942 31.68 ;
      RECT 6.458 0 7.042 31.68 ;
      RECT 5.558 0 6.142 31.68 ;
      RECT 4.658 0 5.242 31.68 ;
      RECT 3.758 0 4.342 31.68 ;
      RECT 2.858 0 3.442 31.68 ;
      RECT 1.958 0 2.542 31.68 ;
      RECT 1.058 0 1.642 31.68 ;
      RECT 0.08 0 0.742 31.68 ;
      RECT 13.658 26.52 14.242 28.68 ;
      RECT 13.658 25.8 14.064 26.52 ;
      RECT 12.848 27.24 13.342 27.96 ;
      RECT 12.758 25.8 13.342 27.24 ;
      RECT 12.758 25.08 13.252 25.8 ;
      RECT 12.036 26.52 12.442 27.24 ;
      RECT 11.858 24.36 12.442 26.52 ;
      RECT 10.058 22.92 10.642 25.8 ;
      RECT 10.492 21.48 10.642 22.92 ;
      RECT 10.058 18 10.642 21.48 ;
      RECT 14.092 24.36 14.242 25.08 ;
      RECT 13.658 22.2 14.242 24.36 ;
      RECT 13.658 21.48 13.808 22.2 ;
      RECT 12.758 21.48 13.342 23.64 ;
      RECT 12.758 20.76 13.164 21.48 ;
      RECT 11.858 20.76 12.442 22.92 ;
      RECT 12.036 20.04 12.442 20.76 ;
      RECT 10.958 18 11.542 22.2 ;
      RECT 11.048 16.56 11.542 18 ;
      RECT 10.958 14.52 11.542 16.56 ;
      RECT 13.836 20.04 14.242 20.76 ;
      RECT 13.658 16.08 14.242 20.04 ;
      RECT 13.192 19.32 13.342 20.04 ;
      RECT 12.848 18.6 13.342 19.32 ;
      RECT 12.758 16.08 13.342 18.6 ;
      RECT 11.858 18.6 12.008 19.32 ;
      RECT 11.858 16.08 12.442 18.6 ;
      RECT 14.558 13.8 15.142 16.56 ;
      RECT 14.736 12.36 15.142 13.8 ;
      RECT 14.648 11.64 15.142 12.36 ;
      RECT 14.558 9.48 15.142 11.64 ;
      RECT 14.736 8.04 15.142 9.48 ;
      RECT 14.558 5.16 15.142 8.04 ;
      RECT 14.736 3.72 15.142 5.16 ;
      RECT 14.558 0 15.142 3.72 ;
      RECT 10.058 13.8 10.642 16.56 ;
      RECT 10.492 12.36 10.642 13.8 ;
      RECT 10.058 10.2 10.642 12.36 ;
      RECT 10.058 9.48 10.552 10.2 ;
      RECT 10.236 8.76 10.552 9.48 ;
      RECT 10.236 8.04 10.642 8.76 ;
      RECT 10.058 5.88 10.642 8.04 ;
      RECT 10.058 5.16 10.208 5.88 ;
      RECT 10.148 4.44 10.208 5.16 ;
      RECT 10.148 3.72 10.642 4.44 ;
      RECT 10.058 1.56 10.642 3.72 ;
      RECT 13.658 13.08 14.242 14.64 ;
      RECT 13.658 12.36 13.808 13.08 ;
      RECT 12.758 12.36 13.342 14.64 ;
      RECT 12.758 11.64 13.164 12.36 ;
      RECT 11.858 11.64 12.442 14.64 ;
      RECT 11.858 10.92 12.352 11.64 ;
      RECT 10.958 10.2 11.542 13.08 ;
      RECT 11.392 8.76 11.542 10.2 ;
      RECT 10.958 6.6 11.542 8.76 ;
      RECT 10.958 5.88 11.452 6.6 ;
      RECT 11.048 5.16 11.452 5.88 ;
      RECT 11.048 4.44 11.542 5.16 ;
      RECT 10.958 2.28 11.542 4.44 ;
      RECT 10.958 0.84 11.364 2.28 ;
      RECT 10.958 0 11.542 0.84 ;
      RECT 13.836 10.92 14.242 11.64 ;
      RECT 13.658 8.76 14.242 10.92 ;
      RECT 13.192 10.2 13.342 10.92 ;
      RECT 12.758 8.04 13.342 10.2 ;
      RECT 12.758 7.32 12.908 8.04 ;
      RECT 11.858 7.32 12.442 9.48 ;
      RECT 11.858 6.6 12.264 7.32 ;
      RECT 13.748 6.6 14.242 7.32 ;
      RECT 13.658 5.16 14.242 6.6 ;
      RECT 13.658 4.44 14.152 5.16 ;
      RECT 12.936 5.88 13.342 6.6 ;
      RECT 12.758 3.72 13.342 5.88 ;
      RECT 12.292 5.16 12.442 5.88 ;
      RECT 11.858 3 12.442 5.16 ;
      RECT 11.858 2.28 12.008 3 ;
      RECT 13.658 0 14.242 3 ;
      RECT 12.848 1.56 13.342 2.28 ;
      RECT 12.758 0 13.342 1.56 ;
      RECT 12.036 0.84 12.442 1.56 ;
      RECT 11.858 0 12.442 0.84 ;
      RECT 10.058 0 10.642 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 30.6 31.678 ;
    LAYER m1 ;
      RECT 0 0 30.6 31.68 ;
    LAYER m2 ;
      RECT 0 0.015 30.6 31.665 ;
    LAYER m3 ;
      RECT 0.015 0 30.585 31.68 ;
    LAYER m4 ;
      RECT 0 0.02 30.6 31.66 ;
    LAYER m5 ;
      RECT 0.012 0 30.588 31.68 ;
    LAYER m6 ;
      RECT 0 0.012 30.6 31.668 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf070b144e1r1w0cbbeheaa4acw

END LIBRARY
