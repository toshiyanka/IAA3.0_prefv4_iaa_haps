module ctech_lib_ident (
   input logic a,
   output logic o
);
   d04bfn00ln0c0 ctech_lib_dcszo (.a(a), .o(o));
endmodule
