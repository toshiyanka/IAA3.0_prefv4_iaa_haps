`ifdef INTEL_FPGA
   `include "<>.sv"
`else
 `include "<>.sv"
`endif 

