//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbra : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbra
(
  // Synchronous Clock/Reset
  sosc_25_clk_core,
  sbi_rst_25_core_b,

  // Asynchronous Clock/Reset(s)
  bb_cclk,
  sosc_125_clk_core,

  // Power Well Isolation Input Signals
  eva_present,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  p3_fab_init_idle_exit,
  p3_fab_init_idle_exit_ack,
  p4_fab_init_idle_exit,
  p4_fab_init_idle_exit_ack,
  p5_fab_init_idle_exit,
  p5_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_sosc_25_clk_core,
  visa_vp_sosc_25_clk_core,
  visa_p0_tier1_bb_cclk,
  visa_p0_tier2_bb_cclk,
  visa_p0_ififo_tier1_sosc_25_clk_core,
  visa_p0_ififo_tier2_sosc_25_clk_core,
  visa_p0_efifo_tier1_sosc_25_clk_core,
  visa_p0_efifo_tier2_sosc_25_clk_core,
  visa_p1_tier1_sosc_125_clk_core,
  visa_p1_tier2_sosc_125_clk_core,
  visa_p1_ififo_tier1_sosc_25_clk_core,
  visa_p1_ififo_tier2_sosc_25_clk_core,
  visa_p1_efifo_tier1_sosc_25_clk_core,
  visa_p1_efifo_tier2_sosc_25_clk_core,
  visa_p2_tier1_sosc_25_clk_core,
  visa_p2_tier2_sosc_25_clk_core,
  visa_p3_tier1_sosc_25_clk_core,
  visa_p3_tier2_sosc_25_clk_core,
  visa_p4_tier1_sosc_25_clk_core,
  visa_p4_tier2_sosc_25_clk_core,
  visa_p5_tier1_sosc_25_clk_core,
  visa_p5_tier2_sosc_25_clk_core,


  // Register wires
  dfxa_sbra_cgovrd,
  dfxa_sbra_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  npsb_sbra_side_ism_agent,
  sbra_npsb_side_ism_fabric,
  npsb_sbra_pccup,
  npsb_sbra_npcup,
  sbra_npsb_pcput,
  sbra_npsb_npput,
  sbra_npsb_eom,
  sbra_npsb_payload,
  sbra_npsb_pccup,
  sbra_npsb_npcup,
  npsb_sbra_pcput,
  npsb_sbra_npput,
  npsb_sbra_eom,
  npsb_sbra_payload,

  // Port 1 declarations
  xpsb_sbra_side_ism_agent,
  sbra_xpsb_side_ism_fabric,
  xpsb_sbra_pccup,
  xpsb_sbra_npcup,
  sbra_xpsb_pcput,
  sbra_xpsb_npput,
  sbra_xpsb_eom,
  sbra_xpsb_payload,
  sbra_xpsb_pccup,
  sbra_xpsb_npcup,
  xpsb_sbra_pcput,
  xpsb_sbra_npput,
  xpsb_sbra_eom,
  xpsb_sbra_payload,

  // Port 2 declarations
  ccsb_sbra_side_ism_agent,
  sbra_ccsb_side_ism_fabric,
  ccsb_sbra_pccup,
  ccsb_sbra_npcup,
  sbra_ccsb_pcput,
  sbra_ccsb_npput,
  sbra_ccsb_eom,
  sbra_ccsb_payload,
  sbra_ccsb_pccup,
  sbra_ccsb_npcup,
  ccsb_sbra_pcput,
  ccsb_sbra_npput,
  ccsb_sbra_eom,
  ccsb_sbra_payload,

  // Port 3 declarations
  io_pxp_sbra_side_ism_agent,
  sbra_io_pxp_side_ism_fabric,
  io_pxp_sbra_pccup,
  io_pxp_sbra_npcup,
  sbra_io_pxp_pcput,
  sbra_io_pxp_npput,
  sbra_io_pxp_eom,
  sbra_io_pxp_payload,
  sbra_io_pxp_pccup,
  sbra_io_pxp_npcup,
  io_pxp_sbra_pcput,
  io_pxp_sbra_npput,
  io_pxp_sbra_eom,
  io_pxp_sbra_payload,

  // Port 4 declarations
  io_dmi_sbra_side_ism_agent,
  sbra_io_dmi_side_ism_fabric,
  io_dmi_sbra_pccup,
  io_dmi_sbra_npcup,
  sbra_io_dmi_pcput,
  sbra_io_dmi_npput,
  sbra_io_dmi_eom,
  sbra_io_dmi_payload,
  sbra_io_dmi_pccup,
  sbra_io_dmi_npcup,
  io_dmi_sbra_pcput,
  io_dmi_sbra_npput,
  io_dmi_sbra_eom,
  io_dmi_sbra_payload,

  // Port 5 declarations
  io_st_sbra_side_ism_agent,
  sbra_io_st_side_ism_fabric,
  io_st_sbra_pccup,
  io_st_sbra_npcup,
  sbra_io_st_pcput,
  sbra_io_st_npput,
  sbra_io_st_eom,
  sbra_io_st_payload,
  sbra_io_st_pccup,
  sbra_io_st_npcup,
  io_st_sbra_pcput,
  io_st_sbra_npput,
  io_st_sbra_eom,
  io_st_sbra_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic sosc_25_clk_core;
  input logic sbi_rst_25_core_b;

  // Asynchronous Clock/Reset(s)
  input logic bb_cclk;
  input logic sosc_125_clk_core;

  // Power Well Isolation Input Signals
  input logic eva_present;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic p3_fab_init_idle_exit;
  input logic p3_fab_init_idle_exit_ack;
  output logic p4_fab_init_idle_exit;
  input logic p4_fab_init_idle_exit_ack;
  output logic p5_fab_init_idle_exit;
  input logic p5_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_sosc_25_clk_core;
  output visa_vp  visa_vp_sosc_25_clk_core;
  output visa_port_tier1 visa_p0_tier1_bb_cclk;
  output visa_port_tier2 visa_p0_tier2_bb_cclk;
  output visa_ififo_tier1 visa_p0_ififo_tier1_sosc_25_clk_core;
  output visa_ififo_tier2 visa_p0_ififo_tier2_sosc_25_clk_core;
  output visa_efifo_tier1 visa_p0_efifo_tier1_sosc_25_clk_core;
  output visa_efifo_tier2 visa_p0_efifo_tier2_sosc_25_clk_core;
  output visa_port_tier1 visa_p1_tier1_sosc_125_clk_core;
  output visa_port_tier2 visa_p1_tier2_sosc_125_clk_core;
  output visa_ififo_tier1 visa_p1_ififo_tier1_sosc_25_clk_core;
  output visa_ififo_tier2 visa_p1_ififo_tier2_sosc_25_clk_core;
  output visa_efifo_tier1 visa_p1_efifo_tier1_sosc_25_clk_core;
  output visa_efifo_tier2 visa_p1_efifo_tier2_sosc_25_clk_core;
  output visa_port_tier1 visa_p2_tier1_sosc_25_clk_core;
  output visa_port_tier2 visa_p2_tier2_sosc_25_clk_core;
  output visa_port_tier1 visa_p3_tier1_sosc_25_clk_core;
  output visa_port_tier2 visa_p3_tier2_sosc_25_clk_core;
  output visa_port_tier1 visa_p4_tier1_sosc_25_clk_core;
  output visa_port_tier2 visa_p4_tier2_sosc_25_clk_core;
  output visa_port_tier1 visa_p5_tier1_sosc_25_clk_core;
  output visa_port_tier2 visa_p5_tier2_sosc_25_clk_core;

  // Register wires
  input logic [4:0]  dfxa_sbra_cgovrd;
  input logic [15:0] dfxa_sbra_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic [1:0] fscan_rstbypen;
  input logic [1:0] fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] npsb_sbra_side_ism_agent;
  output logic [2:0] sbra_npsb_side_ism_fabric;
  input logic npsb_sbra_pccup;
  input logic npsb_sbra_npcup;
  output logic sbra_npsb_pcput;
  output logic sbra_npsb_npput;
  output logic sbra_npsb_eom;
  output logic [7:0] sbra_npsb_payload;
  output logic sbra_npsb_pccup;
  output logic sbra_npsb_npcup;
  input logic npsb_sbra_pcput;
  input logic npsb_sbra_npput;
  input logic npsb_sbra_eom;
  input logic [7:0] npsb_sbra_payload;

  // Port 1 declarations
  input logic [2:0] xpsb_sbra_side_ism_agent;
  output logic [2:0] sbra_xpsb_side_ism_fabric;
  input logic xpsb_sbra_pccup;
  input logic xpsb_sbra_npcup;
  output logic sbra_xpsb_pcput;
  output logic sbra_xpsb_npput;
  output logic sbra_xpsb_eom;
  output logic [7:0] sbra_xpsb_payload;
  output logic sbra_xpsb_pccup;
  output logic sbra_xpsb_npcup;
  input logic xpsb_sbra_pcput;
  input logic xpsb_sbra_npput;
  input logic xpsb_sbra_eom;
  input logic [7:0] xpsb_sbra_payload;

  // Port 2 declarations
  input logic [2:0] ccsb_sbra_side_ism_agent;
  output logic [2:0] sbra_ccsb_side_ism_fabric;
  input logic ccsb_sbra_pccup;
  input logic ccsb_sbra_npcup;
  output logic sbra_ccsb_pcput;
  output logic sbra_ccsb_npput;
  output logic sbra_ccsb_eom;
  output logic [7:0] sbra_ccsb_payload;
  output logic sbra_ccsb_pccup;
  output logic sbra_ccsb_npcup;
  input logic ccsb_sbra_pcput;
  input logic ccsb_sbra_npput;
  input logic ccsb_sbra_eom;
  input logic [7:0] ccsb_sbra_payload;

  // Port 3 declarations
  input logic [2:0] io_pxp_sbra_side_ism_agent;
  output logic [2:0] sbra_io_pxp_side_ism_fabric;
  input logic io_pxp_sbra_pccup;
  input logic io_pxp_sbra_npcup;
  output logic sbra_io_pxp_pcput;
  output logic sbra_io_pxp_npput;
  output logic sbra_io_pxp_eom;
  output logic [7:0] sbra_io_pxp_payload;
  output logic sbra_io_pxp_pccup;
  output logic sbra_io_pxp_npcup;
  input logic io_pxp_sbra_pcput;
  input logic io_pxp_sbra_npput;
  input logic io_pxp_sbra_eom;
  input logic [7:0] io_pxp_sbra_payload;

  // Port 4 declarations
  input logic [2:0] io_dmi_sbra_side_ism_agent;
  output logic [2:0] sbra_io_dmi_side_ism_fabric;
  input logic io_dmi_sbra_pccup;
  input logic io_dmi_sbra_npcup;
  output logic sbra_io_dmi_pcput;
  output logic sbra_io_dmi_npput;
  output logic sbra_io_dmi_eom;
  output logic [7:0] sbra_io_dmi_payload;
  output logic sbra_io_dmi_pccup;
  output logic sbra_io_dmi_npcup;
  input logic io_dmi_sbra_pcput;
  input logic io_dmi_sbra_npput;
  input logic io_dmi_sbra_eom;
  input logic [7:0] io_dmi_sbra_payload;

  // Port 5 declarations
  input logic [2:0] io_st_sbra_side_ism_agent;
  output logic [2:0] sbra_io_st_side_ism_fabric;
  input logic io_st_sbra_pccup;
  input logic io_st_sbra_npcup;
  output logic sbra_io_st_pcput;
  output logic sbra_io_st_npput;
  output logic sbra_io_st_eom;
  output logic [7:0] sbra_io_st_payload;
  output logic sbra_io_st_pccup;
  output logic sbra_io_st_npcup;
  input logic io_st_sbra_pcput;
  input logic io_st_sbra_npput;
  input logic io_st_sbra_eom;
  input logic [7:0] io_st_sbra_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbra_sbcportmap;
always_comb sbra_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbra (sbra)                                   SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {   15 { 17'b0_0000_0000_0000_0000 }},   //   254:240      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //   239          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //   238          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   237          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //   236          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //   235          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //   234          SBCPORTMAPTABLE
      {  224 { 17'b0_0000_0000_0000_0000 }},   //   233: 10      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0100 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //     7          SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_0000_0100 }}    //     6:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  5;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              p3_ism_idle;
logic                              p3_cg_inprogress;
logic                              p3_credit_reinit;
logic                              p4_ism_idle;
logic                              p4_cg_inprogress;
logic                              p4_credit_reinit;
logic                              p5_ism_idle;
logic                              p5_cg_inprogress;
logic                              p5_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              eva_present_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = dfxa_sbra_cgctrl[15];
always_comb cfg_clkgatedef    = dfxa_sbra_cgctrl[14];
always_comb cfg_idlecnt       = dfxa_sbra_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = dfxa_sbra_cgovrd[3];
always_comb jta_force_idle    = dfxa_sbra_cgovrd[1];
always_comb jta_force_notidle = dfxa_sbra_cgovrd[0];
always_comb jta_force_creditreq = dfxa_sbra_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

// Asynchronous port signals
logic                              p0_clkgaten;
logic                              p0_clkgatedef;
logic                              p0_clkgate_ovrd;
logic                              p0_force_idle;
logic                              p0_force_notidle;
logic                              p0_force_creditreq;
logic                              p0_clken;
logic                              p0_gated_clk;
logic                              p0_agent_idle;
logic                              p0_eagent_idle;
logic                              p0_port_idle;
logic                              p0_ififo_idle;
logic                              p0_efifo_idle;
logic                              p0_pctrdy;
logic                              p0_pcirdy;
logic             [INTMAXPLDBIT:0] p0_pcdata;
logic                              p0_pceom;
logic                              p0_nptrdy;
logic                              p0_npirdy;
logic                              p0_npfence;
logic             [INTMAXPLDBIT:0] p0_npdata;
logic                              p0_npeom;
logic                              p0_enpstall;
logic                              p0_epctrdy;
logic                              p0_enptrdy;
logic                              p0_epcirdy;
logic                              p0_enpirdy;
logic                              p0_eom;
logic             [INTMAXPLDBIT:0] p0_data;

logic                              p1_clkgaten;
logic                              p1_clkgatedef;
logic                              p1_clkgate_ovrd;
logic                              p1_force_idle;
logic                              p1_force_notidle;
logic                              p1_force_creditreq;
logic                              p1_clken;
logic                              p1_gated_clk;
logic                              p1_agent_idle;
logic                              p1_eagent_idle;
logic                              p1_port_idle;
logic                              p1_ififo_idle;
logic                              p1_efifo_idle;
logic                              p1_pctrdy;
logic                              p1_pcirdy;
logic             [INTMAXPLDBIT:0] p1_pcdata;
logic                              p1_pceom;
logic                              p1_nptrdy;
logic                              p1_npirdy;
logic                              p1_npfence;
logic             [INTMAXPLDBIT:0] p1_npdata;
logic                              p1_npeom;
logic                              p1_enpstall;
logic                              p1_epctrdy;
logic                              p1_enptrdy;
logic                              p1_epcirdy;
logic                              p1_enpirdy;
logic                              p1_eom;
logic             [INTMAXPLDBIT:0] p1_data;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbra_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbra_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// Async clock reset synchronization
//
//------------------------------------------------------------------------------
logic bb_cclk_rst_b, bb_cclk_rst_b_pre;
sbc_doublesync sync_rst_bb_cclk (
  .d     ( 1'b1 ),
  .clr_b ( sbi_rst_25_core_b ),
  .clk   ( bb_cclk ),
  .q     ( bb_cclk_rst_b_pre ));

always_comb bb_cclk_rst_b = fscan_rstbypen[0] ? fscan_byprst_b[0] : bb_cclk_rst_b_pre;

logic sosc_125_clk_core_rst_b, sosc_125_clk_core_rst_b_pre;
sbc_doublesync sync_rst_sosc_125_clk_core (
  .d     ( 1'b1 ),
  .clr_b ( sbi_rst_25_core_b ),
  .clk   ( sosc_125_clk_core ),
  .q     ( sosc_125_clk_core_rst_b_pre ));

always_comb sosc_125_clk_core_rst_b = fscan_rstbypen[1] ? fscan_byprst_b[1] : sosc_125_clk_core_rst_b_pre;


//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( sbi_rst_25_core_b             ),
  .clk                 ( sosc_25_clk_core              ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( sbi_rst_25_core_b             ),
  .clk                 ( sosc_25_clk_core              ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( sbi_rst_25_core_b             ),
  .clk                 ( sosc_25_clk_core              ),
  .q                   ( force_creditreq               )
);

sbc_doublesync sync_p1_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_force_idle                 )
);

sbc_doublesync sync_p1_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_force_notidle              )
);

sbc_doublesync sync_p1_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_force_creditreq            )
);

sbc_doublesync sync_p0_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_force_idle                 )
);

sbc_doublesync sync_p0_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_force_notidle              )
);

sbc_doublesync sync_p0_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_force_creditreq            )
);

//------------------------------------------------------------------------------
//
// Asynchronous port local clock gating
//
//------------------------------------------------------------------------------
// Port 1
sbc_doublesync sync_p1_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_clkgaten                   )
);

sbc_doublesync sync_p1_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_clkgatedef                 )
);

sbc_doublesync sync_p1_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk                 ( sosc_125_clk_core             ),
  .q                   ( p1_clkgate_ovrd               )
);

always_ff @(posedge sosc_125_clk_core or negedge sosc_125_clk_core_rst_b)
  if (~sosc_125_clk_core_rst_b)
    p1_clken <= '1;
  else
    p1_clken <= ~p1_clkgate_ovrd &
      (p1_clkgatedef | ~p1_clkgaten | ~p1_cg_inprogress |
       ((xpsb_sbra_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbra_xpsb_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (xpsb_sbra_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((xpsb_sbra_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbra_xpsb_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p1_clkgate  (
  .en                  ( p1_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( sosc_125_clk_core             ),
  .enclk               ( p1_gated_clk                  )
);

// Port 0
sbc_doublesync sync_p0_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_clkgaten                   )
);

sbc_doublesync sync_p0_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_clkgatedef                 )
);

sbc_doublesync sync_p0_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( bb_cclk_rst_b ),
  .clk                 ( bb_cclk                       ),
  .q                   ( p0_clkgate_ovrd               )
);

always_ff @(posedge bb_cclk or negedge bb_cclk_rst_b)
  if (~bb_cclk_rst_b)
    p0_clken <= '1;
  else
    p0_clken <= ~p0_clkgate_ovrd &
      (p0_clkgatedef | ~p0_clkgaten | ~p0_cg_inprogress |
       ((npsb_sbra_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbra_npsb_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (npsb_sbra_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((npsb_sbra_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbra_npsb_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p0_clkgate  (
  .en                  ( p0_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( bb_cclk                       ),
  .enclk               ( p0_gated_clk                  )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_eva_present (
  .d                   ( eva_present                   ),
  .clr_b               ( sbi_rst_25_core_b             ),
  .clk                 ( sosc_25_clk_core              ),
  .q                   ( eva_present_ff2               )
);


always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          1'b1,
                          eva_present_ff2,
                          1'b1,
                          1'b1
                        };

logic p2_gated_clk;
sbc_clock_gate p2_pwr_clkgate  (
  .en ( endpoint_pwrgd[2] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p2_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p5_ism_idle | ~endpoint_pwrgd[5])
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  &  p1_efifo_idle
                  &  p0_efifo_idle;

// ISM IDLE cross into router clock domain
logic p0_ism_idle_ff2, p0_ism_idle_pre;
always_ff @(posedge bb_cclk or negedge bb_cclk_rst_b)
  if ( ~bb_cclk_rst_b)
    p0_ism_idle_pre <= '1;
  else
    p0_ism_idle_pre <= p0_ism_idle;

sbc_doublesync sync_idle_p0 (
  .d ( p0_ism_idle_pre ),
  .clr_b ( sbi_rst_25_core_b ),
  .clk   ( sosc_25_clk_core ),
  .q     ( p0_ism_idle_ff2 ));

logic p1_ism_idle_ff2, p1_ism_idle_pre;
always_ff @(posedge sosc_125_clk_core or negedge sosc_125_clk_core_rst_b)
  if ( ~sosc_125_clk_core_rst_b)
    p1_ism_idle_pre <= '1;
  else
    p1_ism_idle_pre <= p1_ism_idle;

sbc_doublesync sync_idle_p1 (
  .d ( p1_ism_idle_pre ),
  .clr_b ( sbi_rst_25_core_b ),
  .clk   ( sosc_25_clk_core ),
  .q     ( p1_ism_idle_ff2 ));

// SBR_IDLE signal for PMU
  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle_ff2 &
                  p1_ism_idle_ff2 &
                  p2_ism_idle &
                  p3_ism_idle &
                  p4_ism_idle &
                  p5_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 1'b0,
                 1'b0
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 pcirdy[1],
                 pcirdy[0]
               };
  end

always_comb
  begin
    npdstvld = { 
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 npirdy[1],
                 npirdy[0]
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_sosc_25_clk_core = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( sosc_25_clk_core              ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_sosc_25_clk_core = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0 (Asynchronous port)
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  logic p0_credit_reinit_ff2;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit_ff2 & p0_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle_ff2 & (~agent_idle[0] || ~p0_efifo_idle) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle_ff2 & agent_idle[0] & p0_efifo_idle & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle_ff2 & p0_side_clk_valid & ~p0_fab_init_idle_exit )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle_ff2 )
          p0_side_clk_valid <= '1;
      end

logic p0_side_clk_valid_ff2;
sbc_doublesync sync_p0_clk_valid (
  .d     ( p0_side_clk_valid ),
  .clr_b ( bb_cclk_rst_b ),
  .clk   ( bb_cclk ),
  .q     ( p0_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p0_credit_reinit (
  .d     ( p0_credit_reinit ),
  .set_b ( sbi_rst_25_core_b ),
  .clk   ( sosc_25_clk_core ),
  .q     ( p0_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

logic [15:0] p0_dbgbus_ing;
logic [15:0] p0_dbgbus_egr;
  always_comb
    begin
      visa_p0_tier1_bb_cclk = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_bb_cclk = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
      visa_p0_ififo_tier1_sosc_25_clk_core = { p0_dbgbus_ing[15:14],
                             p0_dbgbus_ing[5:0]};
      visa_p0_ififo_tier2_sosc_25_clk_core = { p0_dbgbus_ing[13:6] };
      visa_p0_efifo_tier1_sosc_25_clk_core = { p0_dbgbus_egr[7:0] };
      visa_p0_efifo_tier2_sosc_25_clk_core = { p0_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( bb_cclk                       ),
  .gated_side_clk      ( p0_gated_clk                  ),
  .side_rst_b ( bb_cclk_rst_b ),
  .side_clk_valid      ( p0_side_clk_valid_ff2         ),
  .side_ism_in         ( npsb_sbra_side_ism_agent      ),
  .side_ism_out        ( sbra_npsb_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( p0_agent_idle                 ),
  .port_idle           ( p0_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbra_npsb_pccup               ),
  .tnpcup              ( sbra_npsb_npcup               ),
  .tpcput              ( npsb_sbra_pcput               ),
  .tnpput              ( npsb_sbra_npput               ),
  .teom                ( npsb_sbra_eom                 ),
  .tpayload            ( npsb_sbra_payload             ),
  .pctrdy              ( p0_pctrdy                     ),
  .pcirdy              ( p0_pcirdy                     ),
  .pcdata              ( p0_pcdata                     ),
  .pceom               ( p0_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p0_nptrdy                     ),
  .npirdy              ( p0_npirdy                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( p0_npdata                     ),
  .npeom               ( p0_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( npsb_sbra_pccup               ),
  .mnpcup              ( npsb_sbra_npcup               ),
  .mpcput              ( sbra_npsb_pcput               ),
  .mnpput              ( sbra_npsb_npput               ),
  .meom                ( sbra_npsb_eom                 ),
  .mpayload            ( sbra_npsb_payload             ),
  .enpstall            ( p0_enpstall                   ),
  .epctrdy             ( p0_epctrdy                    ),
  .enptrdy             ( p0_enptrdy                    ),
  .epcirdy             ( p0_epcirdy                    ),
  .enpirdy             ( p0_enpirdy                    ),
  .data                ( p0_data                       ),
  .eom                 ( p0_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p0_clkgaten                   ),
  .force_idle          ( p0_force_idle                 ),
  .force_notidle       ( p0_force_notidle              ),
  .force_creditreq     ( p0_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress0 (
  .ing_side_clk        ( p0_gated_clk                  ),
  .ing_side_rst_b ( bb_cclk_rst_b ),
  .port_idle           ( p0_port_idle                  ),
  .pcirdy              ( p0_pcirdy                     ),
  .npirdy              ( p0_npirdy                     ),
  .npfence             ( p0_npfence                    ),
  .pceom               ( p0_pceom                      ),
  .pcdata              ( p0_pcdata                     ),
  .npeom               ( p0_npeom                      ),
  .npdata              ( p0_npdata                     ),
  .pctrdy              ( p0_pctrdy                     ),
  .nptrdy              ( p0_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p0_ififo_idle                 ),
  .egr_side_clk        ( sosc_25_clk_core              ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( sbi_rst_25_core_b             ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[0]                     ),
  .enptrdy             ( nptrdy[0]                     ),
  .epcirdy             ( pcirdy[0]                     ),
  .enpirdy             ( npirdy[0]                     ),
  .eom                 ( npeom[0]                      ),
  .data                ( npdata[0]                     ),
  .opceom              ( pceom[0]                      ),
  .opcdata             ( pcdata[0]                     ),
  .agent_idle          ( port_idle[0]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p0_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress0 (
  .ing_side_clk        ( sosc_25_clk_core              ),
  .ing_side_rst_b      ( sbi_rst_25_core_b             ),
  .port_idle           ( agent_idle[0]                 ),
  .pcirdy              ( epcirdy[0]                    ),
  .npirdy              ( enpirdy[0]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[0]                    ),
  .nptrdy              ( enptrdy[0]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p0_efifo_idle                 ),
  .egr_side_clk        ( bb_cclk                       ),
  .gated_egr_side_clk  ( p0_gated_clk                  ),
  .egr_side_rst_b ( bb_cclk_rst_b ),
  .enpstall            ( p0_enpstall                   ),
  .epctrdy             ( p0_epctrdy                    ),
  .enptrdy             ( p0_enptrdy                    ),
  .epcirdy             ( p0_epcirdy                    ),
  .enpirdy             ( p0_enpirdy                    ),
  .eom                 ( p0_eom                        ),
  .data                ( p0_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p0_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p0_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p0_agent_idle  = p0_eagent_idle & p0_ififo_idle;

// Port 1 (Asynchronous port)
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  logic p1_credit_reinit_ff2;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit_ff2 & p1_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & (~agent_idle[1] || ~p1_efifo_idle) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & agent_idle[1] & p1_efifo_idle & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle_ff2 & p1_side_clk_valid & ~p1_fab_init_idle_exit )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle_ff2 )
          p1_side_clk_valid <= '1;
      end

logic p1_side_clk_valid_ff2;
sbc_doublesync sync_p1_clk_valid (
  .d     ( p1_side_clk_valid ),
  .clr_b ( sosc_125_clk_core_rst_b ),
  .clk   ( sosc_125_clk_core ),
  .q     ( p1_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p1_credit_reinit (
  .d     ( p1_credit_reinit ),
  .set_b ( sbi_rst_25_core_b ),
  .clk   ( sosc_25_clk_core ),
  .q     ( p1_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

logic [15:0] p1_dbgbus_ing;
logic [15:0] p1_dbgbus_egr;
  always_comb
    begin
      visa_p1_tier1_sosc_125_clk_core = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_sosc_125_clk_core = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
      visa_p1_ififo_tier1_sosc_25_clk_core = { p1_dbgbus_ing[15:14],
                             p1_dbgbus_ing[5:0]};
      visa_p1_ififo_tier2_sosc_25_clk_core = { p1_dbgbus_ing[13:6] };
      visa_p1_efifo_tier1_sosc_25_clk_core = { p1_dbgbus_egr[7:0] };
      visa_p1_efifo_tier2_sosc_25_clk_core = { p1_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( sosc_125_clk_core             ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b ( sosc_125_clk_core_rst_b ),
  .side_clk_valid      ( p1_side_clk_valid_ff2         ),
  .side_ism_in         ( xpsb_sbra_side_ism_agent      ),
  .side_ism_out        ( sbra_xpsb_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( p1_agent_idle                 ),
  .port_idle           ( p1_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbra_xpsb_pccup               ),
  .tnpcup              ( sbra_xpsb_npcup               ),
  .tpcput              ( xpsb_sbra_pcput               ),
  .tnpput              ( xpsb_sbra_npput               ),
  .teom                ( xpsb_sbra_eom                 ),
  .tpayload            ( xpsb_sbra_payload             ),
  .pctrdy              ( p1_pctrdy                     ),
  .pcirdy              ( p1_pcirdy                     ),
  .pcdata              ( p1_pcdata                     ),
  .pceom               ( p1_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p1_nptrdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( p1_npdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( xpsb_sbra_pccup               ),
  .mnpcup              ( xpsb_sbra_npcup               ),
  .mpcput              ( sbra_xpsb_pcput               ),
  .mnpput              ( sbra_xpsb_npput               ),
  .meom                ( sbra_xpsb_eom                 ),
  .mpayload            ( sbra_xpsb_payload             ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .data                ( p1_data                       ),
  .eom                 ( p1_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p1_clkgaten                   ),
  .force_idle          ( p1_force_idle                 ),
  .force_notidle       ( p1_force_notidle              ),
  .force_creditreq     ( p1_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress1 (
  .ing_side_clk        ( p1_gated_clk                  ),
  .ing_side_rst_b ( sosc_125_clk_core_rst_b ),
  .port_idle           ( p1_port_idle                  ),
  .pcirdy              ( p1_pcirdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .pceom               ( p1_pceom                      ),
  .pcdata              ( p1_pcdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdata              ( p1_npdata                     ),
  .pctrdy              ( p1_pctrdy                     ),
  .nptrdy              ( p1_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p1_ififo_idle                 ),
  .egr_side_clk        ( sosc_25_clk_core              ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( sbi_rst_25_core_b             ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[1]                     ),
  .enptrdy             ( nptrdy[1]                     ),
  .epcirdy             ( pcirdy[1]                     ),
  .enpirdy             ( npirdy[1]                     ),
  .eom                 ( npeom[1]                      ),
  .data                ( npdata[1]                     ),
  .opceom              ( pceom[1]                      ),
  .opcdata             ( pcdata[1]                     ),
  .agent_idle          ( port_idle[1]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p1_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress1 (
  .ing_side_clk        ( sosc_25_clk_core              ),
  .ing_side_rst_b      ( sbi_rst_25_core_b             ),
  .port_idle           ( agent_idle[1]                 ),
  .pcirdy              ( epcirdy[1]                    ),
  .npirdy              ( enpirdy[1]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[1]                    ),
  .nptrdy              ( enptrdy[1]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p1_efifo_idle                 ),
  .egr_side_clk        ( sosc_125_clk_core             ),
  .gated_egr_side_clk  ( p1_gated_clk                  ),
  .egr_side_rst_b ( sosc_125_clk_core_rst_b ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .eom                 ( p1_eom                        ),
  .data                ( p1_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p1_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p1_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p1_agent_idle  = p1_eagent_idle & p1_ififo_idle;

// Port 2
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit & p2_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle & (~agent_idle[2] || ~p2_idle_egress) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle & agent_idle[2] & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle & p2_side_clk_valid )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle )
          p2_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

  always_comb
    begin
      visa_p2_tier1_sosc_25_clk_core = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_sosc_25_clk_core = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( sosc_25_clk_core              ),
  .gated_side_clk      ( p2_gated_clk                  ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( ccsb_sbra_side_ism_agent      ),
  .side_ism_out        ( sbra_ccsb_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .idle_egress         ( p2_idle_egress                ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbra_ccsb_pccup               ),
  .tnpcup              ( sbra_ccsb_npcup               ),
  .tpcput              ( ccsb_sbra_pcput               ),
  .tnpput              ( ccsb_sbra_npput               ),
  .teom                ( ccsb_sbra_eom                 ),
  .tpayload            ( ccsb_sbra_payload             ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( ccsb_sbra_pccup               ),
  .mnpcup              ( ccsb_sbra_npcup               ),
  .mpcput              ( sbra_ccsb_pcput               ),
  .mnpput              ( sbra_ccsb_npput               ),
  .meom                ( sbra_ccsb_eom                 ),
  .mpayload            ( sbra_ccsb_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

// Port 3
logic p3_side_clk_valid, p3_idle_egress, p3_rst_suppress;
  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p3_rst_suppress <= 1'b1;
    else
      p3_rst_suppress <= p3_credit_reinit & p3_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p3_fab_init_idle_exit <= '1;
    else
      if ( ~p3_rst_suppress & (p3_ism_idle & (~agent_idle[3] || ~p3_idle_egress) & ~p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '1;
      else if ( ~p3_rst_suppress & (p3_ism_idle & agent_idle[3] & p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( p3_ism_idle & p3_side_clk_valid )
          p3_side_clk_valid <= '0;
        else if ( (p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack) || ~p3_ism_idle )
          p3_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

  always_comb
    begin
      visa_p3_tier1_sosc_25_clk_core = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_sosc_25_clk_core = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( sosc_25_clk_core              ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( io_pxp_sbra_side_ism_agent    ),
  .side_ism_out        ( sbra_io_pxp_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .idle_egress         ( p3_idle_egress                ),
  .ism_idle            ( p3_ism_idle                   ),
  .credit_reinit       ( p3_credit_reinit              ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbra_io_pxp_pccup             ),
  .tnpcup              ( sbra_io_pxp_npcup             ),
  .tpcput              ( io_pxp_sbra_pcput             ),
  .tnpput              ( io_pxp_sbra_npput             ),
  .teom                ( io_pxp_sbra_eom               ),
  .tpayload            ( io_pxp_sbra_payload           ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( io_pxp_sbra_pccup             ),
  .mnpcup              ( io_pxp_sbra_npcup             ),
  .mpcput              ( sbra_io_pxp_pcput             ),
  .mnpput              ( sbra_io_pxp_npput             ),
  .meom                ( sbra_io_pxp_eom               ),
  .mpayload            ( sbra_io_pxp_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
logic p4_side_clk_valid, p4_idle_egress, p4_rst_suppress;
  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p4_rst_suppress <= 1'b1;
    else
      p4_rst_suppress <= p4_credit_reinit & p4_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p4_fab_init_idle_exit <= '1;
    else
      if ( ~p4_rst_suppress & (p4_ism_idle & (~agent_idle[4] || ~p4_idle_egress) & ~p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '1;
      else if ( ~p4_rst_suppress & (p4_ism_idle & agent_idle[4] & p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( p4_ism_idle & p4_side_clk_valid )
          p4_side_clk_valid <= '0;
        else if ( (p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack) || ~p4_ism_idle )
          p4_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

  always_comb
    begin
      visa_p4_tier1_sosc_25_clk_core = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_sosc_25_clk_core = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( sosc_25_clk_core              ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( io_dmi_sbra_side_ism_agent    ),
  .side_ism_out        ( sbra_io_dmi_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .idle_egress         ( p4_idle_egress                ),
  .ism_idle            ( p4_ism_idle                   ),
  .credit_reinit       ( p4_credit_reinit              ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbra_io_dmi_pccup             ),
  .tnpcup              ( sbra_io_dmi_npcup             ),
  .tpcput              ( io_dmi_sbra_pcput             ),
  .tnpput              ( io_dmi_sbra_npput             ),
  .teom                ( io_dmi_sbra_eom               ),
  .tpayload            ( io_dmi_sbra_payload           ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( io_dmi_sbra_pccup             ),
  .mnpcup              ( io_dmi_sbra_npcup             ),
  .mpcput              ( sbra_io_dmi_pcput             ),
  .mnpput              ( sbra_io_dmi_npput             ),
  .meom                ( sbra_io_dmi_eom               ),
  .mpayload            ( sbra_io_dmi_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

// Port 5
logic p5_side_clk_valid, p5_idle_egress, p5_rst_suppress;
  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p5_rst_suppress <= 1'b1;
    else
      p5_rst_suppress <= p5_credit_reinit & p5_rst_suppress;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if (~sbi_rst_25_core_b)
      p5_fab_init_idle_exit <= '1;
    else
      if ( ~p5_rst_suppress & (p5_ism_idle & (~agent_idle[5] || ~p5_idle_egress) & ~p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '1;
      else if ( ~p5_rst_suppress & (p5_ism_idle & agent_idle[5] & p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '0;

  always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)
    if ( ~sbi_rst_25_core_b )
      p5_side_clk_valid <= 1'b0;
    else
      begin
        if ( p5_ism_idle & p5_side_clk_valid )
          p5_side_clk_valid <= '0;
        else if ( (p5_fab_init_idle_exit & p5_fab_init_idle_exit_ack) || ~p5_ism_idle )
          p5_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p5_dbgbus;

  always_comb
    begin
      visa_p5_tier1_sosc_25_clk_core = { p5_dbgbus[31],
                            p5_dbgbus[27:24],
                            p5_dbgbus[21:19],
                            p5_dbgbus[15:12],
                            p5_dbgbus[7:4] };
      visa_p5_tier2_sosc_25_clk_core = { p5_dbgbus[30:28],
                            p5_dbgbus[23:22],
                            p5_dbgbus[18:16],
                            p5_dbgbus[11:8],
                            p5_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  1                            ),
  .PCQUEUEDEPTH        (  1                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport5 (
  .side_clk            ( sosc_25_clk_core              ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( sbi_rst_25_core_b             ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( io_st_sbra_side_ism_agent     ),
  .side_ism_out        ( sbra_io_st_side_ism_fabric    ),
  .int_pok             ( endpoint_pwrgd[5] ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .idle_egress         ( p5_idle_egress                ),
  .ism_idle            ( p5_ism_idle                   ),
  .credit_reinit       ( p5_credit_reinit              ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbra_io_st_pccup              ),
  .tnpcup              ( sbra_io_st_npcup              ),
  .tpcput              ( io_st_sbra_pcput              ),
  .tnpput              ( io_st_sbra_npput              ),
  .teom                ( io_st_sbra_eom                ),
  .tpayload            ( io_st_sbra_payload            ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( io_st_sbra_pccup              ),
  .mnpcup              ( io_st_sbra_npcup              ),
  .mpcput              ( sbra_io_st_pcput              ),
  .mnpput              ( sbra_io_st_npput              ),
  .meom                ( sbra_io_st_eom                ),
  .mpayload            ( sbra_io_st_payload            ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p5_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbra_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbra_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge sosc_25_clk_core or negedge sbi_rst_25_core_b)

      if (~sbi_rst_25_core_b) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge sosc_25_clk_core) disable iff (sbi_rst_25_core_b !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge sosc_25_clk_core) disable iff (sbi_rst_25_core_b !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 0, bb_cclk, bb_rst_b, 0, , 4ns
ClockReset, 3, iosf_fust_side_clk, iosf_fust_side_rst_b, 0, , 2ns
ClockReset, 4, iosf_idf_side_clk, iosf_idf_side_rst_b, 0, cgc0, 2ns
ClockReset, 5, iosf_swf_side_clk, iosf_swf_side_rst_b, 0, cgc1, 2ns
ClockReset, 1, sosc_125_clk_core, sbi_rst_125_core_b, 0, , 4ns
ClockReset, 2, sosc_25_clk_core, sbi_rst_25_core_b, 0, , 40ns
SyncRouter, ccsb, ccsb,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 2, sbra, sbr1, , , , , , , , , , , , , , , 
RouterAgentPort, ccsb, 0
RouterAgentPort, ccsb, 1
Endpoint, dfxa,1, 1, 4, 0, 3, 3, 1, 2, 3, 3, 
Endpoint, fust,1, 1, 3, 0, 3, 3, 1, 0, 3, 3, 
Endpoint, idf,1, 1, 4, 0, 3, 3, 1, 5, 3, 3, 
Endpoint, io_dmi,0, 1, 2, 0, 1, 1, 1, 235, 3, 3, 
Endpoint, io_pxp,0, 1, 2, 0, 1, 1, 1, 236, 3, 3, 
Endpoint, io_st,0, 1, 2, 0, 1, 1, 1, 234, 3, 3, 
Endpoint, isa,1, 1, 4, 0, 3, 3, 1, 1, 3, 3, 
Endpoint, npsb,0, 1, 0, 0, 1, 1, 1, 239, 3, 3, 
Endpoint, rsp,1, 1, 4, 0, 3, 3, 1, 6, 3, 3, 
SyncRouter, sbr1, sbr1,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 9, ccsb, fust, sbr2, isa, dfxa, scu0, scu1, idf, rsp, , , , , , , , 
RouterAgentPort, sbr1, 2
SyncRouter, sbr2, sbr2,2, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 5, 3, sbr1, xut, swf, , , , , , , , , , , , , , 
SyncRouter, sbra, sbra,0, 0, 0, 1, 4, 1, 0, 1, noa, dfxa, 2, 6, npsb, xpsb, ccsb, io_pxp, io_dmi, io_st, , , , , , , , , , , 
Endpoint, scu0,1, 1, 4, 0, 3, 3, 1, 3, 3, 3, 
Endpoint, scu1,3, 1, 4, 0, 3, 3, 1, 4, 3, 3, 
Endpoint, swf,2, 1, 5, 0, 3, 3, 1, 9, 3, 3, 
Endpoint, xpsb,0, 1, 1, 0, 1, 1, 1, 238, 3, 3, 
Endpoint, xut,2, 1, 5, 0, 3, 3, 1, 8, 3, 3, 
AsyncPort, ccsb, 0, 4, 4, 0, 
AsyncPort, sbr1, 1, 4, 4, 0, 
AsyncPort, sbr1, 2, 4, 4, 0, 
AsyncPort, sbra, 0, 2, 2, 0, 
AsyncPort, sbra, 1, 2, 2, 0, 
PowerWell, 0, 
PowerWell, 1, eva_present
PowerWell, 2, crp_sbr1_xu_en
PowerWell, 3, crp_sbr1_scu1_en
*/
//------------------------------------------------------------------------------
