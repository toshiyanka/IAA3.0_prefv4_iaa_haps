module ctech_lib_msff_meta (
   input logic clk,
   input logic d, 
   output logic o
);
   d04hgn20ld0b0 ctech_lib_dcszo (.o(o), .d(d), .clk(clk));
endmodule
