parameter NUMBER_OF_HIER  = 0;
parameter NUMBER_OF_STAPS = 0;
