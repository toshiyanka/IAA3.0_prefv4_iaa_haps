VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf192b080e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf192b080e1r1w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 34.2 BY 41.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 21.48 18.128 22.68 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 19.56 15.128 20.76 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 21.48 13.628 22.68 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 21.48 13.716 22.68 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 21.48 13.972 22.68 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 21.48 14.228 22.68 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 21.48 14.316 22.68 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 21.48 14.528 22.68 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 21.48 15.128 22.68 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 21.48 18.216 22.68 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 21.48 18.472 22.68 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 21.48 18.728 22.68 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 21.48 19.116 22.68 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 19.56 16.416 20.76 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 19.56 16.672 20.76 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 19.56 16.928 20.76 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 19.56 17.016 20.76 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 19.56 17.228 20.76 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.784 19.56 17.828 20.76 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 19.56 17.916 20.76 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 19.56 15.216 20.76 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 19.56 15.772 20.76 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 0.24 15.772 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 23.28 15.772 24.48 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 23.28 16.028 24.48 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 23.28 17.316 24.48 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 23.28 17.572 24.48 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 24 16.416 25.2 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 24 15.428 25.2 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 24 16.928 25.2 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 24 17.016 25.2 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 24.72 15.772 25.92 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 24.72 16.028 25.92 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 1.68 17.316 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 24.72 17.572 25.92 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 24.72 16.672 25.92 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 25.44 15.428 26.64 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 25.44 15.516 26.64 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 25.44 17.228 26.64 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 25.44 17.316 26.64 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 26.16 16.116 27.36 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 26.16 16.328 27.36 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 26.16 16.672 27.36 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 26.16 16.928 27.36 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 1.68 17.572 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 26.88 15.428 28.08 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 26.88 15.516 28.08 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 26.88 17.316 28.08 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 26.88 17.572 28.08 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 27.6 16.116 28.8 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 27.6 16.328 28.8 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 27.6 16.672 28.8 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 27.6 16.928 28.8 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 28.32 15.428 29.52 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 28.32 15.516 29.52 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 2.4 16.116 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 28.32 17.316 29.52 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 28.32 17.572 29.52 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 29.04 16.116 30.24 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 29.04 16.328 30.24 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 29.04 16.672 30.24 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 29.04 16.928 30.24 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 29.76 15.428 30.96 ;
    END
  END wrdatap0[136]
  PIN wrdatap0[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 29.76 15.516 30.96 ;
    END
  END wrdatap0[137]
  PIN wrdatap0[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 29.76 17.316 30.96 ;
    END
  END wrdatap0[138]
  PIN wrdatap0[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 29.76 17.572 30.96 ;
    END
  END wrdatap0[139]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 2.4 16.328 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 30.48 16.116 31.68 ;
    END
  END wrdatap0[140]
  PIN wrdatap0[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 30.48 16.328 31.68 ;
    END
  END wrdatap0[141]
  PIN wrdatap0[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 30.48 16.672 31.68 ;
    END
  END wrdatap0[142]
  PIN wrdatap0[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 30.48 16.928 31.68 ;
    END
  END wrdatap0[143]
  PIN wrdatap0[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 31.2 15.428 32.4 ;
    END
  END wrdatap0[144]
  PIN wrdatap0[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 31.2 15.516 32.4 ;
    END
  END wrdatap0[145]
  PIN wrdatap0[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 31.2 17.316 32.4 ;
    END
  END wrdatap0[146]
  PIN wrdatap0[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 31.2 17.572 32.4 ;
    END
  END wrdatap0[147]
  PIN wrdatap0[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 31.92 16.116 33.12 ;
    END
  END wrdatap0[148]
  PIN wrdatap0[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 31.92 16.328 33.12 ;
    END
  END wrdatap0[149]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 2.4 16.672 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 31.92 16.672 33.12 ;
    END
  END wrdatap0[150]
  PIN wrdatap0[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 31.92 16.928 33.12 ;
    END
  END wrdatap0[151]
  PIN wrdatap0[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 32.64 15.428 33.84 ;
    END
  END wrdatap0[152]
  PIN wrdatap0[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 32.64 15.516 33.84 ;
    END
  END wrdatap0[153]
  PIN wrdatap0[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 32.64 17.316 33.84 ;
    END
  END wrdatap0[154]
  PIN wrdatap0[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 32.64 17.572 33.84 ;
    END
  END wrdatap0[155]
  PIN wrdatap0[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 33.36 16.116 34.56 ;
    END
  END wrdatap0[156]
  PIN wrdatap0[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 33.36 16.328 34.56 ;
    END
  END wrdatap0[157]
  PIN wrdatap0[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 33.36 16.672 34.56 ;
    END
  END wrdatap0[158]
  PIN wrdatap0[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 33.36 16.928 34.56 ;
    END
  END wrdatap0[159]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 2.4 16.928 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 34.08 15.428 35.28 ;
    END
  END wrdatap0[160]
  PIN wrdatap0[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 34.08 15.516 35.28 ;
    END
  END wrdatap0[161]
  PIN wrdatap0[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 34.08 17.316 35.28 ;
    END
  END wrdatap0[162]
  PIN wrdatap0[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 34.08 17.572 35.28 ;
    END
  END wrdatap0[163]
  PIN wrdatap0[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 34.8 16.116 36 ;
    END
  END wrdatap0[164]
  PIN wrdatap0[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 34.8 16.328 36 ;
    END
  END wrdatap0[165]
  PIN wrdatap0[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 34.8 16.672 36 ;
    END
  END wrdatap0[166]
  PIN wrdatap0[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 34.8 16.928 36 ;
    END
  END wrdatap0[167]
  PIN wrdatap0[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 35.52 15.428 36.72 ;
    END
  END wrdatap0[168]
  PIN wrdatap0[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 35.52 15.516 36.72 ;
    END
  END wrdatap0[169]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 3.12 15.428 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 35.52 17.316 36.72 ;
    END
  END wrdatap0[170]
  PIN wrdatap0[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 35.52 17.572 36.72 ;
    END
  END wrdatap0[171]
  PIN wrdatap0[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 36.24 16.116 37.44 ;
    END
  END wrdatap0[172]
  PIN wrdatap0[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 36.24 16.328 37.44 ;
    END
  END wrdatap0[173]
  PIN wrdatap0[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 36.24 16.672 37.44 ;
    END
  END wrdatap0[174]
  PIN wrdatap0[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 36.24 16.928 37.44 ;
    END
  END wrdatap0[175]
  PIN wrdatap0[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 36.96 15.428 38.16 ;
    END
  END wrdatap0[176]
  PIN wrdatap0[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 36.96 15.516 38.16 ;
    END
  END wrdatap0[177]
  PIN wrdatap0[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 36.96 17.316 38.16 ;
    END
  END wrdatap0[178]
  PIN wrdatap0[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 36.96 17.572 38.16 ;
    END
  END wrdatap0[179]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 3.12 15.516 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 37.68 16.116 38.88 ;
    END
  END wrdatap0[180]
  PIN wrdatap0[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 37.68 16.328 38.88 ;
    END
  END wrdatap0[181]
  PIN wrdatap0[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 37.68 16.672 38.88 ;
    END
  END wrdatap0[182]
  PIN wrdatap0[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 37.68 16.928 38.88 ;
    END
  END wrdatap0[183]
  PIN wrdatap0[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 38.4 15.428 39.6 ;
    END
  END wrdatap0[184]
  PIN wrdatap0[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 38.4 15.516 39.6 ;
    END
  END wrdatap0[185]
  PIN wrdatap0[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 38.4 17.316 39.6 ;
    END
  END wrdatap0[186]
  PIN wrdatap0[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 38.4 17.572 39.6 ;
    END
  END wrdatap0[187]
  PIN wrdatap0[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 39.12 16.116 40.32 ;
    END
  END wrdatap0[188]
  PIN wrdatap0[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 39.12 16.328 40.32 ;
    END
  END wrdatap0[189]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 3.12 17.316 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 39.12 16.672 40.32 ;
    END
  END wrdatap0[190]
  PIN wrdatap0[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 39.12 16.928 40.32 ;
    END
  END wrdatap0[191]
  PIN wrdatap0[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 39.84 15.428 41.04 ;
    END
  END wrdatap0[192]
  PIN wrdatap0[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 39.84 15.516 41.04 ;
    END
  END wrdatap0[193]
  PIN wrdatap0[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 39.84 17.316 41.04 ;
    END
  END wrdatap0[194]
  PIN wrdatap0[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 39.84 17.572 41.04 ;
    END
  END wrdatap0[195]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 3.12 17.572 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 0.24 16.028 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 3.84 16.116 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 3.84 16.328 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 3.84 16.672 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 3.84 16.928 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.56 15.428 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 4.56 15.516 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 4.56 17.316 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 4.56 17.572 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 5.28 16.116 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 5.28 16.328 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 0.24 17.316 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 5.28 16.672 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 5.28 16.928 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6 15.428 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 6 15.516 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 6 17.316 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 6 17.572 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 6.72 16.116 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 6.72 16.328 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 6.72 16.672 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 6.72 16.928 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 0.24 17.572 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 7.44 15.428 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 7.44 15.516 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 7.44 17.316 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 7.44 17.572 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 8.16 16.116 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 8.16 16.328 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 8.16 16.672 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 8.16 16.928 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.88 15.428 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 8.88 15.516 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 0.96 16.116 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 8.88 17.316 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 8.88 17.572 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 9.6 16.116 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 9.6 16.328 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 9.6 16.672 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 9.6 16.928 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 10.32 15.428 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 10.32 15.516 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 10.32 17.316 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 10.32 17.572 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 0.96 16.328 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 11.04 16.116 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 11.04 16.328 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 11.04 16.672 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 11.04 16.928 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 11.76 15.428 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 11.76 15.516 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 11.76 17.316 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 11.76 17.572 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 12.48 16.116 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 12.48 16.328 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 0.96 16.672 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 12.48 16.672 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 12.48 16.928 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 13.2 15.428 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 13.2 15.516 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 13.2 17.316 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 13.2 17.572 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 13.92 16.116 15.12 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 13.92 16.328 15.12 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 13.92 16.672 15.12 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 13.92 16.928 15.12 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 0.96 16.928 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 14.64 15.428 15.84 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 14.64 15.516 15.84 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 14.64 17.316 15.84 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 14.64 17.572 15.84 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 15.36 16.116 16.56 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 15.36 16.328 16.56 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 15.36 16.672 16.56 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 15.36 16.928 16.56 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 16.08 15.428 17.28 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 16.08 15.516 17.28 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 1.68 15.428 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 16.08 17.316 17.28 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 16.08 17.572 17.28 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 16.8 16.116 18 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 16.8 16.328 18 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 16.8 16.672 18 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 16.8 16.928 18 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 17.52 15.428 18.72 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 17.52 15.516 18.72 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 17.52 17.316 18.72 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 17.52 17.572 18.72 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 1.68 15.516 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 19.56 16.116 20.76 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 19.56 16.328 20.76 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 19.56 16.028 20.76 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 0.24 13.628 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.28 14.616 24.48 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 23.28 14.872 24.48 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.784 23.28 17.828 24.48 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 23.28 17.916 24.48 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 24 13.972 25.2 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 24 14.228 25.2 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 24 18.728 25.2 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 24 18.816 25.2 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 24.72 14.872 25.92 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 24.72 13.628 25.92 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 1.68 18.816 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 24.72 17.916 25.92 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 24.72 18.128 25.92 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 25.44 14.316 26.64 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 25.44 14.528 26.64 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 25.44 18.816 26.64 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 25.44 19.028 26.64 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 26.16 13.628 27.36 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 26.16 13.716 27.36 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 26.16 18.128 27.36 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 26.16 18.216 27.36 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 1.68 19.028 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 26.88 14.616 28.08 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 26.88 14.872 28.08 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.88 18.816 28.08 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.88 19.028 28.08 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 27.6 13.628 28.8 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 27.6 13.716 28.8 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 27.6 18.128 28.8 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 27.6 18.216 28.8 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 28.32 14.616 29.52 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 28.32 14.872 29.52 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 2.4 13.628 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 28.32 18.816 29.52 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 28.32 19.028 29.52 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 29.04 13.628 30.24 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 29.04 13.716 30.24 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 29.04 18.128 30.24 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 29.04 18.216 30.24 ;
    END
  END rddatap0[135]
  PIN rddatap0[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 29.76 14.616 30.96 ;
    END
  END rddatap0[136]
  PIN rddatap0[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 29.76 14.872 30.96 ;
    END
  END rddatap0[137]
  PIN rddatap0[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 29.76 18.816 30.96 ;
    END
  END rddatap0[138]
  PIN rddatap0[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 29.76 19.028 30.96 ;
    END
  END rddatap0[139]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 2.4 13.716 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 30.48 13.628 31.68 ;
    END
  END rddatap0[140]
  PIN rddatap0[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 30.48 13.716 31.68 ;
    END
  END rddatap0[141]
  PIN rddatap0[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 30.48 18.128 31.68 ;
    END
  END rddatap0[142]
  PIN rddatap0[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 30.48 18.216 31.68 ;
    END
  END rddatap0[143]
  PIN rddatap0[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 31.2 14.616 32.4 ;
    END
  END rddatap0[144]
  PIN rddatap0[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 31.2 14.872 32.4 ;
    END
  END rddatap0[145]
  PIN rddatap0[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 31.2 18.816 32.4 ;
    END
  END rddatap0[146]
  PIN rddatap0[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 31.2 19.028 32.4 ;
    END
  END rddatap0[147]
  PIN rddatap0[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 31.92 13.628 33.12 ;
    END
  END rddatap0[148]
  PIN rddatap0[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 31.92 13.716 33.12 ;
    END
  END rddatap0[149]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 2.4 18.128 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 31.92 18.128 33.12 ;
    END
  END rddatap0[150]
  PIN rddatap0[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 31.92 18.216 33.12 ;
    END
  END rddatap0[151]
  PIN rddatap0[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 32.64 14.616 33.84 ;
    END
  END rddatap0[152]
  PIN rddatap0[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 32.64 14.872 33.84 ;
    END
  END rddatap0[153]
  PIN rddatap0[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 32.64 18.816 33.84 ;
    END
  END rddatap0[154]
  PIN rddatap0[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 32.64 19.028 33.84 ;
    END
  END rddatap0[155]
  PIN rddatap0[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 33.36 13.628 34.56 ;
    END
  END rddatap0[156]
  PIN rddatap0[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 33.36 13.716 34.56 ;
    END
  END rddatap0[157]
  PIN rddatap0[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 33.36 18.128 34.56 ;
    END
  END rddatap0[158]
  PIN rddatap0[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 33.36 18.216 34.56 ;
    END
  END rddatap0[159]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 2.4 18.216 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 34.08 14.616 35.28 ;
    END
  END rddatap0[160]
  PIN rddatap0[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 34.08 14.872 35.28 ;
    END
  END rddatap0[161]
  PIN rddatap0[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 34.08 18.816 35.28 ;
    END
  END rddatap0[162]
  PIN rddatap0[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 34.08 19.028 35.28 ;
    END
  END rddatap0[163]
  PIN rddatap0[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 34.8 13.628 36 ;
    END
  END rddatap0[164]
  PIN rddatap0[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 34.8 13.716 36 ;
    END
  END rddatap0[165]
  PIN rddatap0[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 34.8 18.128 36 ;
    END
  END rddatap0[166]
  PIN rddatap0[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 34.8 18.216 36 ;
    END
  END rddatap0[167]
  PIN rddatap0[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 35.52 14.616 36.72 ;
    END
  END rddatap0[168]
  PIN rddatap0[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 35.52 14.872 36.72 ;
    END
  END rddatap0[169]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.12 14.616 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 35.52 18.816 36.72 ;
    END
  END rddatap0[170]
  PIN rddatap0[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 35.52 19.028 36.72 ;
    END
  END rddatap0[171]
  PIN rddatap0[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 36.24 13.628 37.44 ;
    END
  END rddatap0[172]
  PIN rddatap0[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 36.24 13.716 37.44 ;
    END
  END rddatap0[173]
  PIN rddatap0[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 36.24 18.128 37.44 ;
    END
  END rddatap0[174]
  PIN rddatap0[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 36.24 18.216 37.44 ;
    END
  END rddatap0[175]
  PIN rddatap0[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 36.96 14.616 38.16 ;
    END
  END rddatap0[176]
  PIN rddatap0[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 36.96 14.872 38.16 ;
    END
  END rddatap0[177]
  PIN rddatap0[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 36.96 18.816 38.16 ;
    END
  END rddatap0[178]
  PIN rddatap0[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 36.96 19.028 38.16 ;
    END
  END rddatap0[179]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 3.12 14.872 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 37.68 13.628 38.88 ;
    END
  END rddatap0[180]
  PIN rddatap0[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 37.68 13.716 38.88 ;
    END
  END rddatap0[181]
  PIN rddatap0[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 37.68 18.128 38.88 ;
    END
  END rddatap0[182]
  PIN rddatap0[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 37.68 18.216 38.88 ;
    END
  END rddatap0[183]
  PIN rddatap0[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 38.4 14.616 39.6 ;
    END
  END rddatap0[184]
  PIN rddatap0[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 38.4 14.872 39.6 ;
    END
  END rddatap0[185]
  PIN rddatap0[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 38.4 18.816 39.6 ;
    END
  END rddatap0[186]
  PIN rddatap0[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 38.4 19.028 39.6 ;
    END
  END rddatap0[187]
  PIN rddatap0[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 39.12 13.628 40.32 ;
    END
  END rddatap0[188]
  PIN rddatap0[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 39.12 13.716 40.32 ;
    END
  END rddatap0[189]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 3.12 18.816 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 39.12 18.128 40.32 ;
    END
  END rddatap0[190]
  PIN rddatap0[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 39.12 18.216 40.32 ;
    END
  END rddatap0[191]
  PIN rddatap0[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 39.84 14.616 41.04 ;
    END
  END rddatap0[192]
  PIN rddatap0[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 39.84 14.872 41.04 ;
    END
  END rddatap0[193]
  PIN rddatap0[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 39.84 18.816 41.04 ;
    END
  END rddatap0[194]
  PIN rddatap0[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 39.84 19.028 41.04 ;
    END
  END rddatap0[195]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 3.12 19.028 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.24 13.716 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 3.84 13.628 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.84 13.716 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 3.84 18.128 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 3.84 18.216 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 4.56 14.616 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 4.56 14.872 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 4.56 18.816 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 4.56 19.028 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 5.28 13.628 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 5.28 13.716 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 5.28 18.128 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 5.28 18.216 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6 14.616 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 6 14.872 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 6 18.816 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 6 19.028 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 6.72 13.628 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 6.72 13.716 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 6.72 18.128 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 6.72 18.216 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 7.44 14.616 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 7.44 14.872 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 7.44 18.816 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 7.44 19.028 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 8.16 13.628 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 8.16 13.716 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 8.16 18.128 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 8.16 18.216 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.88 14.616 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 8.88 14.872 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.96 13.972 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.88 18.816 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.88 19.028 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 9.6 13.628 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 9.6 13.716 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 9.6 18.128 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 9.6 18.216 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 10.32 14.616 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 10.32 14.872 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 10.32 18.816 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 10.32 19.028 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 0.96 14.228 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.04 13.628 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 11.04 13.716 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 11.04 18.128 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 11.04 18.216 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 11.76 14.616 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 11.76 14.872 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 11.76 18.816 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 11.76 19.028 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 12.48 13.628 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 12.48 13.716 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 0.96 18.128 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 12.48 18.128 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 12.48 18.216 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 13.2 14.616 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 13.2 14.872 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 13.2 18.816 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 13.2 19.028 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 13.92 13.628 15.12 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 13.92 13.716 15.12 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 13.92 18.128 15.12 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 13.92 18.216 15.12 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 0.96 18.216 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 14.64 14.616 15.84 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 14.64 14.872 15.84 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 14.64 18.816 15.84 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 14.64 19.028 15.84 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 15.36 13.628 16.56 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 15.36 13.716 16.56 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 15.36 18.128 16.56 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 15.36 18.216 16.56 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 16.08 14.616 17.28 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 16.08 14.872 17.28 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 1.68 14.616 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 16.08 18.816 17.28 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 16.08 19.028 17.28 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 16.8 13.628 18 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 16.8 13.716 18 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 16.8 18.128 18 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 16.8 18.216 18 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 17.52 14.616 18.72 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 17.52 14.872 18.72 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 17.52 18.816 18.72 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 17.52 19.028 18.72 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 1.68 14.872 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 41.22 ;
        RECT 2.662 0.06 2.738 41.22 ;
        RECT 4.462 0.06 4.538 41.22 ;
        RECT 6.262 0.06 6.338 41.22 ;
        RECT 8.062 0.06 8.138 41.22 ;
        RECT 9.862 0.06 9.938 41.22 ;
        RECT 11.662 0.06 11.738 41.22 ;
        RECT 13.462 0.06 13.538 41.22 ;
        RECT 15.262 0.06 15.338 41.22 ;
        RECT 17.062 0.06 17.138 41.22 ;
        RECT 18.862 0.06 18.938 41.22 ;
        RECT 20.662 0.06 20.738 41.22 ;
        RECT 22.462 0.06 22.538 41.22 ;
        RECT 24.262 0.06 24.338 41.22 ;
        RECT 26.062 0.06 26.138 41.22 ;
        RECT 27.862 0.06 27.938 41.22 ;
        RECT 29.662 0.06 29.738 41.22 ;
        RECT 31.462 0.06 31.538 41.22 ;
        RECT 33.262 0.06 33.338 41.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 41.22 ;
        RECT 3.562 0.06 3.638 41.22 ;
        RECT 5.362 0.06 5.438 41.22 ;
        RECT 7.162 0.06 7.238 41.22 ;
        RECT 8.962 0.06 9.038 41.22 ;
        RECT 10.762 0.06 10.838 41.22 ;
        RECT 12.562 0.06 12.638 41.22 ;
        RECT 14.362 0.06 14.438 41.22 ;
        RECT 16.162 0.06 16.238 41.22 ;
        RECT 17.962 0.06 18.038 41.22 ;
        RECT 19.762 0.06 19.838 41.22 ;
        RECT 21.562 0.06 21.638 41.22 ;
        RECT 23.362 0.06 23.438 41.22 ;
        RECT 25.162 0.06 25.238 41.22 ;
        RECT 26.962 0.06 27.038 41.22 ;
        RECT 28.762 0.06 28.838 41.22 ;
        RECT 30.562 0.06 30.638 41.22 ;
        RECT 32.362 0.06 32.438 41.22 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 34.216 41.294 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 34.22 41.3 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 34.2705 41.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 34.235 41.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 34.27 41.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 34.259 41.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 34.29 41.342 ;
    LAYER m7 SPACING 0 ;
      RECT 33.338 41.34 34.24 41.4 ;
      RECT 33.338 -0.06 34.292 41.34 ;
      RECT 33.338 -0.12 34.24 -0.06 ;
      RECT 32.438 -0.12 33.262 41.4 ;
      RECT 31.538 -0.12 32.362 41.4 ;
      RECT 30.638 -0.12 31.462 41.4 ;
      RECT 29.738 -0.12 30.562 41.4 ;
      RECT 28.838 -0.12 29.662 41.4 ;
      RECT 27.938 -0.12 28.762 41.4 ;
      RECT 27.038 -0.12 27.862 41.4 ;
      RECT 26.138 -0.12 26.962 41.4 ;
      RECT 25.238 -0.12 26.062 41.4 ;
      RECT 24.338 -0.12 25.162 41.4 ;
      RECT 23.438 -0.12 24.262 41.4 ;
      RECT 22.538 -0.12 23.362 41.4 ;
      RECT 21.638 -0.12 22.462 41.4 ;
      RECT 20.738 -0.12 21.562 41.4 ;
      RECT 19.838 -0.12 20.662 41.4 ;
      RECT 18.938 41.04 19.762 41.4 ;
      RECT 18.938 39.84 18.984 41.04 ;
      RECT 19.028 39.84 19.762 41.04 ;
      RECT 18.938 39.6 19.762 39.84 ;
      RECT 18.938 38.4 18.984 39.6 ;
      RECT 19.028 38.4 19.762 39.6 ;
      RECT 18.938 38.16 19.762 38.4 ;
      RECT 18.938 36.96 18.984 38.16 ;
      RECT 19.028 36.96 19.762 38.16 ;
      RECT 18.938 36.72 19.762 36.96 ;
      RECT 18.938 35.52 18.984 36.72 ;
      RECT 19.028 35.52 19.762 36.72 ;
      RECT 18.938 35.28 19.762 35.52 ;
      RECT 18.938 34.08 18.984 35.28 ;
      RECT 19.028 34.08 19.762 35.28 ;
      RECT 18.938 33.84 19.762 34.08 ;
      RECT 18.938 32.64 18.984 33.84 ;
      RECT 19.028 32.64 19.762 33.84 ;
      RECT 18.938 32.4 19.762 32.64 ;
      RECT 18.938 31.2 18.984 32.4 ;
      RECT 19.028 31.2 19.762 32.4 ;
      RECT 18.938 30.96 19.762 31.2 ;
      RECT 18.938 29.76 18.984 30.96 ;
      RECT 19.028 29.76 19.762 30.96 ;
      RECT 18.938 29.52 19.762 29.76 ;
      RECT 18.938 28.32 18.984 29.52 ;
      RECT 19.028 28.32 19.762 29.52 ;
      RECT 18.938 28.08 19.762 28.32 ;
      RECT 18.938 26.88 18.984 28.08 ;
      RECT 19.028 26.88 19.762 28.08 ;
      RECT 18.938 26.64 19.762 26.88 ;
      RECT 18.938 25.44 18.984 26.64 ;
      RECT 19.028 25.44 19.762 26.64 ;
      RECT 18.938 22.68 19.762 25.44 ;
      RECT 18.938 21.48 19.072 22.68 ;
      RECT 19.116 21.48 19.762 22.68 ;
      RECT 18.938 18.72 19.762 21.48 ;
      RECT 18.938 17.52 18.984 18.72 ;
      RECT 19.028 17.52 19.762 18.72 ;
      RECT 18.938 17.28 19.762 17.52 ;
      RECT 18.938 16.08 18.984 17.28 ;
      RECT 19.028 16.08 19.762 17.28 ;
      RECT 18.938 15.84 19.762 16.08 ;
      RECT 18.938 14.64 18.984 15.84 ;
      RECT 19.028 14.64 19.762 15.84 ;
      RECT 18.938 14.4 19.762 14.64 ;
      RECT 18.938 13.2 18.984 14.4 ;
      RECT 19.028 13.2 19.762 14.4 ;
      RECT 18.938 12.96 19.762 13.2 ;
      RECT 18.938 11.76 18.984 12.96 ;
      RECT 19.028 11.76 19.762 12.96 ;
      RECT 18.938 11.52 19.762 11.76 ;
      RECT 18.938 10.32 18.984 11.52 ;
      RECT 19.028 10.32 19.762 11.52 ;
      RECT 18.938 10.08 19.762 10.32 ;
      RECT 18.938 8.88 18.984 10.08 ;
      RECT 19.028 8.88 19.762 10.08 ;
      RECT 18.938 8.64 19.762 8.88 ;
      RECT 18.938 7.44 18.984 8.64 ;
      RECT 19.028 7.44 19.762 8.64 ;
      RECT 18.938 7.2 19.762 7.44 ;
      RECT 18.938 6 18.984 7.2 ;
      RECT 19.028 6 19.762 7.2 ;
      RECT 18.938 5.76 19.762 6 ;
      RECT 18.938 4.56 18.984 5.76 ;
      RECT 19.028 4.56 19.762 5.76 ;
      RECT 18.938 4.32 19.762 4.56 ;
      RECT 18.938 3.12 18.984 4.32 ;
      RECT 19.028 3.12 19.762 4.32 ;
      RECT 18.938 2.88 19.762 3.12 ;
      RECT 18.938 1.68 18.984 2.88 ;
      RECT 19.028 1.68 19.762 2.88 ;
      RECT 18.938 1.44 19.762 1.68 ;
      RECT 18.938 0.24 18.984 1.44 ;
      RECT 19.028 0.24 19.762 1.44 ;
      RECT 18.938 -0.12 19.762 0.24 ;
      RECT 18.038 41.04 18.862 41.4 ;
      RECT 18.038 40.32 18.772 41.04 ;
      RECT 18.816 39.84 18.862 41.04 ;
      RECT 18.216 39.84 18.772 40.32 ;
      RECT 18.216 39.6 18.862 39.84 ;
      RECT 18.038 39.12 18.084 40.32 ;
      RECT 18.128 39.12 18.172 40.32 ;
      RECT 18.216 39.12 18.772 39.6 ;
      RECT 18.038 38.88 18.772 39.12 ;
      RECT 18.816 38.4 18.862 39.6 ;
      RECT 18.216 38.4 18.772 38.88 ;
      RECT 18.216 38.16 18.862 38.4 ;
      RECT 18.038 37.68 18.084 38.88 ;
      RECT 18.128 37.68 18.172 38.88 ;
      RECT 18.216 37.68 18.772 38.16 ;
      RECT 18.038 37.44 18.772 37.68 ;
      RECT 18.816 36.96 18.862 38.16 ;
      RECT 18.216 36.96 18.772 37.44 ;
      RECT 18.216 36.72 18.862 36.96 ;
      RECT 18.038 36.24 18.084 37.44 ;
      RECT 18.128 36.24 18.172 37.44 ;
      RECT 18.216 36.24 18.772 36.72 ;
      RECT 18.038 36 18.772 36.24 ;
      RECT 18.816 35.52 18.862 36.72 ;
      RECT 18.216 35.52 18.772 36 ;
      RECT 18.216 35.28 18.862 35.52 ;
      RECT 18.038 34.8 18.084 36 ;
      RECT 18.128 34.8 18.172 36 ;
      RECT 18.216 34.8 18.772 35.28 ;
      RECT 18.038 34.56 18.772 34.8 ;
      RECT 18.816 34.08 18.862 35.28 ;
      RECT 18.216 34.08 18.772 34.56 ;
      RECT 18.216 33.84 18.862 34.08 ;
      RECT 18.038 33.36 18.084 34.56 ;
      RECT 18.128 33.36 18.172 34.56 ;
      RECT 18.216 33.36 18.772 33.84 ;
      RECT 18.038 33.12 18.772 33.36 ;
      RECT 18.816 32.64 18.862 33.84 ;
      RECT 18.216 32.64 18.772 33.12 ;
      RECT 18.216 32.4 18.862 32.64 ;
      RECT 18.038 31.92 18.084 33.12 ;
      RECT 18.128 31.92 18.172 33.12 ;
      RECT 18.216 31.92 18.772 32.4 ;
      RECT 18.038 31.68 18.772 31.92 ;
      RECT 18.816 31.2 18.862 32.4 ;
      RECT 18.216 31.2 18.772 31.68 ;
      RECT 18.216 30.96 18.862 31.2 ;
      RECT 18.038 30.48 18.084 31.68 ;
      RECT 18.128 30.48 18.172 31.68 ;
      RECT 18.216 30.48 18.772 30.96 ;
      RECT 18.038 30.24 18.772 30.48 ;
      RECT 18.816 29.76 18.862 30.96 ;
      RECT 18.216 29.76 18.772 30.24 ;
      RECT 18.216 29.52 18.862 29.76 ;
      RECT 18.038 29.04 18.084 30.24 ;
      RECT 18.128 29.04 18.172 30.24 ;
      RECT 18.216 29.04 18.772 29.52 ;
      RECT 18.038 28.8 18.772 29.04 ;
      RECT 18.816 28.32 18.862 29.52 ;
      RECT 18.216 28.32 18.772 28.8 ;
      RECT 18.216 28.08 18.862 28.32 ;
      RECT 18.038 27.6 18.084 28.8 ;
      RECT 18.128 27.6 18.172 28.8 ;
      RECT 18.216 27.6 18.772 28.08 ;
      RECT 18.038 27.36 18.772 27.6 ;
      RECT 18.816 26.88 18.862 28.08 ;
      RECT 18.216 26.88 18.772 27.36 ;
      RECT 18.216 26.64 18.862 26.88 ;
      RECT 18.038 26.16 18.084 27.36 ;
      RECT 18.128 26.16 18.172 27.36 ;
      RECT 18.216 26.16 18.772 26.64 ;
      RECT 18.038 25.92 18.772 26.16 ;
      RECT 18.816 25.44 18.862 26.64 ;
      RECT 18.128 25.44 18.772 25.92 ;
      RECT 18.128 25.2 18.862 25.44 ;
      RECT 18.038 24.72 18.084 25.92 ;
      RECT 18.128 24.72 18.684 25.2 ;
      RECT 18.728 24 18.772 25.2 ;
      RECT 18.816 24 18.862 25.2 ;
      RECT 18.038 24 18.684 24.72 ;
      RECT 18.038 22.68 18.862 24 ;
      RECT 18.038 21.48 18.084 22.68 ;
      RECT 18.128 21.48 18.172 22.68 ;
      RECT 18.216 21.48 18.428 22.68 ;
      RECT 18.472 21.48 18.684 22.68 ;
      RECT 18.728 21.48 18.862 22.68 ;
      RECT 18.038 18.72 18.862 21.48 ;
      RECT 18.038 18 18.772 18.72 ;
      RECT 18.816 17.52 18.862 18.72 ;
      RECT 18.216 17.52 18.772 18 ;
      RECT 18.216 17.28 18.862 17.52 ;
      RECT 18.038 16.8 18.084 18 ;
      RECT 18.128 16.8 18.172 18 ;
      RECT 18.216 16.8 18.772 17.28 ;
      RECT 18.038 16.56 18.772 16.8 ;
      RECT 18.816 16.08 18.862 17.28 ;
      RECT 18.216 16.08 18.772 16.56 ;
      RECT 18.216 15.84 18.862 16.08 ;
      RECT 18.038 15.36 18.084 16.56 ;
      RECT 18.128 15.36 18.172 16.56 ;
      RECT 18.216 15.36 18.772 15.84 ;
      RECT 18.038 15.12 18.772 15.36 ;
      RECT 18.816 14.64 18.862 15.84 ;
      RECT 18.216 14.64 18.772 15.12 ;
      RECT 18.216 14.4 18.862 14.64 ;
      RECT 18.038 13.92 18.084 15.12 ;
      RECT 18.128 13.92 18.172 15.12 ;
      RECT 18.216 13.92 18.772 14.4 ;
      RECT 18.038 13.68 18.772 13.92 ;
      RECT 18.816 13.2 18.862 14.4 ;
      RECT 18.216 13.2 18.772 13.68 ;
      RECT 18.216 12.96 18.862 13.2 ;
      RECT 18.038 12.48 18.084 13.68 ;
      RECT 18.128 12.48 18.172 13.68 ;
      RECT 18.216 12.48 18.772 12.96 ;
      RECT 18.038 12.24 18.772 12.48 ;
      RECT 18.816 11.76 18.862 12.96 ;
      RECT 18.216 11.76 18.772 12.24 ;
      RECT 18.216 11.52 18.862 11.76 ;
      RECT 18.038 11.04 18.084 12.24 ;
      RECT 18.128 11.04 18.172 12.24 ;
      RECT 18.216 11.04 18.772 11.52 ;
      RECT 18.038 10.8 18.772 11.04 ;
      RECT 18.816 10.32 18.862 11.52 ;
      RECT 18.216 10.32 18.772 10.8 ;
      RECT 18.216 10.08 18.862 10.32 ;
      RECT 18.038 9.6 18.084 10.8 ;
      RECT 18.128 9.6 18.172 10.8 ;
      RECT 18.216 9.6 18.772 10.08 ;
      RECT 18.038 9.36 18.772 9.6 ;
      RECT 18.816 8.88 18.862 10.08 ;
      RECT 18.216 8.88 18.772 9.36 ;
      RECT 18.216 8.64 18.862 8.88 ;
      RECT 18.038 8.16 18.084 9.36 ;
      RECT 18.128 8.16 18.172 9.36 ;
      RECT 18.216 8.16 18.772 8.64 ;
      RECT 18.038 7.92 18.772 8.16 ;
      RECT 18.816 7.44 18.862 8.64 ;
      RECT 18.216 7.44 18.772 7.92 ;
      RECT 18.216 7.2 18.862 7.44 ;
      RECT 18.038 6.72 18.084 7.92 ;
      RECT 18.128 6.72 18.172 7.92 ;
      RECT 18.216 6.72 18.772 7.2 ;
      RECT 18.038 6.48 18.772 6.72 ;
      RECT 18.816 6 18.862 7.2 ;
      RECT 18.216 6 18.772 6.48 ;
      RECT 18.216 5.76 18.862 6 ;
      RECT 18.038 5.28 18.084 6.48 ;
      RECT 18.128 5.28 18.172 6.48 ;
      RECT 18.216 5.28 18.772 5.76 ;
      RECT 18.038 5.04 18.772 5.28 ;
      RECT 18.816 4.56 18.862 5.76 ;
      RECT 18.216 4.56 18.772 5.04 ;
      RECT 18.216 4.32 18.862 4.56 ;
      RECT 18.038 3.84 18.084 5.04 ;
      RECT 18.128 3.84 18.172 5.04 ;
      RECT 18.216 3.84 18.772 4.32 ;
      RECT 18.038 3.6 18.772 3.84 ;
      RECT 18.816 3.12 18.862 4.32 ;
      RECT 18.216 3.12 18.772 3.6 ;
      RECT 18.216 2.88 18.862 3.12 ;
      RECT 18.038 2.4 18.084 3.6 ;
      RECT 18.128 2.4 18.172 3.6 ;
      RECT 18.216 2.4 18.772 2.88 ;
      RECT 18.038 2.16 18.772 2.4 ;
      RECT 18.816 1.68 18.862 2.88 ;
      RECT 18.216 1.68 18.772 2.16 ;
      RECT 18.216 1.44 18.862 1.68 ;
      RECT 18.038 0.96 18.084 2.16 ;
      RECT 18.128 0.96 18.172 2.16 ;
      RECT 18.216 0.96 18.772 1.44 ;
      RECT 18.816 0.24 18.862 1.44 ;
      RECT 18.038 0.24 18.772 0.96 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 41.04 17.962 41.4 ;
      RECT 17.138 39.84 17.272 41.04 ;
      RECT 17.316 39.84 17.528 41.04 ;
      RECT 17.572 39.84 17.962 41.04 ;
      RECT 17.138 39.6 17.962 39.84 ;
      RECT 17.138 38.4 17.272 39.6 ;
      RECT 17.316 38.4 17.528 39.6 ;
      RECT 17.572 38.4 17.962 39.6 ;
      RECT 17.138 38.16 17.962 38.4 ;
      RECT 17.138 36.96 17.272 38.16 ;
      RECT 17.316 36.96 17.528 38.16 ;
      RECT 17.572 36.96 17.962 38.16 ;
      RECT 17.138 36.72 17.962 36.96 ;
      RECT 17.138 35.52 17.272 36.72 ;
      RECT 17.316 35.52 17.528 36.72 ;
      RECT 17.572 35.52 17.962 36.72 ;
      RECT 17.138 35.28 17.962 35.52 ;
      RECT 17.138 34.08 17.272 35.28 ;
      RECT 17.316 34.08 17.528 35.28 ;
      RECT 17.572 34.08 17.962 35.28 ;
      RECT 17.138 33.84 17.962 34.08 ;
      RECT 17.138 32.64 17.272 33.84 ;
      RECT 17.316 32.64 17.528 33.84 ;
      RECT 17.572 32.64 17.962 33.84 ;
      RECT 17.138 32.4 17.962 32.64 ;
      RECT 17.138 31.2 17.272 32.4 ;
      RECT 17.316 31.2 17.528 32.4 ;
      RECT 17.572 31.2 17.962 32.4 ;
      RECT 17.138 30.96 17.962 31.2 ;
      RECT 17.138 29.76 17.272 30.96 ;
      RECT 17.316 29.76 17.528 30.96 ;
      RECT 17.572 29.76 17.962 30.96 ;
      RECT 17.138 29.52 17.962 29.76 ;
      RECT 17.138 28.32 17.272 29.52 ;
      RECT 17.316 28.32 17.528 29.52 ;
      RECT 17.572 28.32 17.962 29.52 ;
      RECT 17.138 28.08 17.962 28.32 ;
      RECT 17.138 26.88 17.272 28.08 ;
      RECT 17.316 26.88 17.528 28.08 ;
      RECT 17.572 26.88 17.962 28.08 ;
      RECT 17.138 26.64 17.962 26.88 ;
      RECT 17.316 25.92 17.962 26.64 ;
      RECT 17.138 25.44 17.184 26.64 ;
      RECT 17.228 25.44 17.272 26.64 ;
      RECT 17.316 25.44 17.528 25.92 ;
      RECT 17.572 24.72 17.872 25.92 ;
      RECT 17.916 24.72 17.962 25.92 ;
      RECT 17.138 24.72 17.528 25.44 ;
      RECT 17.138 24.48 17.962 24.72 ;
      RECT 17.138 23.28 17.272 24.48 ;
      RECT 17.316 23.28 17.528 24.48 ;
      RECT 17.572 23.28 17.784 24.48 ;
      RECT 17.828 23.28 17.872 24.48 ;
      RECT 17.916 23.28 17.962 24.48 ;
      RECT 17.138 20.76 17.962 23.28 ;
      RECT 17.138 19.56 17.184 20.76 ;
      RECT 17.228 19.56 17.784 20.76 ;
      RECT 17.828 19.56 17.872 20.76 ;
      RECT 17.916 19.56 17.962 20.76 ;
      RECT 17.138 18.72 17.962 19.56 ;
      RECT 17.138 17.52 17.272 18.72 ;
      RECT 17.316 17.52 17.528 18.72 ;
      RECT 17.572 17.52 17.962 18.72 ;
      RECT 17.138 17.28 17.962 17.52 ;
      RECT 17.138 16.08 17.272 17.28 ;
      RECT 17.316 16.08 17.528 17.28 ;
      RECT 17.572 16.08 17.962 17.28 ;
      RECT 17.138 15.84 17.962 16.08 ;
      RECT 17.138 14.64 17.272 15.84 ;
      RECT 17.316 14.64 17.528 15.84 ;
      RECT 17.572 14.64 17.962 15.84 ;
      RECT 17.138 14.4 17.962 14.64 ;
      RECT 17.138 13.2 17.272 14.4 ;
      RECT 17.316 13.2 17.528 14.4 ;
      RECT 17.572 13.2 17.962 14.4 ;
      RECT 17.138 12.96 17.962 13.2 ;
      RECT 17.138 11.76 17.272 12.96 ;
      RECT 17.316 11.76 17.528 12.96 ;
      RECT 17.572 11.76 17.962 12.96 ;
      RECT 17.138 11.52 17.962 11.76 ;
      RECT 17.138 10.32 17.272 11.52 ;
      RECT 17.316 10.32 17.528 11.52 ;
      RECT 17.572 10.32 17.962 11.52 ;
      RECT 17.138 10.08 17.962 10.32 ;
      RECT 17.138 8.88 17.272 10.08 ;
      RECT 17.316 8.88 17.528 10.08 ;
      RECT 17.572 8.88 17.962 10.08 ;
      RECT 17.138 8.64 17.962 8.88 ;
      RECT 17.138 7.44 17.272 8.64 ;
      RECT 17.316 7.44 17.528 8.64 ;
      RECT 17.572 7.44 17.962 8.64 ;
      RECT 17.138 7.2 17.962 7.44 ;
      RECT 17.138 6 17.272 7.2 ;
      RECT 17.316 6 17.528 7.2 ;
      RECT 17.572 6 17.962 7.2 ;
      RECT 17.138 5.76 17.962 6 ;
      RECT 17.138 4.56 17.272 5.76 ;
      RECT 17.316 4.56 17.528 5.76 ;
      RECT 17.572 4.56 17.962 5.76 ;
      RECT 17.138 4.32 17.962 4.56 ;
      RECT 17.138 3.12 17.272 4.32 ;
      RECT 17.316 3.12 17.528 4.32 ;
      RECT 17.572 3.12 17.962 4.32 ;
      RECT 17.138 2.88 17.962 3.12 ;
      RECT 17.138 1.68 17.272 2.88 ;
      RECT 17.316 1.68 17.528 2.88 ;
      RECT 17.572 1.68 17.962 2.88 ;
      RECT 17.138 1.44 17.962 1.68 ;
      RECT 17.138 0.24 17.272 1.44 ;
      RECT 17.316 0.24 17.528 1.44 ;
      RECT 17.572 0.24 17.962 1.44 ;
      RECT 17.138 -0.12 17.962 0.24 ;
      RECT 16.238 40.32 17.062 41.4 ;
      RECT 16.238 39.12 16.284 40.32 ;
      RECT 16.328 39.12 16.628 40.32 ;
      RECT 16.672 39.12 16.884 40.32 ;
      RECT 16.928 39.12 17.062 40.32 ;
      RECT 16.238 38.88 17.062 39.12 ;
      RECT 16.238 37.68 16.284 38.88 ;
      RECT 16.328 37.68 16.628 38.88 ;
      RECT 16.672 37.68 16.884 38.88 ;
      RECT 16.928 37.68 17.062 38.88 ;
      RECT 16.238 37.44 17.062 37.68 ;
      RECT 16.238 36.24 16.284 37.44 ;
      RECT 16.328 36.24 16.628 37.44 ;
      RECT 16.672 36.24 16.884 37.44 ;
      RECT 16.928 36.24 17.062 37.44 ;
      RECT 16.238 36 17.062 36.24 ;
      RECT 16.238 34.8 16.284 36 ;
      RECT 16.328 34.8 16.628 36 ;
      RECT 16.672 34.8 16.884 36 ;
      RECT 16.928 34.8 17.062 36 ;
      RECT 16.238 34.56 17.062 34.8 ;
      RECT 16.238 33.36 16.284 34.56 ;
      RECT 16.328 33.36 16.628 34.56 ;
      RECT 16.672 33.36 16.884 34.56 ;
      RECT 16.928 33.36 17.062 34.56 ;
      RECT 16.238 33.12 17.062 33.36 ;
      RECT 16.238 31.92 16.284 33.12 ;
      RECT 16.328 31.92 16.628 33.12 ;
      RECT 16.672 31.92 16.884 33.12 ;
      RECT 16.928 31.92 17.062 33.12 ;
      RECT 16.238 31.68 17.062 31.92 ;
      RECT 16.238 30.48 16.284 31.68 ;
      RECT 16.328 30.48 16.628 31.68 ;
      RECT 16.672 30.48 16.884 31.68 ;
      RECT 16.928 30.48 17.062 31.68 ;
      RECT 16.238 30.24 17.062 30.48 ;
      RECT 16.238 29.04 16.284 30.24 ;
      RECT 16.328 29.04 16.628 30.24 ;
      RECT 16.672 29.04 16.884 30.24 ;
      RECT 16.928 29.04 17.062 30.24 ;
      RECT 16.238 28.8 17.062 29.04 ;
      RECT 16.238 27.6 16.284 28.8 ;
      RECT 16.328 27.6 16.628 28.8 ;
      RECT 16.672 27.6 16.884 28.8 ;
      RECT 16.928 27.6 17.062 28.8 ;
      RECT 16.238 27.36 17.062 27.6 ;
      RECT 16.238 26.16 16.284 27.36 ;
      RECT 16.328 26.16 16.628 27.36 ;
      RECT 16.672 26.16 16.884 27.36 ;
      RECT 16.928 26.16 17.062 27.36 ;
      RECT 16.238 25.92 17.062 26.16 ;
      RECT 16.238 25.2 16.628 25.92 ;
      RECT 16.672 25.2 17.062 25.92 ;
      RECT 16.416 24.72 16.628 25.2 ;
      RECT 16.672 24.72 16.884 25.2 ;
      RECT 16.238 24 16.372 25.2 ;
      RECT 16.928 24 16.972 25.2 ;
      RECT 17.016 24 17.062 25.2 ;
      RECT 16.416 24 16.884 24.72 ;
      RECT 16.238 20.76 17.062 24 ;
      RECT 16.238 19.56 16.284 20.76 ;
      RECT 16.328 19.56 16.372 20.76 ;
      RECT 16.416 19.56 16.628 20.76 ;
      RECT 16.672 19.56 16.884 20.76 ;
      RECT 16.928 19.56 16.972 20.76 ;
      RECT 17.016 19.56 17.062 20.76 ;
      RECT 16.238 18 17.062 19.56 ;
      RECT 16.238 16.8 16.284 18 ;
      RECT 16.328 16.8 16.628 18 ;
      RECT 16.672 16.8 16.884 18 ;
      RECT 16.928 16.8 17.062 18 ;
      RECT 16.238 16.56 17.062 16.8 ;
      RECT 16.238 15.36 16.284 16.56 ;
      RECT 16.328 15.36 16.628 16.56 ;
      RECT 16.672 15.36 16.884 16.56 ;
      RECT 16.928 15.36 17.062 16.56 ;
      RECT 16.238 15.12 17.062 15.36 ;
      RECT 16.238 13.92 16.284 15.12 ;
      RECT 16.328 13.92 16.628 15.12 ;
      RECT 16.672 13.92 16.884 15.12 ;
      RECT 16.928 13.92 17.062 15.12 ;
      RECT 16.238 13.68 17.062 13.92 ;
      RECT 16.238 12.48 16.284 13.68 ;
      RECT 16.328 12.48 16.628 13.68 ;
      RECT 16.672 12.48 16.884 13.68 ;
      RECT 16.928 12.48 17.062 13.68 ;
      RECT 16.238 12.24 17.062 12.48 ;
      RECT 16.238 11.04 16.284 12.24 ;
      RECT 16.328 11.04 16.628 12.24 ;
      RECT 16.672 11.04 16.884 12.24 ;
      RECT 16.928 11.04 17.062 12.24 ;
      RECT 16.238 10.8 17.062 11.04 ;
      RECT 16.238 9.6 16.284 10.8 ;
      RECT 16.328 9.6 16.628 10.8 ;
      RECT 16.672 9.6 16.884 10.8 ;
      RECT 16.928 9.6 17.062 10.8 ;
      RECT 16.238 9.36 17.062 9.6 ;
      RECT 16.238 8.16 16.284 9.36 ;
      RECT 16.328 8.16 16.628 9.36 ;
      RECT 16.672 8.16 16.884 9.36 ;
      RECT 16.928 8.16 17.062 9.36 ;
      RECT 16.238 7.92 17.062 8.16 ;
      RECT 16.238 6.72 16.284 7.92 ;
      RECT 16.328 6.72 16.628 7.92 ;
      RECT 16.672 6.72 16.884 7.92 ;
      RECT 16.928 6.72 17.062 7.92 ;
      RECT 16.238 6.48 17.062 6.72 ;
      RECT 16.238 5.28 16.284 6.48 ;
      RECT 16.328 5.28 16.628 6.48 ;
      RECT 16.672 5.28 16.884 6.48 ;
      RECT 16.928 5.28 17.062 6.48 ;
      RECT 16.238 5.04 17.062 5.28 ;
      RECT 16.238 3.84 16.284 5.04 ;
      RECT 16.328 3.84 16.628 5.04 ;
      RECT 16.672 3.84 16.884 5.04 ;
      RECT 16.928 3.84 17.062 5.04 ;
      RECT 16.238 3.6 17.062 3.84 ;
      RECT 16.238 2.4 16.284 3.6 ;
      RECT 16.328 2.4 16.628 3.6 ;
      RECT 16.672 2.4 16.884 3.6 ;
      RECT 16.928 2.4 17.062 3.6 ;
      RECT 16.238 2.16 17.062 2.4 ;
      RECT 16.238 0.96 16.284 2.16 ;
      RECT 16.328 0.96 16.628 2.16 ;
      RECT 16.672 0.96 16.884 2.16 ;
      RECT 16.928 0.96 17.062 2.16 ;
      RECT 16.238 -0.12 17.062 0.96 ;
      RECT 15.338 41.04 16.162 41.4 ;
      RECT 15.516 40.32 16.162 41.04 ;
      RECT 15.338 39.84 15.384 41.04 ;
      RECT 15.428 39.84 15.472 41.04 ;
      RECT 15.516 39.84 16.072 40.32 ;
      RECT 15.338 39.6 16.072 39.84 ;
      RECT 16.116 39.12 16.162 40.32 ;
      RECT 15.516 39.12 16.072 39.6 ;
      RECT 15.516 38.88 16.162 39.12 ;
      RECT 15.338 38.4 15.384 39.6 ;
      RECT 15.428 38.4 15.472 39.6 ;
      RECT 15.516 38.4 16.072 38.88 ;
      RECT 15.338 38.16 16.072 38.4 ;
      RECT 16.116 37.68 16.162 38.88 ;
      RECT 15.516 37.68 16.072 38.16 ;
      RECT 15.516 37.44 16.162 37.68 ;
      RECT 15.338 36.96 15.384 38.16 ;
      RECT 15.428 36.96 15.472 38.16 ;
      RECT 15.516 36.96 16.072 37.44 ;
      RECT 15.338 36.72 16.072 36.96 ;
      RECT 16.116 36.24 16.162 37.44 ;
      RECT 15.516 36.24 16.072 36.72 ;
      RECT 15.516 36 16.162 36.24 ;
      RECT 15.338 35.52 15.384 36.72 ;
      RECT 15.428 35.52 15.472 36.72 ;
      RECT 15.516 35.52 16.072 36 ;
      RECT 15.338 35.28 16.072 35.52 ;
      RECT 16.116 34.8 16.162 36 ;
      RECT 15.516 34.8 16.072 35.28 ;
      RECT 15.516 34.56 16.162 34.8 ;
      RECT 15.338 34.08 15.384 35.28 ;
      RECT 15.428 34.08 15.472 35.28 ;
      RECT 15.516 34.08 16.072 34.56 ;
      RECT 15.338 33.84 16.072 34.08 ;
      RECT 16.116 33.36 16.162 34.56 ;
      RECT 15.516 33.36 16.072 33.84 ;
      RECT 15.516 33.12 16.162 33.36 ;
      RECT 15.338 32.64 15.384 33.84 ;
      RECT 15.428 32.64 15.472 33.84 ;
      RECT 15.516 32.64 16.072 33.12 ;
      RECT 15.338 32.4 16.072 32.64 ;
      RECT 16.116 31.92 16.162 33.12 ;
      RECT 15.516 31.92 16.072 32.4 ;
      RECT 15.516 31.68 16.162 31.92 ;
      RECT 15.338 31.2 15.384 32.4 ;
      RECT 15.428 31.2 15.472 32.4 ;
      RECT 15.516 31.2 16.072 31.68 ;
      RECT 15.338 30.96 16.072 31.2 ;
      RECT 16.116 30.48 16.162 31.68 ;
      RECT 15.516 30.48 16.072 30.96 ;
      RECT 15.516 30.24 16.162 30.48 ;
      RECT 15.338 29.76 15.384 30.96 ;
      RECT 15.428 29.76 15.472 30.96 ;
      RECT 15.516 29.76 16.072 30.24 ;
      RECT 15.338 29.52 16.072 29.76 ;
      RECT 16.116 29.04 16.162 30.24 ;
      RECT 15.516 29.04 16.072 29.52 ;
      RECT 15.516 28.8 16.162 29.04 ;
      RECT 15.338 28.32 15.384 29.52 ;
      RECT 15.428 28.32 15.472 29.52 ;
      RECT 15.516 28.32 16.072 28.8 ;
      RECT 15.338 28.08 16.072 28.32 ;
      RECT 16.116 27.6 16.162 28.8 ;
      RECT 15.516 27.6 16.072 28.08 ;
      RECT 15.516 27.36 16.162 27.6 ;
      RECT 15.338 26.88 15.384 28.08 ;
      RECT 15.428 26.88 15.472 28.08 ;
      RECT 15.516 26.88 16.072 27.36 ;
      RECT 15.338 26.64 16.072 26.88 ;
      RECT 16.116 26.16 16.162 27.36 ;
      RECT 15.516 26.16 16.072 26.64 ;
      RECT 15.516 25.92 16.162 26.16 ;
      RECT 15.338 25.44 15.384 26.64 ;
      RECT 15.428 25.44 15.472 26.64 ;
      RECT 15.516 25.44 15.728 25.92 ;
      RECT 15.338 25.2 15.728 25.44 ;
      RECT 15.772 24.72 15.984 25.92 ;
      RECT 16.028 24.72 16.162 25.92 ;
      RECT 15.428 24.72 15.728 25.2 ;
      RECT 15.428 24.48 16.162 24.72 ;
      RECT 15.338 24 15.384 25.2 ;
      RECT 15.428 24 15.728 24.48 ;
      RECT 15.772 23.28 15.984 24.48 ;
      RECT 16.028 23.28 16.162 24.48 ;
      RECT 15.338 23.28 15.728 24 ;
      RECT 15.338 20.76 16.162 23.28 ;
      RECT 15.338 19.56 15.728 20.76 ;
      RECT 15.772 19.56 15.984 20.76 ;
      RECT 16.028 19.56 16.072 20.76 ;
      RECT 16.116 19.56 16.162 20.76 ;
      RECT 15.338 18.72 16.162 19.56 ;
      RECT 15.516 18 16.162 18.72 ;
      RECT 15.338 17.52 15.384 18.72 ;
      RECT 15.428 17.52 15.472 18.72 ;
      RECT 15.516 17.52 16.072 18 ;
      RECT 15.338 17.28 16.072 17.52 ;
      RECT 16.116 16.8 16.162 18 ;
      RECT 15.516 16.8 16.072 17.28 ;
      RECT 15.516 16.56 16.162 16.8 ;
      RECT 15.338 16.08 15.384 17.28 ;
      RECT 15.428 16.08 15.472 17.28 ;
      RECT 15.516 16.08 16.072 16.56 ;
      RECT 15.338 15.84 16.072 16.08 ;
      RECT 16.116 15.36 16.162 16.56 ;
      RECT 15.516 15.36 16.072 15.84 ;
      RECT 15.516 15.12 16.162 15.36 ;
      RECT 15.338 14.64 15.384 15.84 ;
      RECT 15.428 14.64 15.472 15.84 ;
      RECT 15.516 14.64 16.072 15.12 ;
      RECT 15.338 14.4 16.072 14.64 ;
      RECT 16.116 13.92 16.162 15.12 ;
      RECT 15.516 13.92 16.072 14.4 ;
      RECT 15.516 13.68 16.162 13.92 ;
      RECT 15.338 13.2 15.384 14.4 ;
      RECT 15.428 13.2 15.472 14.4 ;
      RECT 15.516 13.2 16.072 13.68 ;
      RECT 15.338 12.96 16.072 13.2 ;
      RECT 16.116 12.48 16.162 13.68 ;
      RECT 15.516 12.48 16.072 12.96 ;
      RECT 15.516 12.24 16.162 12.48 ;
      RECT 15.338 11.76 15.384 12.96 ;
      RECT 15.428 11.76 15.472 12.96 ;
      RECT 15.516 11.76 16.072 12.24 ;
      RECT 15.338 11.52 16.072 11.76 ;
      RECT 16.116 11.04 16.162 12.24 ;
      RECT 15.516 11.04 16.072 11.52 ;
      RECT 15.516 10.8 16.162 11.04 ;
      RECT 15.338 10.32 15.384 11.52 ;
      RECT 15.428 10.32 15.472 11.52 ;
      RECT 15.516 10.32 16.072 10.8 ;
      RECT 15.338 10.08 16.072 10.32 ;
      RECT 16.116 9.6 16.162 10.8 ;
      RECT 15.516 9.6 16.072 10.08 ;
      RECT 15.516 9.36 16.162 9.6 ;
      RECT 15.338 8.88 15.384 10.08 ;
      RECT 15.428 8.88 15.472 10.08 ;
      RECT 15.516 8.88 16.072 9.36 ;
      RECT 15.338 8.64 16.072 8.88 ;
      RECT 16.116 8.16 16.162 9.36 ;
      RECT 15.516 8.16 16.072 8.64 ;
      RECT 15.516 7.92 16.162 8.16 ;
      RECT 15.338 7.44 15.384 8.64 ;
      RECT 15.428 7.44 15.472 8.64 ;
      RECT 15.516 7.44 16.072 7.92 ;
      RECT 15.338 7.2 16.072 7.44 ;
      RECT 16.116 6.72 16.162 7.92 ;
      RECT 15.516 6.72 16.072 7.2 ;
      RECT 15.516 6.48 16.162 6.72 ;
      RECT 15.338 6 15.384 7.2 ;
      RECT 15.428 6 15.472 7.2 ;
      RECT 15.516 6 16.072 6.48 ;
      RECT 15.338 5.76 16.072 6 ;
      RECT 16.116 5.28 16.162 6.48 ;
      RECT 15.516 5.28 16.072 5.76 ;
      RECT 15.516 5.04 16.162 5.28 ;
      RECT 15.338 4.56 15.384 5.76 ;
      RECT 15.428 4.56 15.472 5.76 ;
      RECT 15.516 4.56 16.072 5.04 ;
      RECT 15.338 4.32 16.072 4.56 ;
      RECT 16.116 3.84 16.162 5.04 ;
      RECT 15.516 3.84 16.072 4.32 ;
      RECT 15.516 3.6 16.162 3.84 ;
      RECT 15.338 3.12 15.384 4.32 ;
      RECT 15.428 3.12 15.472 4.32 ;
      RECT 15.516 3.12 16.072 3.6 ;
      RECT 15.338 2.88 16.072 3.12 ;
      RECT 16.116 2.4 16.162 3.6 ;
      RECT 15.516 2.4 16.072 2.88 ;
      RECT 15.516 2.16 16.162 2.4 ;
      RECT 15.338 1.68 15.384 2.88 ;
      RECT 15.428 1.68 15.472 2.88 ;
      RECT 15.516 1.68 16.072 2.16 ;
      RECT 15.338 1.44 16.072 1.68 ;
      RECT 16.116 0.96 16.162 2.16 ;
      RECT 16.028 0.96 16.072 1.44 ;
      RECT 15.338 0.24 15.728 1.44 ;
      RECT 15.772 0.24 15.984 1.44 ;
      RECT 16.028 0.24 16.162 0.96 ;
      RECT 15.338 -0.12 16.162 0.24 ;
      RECT 14.438 41.04 15.262 41.4 ;
      RECT 14.438 39.84 14.572 41.04 ;
      RECT 14.616 39.84 14.828 41.04 ;
      RECT 14.872 39.84 15.262 41.04 ;
      RECT 14.438 39.6 15.262 39.84 ;
      RECT 14.438 38.4 14.572 39.6 ;
      RECT 14.616 38.4 14.828 39.6 ;
      RECT 14.872 38.4 15.262 39.6 ;
      RECT 14.438 38.16 15.262 38.4 ;
      RECT 14.438 36.96 14.572 38.16 ;
      RECT 14.616 36.96 14.828 38.16 ;
      RECT 14.872 36.96 15.262 38.16 ;
      RECT 14.438 36.72 15.262 36.96 ;
      RECT 14.438 35.52 14.572 36.72 ;
      RECT 14.616 35.52 14.828 36.72 ;
      RECT 14.872 35.52 15.262 36.72 ;
      RECT 14.438 35.28 15.262 35.52 ;
      RECT 14.438 34.08 14.572 35.28 ;
      RECT 14.616 34.08 14.828 35.28 ;
      RECT 14.872 34.08 15.262 35.28 ;
      RECT 14.438 33.84 15.262 34.08 ;
      RECT 14.438 32.64 14.572 33.84 ;
      RECT 14.616 32.64 14.828 33.84 ;
      RECT 14.872 32.64 15.262 33.84 ;
      RECT 14.438 32.4 15.262 32.64 ;
      RECT 14.438 31.2 14.572 32.4 ;
      RECT 14.616 31.2 14.828 32.4 ;
      RECT 14.872 31.2 15.262 32.4 ;
      RECT 14.438 30.96 15.262 31.2 ;
      RECT 14.438 29.76 14.572 30.96 ;
      RECT 14.616 29.76 14.828 30.96 ;
      RECT 14.872 29.76 15.262 30.96 ;
      RECT 14.438 29.52 15.262 29.76 ;
      RECT 14.438 28.32 14.572 29.52 ;
      RECT 14.616 28.32 14.828 29.52 ;
      RECT 14.872 28.32 15.262 29.52 ;
      RECT 14.438 28.08 15.262 28.32 ;
      RECT 14.438 26.88 14.572 28.08 ;
      RECT 14.616 26.88 14.828 28.08 ;
      RECT 14.872 26.88 15.262 28.08 ;
      RECT 14.438 26.64 15.262 26.88 ;
      RECT 14.528 25.92 15.262 26.64 ;
      RECT 14.438 25.44 14.484 26.64 ;
      RECT 14.528 25.44 14.828 25.92 ;
      RECT 14.872 24.72 15.262 25.92 ;
      RECT 14.438 24.72 14.828 25.44 ;
      RECT 14.438 24.48 15.262 24.72 ;
      RECT 14.438 23.28 14.572 24.48 ;
      RECT 14.616 23.28 14.828 24.48 ;
      RECT 14.872 23.28 15.262 24.48 ;
      RECT 14.438 22.68 15.262 23.28 ;
      RECT 14.438 21.48 14.484 22.68 ;
      RECT 14.528 21.48 15.084 22.68 ;
      RECT 15.128 21.48 15.262 22.68 ;
      RECT 14.438 20.76 15.262 21.48 ;
      RECT 14.438 19.56 15.084 20.76 ;
      RECT 15.128 19.56 15.172 20.76 ;
      RECT 15.216 19.56 15.262 20.76 ;
      RECT 14.438 18.72 15.262 19.56 ;
      RECT 14.438 17.52 14.572 18.72 ;
      RECT 14.616 17.52 14.828 18.72 ;
      RECT 14.872 17.52 15.262 18.72 ;
      RECT 14.438 17.28 15.262 17.52 ;
      RECT 14.438 16.08 14.572 17.28 ;
      RECT 14.616 16.08 14.828 17.28 ;
      RECT 14.872 16.08 15.262 17.28 ;
      RECT 14.438 15.84 15.262 16.08 ;
      RECT 14.438 14.64 14.572 15.84 ;
      RECT 14.616 14.64 14.828 15.84 ;
      RECT 14.872 14.64 15.262 15.84 ;
      RECT 14.438 14.4 15.262 14.64 ;
      RECT 14.438 13.2 14.572 14.4 ;
      RECT 14.616 13.2 14.828 14.4 ;
      RECT 14.872 13.2 15.262 14.4 ;
      RECT 14.438 12.96 15.262 13.2 ;
      RECT 14.438 11.76 14.572 12.96 ;
      RECT 14.616 11.76 14.828 12.96 ;
      RECT 14.872 11.76 15.262 12.96 ;
      RECT 14.438 11.52 15.262 11.76 ;
      RECT 14.438 10.32 14.572 11.52 ;
      RECT 14.616 10.32 14.828 11.52 ;
      RECT 14.872 10.32 15.262 11.52 ;
      RECT 14.438 10.08 15.262 10.32 ;
      RECT 14.438 8.88 14.572 10.08 ;
      RECT 14.616 8.88 14.828 10.08 ;
      RECT 14.872 8.88 15.262 10.08 ;
      RECT 14.438 8.64 15.262 8.88 ;
      RECT 14.438 7.44 14.572 8.64 ;
      RECT 14.616 7.44 14.828 8.64 ;
      RECT 14.872 7.44 15.262 8.64 ;
      RECT 14.438 7.2 15.262 7.44 ;
      RECT 14.438 6 14.572 7.2 ;
      RECT 14.616 6 14.828 7.2 ;
      RECT 14.872 6 15.262 7.2 ;
      RECT 14.438 5.76 15.262 6 ;
      RECT 14.438 4.56 14.572 5.76 ;
      RECT 14.616 4.56 14.828 5.76 ;
      RECT 14.872 4.56 15.262 5.76 ;
      RECT 14.438 4.32 15.262 4.56 ;
      RECT 14.438 3.12 14.572 4.32 ;
      RECT 14.616 3.12 14.828 4.32 ;
      RECT 14.872 3.12 15.262 4.32 ;
      RECT 14.438 2.88 15.262 3.12 ;
      RECT 14.438 1.68 14.572 2.88 ;
      RECT 14.616 1.68 14.828 2.88 ;
      RECT 14.872 1.68 15.262 2.88 ;
      RECT 14.438 -0.12 15.262 1.68 ;
      RECT 13.538 40.32 14.362 41.4 ;
      RECT 13.538 39.12 13.584 40.32 ;
      RECT 13.628 39.12 13.672 40.32 ;
      RECT 13.716 39.12 14.362 40.32 ;
      RECT 13.538 38.88 14.362 39.12 ;
      RECT 13.538 37.68 13.584 38.88 ;
      RECT 13.628 37.68 13.672 38.88 ;
      RECT 13.716 37.68 14.362 38.88 ;
      RECT 13.538 37.44 14.362 37.68 ;
      RECT 13.538 36.24 13.584 37.44 ;
      RECT 13.628 36.24 13.672 37.44 ;
      RECT 13.716 36.24 14.362 37.44 ;
      RECT 13.538 36 14.362 36.24 ;
      RECT 13.538 34.8 13.584 36 ;
      RECT 13.628 34.8 13.672 36 ;
      RECT 13.716 34.8 14.362 36 ;
      RECT 13.538 34.56 14.362 34.8 ;
      RECT 13.538 33.36 13.584 34.56 ;
      RECT 13.628 33.36 13.672 34.56 ;
      RECT 13.716 33.36 14.362 34.56 ;
      RECT 13.538 33.12 14.362 33.36 ;
      RECT 13.538 31.92 13.584 33.12 ;
      RECT 13.628 31.92 13.672 33.12 ;
      RECT 13.716 31.92 14.362 33.12 ;
      RECT 13.538 31.68 14.362 31.92 ;
      RECT 13.538 30.48 13.584 31.68 ;
      RECT 13.628 30.48 13.672 31.68 ;
      RECT 13.716 30.48 14.362 31.68 ;
      RECT 13.538 30.24 14.362 30.48 ;
      RECT 13.538 29.04 13.584 30.24 ;
      RECT 13.628 29.04 13.672 30.24 ;
      RECT 13.716 29.04 14.362 30.24 ;
      RECT 13.538 28.8 14.362 29.04 ;
      RECT 13.538 27.6 13.584 28.8 ;
      RECT 13.628 27.6 13.672 28.8 ;
      RECT 13.716 27.6 14.362 28.8 ;
      RECT 13.538 27.36 14.362 27.6 ;
      RECT 13.716 26.64 14.362 27.36 ;
      RECT 13.538 26.16 13.584 27.36 ;
      RECT 13.628 26.16 13.672 27.36 ;
      RECT 13.716 26.16 14.272 26.64 ;
      RECT 13.538 25.92 14.272 26.16 ;
      RECT 14.316 25.44 14.362 26.64 ;
      RECT 13.628 25.44 14.272 25.92 ;
      RECT 13.628 25.2 14.362 25.44 ;
      RECT 13.538 24.72 13.584 25.92 ;
      RECT 13.628 24.72 13.928 25.2 ;
      RECT 13.972 24 14.184 25.2 ;
      RECT 14.228 24 14.362 25.2 ;
      RECT 13.538 24 13.928 24.72 ;
      RECT 13.538 22.68 14.362 24 ;
      RECT 13.538 21.48 13.584 22.68 ;
      RECT 13.628 21.48 13.672 22.68 ;
      RECT 13.716 21.48 13.928 22.68 ;
      RECT 13.972 21.48 14.184 22.68 ;
      RECT 14.228 21.48 14.272 22.68 ;
      RECT 14.316 21.48 14.362 22.68 ;
      RECT 13.538 18 14.362 21.48 ;
      RECT 13.538 16.8 13.584 18 ;
      RECT 13.628 16.8 13.672 18 ;
      RECT 13.716 16.8 14.362 18 ;
      RECT 13.538 16.56 14.362 16.8 ;
      RECT 13.538 15.36 13.584 16.56 ;
      RECT 13.628 15.36 13.672 16.56 ;
      RECT 13.716 15.36 14.362 16.56 ;
      RECT 13.538 15.12 14.362 15.36 ;
      RECT 13.538 13.92 13.584 15.12 ;
      RECT 13.628 13.92 13.672 15.12 ;
      RECT 13.716 13.92 14.362 15.12 ;
      RECT 13.538 13.68 14.362 13.92 ;
      RECT 13.538 12.48 13.584 13.68 ;
      RECT 13.628 12.48 13.672 13.68 ;
      RECT 13.716 12.48 14.362 13.68 ;
      RECT 13.538 12.24 14.362 12.48 ;
      RECT 13.538 11.04 13.584 12.24 ;
      RECT 13.628 11.04 13.672 12.24 ;
      RECT 13.716 11.04 14.362 12.24 ;
      RECT 13.538 10.8 14.362 11.04 ;
      RECT 13.538 9.6 13.584 10.8 ;
      RECT 13.628 9.6 13.672 10.8 ;
      RECT 13.716 9.6 14.362 10.8 ;
      RECT 13.538 9.36 14.362 9.6 ;
      RECT 13.538 8.16 13.584 9.36 ;
      RECT 13.628 8.16 13.672 9.36 ;
      RECT 13.716 8.16 14.362 9.36 ;
      RECT 13.538 7.92 14.362 8.16 ;
      RECT 13.538 6.72 13.584 7.92 ;
      RECT 13.628 6.72 13.672 7.92 ;
      RECT 13.716 6.72 14.362 7.92 ;
      RECT 13.538 6.48 14.362 6.72 ;
      RECT 13.538 5.28 13.584 6.48 ;
      RECT 13.628 5.28 13.672 6.48 ;
      RECT 13.716 5.28 14.362 6.48 ;
      RECT 13.538 5.04 14.362 5.28 ;
      RECT 13.538 3.84 13.584 5.04 ;
      RECT 13.628 3.84 13.672 5.04 ;
      RECT 13.716 3.84 14.362 5.04 ;
      RECT 13.538 3.6 14.362 3.84 ;
      RECT 13.538 2.4 13.584 3.6 ;
      RECT 13.628 2.4 13.672 3.6 ;
      RECT 13.716 2.4 14.362 3.6 ;
      RECT 13.538 2.16 14.362 2.4 ;
      RECT 13.538 1.44 13.928 2.16 ;
      RECT 13.972 0.96 14.184 2.16 ;
      RECT 14.228 0.96 14.362 2.16 ;
      RECT 13.716 0.96 13.928 1.44 ;
      RECT 13.538 0.24 13.584 1.44 ;
      RECT 13.628 0.24 13.672 1.44 ;
      RECT 13.716 0.24 14.362 0.96 ;
      RECT 13.538 -0.12 14.362 0.24 ;
      RECT 12.638 -0.12 13.462 41.4 ;
      RECT 11.738 -0.12 12.562 41.4 ;
      RECT 10.838 -0.12 11.662 41.4 ;
      RECT 9.938 -0.12 10.762 41.4 ;
      RECT 9.038 -0.12 9.862 41.4 ;
      RECT 8.138 -0.12 8.962 41.4 ;
      RECT 7.238 -0.12 8.062 41.4 ;
      RECT 6.338 -0.12 7.162 41.4 ;
      RECT 5.438 -0.12 6.262 41.4 ;
      RECT 4.538 -0.12 5.362 41.4 ;
      RECT 3.638 -0.12 4.462 41.4 ;
      RECT 2.738 -0.12 3.562 41.4 ;
      RECT 1.838 -0.12 2.662 41.4 ;
      RECT 0.938 -0.12 1.762 41.4 ;
      RECT -0.04 41.34 0.862 41.4 ;
      RECT -0.092 -0.06 0.862 41.34 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 33.458 0 34.12 41.28 ;
      RECT 32.558 0 33.142 41.28 ;
      RECT 31.658 0 32.242 41.28 ;
      RECT 30.758 0 31.342 41.28 ;
      RECT 29.858 0 30.442 41.28 ;
      RECT 28.958 0 29.542 41.28 ;
      RECT 28.058 0 28.642 41.28 ;
      RECT 27.158 0 27.742 41.28 ;
      RECT 26.258 0 26.842 41.28 ;
      RECT 25.358 0 25.942 41.28 ;
      RECT 24.458 0 25.042 41.28 ;
      RECT 23.558 0 24.142 41.28 ;
      RECT 22.658 0 23.242 41.28 ;
      RECT 21.758 0 22.342 41.28 ;
      RECT 20.858 0 21.442 41.28 ;
      RECT 19.958 0 20.542 41.28 ;
      RECT 19.058 41.16 19.642 41.28 ;
      RECT 19.148 25.32 19.642 41.16 ;
      RECT 19.058 22.8 19.642 25.32 ;
      RECT 19.236 21.36 19.642 22.8 ;
      RECT 19.058 18.84 19.642 21.36 ;
      RECT 19.148 0.12 19.642 18.84 ;
      RECT 19.058 0 19.642 0.12 ;
      RECT 18.158 41.16 18.742 41.28 ;
      RECT 18.158 40.44 18.652 41.16 ;
      RECT 18.336 26.04 18.652 40.44 ;
      RECT 18.248 25.32 18.652 26.04 ;
      RECT 18.248 24.6 18.564 25.32 ;
      RECT 18.158 23.88 18.564 24.6 ;
      RECT 18.158 22.8 18.742 23.88 ;
      RECT 17.258 41.16 17.842 41.28 ;
      RECT 17.692 26.76 17.842 41.16 ;
      RECT 17.436 26.04 17.842 26.76 ;
      RECT 17.692 24.6 17.752 26.04 ;
      RECT 16.358 40.44 16.942 41.28 ;
      RECT 16.448 26.04 16.508 40.44 ;
      RECT 16.358 25.32 16.508 26.04 ;
      RECT 15.458 41.16 16.042 41.28 ;
      RECT 15.636 40.44 16.042 41.16 ;
      RECT 15.636 26.04 15.952 40.44 ;
      RECT 14.558 41.16 15.142 41.28 ;
      RECT 14.992 26.76 15.142 41.16 ;
      RECT 14.648 26.04 15.142 26.76 ;
      RECT 14.648 25.32 14.708 26.04 ;
      RECT 14.558 24.6 14.708 25.32 ;
      RECT 14.992 23.16 15.142 26.04 ;
      RECT 14.558 22.8 15.142 23.16 ;
      RECT 14.648 21.36 14.964 22.8 ;
      RECT 14.558 20.88 15.142 21.36 ;
      RECT 14.558 19.44 14.964 20.88 ;
      RECT 14.558 18.84 15.142 19.44 ;
      RECT 14.992 1.56 15.142 18.84 ;
      RECT 14.558 0 15.142 1.56 ;
      RECT 13.658 40.44 14.242 41.28 ;
      RECT 13.836 26.76 14.242 40.44 ;
      RECT 13.836 26.04 14.152 26.76 ;
      RECT 13.748 25.32 14.152 26.04 ;
      RECT 13.748 24.6 13.808 25.32 ;
      RECT 13.658 23.88 13.808 24.6 ;
      RECT 13.658 22.8 14.242 23.88 ;
      RECT 12.758 0 13.342 41.28 ;
      RECT 11.858 0 12.442 41.28 ;
      RECT 10.958 0 11.542 41.28 ;
      RECT 10.058 0 10.642 41.28 ;
      RECT 9.158 0 9.742 41.28 ;
      RECT 8.258 0 8.842 41.28 ;
      RECT 7.358 0 7.942 41.28 ;
      RECT 6.458 0 7.042 41.28 ;
      RECT 5.558 0 6.142 41.28 ;
      RECT 4.658 0 5.242 41.28 ;
      RECT 3.758 0 4.342 41.28 ;
      RECT 2.858 0 3.442 41.28 ;
      RECT 1.958 0 2.542 41.28 ;
      RECT 1.058 0 1.642 41.28 ;
      RECT 0.08 0 0.742 41.28 ;
      RECT 16.792 25.32 16.942 26.04 ;
      RECT 17.258 24.6 17.408 25.32 ;
      RECT 15.548 23.88 15.608 25.32 ;
      RECT 15.458 23.16 15.608 23.88 ;
      RECT 15.458 20.88 16.042 23.16 ;
      RECT 15.458 19.44 15.608 20.88 ;
      RECT 15.458 18.84 16.042 19.44 ;
      RECT 15.636 18.12 16.042 18.84 ;
      RECT 15.636 1.56 15.952 18.12 ;
      RECT 16.536 23.88 16.764 24.6 ;
      RECT 16.358 20.88 16.942 23.88 ;
      RECT 17.258 20.88 17.842 23.16 ;
      RECT 17.348 19.44 17.664 20.88 ;
      RECT 17.258 18.84 17.842 19.44 ;
      RECT 17.692 0.12 17.842 18.84 ;
      RECT 17.258 0 17.842 0.12 ;
      RECT 18.158 18.84 18.742 21.36 ;
      RECT 18.158 18.12 18.652 18.84 ;
      RECT 18.336 0.84 18.652 18.12 ;
      RECT 18.158 0.12 18.652 0.84 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 13.658 18.12 14.242 21.36 ;
      RECT 13.836 2.28 14.242 18.12 ;
      RECT 16.358 18.12 16.942 19.44 ;
      RECT 16.448 0.84 16.508 18.12 ;
      RECT 16.358 0 16.942 0.84 ;
      RECT 13.658 1.56 13.808 2.28 ;
      RECT 15.458 0.12 15.608 1.56 ;
      RECT 15.458 0 16.042 0.12 ;
      RECT 13.836 0.12 14.242 0.84 ;
      RECT 13.658 0 14.242 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 34.2 41.278 ;
    LAYER m1 ;
      RECT 0 0 34.2 41.28 ;
    LAYER m2 ;
      RECT 0 0.015 34.2 41.265 ;
    LAYER m3 ;
      RECT 0.015 0 34.185 41.28 ;
    LAYER m4 ;
      RECT 0 0.02 34.2 41.26 ;
    LAYER m5 ;
      RECT 0.012 0 34.188 41.28 ;
    LAYER m6 ;
      RECT 0 0.012 34.2 41.268 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf192b080e1r1w0cbbehbaa4acw

END LIBRARY
