//-----------------------------------------------------------------
// Intel Proprietary -- Copyright 2011 Intel -- All rights reserved 
//-----------------------------------------------------------------
// Author       : rravindr
// Date Created : 2014-10-30 
//-----------------------------------------------------------------
// Description:
// ccu_vc_test_pkg package definition
//------------------------------------------------------------------

/**
 * TODO: Add package description
 */
package ccu_vc_test_pkg;
   //------------------------------------------
   // Needed Packages 
   //------------------------------------------
   // OVM
   import ovm_pkg::*;
   `include "ovm_macros.svh"

   // Saola
   import sla_pkg::*;
   `include "sla_macros.svh"

   import ccu_vc_pkg::*;
   import ccu_vc_env_pkg::*;
   
   //------------------------------------------
   // Classes definitions 
   //------------------------------------------
   `include "ccu_vc_test.svh"
   `include "ccu_vc_test_rand_dly.svh"
   `include "test01.svh"
   `include "test02.svh"
   `include "test03.svh"
   `include "test04.svh"
   `include "test05.svh"
   `include "test06.svh"
   `include "test07.svh"
   `include "test08.svh"
   `include "test09.svh"
   `include "test10.svh"
   `include "test11.svh"
   `include "test12.svh"
   `include "test13.svh"
   `include "test14.svh"
   `include "test15.svh"
   `include "test16.svh"
   `include "test17.svh"
endpackage :ccu_vc_test_pkg

