VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf124b064e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf124b064e1r1w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 27 BY 28.8 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 14.76 13.972 15.96 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 12.84 11.016 14.04 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 14.76 15.216 15.96 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 14.76 15.428 15.96 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 14.76 15.516 15.96 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 14.76 10.372 15.96 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 14.76 10.628 15.96 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 14.76 10.716 15.96 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 14.76 14.228 15.96 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 14.76 14.316 15.96 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 14.76 14.872 15.96 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 14.76 15.128 15.96 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 12.84 12.172 14.04 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 12.84 12.428 14.04 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 12.84 12.816 14.04 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 12.84 13.416 14.04 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 12.84 13.628 14.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 12.84 13.716 14.04 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 12.84 11.272 14.04 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 12.84 11.528 14.04 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 0.24 12.172 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 23.04 11.828 24.24 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 23.04 11.916 24.24 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 23.04 13.716 24.24 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 23.04 13.972 24.24 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 23.76 12.516 24.96 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 23.76 12.728 24.96 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 23.76 13.072 24.96 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 23.76 13.328 24.96 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 24.48 11.828 25.68 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 24.48 11.916 25.68 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 1.68 13.716 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 24.48 13.716 25.68 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 24.48 13.972 25.68 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 25.2 12.516 26.4 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 25.2 12.728 26.4 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 25.2 13.072 26.4 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 25.2 13.328 26.4 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 25.92 11.828 27.12 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 25.92 11.916 27.12 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 25.92 13.716 27.12 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 25.92 13.972 27.12 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 1.68 13.972 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 26.64 12.516 27.84 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 26.64 12.728 27.84 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 26.64 13.072 27.84 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 26.64 13.328 27.84 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 27.36 11.828 28.56 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 27.36 11.916 28.56 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 27.36 13.716 28.56 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 27.36 13.972 28.56 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 2.4 12.516 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 2.4 12.728 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 2.4 13.072 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 2.4 13.328 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 3.12 11.828 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 3.12 11.916 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.12 13.716 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.12 13.972 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 0.24 12.428 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 3.84 12.516 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 3.84 12.728 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 3.84 13.072 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 3.84 13.328 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 4.56 11.828 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 4.56 11.916 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 4.56 13.716 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 4.56 13.972 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 5.28 12.516 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 5.28 12.728 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.24 13.716 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 5.28 13.072 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 5.28 13.328 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 6 11.828 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 6 11.916 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 6 13.716 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 6 13.972 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 6.72 12.516 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 6.72 12.728 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 6.72 13.072 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 6.72 13.328 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.24 13.972 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 7.44 11.828 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 7.44 11.916 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 7.44 13.716 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 7.44 13.972 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 8.16 12.516 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 8.16 12.728 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 8.16 13.072 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 8.16 13.328 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 8.88 11.828 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 8.88 11.916 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 0.96 12.516 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 8.88 13.716 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 8.88 13.972 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 9.6 12.516 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 9.6 12.728 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 9.6 13.072 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 9.6 13.328 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 10.32 11.828 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 10.32 11.916 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 10.32 13.716 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 10.32 13.972 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 0.96 12.728 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 11.04 12.516 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 11.04 12.728 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 11.04 13.072 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 11.04 13.328 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 16.56 12.728 17.76 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 16.56 12.816 17.76 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 16.56 13.072 17.76 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 16.56 13.328 17.76 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 17.28 12.516 18.48 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 17.28 11.828 18.48 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 0.96 13.072 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 17.28 13.628 18.48 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 17.28 13.716 18.48 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 18 12.172 19.2 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 18 12.428 19.2 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 18 13.972 19.2 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 18 13.072 19.2 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 18.72 11.828 19.92 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 18.72 11.916 19.92 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 18.72 13.628 19.92 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 18.72 13.716 19.92 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 0.96 13.328 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 19.44 12.516 20.64 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 19.44 12.728 20.64 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 19.44 13.072 20.64 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 19.44 13.328 20.64 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 20.16 11.828 21.36 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 20.16 11.916 21.36 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 20.16 13.716 21.36 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 20.16 13.972 21.36 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 20.88 12.516 22.08 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 20.88 12.728 22.08 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 1.68 11.828 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 20.88 13.072 22.08 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 20.88 13.328 22.08 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 21.6 11.828 22.8 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 21.6 11.916 22.8 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 21.6 13.716 22.8 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 21.6 13.972 22.8 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 22.32 12.516 23.52 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 22.32 12.728 23.52 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 22.32 13.072 23.52 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 22.32 13.328 23.52 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 1.68 11.916 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 12.84 11.828 14.04 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 12.84 11.916 14.04 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 12.84 11.616 14.04 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 23.04 11.016 24.24 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 23.04 11.272 24.24 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 23.04 15.216 24.24 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 23.04 15.428 24.24 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 23.76 10.028 24.96 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 23.76 10.116 24.96 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 23.76 14.528 24.96 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.76 14.616 24.96 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 24.48 11.016 25.68 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 24.48 11.272 25.68 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 1.68 15.216 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 24.48 15.216 25.68 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 24.48 15.428 25.68 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 25.2 10.028 26.4 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 25.2 10.116 26.4 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 25.2 14.528 26.4 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 25.2 14.616 26.4 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 25.92 11.016 27.12 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 25.92 11.272 27.12 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 25.92 15.216 27.12 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 25.92 15.428 27.12 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 1.68 15.428 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 26.64 10.028 27.84 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 26.64 10.116 27.84 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 26.64 14.528 27.84 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 26.64 14.616 27.84 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 27.36 11.016 28.56 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 27.36 11.272 28.56 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 27.36 15.216 28.56 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 27.36 15.428 28.56 ;
    END
  END rddatap0[127]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 2.4 10.028 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 2.4 10.116 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 2.4 14.528 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 2.4 14.616 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 3.12 11.016 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 3.12 11.272 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 3.12 15.216 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 3.12 15.428 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 3.84 10.028 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 3.84 10.116 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 3.84 14.528 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.84 14.616 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 4.56 11.016 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 4.56 11.272 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 4.56 15.216 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.56 15.428 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 5.28 10.028 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 5.28 10.116 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 0.24 15.216 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 5.28 14.528 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 5.28 14.616 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 6 11.016 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 6 11.272 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 6 15.216 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6 15.428 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 6.72 10.028 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 6.72 10.116 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 6.72 14.528 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6.72 14.616 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 0.24 15.428 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 7.44 11.016 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 7.44 11.272 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 7.44 15.216 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 7.44 15.428 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 8.16 10.028 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.16 10.116 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 8.16 14.528 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.16 14.616 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 8.88 11.016 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 8.88 11.272 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.96 10.372 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 8.88 15.216 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.88 15.428 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 9.6 10.028 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 9.6 10.116 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 9.6 14.528 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 9.6 14.616 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 10.32 11.016 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 10.32 11.272 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 10.32 15.216 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 10.32 15.428 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 0.96 10.628 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 11.04 10.028 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 11.04 10.116 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 11.04 14.528 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 11.04 14.616 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 16.56 11.016 17.76 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 16.56 11.272 17.76 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 16.56 14.528 17.76 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 16.56 14.616 17.76 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 17.28 10.372 18.48 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 17.28 10.628 18.48 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 0.96 14.528 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 17.28 15.128 18.48 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 17.28 15.216 18.48 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 18 11.272 19.2 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 18 10.028 19.2 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 18 14.316 19.2 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 18 14.528 19.2 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 18.72 10.716 19.92 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 18.72 10.928 19.92 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 18.72 15.216 19.92 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 18.72 15.428 19.92 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 0.96 14.616 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 19.44 10.028 20.64 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 19.44 10.116 20.64 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 19.44 14.528 20.64 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 19.44 14.616 20.64 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 20.16 11.016 21.36 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 20.16 11.272 21.36 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 20.16 15.216 21.36 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 20.16 15.428 21.36 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 20.88 10.028 22.08 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 20.88 10.116 22.08 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 1.68 11.016 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 20.88 14.528 22.08 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 20.88 14.616 22.08 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 21.6 11.016 22.8 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 21.6 11.272 22.8 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 21.6 15.216 22.8 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 21.6 15.428 22.8 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 22.32 10.028 23.52 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 22.32 10.116 23.52 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 22.32 14.528 23.52 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 22.32 14.616 23.52 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 1.68 11.272 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 28.74 ;
        RECT 2.662 0.06 2.738 28.74 ;
        RECT 4.462 0.06 4.538 28.74 ;
        RECT 6.262 0.06 6.338 28.74 ;
        RECT 8.062 0.06 8.138 28.74 ;
        RECT 9.862 0.06 9.938 28.74 ;
        RECT 11.662 0.06 11.738 28.74 ;
        RECT 13.462 0.06 13.538 28.74 ;
        RECT 15.262 0.06 15.338 28.74 ;
        RECT 17.062 0.06 17.138 28.74 ;
        RECT 18.862 0.06 18.938 28.74 ;
        RECT 20.662 0.06 20.738 28.74 ;
        RECT 22.462 0.06 22.538 28.74 ;
        RECT 24.262 0.06 24.338 28.74 ;
        RECT 26.062 0.06 26.138 28.74 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 28.74 ;
        RECT 3.562 0.06 3.638 28.74 ;
        RECT 5.362 0.06 5.438 28.74 ;
        RECT 7.162 0.06 7.238 28.74 ;
        RECT 8.962 0.06 9.038 28.74 ;
        RECT 10.762 0.06 10.838 28.74 ;
        RECT 12.562 0.06 12.638 28.74 ;
        RECT 14.362 0.06 14.438 28.74 ;
        RECT 16.162 0.06 16.238 28.74 ;
        RECT 17.962 0.06 18.038 28.74 ;
        RECT 19.762 0.06 19.838 28.74 ;
        RECT 21.562 0.06 21.638 28.74 ;
        RECT 23.362 0.06 23.438 28.74 ;
        RECT 25.162 0.06 25.238 28.74 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 27.016 28.814 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 27.02 28.82 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 27.0705 28.838 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 27.035 28.87 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 27.07 28.838 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 27.059 28.89 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 27.09 28.862 ;
    LAYER m7 SPACING 0 ;
      RECT 26.138 28.86 27.04 28.92 ;
      RECT 26.138 -0.06 27.092 28.86 ;
      RECT 26.138 -0.12 27.04 -0.06 ;
      RECT 25.238 -0.12 26.062 28.92 ;
      RECT 24.338 -0.12 25.162 28.92 ;
      RECT 23.438 -0.12 24.262 28.92 ;
      RECT 22.538 -0.12 23.362 28.92 ;
      RECT 21.638 -0.12 22.462 28.92 ;
      RECT 20.738 -0.12 21.562 28.92 ;
      RECT 19.838 -0.12 20.662 28.92 ;
      RECT 18.938 -0.12 19.762 28.92 ;
      RECT 18.038 -0.12 18.862 28.92 ;
      RECT 17.138 -0.12 17.962 28.92 ;
      RECT 16.238 -0.12 17.062 28.92 ;
      RECT 15.338 28.56 16.162 28.92 ;
      RECT 15.338 27.36 15.384 28.56 ;
      RECT 15.428 27.36 16.162 28.56 ;
      RECT 15.338 27.12 16.162 27.36 ;
      RECT 15.338 25.92 15.384 27.12 ;
      RECT 15.428 25.92 16.162 27.12 ;
      RECT 15.338 25.68 16.162 25.92 ;
      RECT 15.338 24.48 15.384 25.68 ;
      RECT 15.428 24.48 16.162 25.68 ;
      RECT 15.338 24.24 16.162 24.48 ;
      RECT 15.338 23.04 15.384 24.24 ;
      RECT 15.428 23.04 16.162 24.24 ;
      RECT 15.338 22.8 16.162 23.04 ;
      RECT 15.338 21.6 15.384 22.8 ;
      RECT 15.428 21.6 16.162 22.8 ;
      RECT 15.338 21.36 16.162 21.6 ;
      RECT 15.338 20.16 15.384 21.36 ;
      RECT 15.428 20.16 16.162 21.36 ;
      RECT 15.338 19.92 16.162 20.16 ;
      RECT 15.338 18.72 15.384 19.92 ;
      RECT 15.428 18.72 16.162 19.92 ;
      RECT 15.338 15.96 16.162 18.72 ;
      RECT 15.338 14.76 15.384 15.96 ;
      RECT 15.428 14.76 15.472 15.96 ;
      RECT 15.516 14.76 16.162 15.96 ;
      RECT 15.338 11.52 16.162 14.76 ;
      RECT 15.338 10.32 15.384 11.52 ;
      RECT 15.428 10.32 16.162 11.52 ;
      RECT 15.338 10.08 16.162 10.32 ;
      RECT 15.338 8.88 15.384 10.08 ;
      RECT 15.428 8.88 16.162 10.08 ;
      RECT 15.338 8.64 16.162 8.88 ;
      RECT 15.338 7.44 15.384 8.64 ;
      RECT 15.428 7.44 16.162 8.64 ;
      RECT 15.338 7.2 16.162 7.44 ;
      RECT 15.338 6 15.384 7.2 ;
      RECT 15.428 6 16.162 7.2 ;
      RECT 15.338 5.76 16.162 6 ;
      RECT 15.338 4.56 15.384 5.76 ;
      RECT 15.428 4.56 16.162 5.76 ;
      RECT 15.338 4.32 16.162 4.56 ;
      RECT 15.338 3.12 15.384 4.32 ;
      RECT 15.428 3.12 16.162 4.32 ;
      RECT 15.338 2.88 16.162 3.12 ;
      RECT 15.338 1.68 15.384 2.88 ;
      RECT 15.428 1.68 16.162 2.88 ;
      RECT 15.338 1.44 16.162 1.68 ;
      RECT 15.338 0.24 15.384 1.44 ;
      RECT 15.428 0.24 16.162 1.44 ;
      RECT 15.338 -0.12 16.162 0.24 ;
      RECT 14.438 28.56 15.262 28.92 ;
      RECT 14.438 27.84 15.172 28.56 ;
      RECT 15.216 27.36 15.262 28.56 ;
      RECT 14.616 27.36 15.172 27.84 ;
      RECT 14.616 27.12 15.262 27.36 ;
      RECT 14.438 26.64 14.484 27.84 ;
      RECT 14.528 26.64 14.572 27.84 ;
      RECT 14.616 26.64 15.172 27.12 ;
      RECT 14.438 26.4 15.172 26.64 ;
      RECT 15.216 25.92 15.262 27.12 ;
      RECT 14.616 25.92 15.172 26.4 ;
      RECT 14.616 25.68 15.262 25.92 ;
      RECT 14.438 25.2 14.484 26.4 ;
      RECT 14.528 25.2 14.572 26.4 ;
      RECT 14.616 25.2 15.172 25.68 ;
      RECT 14.438 24.96 15.172 25.2 ;
      RECT 15.216 24.48 15.262 25.68 ;
      RECT 14.616 24.48 15.172 24.96 ;
      RECT 14.616 24.24 15.262 24.48 ;
      RECT 14.438 23.76 14.484 24.96 ;
      RECT 14.528 23.76 14.572 24.96 ;
      RECT 14.616 23.76 15.172 24.24 ;
      RECT 14.438 23.52 15.172 23.76 ;
      RECT 15.216 23.04 15.262 24.24 ;
      RECT 14.616 23.04 15.172 23.52 ;
      RECT 14.616 22.8 15.262 23.04 ;
      RECT 14.438 22.32 14.484 23.52 ;
      RECT 14.528 22.32 14.572 23.52 ;
      RECT 14.616 22.32 15.172 22.8 ;
      RECT 14.438 22.08 15.172 22.32 ;
      RECT 15.216 21.6 15.262 22.8 ;
      RECT 14.616 21.6 15.172 22.08 ;
      RECT 14.616 21.36 15.262 21.6 ;
      RECT 14.438 20.88 14.484 22.08 ;
      RECT 14.528 20.88 14.572 22.08 ;
      RECT 14.616 20.88 15.172 21.36 ;
      RECT 14.438 20.64 15.172 20.88 ;
      RECT 15.216 20.16 15.262 21.36 ;
      RECT 14.616 20.16 15.172 20.64 ;
      RECT 14.616 19.92 15.262 20.16 ;
      RECT 14.438 19.44 14.484 20.64 ;
      RECT 14.528 19.44 14.572 20.64 ;
      RECT 14.616 19.44 15.172 19.92 ;
      RECT 14.438 19.2 15.172 19.44 ;
      RECT 15.216 18.72 15.262 19.92 ;
      RECT 14.528 18.72 15.172 19.2 ;
      RECT 14.528 18.48 15.262 18.72 ;
      RECT 14.438 18 14.484 19.2 ;
      RECT 14.528 18 15.084 18.48 ;
      RECT 14.438 17.76 15.084 18 ;
      RECT 15.128 17.28 15.172 18.48 ;
      RECT 15.216 17.28 15.262 18.48 ;
      RECT 14.616 17.28 15.084 17.76 ;
      RECT 14.438 16.56 14.484 17.76 ;
      RECT 14.528 16.56 14.572 17.76 ;
      RECT 14.616 16.56 15.262 17.28 ;
      RECT 14.438 15.96 15.262 16.56 ;
      RECT 14.438 14.76 14.828 15.96 ;
      RECT 14.872 14.76 15.084 15.96 ;
      RECT 15.128 14.76 15.172 15.96 ;
      RECT 15.216 14.76 15.262 15.96 ;
      RECT 14.438 12.24 15.262 14.76 ;
      RECT 14.616 11.52 15.262 12.24 ;
      RECT 14.438 11.04 14.484 12.24 ;
      RECT 14.528 11.04 14.572 12.24 ;
      RECT 14.616 11.04 15.172 11.52 ;
      RECT 14.438 10.8 15.172 11.04 ;
      RECT 15.216 10.32 15.262 11.52 ;
      RECT 14.616 10.32 15.172 10.8 ;
      RECT 14.616 10.08 15.262 10.32 ;
      RECT 14.438 9.6 14.484 10.8 ;
      RECT 14.528 9.6 14.572 10.8 ;
      RECT 14.616 9.6 15.172 10.08 ;
      RECT 14.438 9.36 15.172 9.6 ;
      RECT 15.216 8.88 15.262 10.08 ;
      RECT 14.616 8.88 15.172 9.36 ;
      RECT 14.616 8.64 15.262 8.88 ;
      RECT 14.438 8.16 14.484 9.36 ;
      RECT 14.528 8.16 14.572 9.36 ;
      RECT 14.616 8.16 15.172 8.64 ;
      RECT 14.438 7.92 15.172 8.16 ;
      RECT 15.216 7.44 15.262 8.64 ;
      RECT 14.616 7.44 15.172 7.92 ;
      RECT 14.616 7.2 15.262 7.44 ;
      RECT 14.438 6.72 14.484 7.92 ;
      RECT 14.528 6.72 14.572 7.92 ;
      RECT 14.616 6.72 15.172 7.2 ;
      RECT 14.438 6.48 15.172 6.72 ;
      RECT 15.216 6 15.262 7.2 ;
      RECT 14.616 6 15.172 6.48 ;
      RECT 14.616 5.76 15.262 6 ;
      RECT 14.438 5.28 14.484 6.48 ;
      RECT 14.528 5.28 14.572 6.48 ;
      RECT 14.616 5.28 15.172 5.76 ;
      RECT 14.438 5.04 15.172 5.28 ;
      RECT 15.216 4.56 15.262 5.76 ;
      RECT 14.616 4.56 15.172 5.04 ;
      RECT 14.616 4.32 15.262 4.56 ;
      RECT 14.438 3.84 14.484 5.04 ;
      RECT 14.528 3.84 14.572 5.04 ;
      RECT 14.616 3.84 15.172 4.32 ;
      RECT 14.438 3.6 15.172 3.84 ;
      RECT 15.216 3.12 15.262 4.32 ;
      RECT 14.616 3.12 15.172 3.6 ;
      RECT 14.616 2.88 15.262 3.12 ;
      RECT 14.438 2.4 14.484 3.6 ;
      RECT 14.528 2.4 14.572 3.6 ;
      RECT 14.616 2.4 15.172 2.88 ;
      RECT 14.438 2.16 15.172 2.4 ;
      RECT 15.216 1.68 15.262 2.88 ;
      RECT 14.616 1.68 15.172 2.16 ;
      RECT 14.616 1.44 15.262 1.68 ;
      RECT 14.438 0.96 14.484 2.16 ;
      RECT 14.528 0.96 14.572 2.16 ;
      RECT 14.616 0.96 15.172 1.44 ;
      RECT 15.216 0.24 15.262 1.44 ;
      RECT 14.438 0.24 15.172 0.96 ;
      RECT 14.438 -0.12 15.262 0.24 ;
      RECT 13.538 28.56 14.362 28.92 ;
      RECT 13.538 27.36 13.672 28.56 ;
      RECT 13.716 27.36 13.928 28.56 ;
      RECT 13.972 27.36 14.362 28.56 ;
      RECT 13.538 27.12 14.362 27.36 ;
      RECT 13.538 25.92 13.672 27.12 ;
      RECT 13.716 25.92 13.928 27.12 ;
      RECT 13.972 25.92 14.362 27.12 ;
      RECT 13.538 25.68 14.362 25.92 ;
      RECT 13.538 24.48 13.672 25.68 ;
      RECT 13.716 24.48 13.928 25.68 ;
      RECT 13.972 24.48 14.362 25.68 ;
      RECT 13.538 24.24 14.362 24.48 ;
      RECT 13.538 23.04 13.672 24.24 ;
      RECT 13.716 23.04 13.928 24.24 ;
      RECT 13.972 23.04 14.362 24.24 ;
      RECT 13.538 22.8 14.362 23.04 ;
      RECT 13.538 21.6 13.672 22.8 ;
      RECT 13.716 21.6 13.928 22.8 ;
      RECT 13.972 21.6 14.362 22.8 ;
      RECT 13.538 21.36 14.362 21.6 ;
      RECT 13.538 20.16 13.672 21.36 ;
      RECT 13.716 20.16 13.928 21.36 ;
      RECT 13.972 20.16 14.362 21.36 ;
      RECT 13.538 19.92 14.362 20.16 ;
      RECT 13.716 19.2 14.362 19.92 ;
      RECT 13.538 18.72 13.584 19.92 ;
      RECT 13.628 18.72 13.672 19.92 ;
      RECT 13.716 18.72 13.928 19.2 ;
      RECT 13.538 18.48 13.928 18.72 ;
      RECT 13.972 18 14.272 19.2 ;
      RECT 14.316 18 14.362 19.2 ;
      RECT 13.716 18 13.928 18.48 ;
      RECT 13.538 17.28 13.584 18.48 ;
      RECT 13.628 17.28 13.672 18.48 ;
      RECT 13.716 17.28 14.362 18 ;
      RECT 13.538 15.96 14.362 17.28 ;
      RECT 13.538 14.76 13.928 15.96 ;
      RECT 13.972 14.76 14.184 15.96 ;
      RECT 14.228 14.76 14.272 15.96 ;
      RECT 14.316 14.76 14.362 15.96 ;
      RECT 13.538 14.04 14.362 14.76 ;
      RECT 13.538 12.84 13.584 14.04 ;
      RECT 13.628 12.84 13.672 14.04 ;
      RECT 13.716 12.84 14.362 14.04 ;
      RECT 13.538 11.52 14.362 12.84 ;
      RECT 13.538 10.32 13.672 11.52 ;
      RECT 13.716 10.32 13.928 11.52 ;
      RECT 13.972 10.32 14.362 11.52 ;
      RECT 13.538 10.08 14.362 10.32 ;
      RECT 13.538 8.88 13.672 10.08 ;
      RECT 13.716 8.88 13.928 10.08 ;
      RECT 13.972 8.88 14.362 10.08 ;
      RECT 13.538 8.64 14.362 8.88 ;
      RECT 13.538 7.44 13.672 8.64 ;
      RECT 13.716 7.44 13.928 8.64 ;
      RECT 13.972 7.44 14.362 8.64 ;
      RECT 13.538 7.2 14.362 7.44 ;
      RECT 13.538 6 13.672 7.2 ;
      RECT 13.716 6 13.928 7.2 ;
      RECT 13.972 6 14.362 7.2 ;
      RECT 13.538 5.76 14.362 6 ;
      RECT 13.538 4.56 13.672 5.76 ;
      RECT 13.716 4.56 13.928 5.76 ;
      RECT 13.972 4.56 14.362 5.76 ;
      RECT 13.538 4.32 14.362 4.56 ;
      RECT 13.538 3.12 13.672 4.32 ;
      RECT 13.716 3.12 13.928 4.32 ;
      RECT 13.972 3.12 14.362 4.32 ;
      RECT 13.538 2.88 14.362 3.12 ;
      RECT 13.538 1.68 13.672 2.88 ;
      RECT 13.716 1.68 13.928 2.88 ;
      RECT 13.972 1.68 14.362 2.88 ;
      RECT 13.538 1.44 14.362 1.68 ;
      RECT 13.538 0.24 13.672 1.44 ;
      RECT 13.716 0.24 13.928 1.44 ;
      RECT 13.972 0.24 14.362 1.44 ;
      RECT 13.538 -0.12 14.362 0.24 ;
      RECT 12.638 27.84 13.462 28.92 ;
      RECT 12.638 26.64 12.684 27.84 ;
      RECT 12.728 26.64 13.028 27.84 ;
      RECT 13.072 26.64 13.284 27.84 ;
      RECT 13.328 26.64 13.462 27.84 ;
      RECT 12.638 26.4 13.462 26.64 ;
      RECT 12.638 25.2 12.684 26.4 ;
      RECT 12.728 25.2 13.028 26.4 ;
      RECT 13.072 25.2 13.284 26.4 ;
      RECT 13.328 25.2 13.462 26.4 ;
      RECT 12.638 24.96 13.462 25.2 ;
      RECT 12.638 23.76 12.684 24.96 ;
      RECT 12.728 23.76 13.028 24.96 ;
      RECT 13.072 23.76 13.284 24.96 ;
      RECT 13.328 23.76 13.462 24.96 ;
      RECT 12.638 23.52 13.462 23.76 ;
      RECT 12.638 22.32 12.684 23.52 ;
      RECT 12.728 22.32 13.028 23.52 ;
      RECT 13.072 22.32 13.284 23.52 ;
      RECT 13.328 22.32 13.462 23.52 ;
      RECT 12.638 22.08 13.462 22.32 ;
      RECT 12.638 20.88 12.684 22.08 ;
      RECT 12.728 20.88 13.028 22.08 ;
      RECT 13.072 20.88 13.284 22.08 ;
      RECT 13.328 20.88 13.462 22.08 ;
      RECT 12.638 20.64 13.462 20.88 ;
      RECT 12.638 19.44 12.684 20.64 ;
      RECT 12.728 19.44 13.028 20.64 ;
      RECT 13.072 19.44 13.284 20.64 ;
      RECT 13.328 19.44 13.462 20.64 ;
      RECT 12.638 19.2 13.462 19.44 ;
      RECT 12.638 18 13.028 19.2 ;
      RECT 13.072 18 13.462 19.2 ;
      RECT 12.638 17.76 13.462 18 ;
      RECT 12.638 16.56 12.684 17.76 ;
      RECT 12.728 16.56 12.772 17.76 ;
      RECT 12.816 16.56 13.028 17.76 ;
      RECT 13.072 16.56 13.284 17.76 ;
      RECT 13.328 16.56 13.462 17.76 ;
      RECT 12.638 14.04 13.462 16.56 ;
      RECT 12.638 12.84 12.772 14.04 ;
      RECT 12.816 12.84 13.372 14.04 ;
      RECT 13.416 12.84 13.462 14.04 ;
      RECT 12.638 12.24 13.462 12.84 ;
      RECT 12.638 11.04 12.684 12.24 ;
      RECT 12.728 11.04 13.028 12.24 ;
      RECT 13.072 11.04 13.284 12.24 ;
      RECT 13.328 11.04 13.462 12.24 ;
      RECT 12.638 10.8 13.462 11.04 ;
      RECT 12.638 9.6 12.684 10.8 ;
      RECT 12.728 9.6 13.028 10.8 ;
      RECT 13.072 9.6 13.284 10.8 ;
      RECT 13.328 9.6 13.462 10.8 ;
      RECT 12.638 9.36 13.462 9.6 ;
      RECT 12.638 8.16 12.684 9.36 ;
      RECT 12.728 8.16 13.028 9.36 ;
      RECT 13.072 8.16 13.284 9.36 ;
      RECT 13.328 8.16 13.462 9.36 ;
      RECT 12.638 7.92 13.462 8.16 ;
      RECT 12.638 6.72 12.684 7.92 ;
      RECT 12.728 6.72 13.028 7.92 ;
      RECT 13.072 6.72 13.284 7.92 ;
      RECT 13.328 6.72 13.462 7.92 ;
      RECT 12.638 6.48 13.462 6.72 ;
      RECT 12.638 5.28 12.684 6.48 ;
      RECT 12.728 5.28 13.028 6.48 ;
      RECT 13.072 5.28 13.284 6.48 ;
      RECT 13.328 5.28 13.462 6.48 ;
      RECT 12.638 5.04 13.462 5.28 ;
      RECT 12.638 3.84 12.684 5.04 ;
      RECT 12.728 3.84 13.028 5.04 ;
      RECT 13.072 3.84 13.284 5.04 ;
      RECT 13.328 3.84 13.462 5.04 ;
      RECT 12.638 3.6 13.462 3.84 ;
      RECT 12.638 2.4 12.684 3.6 ;
      RECT 12.728 2.4 13.028 3.6 ;
      RECT 13.072 2.4 13.284 3.6 ;
      RECT 13.328 2.4 13.462 3.6 ;
      RECT 12.638 2.16 13.462 2.4 ;
      RECT 12.638 0.96 12.684 2.16 ;
      RECT 12.728 0.96 13.028 2.16 ;
      RECT 13.072 0.96 13.284 2.16 ;
      RECT 13.328 0.96 13.462 2.16 ;
      RECT 12.638 -0.12 13.462 0.96 ;
      RECT 11.738 28.56 12.562 28.92 ;
      RECT 11.916 27.84 12.562 28.56 ;
      RECT 11.738 27.36 11.784 28.56 ;
      RECT 11.828 27.36 11.872 28.56 ;
      RECT 11.916 27.36 12.472 27.84 ;
      RECT 11.738 27.12 12.472 27.36 ;
      RECT 12.516 26.64 12.562 27.84 ;
      RECT 11.916 26.64 12.472 27.12 ;
      RECT 11.916 26.4 12.562 26.64 ;
      RECT 11.738 25.92 11.784 27.12 ;
      RECT 11.828 25.92 11.872 27.12 ;
      RECT 11.916 25.92 12.472 26.4 ;
      RECT 11.738 25.68 12.472 25.92 ;
      RECT 12.516 25.2 12.562 26.4 ;
      RECT 11.916 25.2 12.472 25.68 ;
      RECT 11.916 24.96 12.562 25.2 ;
      RECT 11.738 24.48 11.784 25.68 ;
      RECT 11.828 24.48 11.872 25.68 ;
      RECT 11.916 24.48 12.472 24.96 ;
      RECT 11.738 24.24 12.472 24.48 ;
      RECT 12.516 23.76 12.562 24.96 ;
      RECT 11.916 23.76 12.472 24.24 ;
      RECT 11.916 23.52 12.562 23.76 ;
      RECT 11.738 23.04 11.784 24.24 ;
      RECT 11.828 23.04 11.872 24.24 ;
      RECT 11.916 23.04 12.472 23.52 ;
      RECT 11.738 22.8 12.472 23.04 ;
      RECT 12.516 22.32 12.562 23.52 ;
      RECT 11.916 22.32 12.472 22.8 ;
      RECT 11.916 22.08 12.562 22.32 ;
      RECT 11.738 21.6 11.784 22.8 ;
      RECT 11.828 21.6 11.872 22.8 ;
      RECT 11.916 21.6 12.472 22.08 ;
      RECT 11.738 21.36 12.472 21.6 ;
      RECT 12.516 20.88 12.562 22.08 ;
      RECT 11.916 20.88 12.472 21.36 ;
      RECT 11.916 20.64 12.562 20.88 ;
      RECT 11.738 20.16 11.784 21.36 ;
      RECT 11.828 20.16 11.872 21.36 ;
      RECT 11.916 20.16 12.472 20.64 ;
      RECT 11.738 19.92 12.472 20.16 ;
      RECT 12.516 19.44 12.562 20.64 ;
      RECT 11.916 19.44 12.472 19.92 ;
      RECT 11.916 19.2 12.562 19.44 ;
      RECT 11.738 18.72 11.784 19.92 ;
      RECT 11.828 18.72 11.872 19.92 ;
      RECT 11.916 18.72 12.128 19.2 ;
      RECT 12.428 18.48 12.562 19.2 ;
      RECT 11.738 18.48 12.128 18.72 ;
      RECT 12.172 18 12.384 19.2 ;
      RECT 11.828 18 12.128 18.48 ;
      RECT 12.428 18 12.472 18.48 ;
      RECT 11.738 17.28 11.784 18.48 ;
      RECT 12.516 17.28 12.562 18.48 ;
      RECT 11.828 17.28 12.472 18 ;
      RECT 11.738 14.04 12.562 17.28 ;
      RECT 11.738 12.84 11.784 14.04 ;
      RECT 11.828 12.84 11.872 14.04 ;
      RECT 11.916 12.84 12.128 14.04 ;
      RECT 12.172 12.84 12.384 14.04 ;
      RECT 12.428 12.84 12.562 14.04 ;
      RECT 11.738 12.24 12.562 12.84 ;
      RECT 11.738 11.52 12.472 12.24 ;
      RECT 12.516 11.04 12.562 12.24 ;
      RECT 11.916 11.04 12.472 11.52 ;
      RECT 11.916 10.8 12.562 11.04 ;
      RECT 11.738 10.32 11.784 11.52 ;
      RECT 11.828 10.32 11.872 11.52 ;
      RECT 11.916 10.32 12.472 10.8 ;
      RECT 11.738 10.08 12.472 10.32 ;
      RECT 12.516 9.6 12.562 10.8 ;
      RECT 11.916 9.6 12.472 10.08 ;
      RECT 11.916 9.36 12.562 9.6 ;
      RECT 11.738 8.88 11.784 10.08 ;
      RECT 11.828 8.88 11.872 10.08 ;
      RECT 11.916 8.88 12.472 9.36 ;
      RECT 11.738 8.64 12.472 8.88 ;
      RECT 12.516 8.16 12.562 9.36 ;
      RECT 11.916 8.16 12.472 8.64 ;
      RECT 11.916 7.92 12.562 8.16 ;
      RECT 11.738 7.44 11.784 8.64 ;
      RECT 11.828 7.44 11.872 8.64 ;
      RECT 11.916 7.44 12.472 7.92 ;
      RECT 11.738 7.2 12.472 7.44 ;
      RECT 12.516 6.72 12.562 7.92 ;
      RECT 11.916 6.72 12.472 7.2 ;
      RECT 11.916 6.48 12.562 6.72 ;
      RECT 11.738 6 11.784 7.2 ;
      RECT 11.828 6 11.872 7.2 ;
      RECT 11.916 6 12.472 6.48 ;
      RECT 11.738 5.76 12.472 6 ;
      RECT 12.516 5.28 12.562 6.48 ;
      RECT 11.916 5.28 12.472 5.76 ;
      RECT 11.916 5.04 12.562 5.28 ;
      RECT 11.738 4.56 11.784 5.76 ;
      RECT 11.828 4.56 11.872 5.76 ;
      RECT 11.916 4.56 12.472 5.04 ;
      RECT 11.738 4.32 12.472 4.56 ;
      RECT 12.516 3.84 12.562 5.04 ;
      RECT 11.916 3.84 12.472 4.32 ;
      RECT 11.916 3.6 12.562 3.84 ;
      RECT 11.738 3.12 11.784 4.32 ;
      RECT 11.828 3.12 11.872 4.32 ;
      RECT 11.916 3.12 12.472 3.6 ;
      RECT 11.738 2.88 12.472 3.12 ;
      RECT 12.516 2.4 12.562 3.6 ;
      RECT 11.916 2.4 12.472 2.88 ;
      RECT 11.916 2.16 12.562 2.4 ;
      RECT 11.738 1.68 11.784 2.88 ;
      RECT 11.828 1.68 11.872 2.88 ;
      RECT 11.916 1.68 12.472 2.16 ;
      RECT 11.738 1.44 12.472 1.68 ;
      RECT 12.516 0.96 12.562 2.16 ;
      RECT 12.428 0.96 12.472 1.44 ;
      RECT 11.738 0.24 12.128 1.44 ;
      RECT 12.172 0.24 12.384 1.44 ;
      RECT 12.428 0.24 12.562 0.96 ;
      RECT 11.738 -0.12 12.562 0.24 ;
      RECT 10.838 28.56 11.662 28.92 ;
      RECT 10.838 27.36 10.972 28.56 ;
      RECT 11.016 27.36 11.228 28.56 ;
      RECT 11.272 27.36 11.662 28.56 ;
      RECT 10.838 27.12 11.662 27.36 ;
      RECT 10.838 25.92 10.972 27.12 ;
      RECT 11.016 25.92 11.228 27.12 ;
      RECT 11.272 25.92 11.662 27.12 ;
      RECT 10.838 25.68 11.662 25.92 ;
      RECT 10.838 24.48 10.972 25.68 ;
      RECT 11.016 24.48 11.228 25.68 ;
      RECT 11.272 24.48 11.662 25.68 ;
      RECT 10.838 24.24 11.662 24.48 ;
      RECT 10.838 23.04 10.972 24.24 ;
      RECT 11.016 23.04 11.228 24.24 ;
      RECT 11.272 23.04 11.662 24.24 ;
      RECT 10.838 22.8 11.662 23.04 ;
      RECT 10.838 21.6 10.972 22.8 ;
      RECT 11.016 21.6 11.228 22.8 ;
      RECT 11.272 21.6 11.662 22.8 ;
      RECT 10.838 21.36 11.662 21.6 ;
      RECT 10.838 20.16 10.972 21.36 ;
      RECT 11.016 20.16 11.228 21.36 ;
      RECT 11.272 20.16 11.662 21.36 ;
      RECT 10.838 19.92 11.662 20.16 ;
      RECT 10.928 19.2 11.662 19.92 ;
      RECT 10.838 18.72 10.884 19.92 ;
      RECT 10.928 18.72 11.228 19.2 ;
      RECT 11.272 18 11.662 19.2 ;
      RECT 10.838 18 11.228 18.72 ;
      RECT 10.838 17.76 11.662 18 ;
      RECT 10.838 16.56 10.972 17.76 ;
      RECT 11.016 16.56 11.228 17.76 ;
      RECT 11.272 16.56 11.662 17.76 ;
      RECT 10.838 14.04 11.662 16.56 ;
      RECT 10.838 12.84 10.972 14.04 ;
      RECT 11.016 12.84 11.228 14.04 ;
      RECT 11.272 12.84 11.484 14.04 ;
      RECT 11.528 12.84 11.572 14.04 ;
      RECT 11.616 12.84 11.662 14.04 ;
      RECT 10.838 11.52 11.662 12.84 ;
      RECT 10.838 10.32 10.972 11.52 ;
      RECT 11.016 10.32 11.228 11.52 ;
      RECT 11.272 10.32 11.662 11.52 ;
      RECT 10.838 10.08 11.662 10.32 ;
      RECT 10.838 8.88 10.972 10.08 ;
      RECT 11.016 8.88 11.228 10.08 ;
      RECT 11.272 8.88 11.662 10.08 ;
      RECT 10.838 8.64 11.662 8.88 ;
      RECT 10.838 7.44 10.972 8.64 ;
      RECT 11.016 7.44 11.228 8.64 ;
      RECT 11.272 7.44 11.662 8.64 ;
      RECT 10.838 7.2 11.662 7.44 ;
      RECT 10.838 6 10.972 7.2 ;
      RECT 11.016 6 11.228 7.2 ;
      RECT 11.272 6 11.662 7.2 ;
      RECT 10.838 5.76 11.662 6 ;
      RECT 10.838 4.56 10.972 5.76 ;
      RECT 11.016 4.56 11.228 5.76 ;
      RECT 11.272 4.56 11.662 5.76 ;
      RECT 10.838 4.32 11.662 4.56 ;
      RECT 10.838 3.12 10.972 4.32 ;
      RECT 11.016 3.12 11.228 4.32 ;
      RECT 11.272 3.12 11.662 4.32 ;
      RECT 10.838 2.88 11.662 3.12 ;
      RECT 10.838 1.68 10.972 2.88 ;
      RECT 11.016 1.68 11.228 2.88 ;
      RECT 11.272 1.68 11.662 2.88 ;
      RECT 10.838 -0.12 11.662 1.68 ;
      RECT 9.938 27.84 10.762 28.92 ;
      RECT 9.938 26.64 9.984 27.84 ;
      RECT 10.028 26.64 10.072 27.84 ;
      RECT 10.116 26.64 10.762 27.84 ;
      RECT 9.938 26.4 10.762 26.64 ;
      RECT 9.938 25.2 9.984 26.4 ;
      RECT 10.028 25.2 10.072 26.4 ;
      RECT 10.116 25.2 10.762 26.4 ;
      RECT 9.938 24.96 10.762 25.2 ;
      RECT 9.938 23.76 9.984 24.96 ;
      RECT 10.028 23.76 10.072 24.96 ;
      RECT 10.116 23.76 10.762 24.96 ;
      RECT 9.938 23.52 10.762 23.76 ;
      RECT 9.938 22.32 9.984 23.52 ;
      RECT 10.028 22.32 10.072 23.52 ;
      RECT 10.116 22.32 10.762 23.52 ;
      RECT 9.938 22.08 10.762 22.32 ;
      RECT 9.938 20.88 9.984 22.08 ;
      RECT 10.028 20.88 10.072 22.08 ;
      RECT 10.116 20.88 10.762 22.08 ;
      RECT 9.938 20.64 10.762 20.88 ;
      RECT 10.116 19.92 10.762 20.64 ;
      RECT 9.938 19.44 9.984 20.64 ;
      RECT 10.028 19.44 10.072 20.64 ;
      RECT 10.116 19.44 10.672 19.92 ;
      RECT 9.938 19.2 10.672 19.44 ;
      RECT 10.716 18.72 10.762 19.92 ;
      RECT 10.028 18.72 10.672 19.2 ;
      RECT 10.028 18.48 10.762 18.72 ;
      RECT 9.938 18 9.984 19.2 ;
      RECT 10.028 18 10.328 18.48 ;
      RECT 10.372 17.28 10.584 18.48 ;
      RECT 10.628 17.28 10.762 18.48 ;
      RECT 9.938 17.28 10.328 18 ;
      RECT 9.938 15.96 10.762 17.28 ;
      RECT 9.938 14.76 10.328 15.96 ;
      RECT 10.372 14.76 10.584 15.96 ;
      RECT 10.628 14.76 10.672 15.96 ;
      RECT 10.716 14.76 10.762 15.96 ;
      RECT 9.938 12.24 10.762 14.76 ;
      RECT 9.938 11.04 9.984 12.24 ;
      RECT 10.028 11.04 10.072 12.24 ;
      RECT 10.116 11.04 10.762 12.24 ;
      RECT 9.938 10.8 10.762 11.04 ;
      RECT 9.938 9.6 9.984 10.8 ;
      RECT 10.028 9.6 10.072 10.8 ;
      RECT 10.116 9.6 10.762 10.8 ;
      RECT 9.938 9.36 10.762 9.6 ;
      RECT 9.938 8.16 9.984 9.36 ;
      RECT 10.028 8.16 10.072 9.36 ;
      RECT 10.116 8.16 10.762 9.36 ;
      RECT 9.938 7.92 10.762 8.16 ;
      RECT 9.938 6.72 9.984 7.92 ;
      RECT 10.028 6.72 10.072 7.92 ;
      RECT 10.116 6.72 10.762 7.92 ;
      RECT 9.938 6.48 10.762 6.72 ;
      RECT 9.938 5.28 9.984 6.48 ;
      RECT 10.028 5.28 10.072 6.48 ;
      RECT 10.116 5.28 10.762 6.48 ;
      RECT 9.938 5.04 10.762 5.28 ;
      RECT 9.938 3.84 9.984 5.04 ;
      RECT 10.028 3.84 10.072 5.04 ;
      RECT 10.116 3.84 10.762 5.04 ;
      RECT 9.938 3.6 10.762 3.84 ;
      RECT 9.938 2.4 9.984 3.6 ;
      RECT 10.028 2.4 10.072 3.6 ;
      RECT 10.116 2.4 10.762 3.6 ;
      RECT 9.938 2.16 10.762 2.4 ;
      RECT 9.938 1.44 10.328 2.16 ;
      RECT 10.372 0.96 10.584 2.16 ;
      RECT 10.628 0.96 10.762 2.16 ;
      RECT 10.116 0.96 10.328 1.44 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.762 0.96 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 28.92 ;
      RECT 8.138 -0.12 8.962 28.92 ;
      RECT 7.238 -0.12 8.062 28.92 ;
      RECT 6.338 -0.12 7.162 28.92 ;
      RECT 5.438 -0.12 6.262 28.92 ;
      RECT 4.538 -0.12 5.362 28.92 ;
      RECT 3.638 -0.12 4.462 28.92 ;
      RECT 2.738 -0.12 3.562 28.92 ;
      RECT 1.838 -0.12 2.662 28.92 ;
      RECT 0.938 -0.12 1.762 28.92 ;
      RECT -0.04 28.86 0.862 28.92 ;
      RECT -0.092 -0.06 0.862 28.86 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 26.258 0 26.92 28.8 ;
      RECT 25.358 0 25.942 28.8 ;
      RECT 24.458 0 25.042 28.8 ;
      RECT 23.558 0 24.142 28.8 ;
      RECT 22.658 0 23.242 28.8 ;
      RECT 21.758 0 22.342 28.8 ;
      RECT 20.858 0 21.442 28.8 ;
      RECT 19.958 0 20.542 28.8 ;
      RECT 19.058 0 19.642 28.8 ;
      RECT 18.158 0 18.742 28.8 ;
      RECT 17.258 0 17.842 28.8 ;
      RECT 16.358 0 16.942 28.8 ;
      RECT 15.458 28.68 16.042 28.8 ;
      RECT 15.548 18.6 16.042 28.68 ;
      RECT 15.458 16.08 16.042 18.6 ;
      RECT 15.636 14.64 16.042 16.08 ;
      RECT 15.458 11.64 16.042 14.64 ;
      RECT 15.548 0.12 16.042 11.64 ;
      RECT 15.458 0 16.042 0.12 ;
      RECT 14.558 28.68 15.142 28.8 ;
      RECT 14.558 27.96 15.052 28.68 ;
      RECT 14.736 19.32 15.052 27.96 ;
      RECT 14.648 18.6 15.052 19.32 ;
      RECT 14.648 17.88 14.964 18.6 ;
      RECT 14.736 17.16 14.964 17.88 ;
      RECT 14.736 16.44 15.142 17.16 ;
      RECT 14.558 16.08 15.142 16.44 ;
      RECT 14.558 14.64 14.708 16.08 ;
      RECT 14.558 12.36 15.142 14.64 ;
      RECT 14.736 11.64 15.142 12.36 ;
      RECT 14.736 0.84 15.052 11.64 ;
      RECT 14.558 0.12 15.052 0.84 ;
      RECT 14.558 0 15.142 0.12 ;
      RECT 13.658 28.68 14.242 28.8 ;
      RECT 14.092 20.04 14.242 28.68 ;
      RECT 13.836 19.32 14.242 20.04 ;
      RECT 14.092 17.88 14.152 19.32 ;
      RECT 13.836 17.16 14.242 17.88 ;
      RECT 13.658 16.08 14.242 17.16 ;
      RECT 13.658 14.64 13.808 16.08 ;
      RECT 13.658 14.16 14.242 14.64 ;
      RECT 13.836 12.72 14.242 14.16 ;
      RECT 13.658 11.64 14.242 12.72 ;
      RECT 14.092 0.12 14.242 11.64 ;
      RECT 13.658 0 14.242 0.12 ;
      RECT 12.758 27.96 13.342 28.8 ;
      RECT 12.848 19.32 12.908 27.96 ;
      RECT 12.758 17.88 12.908 19.32 ;
      RECT 11.858 28.68 12.442 28.8 ;
      RECT 12.036 27.96 12.442 28.68 ;
      RECT 12.036 19.32 12.352 27.96 ;
      RECT 10.958 28.68 11.542 28.8 ;
      RECT 11.392 20.04 11.542 28.68 ;
      RECT 11.048 19.32 11.542 20.04 ;
      RECT 11.048 18.6 11.108 19.32 ;
      RECT 10.958 17.88 11.108 18.6 ;
      RECT 11.392 16.44 11.542 19.32 ;
      RECT 10.958 14.16 11.542 16.44 ;
      RECT 10.058 27.96 10.642 28.8 ;
      RECT 10.236 20.04 10.642 27.96 ;
      RECT 10.236 19.32 10.552 20.04 ;
      RECT 10.148 18.6 10.552 19.32 ;
      RECT 10.148 17.88 10.208 18.6 ;
      RECT 10.058 17.16 10.208 17.88 ;
      RECT 10.058 16.08 10.642 17.16 ;
      RECT 10.058 14.64 10.208 16.08 ;
      RECT 10.058 12.36 10.642 14.64 ;
      RECT 10.236 2.28 10.642 12.36 ;
      RECT 9.158 0 9.742 28.8 ;
      RECT 8.258 0 8.842 28.8 ;
      RECT 7.358 0 7.942 28.8 ;
      RECT 6.458 0 7.042 28.8 ;
      RECT 5.558 0 6.142 28.8 ;
      RECT 4.658 0 5.242 28.8 ;
      RECT 3.758 0 4.342 28.8 ;
      RECT 2.858 0 3.442 28.8 ;
      RECT 1.958 0 2.542 28.8 ;
      RECT 1.058 0 1.642 28.8 ;
      RECT 0.08 0 0.742 28.8 ;
      RECT 13.192 17.88 13.342 19.32 ;
      RECT 11.948 17.88 12.008 18.6 ;
      RECT 11.948 17.16 12.352 17.88 ;
      RECT 11.858 14.16 12.442 17.16 ;
      RECT 12.758 14.16 13.342 16.44 ;
      RECT 12.936 12.72 13.252 14.16 ;
      RECT 12.758 12.36 13.342 12.72 ;
      RECT 12.848 0.84 12.908 12.36 ;
      RECT 12.758 0 13.342 0.84 ;
      RECT 11.858 12.36 12.442 12.72 ;
      RECT 11.858 11.64 12.352 12.36 ;
      RECT 12.036 1.56 12.352 11.64 ;
      RECT 10.958 11.64 11.542 12.72 ;
      RECT 11.392 1.56 11.542 11.64 ;
      RECT 10.958 0 11.542 1.56 ;
      RECT 10.058 1.56 10.208 2.28 ;
      RECT 11.858 0.12 12.008 1.56 ;
      RECT 11.858 0 12.442 0.12 ;
      RECT 10.236 0.12 10.642 0.84 ;
      RECT 10.058 0 10.642 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 27 28.798 ;
    LAYER m1 ;
      RECT 0 0 27 28.8 ;
    LAYER m2 ;
      RECT 0 0.015 27 28.785 ;
    LAYER m3 ;
      RECT 0.015 0 26.985 28.8 ;
    LAYER m4 ;
      RECT 0 0.02 27 28.78 ;
    LAYER m5 ;
      RECT 0.012 0 26.988 28.8 ;
    LAYER m6 ;
      RECT 0 0.012 27 28.788 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf124b064e1r1w0cbbehbaa4acw

END LIBRARY
