#############################################################################################
## Intel Confidential                                                                      ##
#############################################################################################
## Copyright 2023 Intel Corporation. The information contained herein is the proprietary   ##
## and confidential information of Intel or its licensors, and is supplied subject to, and ##
## may be used only in accordance with, previously executed agreements with Intel.         ##
## EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING: (1) ALL MATERIALS FURNISHED BY INTEL      ##
## HEREUNDER ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY KIND; (2) INTEL SPECIFICALLY     ##
## DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS FOR A PARTICULAR PURPOSE OR          ##
## MERCHANTABILITY; AND (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF       ##
## SUBSTITUTES, LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR FOR ANY OTHER SPECIAL,       ##
## CONSEQUENTIAL OR INCIDENTAL DAMAGES, HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY,    ##
## CONTRACT, TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                              ##
#############################################################################################
#############################################################################################
##                                                                                         ##
##  Vendor:                Intel Corporation                                               ##
##  Product:               c764hduspsr                                                     ##
##  Version:               r1.0.0                                                          ##
##  Technology:            p1276.4                                                         ##
##  Celltype:              MemoryIP                                                        ##
##  IP Owner:              Intel CMO                                                       ##
##  Creation Time:         Tue Mar 28 2023 19:06:49                                        ##
##  Memory Name:           ip764hduspsr2048x39m8b2s0r2p0d0                                 ##
##  Memory Name Generated: ip764hduspsr2048x39m8b2s0r2p0d0                                 ##
##                                                                                         ##
#############################################################################################

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 4000 ;
END UNITS
SITE ip764hduspsr2048x39m8b2s0r2p0d0
  SIZE 36.3 by 105.12 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END ip764hduspsr2048x39m8b2s0r2p0d0


MACRO ip764hduspsr2048x39m8b2s0r2p0d0
     FIXEDMASK ;
     FOREIGN ip764hduspsr2048x39m8b2s0r2p0d0 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 36.3 by 105.12 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE ip764hduspsr2048x39m8b2s0r2p0d0 ;
     PIN q[0]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 0.62 17.176 1.78 ;
               LAYER v4 ;
               RECT 17.136 1.329 17.176 1.365 ;
          END
     END q[0]
     PIN din[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 0.62 17.452 1.78 ;
               LAYER v4 ;
               RECT 17.412 1.558 17.452 1.594 ;
          END
     END din[0]
     PIN q[1]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 3.02 17.176 4.18 ;
               LAYER v4 ;
               RECT 17.136 3.729 17.176 3.765 ;
          END
     END q[1]
     PIN din[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 3.02 17.452 4.18 ;
               LAYER v4 ;
               RECT 17.412 3.958 17.452 3.994 ;
          END
     END din[1]
     PIN q[2]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 5.42 17.176 6.58 ;
               LAYER v4 ;
               RECT 17.136 6.129 17.176 6.165 ;
          END
     END q[2]
     PIN din[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 5.42 17.452 6.58 ;
               LAYER v4 ;
               RECT 17.412 6.358 17.452 6.394 ;
          END
     END din[2]
     PIN q[3]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 7.82 17.176 8.98 ;
               LAYER v4 ;
               RECT 17.136 8.529 17.176 8.565 ;
          END
     END q[3]
     PIN din[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 7.82 17.452 8.98 ;
               LAYER v4 ;
               RECT 17.412 8.758 17.452 8.794 ;
          END
     END din[3]
     PIN q[4]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 10.22 17.176 11.38 ;
               LAYER v4 ;
               RECT 17.136 10.929 17.176 10.965 ;
          END
     END q[4]
     PIN din[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 10.22 17.452 11.38 ;
               LAYER v4 ;
               RECT 17.412 11.158 17.452 11.194 ;
          END
     END din[4]
     PIN q[5]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 12.62 17.176 13.78 ;
               LAYER v4 ;
               RECT 17.136 13.329 17.176 13.365 ;
          END
     END q[5]
     PIN din[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 12.62 17.452 13.78 ;
               LAYER v4 ;
               RECT 17.412 13.558 17.452 13.594 ;
          END
     END din[5]
     PIN q[6]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 15.02 17.176 16.18 ;
               LAYER v4 ;
               RECT 17.136 15.729 17.176 15.765 ;
          END
     END q[6]
     PIN din[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 15.02 17.452 16.18 ;
               LAYER v4 ;
               RECT 17.412 15.958 17.452 15.994 ;
          END
     END din[6]
     PIN q[7]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 17.42 17.176 18.58 ;
               LAYER v4 ;
               RECT 17.136 18.129 17.176 18.165 ;
          END
     END q[7]
     PIN din[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 17.42 17.452 18.58 ;
               LAYER v4 ;
               RECT 17.412 18.358 17.452 18.394 ;
          END
     END din[7]
     PIN q[8]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 19.82 17.176 20.98 ;
               LAYER v4 ;
               RECT 17.136 20.529 17.176 20.565 ;
          END
     END q[8]
     PIN din[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 19.82 17.452 20.98 ;
               LAYER v4 ;
               RECT 17.412 20.758 17.452 20.794 ;
          END
     END din[8]
     PIN q[9]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 22.22 17.176 23.38 ;
               LAYER v4 ;
               RECT 17.136 22.929 17.176 22.965 ;
          END
     END q[9]
     PIN din[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 22.22 17.452 23.38 ;
               LAYER v4 ;
               RECT 17.412 23.158 17.452 23.194 ;
          END
     END din[9]
     PIN q[10]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 24.62 17.176 25.78 ;
               LAYER v4 ;
               RECT 17.136 25.329 17.176 25.365 ;
          END
     END q[10]
     PIN din[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 24.62 17.452 25.78 ;
               LAYER v4 ;
               RECT 17.412 25.558 17.452 25.594 ;
          END
     END din[10]
     PIN q[11]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 27.02 17.176 28.18 ;
               LAYER v4 ;
               RECT 17.136 27.729 17.176 27.765 ;
          END
     END q[11]
     PIN din[11]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 27.02 17.452 28.18 ;
               LAYER v4 ;
               RECT 17.412 27.958 17.452 27.994 ;
          END
     END din[11]
     PIN q[12]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 29.42 17.176 30.58 ;
               LAYER v4 ;
               RECT 17.136 30.129 17.176 30.165 ;
          END
     END q[12]
     PIN din[12]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 29.42 17.452 30.58 ;
               LAYER v4 ;
               RECT 17.412 30.358 17.452 30.394 ;
          END
     END din[12]
     PIN q[13]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 31.82 17.176 32.98 ;
               LAYER v4 ;
               RECT 17.136 32.529 17.176 32.565 ;
          END
     END q[13]
     PIN din[13]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 31.82 17.452 32.98 ;
               LAYER v4 ;
               RECT 17.412 32.758 17.452 32.794 ;
          END
     END din[13]
     PIN q[14]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 34.22 17.176 35.38 ;
               LAYER v4 ;
               RECT 17.136 34.929 17.176 34.965 ;
          END
     END q[14]
     PIN din[14]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 34.22 17.452 35.38 ;
               LAYER v4 ;
               RECT 17.412 35.158 17.452 35.194 ;
          END
     END din[14]
     PIN q[15]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 36.62 17.176 37.78 ;
               LAYER v4 ;
               RECT 17.136 37.329 17.176 37.365 ;
          END
     END q[15]
     PIN din[15]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 36.62 17.452 37.78 ;
               LAYER v4 ;
               RECT 17.412 37.558 17.452 37.594 ;
          END
     END din[15]
     PIN q[16]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 39.02 17.176 40.18 ;
               LAYER v4 ;
               RECT 17.136 39.729 17.176 39.765 ;
          END
     END q[16]
     PIN din[16]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 39.02 17.452 40.18 ;
               LAYER v4 ;
               RECT 17.412 39.958 17.452 39.994 ;
          END
     END din[16]
     PIN q[17]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 41.42 17.176 42.58 ;
               LAYER v4 ;
               RECT 17.136 42.129 17.176 42.165 ;
          END
     END q[17]
     PIN din[17]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 41.42 17.452 42.58 ;
               LAYER v4 ;
               RECT 17.412 42.358 17.452 42.394 ;
          END
     END din[17]
     PIN q[18]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 43.82 17.176 44.98 ;
               LAYER v4 ;
               RECT 17.136 44.529 17.176 44.565 ;
          END
     END q[18]
     PIN din[18]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 43.82 17.452 44.98 ;
               LAYER v4 ;
               RECT 17.412 44.758 17.452 44.794 ;
          END
     END din[18]
     PIN q[19]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 46.22 17.176 47.38 ;
               LAYER v4 ;
               RECT 17.136 46.929 17.176 46.965 ;
          END
     END q[19]
     PIN din[19]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 46.22 17.452 47.38 ;
               LAYER v4 ;
               RECT 17.412 47.158 17.452 47.194 ;
          END
     END din[19]
     PIN arysleep
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.344 48.98 17.384 49.94 ;
               LAYER v4 ;
               RECT 17.344 49.0005 17.384 49.0365 ;
          END
     END arysleep
     PIN sbc[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.548 48.98 17.588 49.94 ;
               LAYER v4 ;
               RECT 17.548 49.2405 17.588 49.2765 ;
          END
     END sbc[1]
     PIN async_reset
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 48.98 17.656 49.94 ;
               LAYER v4 ;
               RECT 17.616 49.1235 17.656 49.1595 ;
          END
     END async_reset
     PIN sbc[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.284 48.98 18.328 49.94 ;
               LAYER v4 ;
               RECT 18.284 49.062 18.328 49.098 ;
          END
     END sbc[0]
     PIN wen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.272 49.98 17.316 50.94 ;
               LAYER v4 ;
               RECT 17.272 50.5635 17.316 50.5995 ;
          END
     END wen
     PIN adr[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 49.98 17.656 50.94 ;
               LAYER v4 ;
               RECT 17.616 50.2005 17.656 50.2365 ;
          END
     END adr[2]
     PIN adr[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.944 49.98 17.984 50.94 ;
               LAYER v4 ;
               RECT 17.944 50.022 17.984 50.058 ;
          END
     END adr[7]
     PIN redrowen[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.012 49.98 18.052 50.94 ;
               LAYER v4 ;
               RECT 18.012 50.262 18.052 50.298 ;
          END
     END redrowen[1]
     PIN adr[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.284 49.98 18.328 50.94 ;
               LAYER v4 ;
               RECT 18.284 50.742 18.328 50.778 ;
          END
     END adr[5]
     PIN adr[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 50.1 17.176 51.06 ;
               LAYER v4 ;
               RECT 17.136 50.742 17.176 50.778 ;
          END
     END adr[6]
     PIN adr[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.48 50.1 17.52 51.06 ;
               LAYER v4 ;
               RECT 17.48 50.8035 17.52 50.8395 ;
          END
     END adr[3]
     PIN ren
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.064 50.98 17.108 51.94 ;
               LAYER v4 ;
               RECT 17.064 51.222 17.108 51.258 ;
          END
     END ren
     PIN adr[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.272 50.98 17.316 51.94 ;
               LAYER v4 ;
               RECT 17.272 51.0435 17.316 51.0795 ;
          END
     END adr[9]
     PIN adr[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.344 50.98 17.384 51.94 ;
               LAYER v4 ;
               RECT 17.344 51.702 17.384 51.738 ;
          END
     END adr[0]
     PIN adr[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 50.98 17.656 51.94 ;
               LAYER v4 ;
               RECT 17.616 51.1605 17.656 51.1965 ;
          END
     END adr[10]
     PIN stbyp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.012 50.98 18.052 51.94 ;
               LAYER v4 ;
               RECT 18.012 51.462 18.052 51.498 ;
          END
     END stbyp
     PIN adr[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.284 50.98 18.328 51.94 ;
               LAYER v4 ;
               RECT 18.284 51.702 18.328 51.738 ;
          END
     END adr[8]
     PIN adr[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 51.1 17.176 52.06 ;
               LAYER v4 ;
               RECT 17.136 51.702 17.176 51.738 ;
          END
     END adr[4]
     PIN adr[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.48 51.1 17.52 52.06 ;
               LAYER v4 ;
               RECT 17.48 51.4005 17.52 51.4365 ;
          END
     END adr[1]
     PIN wa[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.344 52.65 17.384 53.61 ;
               LAYER v4 ;
               RECT 17.344 53.142 17.384 53.178 ;
          END
     END wa[1]
     PIN redrowen[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 52.65 17.656 53.61 ;
               LAYER v4 ;
               RECT 17.616 52.902 17.656 52.938 ;
          END
     END redrowen[0]
     PIN wpulse[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 53.65 17.176 54.61 ;
               LAYER v4 ;
               RECT 17.136 54.0405 17.176 54.0765 ;
          END
     END wpulse[1]
     PIN wmce[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.344 53.65 17.384 54.61 ;
               LAYER v4 ;
               RECT 17.344 53.6835 17.384 53.7195 ;
          END
     END wmce[1]
     PIN wpulse[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.548 53.65 17.588 54.61 ;
               LAYER v4 ;
               RECT 17.548 54.2805 17.588 54.3165 ;
          END
     END wpulse[0]
     PIN wa[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 53.65 17.656 54.61 ;
               LAYER v4 ;
               RECT 17.616 54.102 17.656 54.138 ;
          END
     END wa[0]
     PIN wpulse[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.944 53.65 17.984 54.61 ;
               LAYER v4 ;
               RECT 17.944 54.0405 17.984 54.0765 ;
          END
     END wpulse[2]
     PIN ra[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.012 53.65 18.052 54.61 ;
               LAYER v4 ;
               RECT 18.012 54.342 18.052 54.378 ;
          END
     END ra[1]
     PIN wa[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.08 53.65 18.12 54.61 ;
               LAYER v4 ;
               RECT 18.08 53.6835 18.12 53.7195 ;
          END
     END wa[2]
     PIN ra[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 18.424 53.65 18.464 54.61 ;
               LAYER v4 ;
               RECT 18.424 54.5205 18.464 54.5565 ;
          END
     END ra[0]
     PIN wmce[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.48 53.77 17.52 54.73 ;
               LAYER v4 ;
               RECT 17.48 54.1635 17.52 54.1995 ;
          END
     END wmce[0]
     PIN mce
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 54.65 17.176 55.61 ;
               LAYER v4 ;
               RECT 17.136 54.822 17.176 54.858 ;
          END
     END mce
     PIN rmce[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.344 54.65 17.384 55.61 ;
               LAYER v4 ;
               RECT 17.344 54.7605 17.384 54.7965 ;
          END
     END rmce[2]
     PIN rmce[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.548 54.65 17.588 55.61 ;
               LAYER v4 ;
               RECT 17.548 55.0005 17.588 55.0365 ;
          END
     END rmce[1]
     PIN rmce[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.616 54.65 17.656 55.61 ;
               LAYER v4 ;
               RECT 17.616 55.302 17.656 55.338 ;
          END
     END rmce[0]
     PIN rmce[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.48 54.77 17.52 55.73 ;
               LAYER v4 ;
               RECT 17.48 55.1235 17.52 55.1595 ;
          END
     END rmce[3]
     PIN q[20]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 56.54 17.176 57.7 ;
               LAYER v4 ;
               RECT 17.136 57.249 17.176 57.285 ;
          END
     END q[20]
     PIN din[20]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 56.54 17.452 57.7 ;
               LAYER v4 ;
               RECT 17.412 57.478 17.452 57.514 ;
          END
     END din[20]
     PIN q[21]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 58.94 17.176 60.1 ;
               LAYER v4 ;
               RECT 17.136 59.649 17.176 59.685 ;
          END
     END q[21]
     PIN din[21]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 58.94 17.452 60.1 ;
               LAYER v4 ;
               RECT 17.412 59.878 17.452 59.914 ;
          END
     END din[21]
     PIN q[22]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 61.34 17.176 62.5 ;
               LAYER v4 ;
               RECT 17.136 62.049 17.176 62.085 ;
          END
     END q[22]
     PIN din[22]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 61.34 17.452 62.5 ;
               LAYER v4 ;
               RECT 17.412 62.278 17.452 62.314 ;
          END
     END din[22]
     PIN q[23]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 63.74 17.176 64.9 ;
               LAYER v4 ;
               RECT 17.136 64.449 17.176 64.485 ;
          END
     END q[23]
     PIN din[23]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 63.74 17.452 64.9 ;
               LAYER v4 ;
               RECT 17.412 64.678 17.452 64.714 ;
          END
     END din[23]
     PIN q[24]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 66.14 17.176 67.3 ;
               LAYER v4 ;
               RECT 17.136 66.849 17.176 66.885 ;
          END
     END q[24]
     PIN din[24]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 66.14 17.452 67.3 ;
               LAYER v4 ;
               RECT 17.412 67.078 17.452 67.114 ;
          END
     END din[24]
     PIN q[25]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 68.54 17.176 69.7 ;
               LAYER v4 ;
               RECT 17.136 69.249 17.176 69.285 ;
          END
     END q[25]
     PIN din[25]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 68.54 17.452 69.7 ;
               LAYER v4 ;
               RECT 17.412 69.478 17.452 69.514 ;
          END
     END din[25]
     PIN q[26]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 70.94 17.176 72.1 ;
               LAYER v4 ;
               RECT 17.136 71.649 17.176 71.685 ;
          END
     END q[26]
     PIN din[26]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 70.94 17.452 72.1 ;
               LAYER v4 ;
               RECT 17.412 71.878 17.452 71.914 ;
          END
     END din[26]
     PIN q[27]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 73.34 17.176 74.5 ;
               LAYER v4 ;
               RECT 17.136 74.049 17.176 74.085 ;
          END
     END q[27]
     PIN din[27]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 73.34 17.452 74.5 ;
               LAYER v4 ;
               RECT 17.412 74.278 17.452 74.314 ;
          END
     END din[27]
     PIN q[28]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 75.74 17.176 76.9 ;
               LAYER v4 ;
               RECT 17.136 76.449 17.176 76.485 ;
          END
     END q[28]
     PIN din[28]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 75.74 17.452 76.9 ;
               LAYER v4 ;
               RECT 17.412 76.678 17.452 76.714 ;
          END
     END din[28]
     PIN q[29]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 78.14 17.176 79.3 ;
               LAYER v4 ;
               RECT 17.136 78.849 17.176 78.885 ;
          END
     END q[29]
     PIN din[29]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 78.14 17.452 79.3 ;
               LAYER v4 ;
               RECT 17.412 79.078 17.452 79.114 ;
          END
     END din[29]
     PIN q[30]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 80.54 17.176 81.7 ;
               LAYER v4 ;
               RECT 17.136 81.249 17.176 81.285 ;
          END
     END q[30]
     PIN din[30]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 80.54 17.452 81.7 ;
               LAYER v4 ;
               RECT 17.412 81.478 17.452 81.514 ;
          END
     END din[30]
     PIN q[31]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 82.94 17.176 84.1 ;
               LAYER v4 ;
               RECT 17.136 83.649 17.176 83.685 ;
          END
     END q[31]
     PIN din[31]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 82.94 17.452 84.1 ;
               LAYER v4 ;
               RECT 17.412 83.878 17.452 83.914 ;
          END
     END din[31]
     PIN q[32]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 85.34 17.176 86.5 ;
               LAYER v4 ;
               RECT 17.136 86.049 17.176 86.085 ;
          END
     END q[32]
     PIN din[32]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 85.34 17.452 86.5 ;
               LAYER v4 ;
               RECT 17.412 86.278 17.452 86.314 ;
          END
     END din[32]
     PIN q[33]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 87.74 17.176 88.9 ;
               LAYER v4 ;
               RECT 17.136 88.449 17.176 88.485 ;
          END
     END q[33]
     PIN din[33]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 87.74 17.452 88.9 ;
               LAYER v4 ;
               RECT 17.412 88.678 17.452 88.714 ;
          END
     END din[33]
     PIN q[34]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 90.14 17.176 91.3 ;
               LAYER v4 ;
               RECT 17.136 90.849 17.176 90.885 ;
          END
     END q[34]
     PIN din[34]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 90.14 17.452 91.3 ;
               LAYER v4 ;
               RECT 17.412 91.078 17.452 91.114 ;
          END
     END din[34]
     PIN q[35]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 92.54 17.176 93.7 ;
               LAYER v4 ;
               RECT 17.136 93.249 17.176 93.285 ;
          END
     END q[35]
     PIN din[35]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 92.54 17.452 93.7 ;
               LAYER v4 ;
               RECT 17.412 93.478 17.452 93.514 ;
          END
     END din[35]
     PIN q[36]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 94.94 17.176 96.1 ;
               LAYER v4 ;
               RECT 17.136 95.649 17.176 95.685 ;
          END
     END q[36]
     PIN din[36]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 94.94 17.452 96.1 ;
               LAYER v4 ;
               RECT 17.412 95.878 17.452 95.914 ;
          END
     END din[36]
     PIN q[37]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 97.34 17.176 98.5 ;
               LAYER v4 ;
               RECT 17.136 98.049 17.176 98.085 ;
          END
     END q[37]
     PIN din[37]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 97.34 17.452 98.5 ;
               LAYER v4 ;
               RECT 17.412 98.278 17.452 98.314 ;
          END
     END din[37]
     PIN q[38]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 99.74 17.176 100.9 ;
               LAYER v4 ;
               RECT 17.136 100.449 17.176 100.485 ;
          END
     END q[38]
     PIN din[38]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 99.74 17.452 100.9 ;
               LAYER v4 ;
               RECT 17.412 100.678 17.452 100.714 ;
          END
     END din[38]
     PIN q[39]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.136 102.14 17.176 103.3 ;
               LAYER v4 ;
               RECT 17.136 102.849 17.176 102.885 ;
          END
     END q[39]
     PIN din[39]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m5 ;
               RECT 17.412 102.14 17.452 103.3 ;
               LAYER v4 ;
               RECT 17.412 103.078 17.452 103.114 ;
          END
     END din[39]
     PIN clk
     DIRECTION input ;
          USE CLOCK ;
          PORT
               LAYER m5 ;
               RECT 17.136 52.65 17.176 53.61 ;
               LAYER v4 ;
               RECT 17.136 53.142 17.176 53.178 ;
          END
     END clk
     PIN vddp
     SHAPE ABUTMENT ;
     DIRECTION input ;
          USE POWER ;
          PORT
               LAYER m5 ;
               RECT 0.654 49.7505 0.706 55.3695 ;
               LAYER v4 ;
               RECT 0.654 49.782 0.706 49.818 ;
               RECT 0.654 50.262 0.706 50.298 ;
               RECT 0.654 50.502 0.706 50.538 ;
               RECT 0.654 50.982 0.706 51.018 ;
               RECT 0.654 51.102 0.706 51.138 ;
               RECT 0.654 51.582 0.706 51.618 ;
               RECT 0.654 52.062 0.706 52.098 ;
               RECT 0.654 52.182 0.706 52.218 ;
               RECT 0.654 52.542 0.706 52.578 ;
               RECT 0.654 52.662 0.706 52.698 ;
               RECT 0.654 52.902 0.706 52.938 ;
               RECT 0.654 53.022 0.706 53.058 ;
               RECT 0.654 53.502 0.706 53.538 ;
               RECT 0.654 53.982 0.706 54.018 ;
               RECT 0.654 54.102 0.706 54.138 ;
               RECT 0.654 54.582 0.706 54.618 ;
               RECT 0.654 54.822 0.706 54.858 ;
               RECT 0.654 55.302 0.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 0.974 0.6 1.026 104.52 ;
               LAYER v4 ;
               RECT 0.974 49.542 1.026 49.578 ;
               RECT 0.974 49.782 1.026 49.818 ;
               RECT 0.974 50.262 1.026 50.298 ;
               RECT 0.974 50.502 1.026 50.538 ;
               RECT 0.974 50.982 1.026 51.018 ;
               RECT 0.974 51.102 1.026 51.138 ;
               RECT 0.974 51.582 1.026 51.618 ;
               RECT 0.974 52.062 1.026 52.098 ;
               RECT 0.974 52.182 1.026 52.218 ;
               RECT 0.974 52.542 1.026 52.578 ;
               RECT 0.974 52.662 1.026 52.698 ;
               RECT 0.974 52.902 1.026 52.938 ;
               RECT 0.974 53.502 1.026 53.538 ;
               RECT 0.974 53.982 1.026 54.018 ;
               RECT 0.974 54.102 1.026 54.138 ;
               RECT 0.974 54.582 1.026 54.618 ;
               RECT 0.974 54.822 1.026 54.858 ;
               RECT 0.974 55.302 1.026 55.338 ;
               RECT 0.974 55.542 1.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 1.454 49.7505 1.506 55.3695 ;
               LAYER v4 ;
               RECT 1.454 49.782 1.506 49.818 ;
               RECT 1.454 50.262 1.506 50.298 ;
               RECT 1.454 50.502 1.506 50.538 ;
               RECT 1.454 50.982 1.506 51.018 ;
               RECT 1.454 51.102 1.506 51.138 ;
               RECT 1.454 51.582 1.506 51.618 ;
               RECT 1.454 52.062 1.506 52.098 ;
               RECT 1.454 52.182 1.506 52.218 ;
               RECT 1.454 52.542 1.506 52.578 ;
               RECT 1.454 52.662 1.506 52.698 ;
               RECT 1.454 52.902 1.506 52.938 ;
               RECT 1.454 53.022 1.506 53.058 ;
               RECT 1.454 53.502 1.506 53.538 ;
               RECT 1.454 53.982 1.506 54.018 ;
               RECT 1.454 54.102 1.506 54.138 ;
               RECT 1.454 54.582 1.506 54.618 ;
               RECT 1.454 54.822 1.506 54.858 ;
               RECT 1.454 55.302 1.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 1.774 0.6 1.826 104.52 ;
               LAYER v4 ;
               RECT 1.774 49.542 1.826 49.578 ;
               RECT 1.774 49.782 1.826 49.818 ;
               RECT 1.774 50.262 1.826 50.298 ;
               RECT 1.774 50.502 1.826 50.538 ;
               RECT 1.774 50.982 1.826 51.018 ;
               RECT 1.774 51.102 1.826 51.138 ;
               RECT 1.774 51.582 1.826 51.618 ;
               RECT 1.774 52.062 1.826 52.098 ;
               RECT 1.774 52.182 1.826 52.218 ;
               RECT 1.774 52.542 1.826 52.578 ;
               RECT 1.774 52.662 1.826 52.698 ;
               RECT 1.774 52.902 1.826 52.938 ;
               RECT 1.774 53.502 1.826 53.538 ;
               RECT 1.774 53.982 1.826 54.018 ;
               RECT 1.774 54.102 1.826 54.138 ;
               RECT 1.774 54.582 1.826 54.618 ;
               RECT 1.774 54.822 1.826 54.858 ;
               RECT 1.774 55.302 1.826 55.338 ;
               RECT 1.774 55.542 1.826 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 10.254 49.7505 10.306 55.3695 ;
               LAYER v4 ;
               RECT 10.254 49.782 10.306 49.818 ;
               RECT 10.254 50.262 10.306 50.298 ;
               RECT 10.254 50.502 10.306 50.538 ;
               RECT 10.254 50.982 10.306 51.018 ;
               RECT 10.254 51.102 10.306 51.138 ;
               RECT 10.254 51.582 10.306 51.618 ;
               RECT 10.254 52.062 10.306 52.098 ;
               RECT 10.254 52.182 10.306 52.218 ;
               RECT 10.254 52.542 10.306 52.578 ;
               RECT 10.254 52.662 10.306 52.698 ;
               RECT 10.254 52.902 10.306 52.938 ;
               RECT 10.254 53.022 10.306 53.058 ;
               RECT 10.254 53.502 10.306 53.538 ;
               RECT 10.254 53.982 10.306 54.018 ;
               RECT 10.254 54.102 10.306 54.138 ;
               RECT 10.254 54.582 10.306 54.618 ;
               RECT 10.254 54.822 10.306 54.858 ;
               RECT 10.254 55.302 10.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 10.574 0.6 10.626 104.52 ;
               LAYER v4 ;
               RECT 10.574 49.542 10.626 49.578 ;
               RECT 10.574 49.782 10.626 49.818 ;
               RECT 10.574 50.262 10.626 50.298 ;
               RECT 10.574 50.502 10.626 50.538 ;
               RECT 10.574 50.982 10.626 51.018 ;
               RECT 10.574 51.102 10.626 51.138 ;
               RECT 10.574 51.582 10.626 51.618 ;
               RECT 10.574 52.062 10.626 52.098 ;
               RECT 10.574 52.182 10.626 52.218 ;
               RECT 10.574 52.542 10.626 52.578 ;
               RECT 10.574 52.662 10.626 52.698 ;
               RECT 10.574 52.902 10.626 52.938 ;
               RECT 10.574 53.502 10.626 53.538 ;
               RECT 10.574 53.982 10.626 54.018 ;
               RECT 10.574 54.102 10.626 54.138 ;
               RECT 10.574 54.582 10.626 54.618 ;
               RECT 10.574 54.822 10.626 54.858 ;
               RECT 10.574 55.302 10.626 55.338 ;
               RECT 10.574 55.542 10.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 11.054 49.7505 11.106 55.3695 ;
               LAYER v4 ;
               RECT 11.054 49.782 11.106 49.818 ;
               RECT 11.054 50.262 11.106 50.298 ;
               RECT 11.054 50.502 11.106 50.538 ;
               RECT 11.054 50.982 11.106 51.018 ;
               RECT 11.054 51.102 11.106 51.138 ;
               RECT 11.054 51.582 11.106 51.618 ;
               RECT 11.054 52.062 11.106 52.098 ;
               RECT 11.054 52.182 11.106 52.218 ;
               RECT 11.054 52.542 11.106 52.578 ;
               RECT 11.054 52.662 11.106 52.698 ;
               RECT 11.054 52.902 11.106 52.938 ;
               RECT 11.054 53.022 11.106 53.058 ;
               RECT 11.054 53.502 11.106 53.538 ;
               RECT 11.054 53.982 11.106 54.018 ;
               RECT 11.054 54.102 11.106 54.138 ;
               RECT 11.054 54.582 11.106 54.618 ;
               RECT 11.054 54.822 11.106 54.858 ;
               RECT 11.054 55.302 11.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 11.374 0.6 11.426 104.52 ;
               LAYER v4 ;
               RECT 11.374 49.542 11.426 49.578 ;
               RECT 11.374 49.782 11.426 49.818 ;
               RECT 11.374 50.262 11.426 50.298 ;
               RECT 11.374 50.502 11.426 50.538 ;
               RECT 11.374 50.982 11.426 51.018 ;
               RECT 11.374 51.102 11.426 51.138 ;
               RECT 11.374 51.582 11.426 51.618 ;
               RECT 11.374 52.062 11.426 52.098 ;
               RECT 11.374 52.182 11.426 52.218 ;
               RECT 11.374 52.542 11.426 52.578 ;
               RECT 11.374 52.662 11.426 52.698 ;
               RECT 11.374 52.902 11.426 52.938 ;
               RECT 11.374 53.502 11.426 53.538 ;
               RECT 11.374 53.982 11.426 54.018 ;
               RECT 11.374 54.102 11.426 54.138 ;
               RECT 11.374 54.582 11.426 54.618 ;
               RECT 11.374 54.822 11.426 54.858 ;
               RECT 11.374 55.302 11.426 55.338 ;
               RECT 11.374 55.542 11.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 11.854 49.7505 11.906 55.3695 ;
               LAYER v4 ;
               RECT 11.854 49.782 11.906 49.818 ;
               RECT 11.854 50.262 11.906 50.298 ;
               RECT 11.854 50.502 11.906 50.538 ;
               RECT 11.854 50.982 11.906 51.018 ;
               RECT 11.854 51.102 11.906 51.138 ;
               RECT 11.854 51.582 11.906 51.618 ;
               RECT 11.854 52.062 11.906 52.098 ;
               RECT 11.854 52.182 11.906 52.218 ;
               RECT 11.854 52.542 11.906 52.578 ;
               RECT 11.854 52.662 11.906 52.698 ;
               RECT 11.854 52.902 11.906 52.938 ;
               RECT 11.854 53.022 11.906 53.058 ;
               RECT 11.854 53.502 11.906 53.538 ;
               RECT 11.854 53.982 11.906 54.018 ;
               RECT 11.854 54.102 11.906 54.138 ;
               RECT 11.854 54.582 11.906 54.618 ;
               RECT 11.854 54.822 11.906 54.858 ;
               RECT 11.854 55.302 11.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 12.174 0.6 12.226 104.52 ;
               LAYER v4 ;
               RECT 12.174 49.542 12.226 49.578 ;
               RECT 12.174 49.782 12.226 49.818 ;
               RECT 12.174 50.262 12.226 50.298 ;
               RECT 12.174 50.502 12.226 50.538 ;
               RECT 12.174 50.982 12.226 51.018 ;
               RECT 12.174 51.102 12.226 51.138 ;
               RECT 12.174 51.582 12.226 51.618 ;
               RECT 12.174 52.062 12.226 52.098 ;
               RECT 12.174 52.182 12.226 52.218 ;
               RECT 12.174 52.542 12.226 52.578 ;
               RECT 12.174 52.662 12.226 52.698 ;
               RECT 12.174 52.902 12.226 52.938 ;
               RECT 12.174 53.502 12.226 53.538 ;
               RECT 12.174 53.982 12.226 54.018 ;
               RECT 12.174 54.102 12.226 54.138 ;
               RECT 12.174 54.582 12.226 54.618 ;
               RECT 12.174 54.822 12.226 54.858 ;
               RECT 12.174 55.302 12.226 55.338 ;
               RECT 12.174 55.542 12.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 12.654 49.7505 12.706 55.3695 ;
               LAYER v4 ;
               RECT 12.654 49.782 12.706 49.818 ;
               RECT 12.654 50.262 12.706 50.298 ;
               RECT 12.654 50.502 12.706 50.538 ;
               RECT 12.654 50.982 12.706 51.018 ;
               RECT 12.654 51.102 12.706 51.138 ;
               RECT 12.654 51.582 12.706 51.618 ;
               RECT 12.654 52.062 12.706 52.098 ;
               RECT 12.654 52.182 12.706 52.218 ;
               RECT 12.654 52.542 12.706 52.578 ;
               RECT 12.654 52.662 12.706 52.698 ;
               RECT 12.654 52.902 12.706 52.938 ;
               RECT 12.654 53.022 12.706 53.058 ;
               RECT 12.654 53.502 12.706 53.538 ;
               RECT 12.654 53.982 12.706 54.018 ;
               RECT 12.654 54.102 12.706 54.138 ;
               RECT 12.654 54.582 12.706 54.618 ;
               RECT 12.654 54.822 12.706 54.858 ;
               RECT 12.654 55.302 12.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 12.974 0.6 13.026 104.52 ;
               LAYER v4 ;
               RECT 12.974 49.542 13.026 49.578 ;
               RECT 12.974 49.782 13.026 49.818 ;
               RECT 12.974 50.262 13.026 50.298 ;
               RECT 12.974 50.502 13.026 50.538 ;
               RECT 12.974 50.982 13.026 51.018 ;
               RECT 12.974 51.102 13.026 51.138 ;
               RECT 12.974 51.582 13.026 51.618 ;
               RECT 12.974 52.062 13.026 52.098 ;
               RECT 12.974 52.182 13.026 52.218 ;
               RECT 12.974 52.542 13.026 52.578 ;
               RECT 12.974 52.662 13.026 52.698 ;
               RECT 12.974 52.902 13.026 52.938 ;
               RECT 12.974 53.502 13.026 53.538 ;
               RECT 12.974 53.982 13.026 54.018 ;
               RECT 12.974 54.102 13.026 54.138 ;
               RECT 12.974 54.582 13.026 54.618 ;
               RECT 12.974 54.822 13.026 54.858 ;
               RECT 12.974 55.302 13.026 55.338 ;
               RECT 12.974 55.542 13.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 14.05 0.5695 14.104 104.5505 ;
               LAYER v4 ;
               RECT 14.05 0.729 14.104 0.765 ;
               RECT 14.05 0.958 14.104 0.994 ;
               RECT 14.05 1.406 14.104 1.442 ;
               RECT 14.05 1.929 14.104 1.965 ;
               RECT 14.05 2.158 14.104 2.194 ;
               RECT 14.05 2.606 14.104 2.642 ;
               RECT 14.05 3.129 14.104 3.165 ;
               RECT 14.05 3.358 14.104 3.394 ;
               RECT 14.05 3.806 14.104 3.842 ;
               RECT 14.05 4.329 14.104 4.365 ;
               RECT 14.05 4.558 14.104 4.594 ;
               RECT 14.05 5.006 14.104 5.042 ;
               RECT 14.05 5.529 14.104 5.565 ;
               RECT 14.05 5.758 14.104 5.794 ;
               RECT 14.05 6.206 14.104 6.242 ;
               RECT 14.05 6.729 14.104 6.765 ;
               RECT 14.05 6.958 14.104 6.994 ;
               RECT 14.05 7.406 14.104 7.442 ;
               RECT 14.05 7.929 14.104 7.965 ;
               RECT 14.05 8.158 14.104 8.194 ;
               RECT 14.05 8.606 14.104 8.642 ;
               RECT 14.05 9.129 14.104 9.165 ;
               RECT 14.05 9.358 14.104 9.394 ;
               RECT 14.05 9.806 14.104 9.842 ;
               RECT 14.05 10.329 14.104 10.365 ;
               RECT 14.05 10.558 14.104 10.594 ;
               RECT 14.05 11.006 14.104 11.042 ;
               RECT 14.05 11.529 14.104 11.565 ;
               RECT 14.05 11.758 14.104 11.794 ;
               RECT 14.05 12.206 14.104 12.242 ;
               RECT 14.05 12.729 14.104 12.765 ;
               RECT 14.05 12.958 14.104 12.994 ;
               RECT 14.05 13.406 14.104 13.442 ;
               RECT 14.05 13.929 14.104 13.965 ;
               RECT 14.05 14.158 14.104 14.194 ;
               RECT 14.05 14.606 14.104 14.642 ;
               RECT 14.05 15.129 14.104 15.165 ;
               RECT 14.05 15.358 14.104 15.394 ;
               RECT 14.05 15.806 14.104 15.842 ;
               RECT 14.05 16.329 14.104 16.365 ;
               RECT 14.05 16.558 14.104 16.594 ;
               RECT 14.05 17.006 14.104 17.042 ;
               RECT 14.05 17.529 14.104 17.565 ;
               RECT 14.05 17.758 14.104 17.794 ;
               RECT 14.05 18.206 14.104 18.242 ;
               RECT 14.05 18.729 14.104 18.765 ;
               RECT 14.05 18.958 14.104 18.994 ;
               RECT 14.05 19.406 14.104 19.442 ;
               RECT 14.05 19.929 14.104 19.965 ;
               RECT 14.05 20.158 14.104 20.194 ;
               RECT 14.05 20.606 14.104 20.642 ;
               RECT 14.05 21.129 14.104 21.165 ;
               RECT 14.05 21.358 14.104 21.394 ;
               RECT 14.05 21.806 14.104 21.842 ;
               RECT 14.05 22.329 14.104 22.365 ;
               RECT 14.05 22.558 14.104 22.594 ;
               RECT 14.05 23.006 14.104 23.042 ;
               RECT 14.05 23.529 14.104 23.565 ;
               RECT 14.05 23.758 14.104 23.794 ;
               RECT 14.05 24.206 14.104 24.242 ;
               RECT 14.05 24.729 14.104 24.765 ;
               RECT 14.05 24.958 14.104 24.994 ;
               RECT 14.05 25.406 14.104 25.442 ;
               RECT 14.05 25.929 14.104 25.965 ;
               RECT 14.05 26.158 14.104 26.194 ;
               RECT 14.05 26.606 14.104 26.642 ;
               RECT 14.05 27.129 14.104 27.165 ;
               RECT 14.05 27.358 14.104 27.394 ;
               RECT 14.05 27.806 14.104 27.842 ;
               RECT 14.05 28.329 14.104 28.365 ;
               RECT 14.05 28.558 14.104 28.594 ;
               RECT 14.05 29.006 14.104 29.042 ;
               RECT 14.05 29.529 14.104 29.565 ;
               RECT 14.05 29.758 14.104 29.794 ;
               RECT 14.05 30.206 14.104 30.242 ;
               RECT 14.05 30.729 14.104 30.765 ;
               RECT 14.05 30.958 14.104 30.994 ;
               RECT 14.05 31.406 14.104 31.442 ;
               RECT 14.05 31.929 14.104 31.965 ;
               RECT 14.05 32.158 14.104 32.194 ;
               RECT 14.05 32.606 14.104 32.642 ;
               RECT 14.05 33.129 14.104 33.165 ;
               RECT 14.05 33.358 14.104 33.394 ;
               RECT 14.05 33.806 14.104 33.842 ;
               RECT 14.05 34.329 14.104 34.365 ;
               RECT 14.05 34.558 14.104 34.594 ;
               RECT 14.05 35.006 14.104 35.042 ;
               RECT 14.05 35.529 14.104 35.565 ;
               RECT 14.05 35.758 14.104 35.794 ;
               RECT 14.05 36.206 14.104 36.242 ;
               RECT 14.05 36.729 14.104 36.765 ;
               RECT 14.05 36.958 14.104 36.994 ;
               RECT 14.05 37.406 14.104 37.442 ;
               RECT 14.05 37.929 14.104 37.965 ;
               RECT 14.05 38.158 14.104 38.194 ;
               RECT 14.05 38.606 14.104 38.642 ;
               RECT 14.05 39.129 14.104 39.165 ;
               RECT 14.05 39.358 14.104 39.394 ;
               RECT 14.05 39.806 14.104 39.842 ;
               RECT 14.05 40.329 14.104 40.365 ;
               RECT 14.05 40.558 14.104 40.594 ;
               RECT 14.05 41.006 14.104 41.042 ;
               RECT 14.05 41.529 14.104 41.565 ;
               RECT 14.05 41.758 14.104 41.794 ;
               RECT 14.05 42.206 14.104 42.242 ;
               RECT 14.05 42.729 14.104 42.765 ;
               RECT 14.05 42.958 14.104 42.994 ;
               RECT 14.05 43.406 14.104 43.442 ;
               RECT 14.05 43.929 14.104 43.965 ;
               RECT 14.05 44.158 14.104 44.194 ;
               RECT 14.05 44.606 14.104 44.642 ;
               RECT 14.05 45.129 14.104 45.165 ;
               RECT 14.05 45.358 14.104 45.394 ;
               RECT 14.05 45.806 14.104 45.842 ;
               RECT 14.05 46.329 14.104 46.365 ;
               RECT 14.05 46.558 14.104 46.594 ;
               RECT 14.05 47.006 14.104 47.042 ;
               RECT 14.05 47.529 14.104 47.565 ;
               RECT 14.05 47.758 14.104 47.794 ;
               RECT 14.05 48.206 14.104 48.242 ;
               RECT 14.05 49.062 14.104 49.098 ;
               RECT 14.05 49.182 14.104 49.218 ;
               RECT 14.05 49.542 14.104 49.578 ;
               RECT 14.05 49.662 14.104 49.698 ;
               RECT 14.05 49.782 14.104 49.818 ;
               RECT 14.05 50.142 14.104 50.178 ;
               RECT 14.05 50.262 14.104 50.298 ;
               RECT 14.05 50.622 14.104 50.658 ;
               RECT 14.05 51.5875 14.104 51.6125 ;
               RECT 14.05 52.062 14.104 52.098 ;
               RECT 14.05 52.182 14.104 52.218 ;
               RECT 14.05 52.542 14.104 52.578 ;
               RECT 14.05 52.902 14.104 52.938 ;
               RECT 14.05 53.022 14.104 53.058 ;
               RECT 14.05 53.502 14.104 53.538 ;
               RECT 14.05 53.9875 14.104 54.0125 ;
               RECT 14.05 54.462 14.104 54.498 ;
               RECT 14.05 54.822 14.104 54.858 ;
               RECT 14.05 54.942 14.104 54.978 ;
               RECT 14.05 55.302 14.104 55.338 ;
               RECT 14.05 55.422 14.104 55.458 ;
               RECT 14.05 55.542 14.104 55.578 ;
               RECT 14.05 55.902 14.104 55.938 ;
               RECT 14.05 56.649 14.104 56.685 ;
               RECT 14.05 56.878 14.104 56.914 ;
               RECT 14.05 57.326 14.104 57.362 ;
               RECT 14.05 57.849 14.104 57.885 ;
               RECT 14.05 58.078 14.104 58.114 ;
               RECT 14.05 58.526 14.104 58.562 ;
               RECT 14.05 59.049 14.104 59.085 ;
               RECT 14.05 59.278 14.104 59.314 ;
               RECT 14.05 59.726 14.104 59.762 ;
               RECT 14.05 60.249 14.104 60.285 ;
               RECT 14.05 60.478 14.104 60.514 ;
               RECT 14.05 60.926 14.104 60.962 ;
               RECT 14.05 61.449 14.104 61.485 ;
               RECT 14.05 61.678 14.104 61.714 ;
               RECT 14.05 62.126 14.104 62.162 ;
               RECT 14.05 62.649 14.104 62.685 ;
               RECT 14.05 62.878 14.104 62.914 ;
               RECT 14.05 63.326 14.104 63.362 ;
               RECT 14.05 63.849 14.104 63.885 ;
               RECT 14.05 64.078 14.104 64.114 ;
               RECT 14.05 64.526 14.104 64.562 ;
               RECT 14.05 65.049 14.104 65.085 ;
               RECT 14.05 65.278 14.104 65.314 ;
               RECT 14.05 65.726 14.104 65.762 ;
               RECT 14.05 66.249 14.104 66.285 ;
               RECT 14.05 66.478 14.104 66.514 ;
               RECT 14.05 66.926 14.104 66.962 ;
               RECT 14.05 67.449 14.104 67.485 ;
               RECT 14.05 67.678 14.104 67.714 ;
               RECT 14.05 68.126 14.104 68.162 ;
               RECT 14.05 68.649 14.104 68.685 ;
               RECT 14.05 68.878 14.104 68.914 ;
               RECT 14.05 69.326 14.104 69.362 ;
               RECT 14.05 69.849 14.104 69.885 ;
               RECT 14.05 70.078 14.104 70.114 ;
               RECT 14.05 70.526 14.104 70.562 ;
               RECT 14.05 71.049 14.104 71.085 ;
               RECT 14.05 71.278 14.104 71.314 ;
               RECT 14.05 71.726 14.104 71.762 ;
               RECT 14.05 72.249 14.104 72.285 ;
               RECT 14.05 72.478 14.104 72.514 ;
               RECT 14.05 72.926 14.104 72.962 ;
               RECT 14.05 73.449 14.104 73.485 ;
               RECT 14.05 73.678 14.104 73.714 ;
               RECT 14.05 74.126 14.104 74.162 ;
               RECT 14.05 74.649 14.104 74.685 ;
               RECT 14.05 74.878 14.104 74.914 ;
               RECT 14.05 75.326 14.104 75.362 ;
               RECT 14.05 75.849 14.104 75.885 ;
               RECT 14.05 76.078 14.104 76.114 ;
               RECT 14.05 76.526 14.104 76.562 ;
               RECT 14.05 77.049 14.104 77.085 ;
               RECT 14.05 77.278 14.104 77.314 ;
               RECT 14.05 77.726 14.104 77.762 ;
               RECT 14.05 78.249 14.104 78.285 ;
               RECT 14.05 78.478 14.104 78.514 ;
               RECT 14.05 78.926 14.104 78.962 ;
               RECT 14.05 79.449 14.104 79.485 ;
               RECT 14.05 79.678 14.104 79.714 ;
               RECT 14.05 80.126 14.104 80.162 ;
               RECT 14.05 80.649 14.104 80.685 ;
               RECT 14.05 80.878 14.104 80.914 ;
               RECT 14.05 81.326 14.104 81.362 ;
               RECT 14.05 81.849 14.104 81.885 ;
               RECT 14.05 82.078 14.104 82.114 ;
               RECT 14.05 82.526 14.104 82.562 ;
               RECT 14.05 83.049 14.104 83.085 ;
               RECT 14.05 83.278 14.104 83.314 ;
               RECT 14.05 83.726 14.104 83.762 ;
               RECT 14.05 84.249 14.104 84.285 ;
               RECT 14.05 84.478 14.104 84.514 ;
               RECT 14.05 84.926 14.104 84.962 ;
               RECT 14.05 85.449 14.104 85.485 ;
               RECT 14.05 85.678 14.104 85.714 ;
               RECT 14.05 86.126 14.104 86.162 ;
               RECT 14.05 86.649 14.104 86.685 ;
               RECT 14.05 86.878 14.104 86.914 ;
               RECT 14.05 87.326 14.104 87.362 ;
               RECT 14.05 87.849 14.104 87.885 ;
               RECT 14.05 88.078 14.104 88.114 ;
               RECT 14.05 88.526 14.104 88.562 ;
               RECT 14.05 89.049 14.104 89.085 ;
               RECT 14.05 89.278 14.104 89.314 ;
               RECT 14.05 89.726 14.104 89.762 ;
               RECT 14.05 90.249 14.104 90.285 ;
               RECT 14.05 90.478 14.104 90.514 ;
               RECT 14.05 90.926 14.104 90.962 ;
               RECT 14.05 91.449 14.104 91.485 ;
               RECT 14.05 91.678 14.104 91.714 ;
               RECT 14.05 92.126 14.104 92.162 ;
               RECT 14.05 92.649 14.104 92.685 ;
               RECT 14.05 92.878 14.104 92.914 ;
               RECT 14.05 93.326 14.104 93.362 ;
               RECT 14.05 93.849 14.104 93.885 ;
               RECT 14.05 94.078 14.104 94.114 ;
               RECT 14.05 94.526 14.104 94.562 ;
               RECT 14.05 95.049 14.104 95.085 ;
               RECT 14.05 95.278 14.104 95.314 ;
               RECT 14.05 95.726 14.104 95.762 ;
               RECT 14.05 96.249 14.104 96.285 ;
               RECT 14.05 96.478 14.104 96.514 ;
               RECT 14.05 96.926 14.104 96.962 ;
               RECT 14.05 97.449 14.104 97.485 ;
               RECT 14.05 97.678 14.104 97.714 ;
               RECT 14.05 98.126 14.104 98.162 ;
               RECT 14.05 98.649 14.104 98.685 ;
               RECT 14.05 98.878 14.104 98.914 ;
               RECT 14.05 99.326 14.104 99.362 ;
               RECT 14.05 99.849 14.104 99.885 ;
               RECT 14.05 100.078 14.104 100.114 ;
               RECT 14.05 100.526 14.104 100.562 ;
               RECT 14.05 101.049 14.104 101.085 ;
               RECT 14.05 101.278 14.104 101.314 ;
               RECT 14.05 101.726 14.104 101.762 ;
               RECT 14.05 102.249 14.104 102.285 ;
               RECT 14.05 102.478 14.104 102.514 ;
               RECT 14.05 102.926 14.104 102.962 ;
               RECT 14.05 103.449 14.104 103.485 ;
               RECT 14.05 103.678 14.104 103.714 ;
               RECT 14.05 104.126 14.104 104.162 ;
          END
          PORT
               LAYER m5 ;
               RECT 14.296 0.5695 14.35 104.5505 ;
               LAYER v4 ;
               RECT 14.296 0.958 14.35 0.994 ;
               RECT 14.296 1.406 14.35 1.442 ;
               RECT 14.296 1.635 14.35 1.671 ;
               RECT 14.296 2.158 14.35 2.194 ;
               RECT 14.296 2.606 14.35 2.642 ;
               RECT 14.296 2.835 14.35 2.871 ;
               RECT 14.296 3.358 14.35 3.394 ;
               RECT 14.296 3.806 14.35 3.842 ;
               RECT 14.296 4.035 14.35 4.071 ;
               RECT 14.296 4.558 14.35 4.594 ;
               RECT 14.296 5.006 14.35 5.042 ;
               RECT 14.296 5.235 14.35 5.271 ;
               RECT 14.296 5.758 14.35 5.794 ;
               RECT 14.296 6.206 14.35 6.242 ;
               RECT 14.296 6.435 14.35 6.471 ;
               RECT 14.296 6.958 14.35 6.994 ;
               RECT 14.296 7.406 14.35 7.442 ;
               RECT 14.296 7.635 14.35 7.671 ;
               RECT 14.296 8.158 14.35 8.194 ;
               RECT 14.296 8.606 14.35 8.642 ;
               RECT 14.296 8.835 14.35 8.871 ;
               RECT 14.296 9.358 14.35 9.394 ;
               RECT 14.296 9.806 14.35 9.842 ;
               RECT 14.296 10.035 14.35 10.071 ;
               RECT 14.296 10.558 14.35 10.594 ;
               RECT 14.296 11.006 14.35 11.042 ;
               RECT 14.296 11.235 14.35 11.271 ;
               RECT 14.296 11.758 14.35 11.794 ;
               RECT 14.296 12.206 14.35 12.242 ;
               RECT 14.296 12.435 14.35 12.471 ;
               RECT 14.296 12.958 14.35 12.994 ;
               RECT 14.296 13.406 14.35 13.442 ;
               RECT 14.296 13.635 14.35 13.671 ;
               RECT 14.296 14.158 14.35 14.194 ;
               RECT 14.296 14.606 14.35 14.642 ;
               RECT 14.296 14.835 14.35 14.871 ;
               RECT 14.296 15.358 14.35 15.394 ;
               RECT 14.296 15.806 14.35 15.842 ;
               RECT 14.296 16.035 14.35 16.071 ;
               RECT 14.296 16.558 14.35 16.594 ;
               RECT 14.296 17.006 14.35 17.042 ;
               RECT 14.296 17.235 14.35 17.271 ;
               RECT 14.296 17.758 14.35 17.794 ;
               RECT 14.296 18.206 14.35 18.242 ;
               RECT 14.296 18.435 14.35 18.471 ;
               RECT 14.296 18.958 14.35 18.994 ;
               RECT 14.296 19.406 14.35 19.442 ;
               RECT 14.296 19.635 14.35 19.671 ;
               RECT 14.296 20.158 14.35 20.194 ;
               RECT 14.296 20.606 14.35 20.642 ;
               RECT 14.296 20.835 14.35 20.871 ;
               RECT 14.296 21.358 14.35 21.394 ;
               RECT 14.296 21.806 14.35 21.842 ;
               RECT 14.296 22.035 14.35 22.071 ;
               RECT 14.296 22.558 14.35 22.594 ;
               RECT 14.296 23.006 14.35 23.042 ;
               RECT 14.296 23.235 14.35 23.271 ;
               RECT 14.296 23.758 14.35 23.794 ;
               RECT 14.296 24.206 14.35 24.242 ;
               RECT 14.296 24.435 14.35 24.471 ;
               RECT 14.296 24.958 14.35 24.994 ;
               RECT 14.296 25.406 14.35 25.442 ;
               RECT 14.296 25.635 14.35 25.671 ;
               RECT 14.296 26.158 14.35 26.194 ;
               RECT 14.296 26.606 14.35 26.642 ;
               RECT 14.296 26.835 14.35 26.871 ;
               RECT 14.296 27.358 14.35 27.394 ;
               RECT 14.296 27.806 14.35 27.842 ;
               RECT 14.296 28.035 14.35 28.071 ;
               RECT 14.296 28.558 14.35 28.594 ;
               RECT 14.296 29.006 14.35 29.042 ;
               RECT 14.296 29.235 14.35 29.271 ;
               RECT 14.296 29.758 14.35 29.794 ;
               RECT 14.296 30.206 14.35 30.242 ;
               RECT 14.296 30.435 14.35 30.471 ;
               RECT 14.296 30.958 14.35 30.994 ;
               RECT 14.296 31.406 14.35 31.442 ;
               RECT 14.296 31.635 14.35 31.671 ;
               RECT 14.296 32.158 14.35 32.194 ;
               RECT 14.296 32.606 14.35 32.642 ;
               RECT 14.296 32.835 14.35 32.871 ;
               RECT 14.296 33.358 14.35 33.394 ;
               RECT 14.296 33.806 14.35 33.842 ;
               RECT 14.296 34.035 14.35 34.071 ;
               RECT 14.296 34.558 14.35 34.594 ;
               RECT 14.296 35.006 14.35 35.042 ;
               RECT 14.296 35.235 14.35 35.271 ;
               RECT 14.296 35.758 14.35 35.794 ;
               RECT 14.296 36.206 14.35 36.242 ;
               RECT 14.296 36.435 14.35 36.471 ;
               RECT 14.296 36.958 14.35 36.994 ;
               RECT 14.296 37.406 14.35 37.442 ;
               RECT 14.296 37.635 14.35 37.671 ;
               RECT 14.296 38.158 14.35 38.194 ;
               RECT 14.296 38.606 14.35 38.642 ;
               RECT 14.296 38.835 14.35 38.871 ;
               RECT 14.296 39.358 14.35 39.394 ;
               RECT 14.296 39.806 14.35 39.842 ;
               RECT 14.296 40.035 14.35 40.071 ;
               RECT 14.296 40.558 14.35 40.594 ;
               RECT 14.296 41.006 14.35 41.042 ;
               RECT 14.296 41.235 14.35 41.271 ;
               RECT 14.296 41.758 14.35 41.794 ;
               RECT 14.296 42.206 14.35 42.242 ;
               RECT 14.296 42.435 14.35 42.471 ;
               RECT 14.296 42.958 14.35 42.994 ;
               RECT 14.296 43.406 14.35 43.442 ;
               RECT 14.296 43.635 14.35 43.671 ;
               RECT 14.296 44.158 14.35 44.194 ;
               RECT 14.296 44.606 14.35 44.642 ;
               RECT 14.296 44.835 14.35 44.871 ;
               RECT 14.296 45.358 14.35 45.394 ;
               RECT 14.296 45.806 14.35 45.842 ;
               RECT 14.296 46.035 14.35 46.071 ;
               RECT 14.296 46.558 14.35 46.594 ;
               RECT 14.296 47.006 14.35 47.042 ;
               RECT 14.296 47.235 14.35 47.271 ;
               RECT 14.296 47.758 14.35 47.794 ;
               RECT 14.296 48.206 14.35 48.242 ;
               RECT 14.296 48.435 14.35 48.471 ;
               RECT 14.296 49.062 14.35 49.098 ;
               RECT 14.296 49.1875 14.35 49.2125 ;
               RECT 14.296 49.542 14.35 49.578 ;
               RECT 14.296 49.662 14.35 49.698 ;
               RECT 14.296 49.782 14.35 49.818 ;
               RECT 14.296 50.142 14.35 50.178 ;
               RECT 14.296 50.262 14.35 50.298 ;
               RECT 14.296 50.622 14.35 50.658 ;
               RECT 14.296 51.102 14.35 51.138 ;
               RECT 14.296 51.582 14.35 51.618 ;
               RECT 14.296 52.062 14.35 52.098 ;
               RECT 14.296 52.182 14.35 52.218 ;
               RECT 14.296 52.542 14.35 52.578 ;
               RECT 14.296 52.902 14.35 52.938 ;
               RECT 14.296 53.022 14.35 53.058 ;
               RECT 14.296 53.5075 14.35 53.5325 ;
               RECT 14.296 53.9875 14.35 54.0125 ;
               RECT 14.296 54.462 14.35 54.498 ;
               RECT 14.296 54.822 14.35 54.858 ;
               RECT 14.296 54.942 14.35 54.978 ;
               RECT 14.296 55.302 14.35 55.338 ;
               RECT 14.296 55.4275 14.35 55.4525 ;
               RECT 14.296 55.542 14.35 55.578 ;
               RECT 14.296 55.902 14.35 55.938 ;
               RECT 14.296 56.878 14.35 56.914 ;
               RECT 14.296 57.326 14.35 57.362 ;
               RECT 14.296 57.555 14.35 57.591 ;
               RECT 14.296 58.078 14.35 58.114 ;
               RECT 14.296 58.526 14.35 58.562 ;
               RECT 14.296 58.755 14.35 58.791 ;
               RECT 14.296 59.278 14.35 59.314 ;
               RECT 14.296 59.726 14.35 59.762 ;
               RECT 14.296 59.955 14.35 59.991 ;
               RECT 14.296 60.478 14.35 60.514 ;
               RECT 14.296 60.926 14.35 60.962 ;
               RECT 14.296 61.155 14.35 61.191 ;
               RECT 14.296 61.678 14.35 61.714 ;
               RECT 14.296 62.126 14.35 62.162 ;
               RECT 14.296 62.355 14.35 62.391 ;
               RECT 14.296 62.878 14.35 62.914 ;
               RECT 14.296 63.326 14.35 63.362 ;
               RECT 14.296 63.555 14.35 63.591 ;
               RECT 14.296 64.078 14.35 64.114 ;
               RECT 14.296 64.526 14.35 64.562 ;
               RECT 14.296 64.755 14.35 64.791 ;
               RECT 14.296 65.278 14.35 65.314 ;
               RECT 14.296 65.726 14.35 65.762 ;
               RECT 14.296 65.955 14.35 65.991 ;
               RECT 14.296 66.478 14.35 66.514 ;
               RECT 14.296 66.926 14.35 66.962 ;
               RECT 14.296 67.155 14.35 67.191 ;
               RECT 14.296 67.678 14.35 67.714 ;
               RECT 14.296 68.126 14.35 68.162 ;
               RECT 14.296 68.355 14.35 68.391 ;
               RECT 14.296 68.878 14.35 68.914 ;
               RECT 14.296 69.326 14.35 69.362 ;
               RECT 14.296 69.555 14.35 69.591 ;
               RECT 14.296 70.078 14.35 70.114 ;
               RECT 14.296 70.526 14.35 70.562 ;
               RECT 14.296 70.755 14.35 70.791 ;
               RECT 14.296 71.278 14.35 71.314 ;
               RECT 14.296 71.726 14.35 71.762 ;
               RECT 14.296 71.955 14.35 71.991 ;
               RECT 14.296 72.478 14.35 72.514 ;
               RECT 14.296 72.926 14.35 72.962 ;
               RECT 14.296 73.155 14.35 73.191 ;
               RECT 14.296 73.678 14.35 73.714 ;
               RECT 14.296 74.126 14.35 74.162 ;
               RECT 14.296 74.355 14.35 74.391 ;
               RECT 14.296 74.878 14.35 74.914 ;
               RECT 14.296 75.326 14.35 75.362 ;
               RECT 14.296 75.555 14.35 75.591 ;
               RECT 14.296 76.078 14.35 76.114 ;
               RECT 14.296 76.526 14.35 76.562 ;
               RECT 14.296 76.755 14.35 76.791 ;
               RECT 14.296 77.278 14.35 77.314 ;
               RECT 14.296 77.726 14.35 77.762 ;
               RECT 14.296 77.955 14.35 77.991 ;
               RECT 14.296 78.478 14.35 78.514 ;
               RECT 14.296 78.926 14.35 78.962 ;
               RECT 14.296 79.155 14.35 79.191 ;
               RECT 14.296 79.678 14.35 79.714 ;
               RECT 14.296 80.126 14.35 80.162 ;
               RECT 14.296 80.355 14.35 80.391 ;
               RECT 14.296 80.878 14.35 80.914 ;
               RECT 14.296 81.326 14.35 81.362 ;
               RECT 14.296 81.555 14.35 81.591 ;
               RECT 14.296 82.078 14.35 82.114 ;
               RECT 14.296 82.526 14.35 82.562 ;
               RECT 14.296 82.755 14.35 82.791 ;
               RECT 14.296 83.278 14.35 83.314 ;
               RECT 14.296 83.726 14.35 83.762 ;
               RECT 14.296 83.955 14.35 83.991 ;
               RECT 14.296 84.478 14.35 84.514 ;
               RECT 14.296 84.926 14.35 84.962 ;
               RECT 14.296 85.155 14.35 85.191 ;
               RECT 14.296 85.678 14.35 85.714 ;
               RECT 14.296 86.126 14.35 86.162 ;
               RECT 14.296 86.355 14.35 86.391 ;
               RECT 14.296 86.878 14.35 86.914 ;
               RECT 14.296 87.326 14.35 87.362 ;
               RECT 14.296 87.555 14.35 87.591 ;
               RECT 14.296 88.078 14.35 88.114 ;
               RECT 14.296 88.526 14.35 88.562 ;
               RECT 14.296 88.755 14.35 88.791 ;
               RECT 14.296 89.278 14.35 89.314 ;
               RECT 14.296 89.726 14.35 89.762 ;
               RECT 14.296 89.955 14.35 89.991 ;
               RECT 14.296 90.478 14.35 90.514 ;
               RECT 14.296 90.926 14.35 90.962 ;
               RECT 14.296 91.155 14.35 91.191 ;
               RECT 14.296 91.678 14.35 91.714 ;
               RECT 14.296 92.126 14.35 92.162 ;
               RECT 14.296 92.355 14.35 92.391 ;
               RECT 14.296 92.878 14.35 92.914 ;
               RECT 14.296 93.326 14.35 93.362 ;
               RECT 14.296 93.555 14.35 93.591 ;
               RECT 14.296 94.078 14.35 94.114 ;
               RECT 14.296 94.526 14.35 94.562 ;
               RECT 14.296 94.755 14.35 94.791 ;
               RECT 14.296 95.278 14.35 95.314 ;
               RECT 14.296 95.726 14.35 95.762 ;
               RECT 14.296 95.955 14.35 95.991 ;
               RECT 14.296 96.478 14.35 96.514 ;
               RECT 14.296 96.926 14.35 96.962 ;
               RECT 14.296 97.155 14.35 97.191 ;
               RECT 14.296 97.678 14.35 97.714 ;
               RECT 14.296 98.126 14.35 98.162 ;
               RECT 14.296 98.355 14.35 98.391 ;
               RECT 14.296 98.878 14.35 98.914 ;
               RECT 14.296 99.326 14.35 99.362 ;
               RECT 14.296 99.555 14.35 99.591 ;
               RECT 14.296 100.078 14.35 100.114 ;
               RECT 14.296 100.526 14.35 100.562 ;
               RECT 14.296 100.755 14.35 100.791 ;
               RECT 14.296 101.278 14.35 101.314 ;
               RECT 14.296 101.726 14.35 101.762 ;
               RECT 14.296 101.955 14.35 101.991 ;
               RECT 14.296 102.478 14.35 102.514 ;
               RECT 14.296 102.926 14.35 102.962 ;
               RECT 14.296 103.155 14.35 103.191 ;
               RECT 14.296 103.678 14.35 103.714 ;
               RECT 14.296 104.126 14.35 104.162 ;
               RECT 14.296 104.355 14.35 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 14.932 0.5695 14.986 104.5505 ;
               LAYER v4 ;
               RECT 14.932 0.729 14.986 0.765 ;
               RECT 14.932 0.958 14.986 0.994 ;
               RECT 14.932 1.406 14.986 1.442 ;
               RECT 14.932 1.635 14.986 1.671 ;
               RECT 14.932 1.929 14.986 1.965 ;
               RECT 14.932 2.158 14.986 2.194 ;
               RECT 14.932 2.606 14.986 2.642 ;
               RECT 14.932 2.835 14.986 2.871 ;
               RECT 14.932 3.129 14.986 3.165 ;
               RECT 14.932 3.358 14.986 3.394 ;
               RECT 14.932 3.806 14.986 3.842 ;
               RECT 14.932 4.035 14.986 4.071 ;
               RECT 14.932 4.329 14.986 4.365 ;
               RECT 14.932 4.558 14.986 4.594 ;
               RECT 14.932 5.006 14.986 5.042 ;
               RECT 14.932 5.235 14.986 5.271 ;
               RECT 14.932 5.529 14.986 5.565 ;
               RECT 14.932 5.758 14.986 5.794 ;
               RECT 14.932 6.206 14.986 6.242 ;
               RECT 14.932 6.435 14.986 6.471 ;
               RECT 14.932 6.729 14.986 6.765 ;
               RECT 14.932 6.958 14.986 6.994 ;
               RECT 14.932 7.406 14.986 7.442 ;
               RECT 14.932 7.635 14.986 7.671 ;
               RECT 14.932 7.929 14.986 7.965 ;
               RECT 14.932 8.158 14.986 8.194 ;
               RECT 14.932 8.606 14.986 8.642 ;
               RECT 14.932 8.835 14.986 8.871 ;
               RECT 14.932 9.129 14.986 9.165 ;
               RECT 14.932 9.358 14.986 9.394 ;
               RECT 14.932 9.806 14.986 9.842 ;
               RECT 14.932 10.035 14.986 10.071 ;
               RECT 14.932 10.329 14.986 10.365 ;
               RECT 14.932 10.558 14.986 10.594 ;
               RECT 14.932 11.006 14.986 11.042 ;
               RECT 14.932 11.235 14.986 11.271 ;
               RECT 14.932 11.529 14.986 11.565 ;
               RECT 14.932 11.758 14.986 11.794 ;
               RECT 14.932 12.206 14.986 12.242 ;
               RECT 14.932 12.435 14.986 12.471 ;
               RECT 14.932 12.729 14.986 12.765 ;
               RECT 14.932 12.958 14.986 12.994 ;
               RECT 14.932 13.406 14.986 13.442 ;
               RECT 14.932 13.635 14.986 13.671 ;
               RECT 14.932 13.929 14.986 13.965 ;
               RECT 14.932 14.158 14.986 14.194 ;
               RECT 14.932 14.606 14.986 14.642 ;
               RECT 14.932 14.835 14.986 14.871 ;
               RECT 14.932 15.129 14.986 15.165 ;
               RECT 14.932 15.358 14.986 15.394 ;
               RECT 14.932 15.806 14.986 15.842 ;
               RECT 14.932 16.035 14.986 16.071 ;
               RECT 14.932 16.329 14.986 16.365 ;
               RECT 14.932 16.558 14.986 16.594 ;
               RECT 14.932 17.006 14.986 17.042 ;
               RECT 14.932 17.235 14.986 17.271 ;
               RECT 14.932 17.529 14.986 17.565 ;
               RECT 14.932 17.758 14.986 17.794 ;
               RECT 14.932 18.206 14.986 18.242 ;
               RECT 14.932 18.435 14.986 18.471 ;
               RECT 14.932 18.729 14.986 18.765 ;
               RECT 14.932 18.958 14.986 18.994 ;
               RECT 14.932 19.406 14.986 19.442 ;
               RECT 14.932 19.635 14.986 19.671 ;
               RECT 14.932 19.929 14.986 19.965 ;
               RECT 14.932 20.158 14.986 20.194 ;
               RECT 14.932 20.606 14.986 20.642 ;
               RECT 14.932 20.835 14.986 20.871 ;
               RECT 14.932 21.129 14.986 21.165 ;
               RECT 14.932 21.358 14.986 21.394 ;
               RECT 14.932 21.806 14.986 21.842 ;
               RECT 14.932 22.035 14.986 22.071 ;
               RECT 14.932 22.329 14.986 22.365 ;
               RECT 14.932 22.558 14.986 22.594 ;
               RECT 14.932 23.006 14.986 23.042 ;
               RECT 14.932 23.235 14.986 23.271 ;
               RECT 14.932 23.529 14.986 23.565 ;
               RECT 14.932 23.758 14.986 23.794 ;
               RECT 14.932 24.206 14.986 24.242 ;
               RECT 14.932 24.435 14.986 24.471 ;
               RECT 14.932 24.729 14.986 24.765 ;
               RECT 14.932 24.958 14.986 24.994 ;
               RECT 14.932 25.406 14.986 25.442 ;
               RECT 14.932 25.635 14.986 25.671 ;
               RECT 14.932 25.929 14.986 25.965 ;
               RECT 14.932 26.158 14.986 26.194 ;
               RECT 14.932 26.606 14.986 26.642 ;
               RECT 14.932 26.835 14.986 26.871 ;
               RECT 14.932 27.129 14.986 27.165 ;
               RECT 14.932 27.358 14.986 27.394 ;
               RECT 14.932 27.806 14.986 27.842 ;
               RECT 14.932 28.035 14.986 28.071 ;
               RECT 14.932 28.329 14.986 28.365 ;
               RECT 14.932 28.558 14.986 28.594 ;
               RECT 14.932 29.006 14.986 29.042 ;
               RECT 14.932 29.235 14.986 29.271 ;
               RECT 14.932 29.529 14.986 29.565 ;
               RECT 14.932 29.758 14.986 29.794 ;
               RECT 14.932 30.206 14.986 30.242 ;
               RECT 14.932 30.435 14.986 30.471 ;
               RECT 14.932 30.729 14.986 30.765 ;
               RECT 14.932 30.958 14.986 30.994 ;
               RECT 14.932 31.406 14.986 31.442 ;
               RECT 14.932 31.635 14.986 31.671 ;
               RECT 14.932 31.929 14.986 31.965 ;
               RECT 14.932 32.158 14.986 32.194 ;
               RECT 14.932 32.606 14.986 32.642 ;
               RECT 14.932 32.835 14.986 32.871 ;
               RECT 14.932 33.129 14.986 33.165 ;
               RECT 14.932 33.358 14.986 33.394 ;
               RECT 14.932 33.806 14.986 33.842 ;
               RECT 14.932 34.035 14.986 34.071 ;
               RECT 14.932 34.329 14.986 34.365 ;
               RECT 14.932 34.558 14.986 34.594 ;
               RECT 14.932 35.006 14.986 35.042 ;
               RECT 14.932 35.235 14.986 35.271 ;
               RECT 14.932 35.529 14.986 35.565 ;
               RECT 14.932 35.758 14.986 35.794 ;
               RECT 14.932 36.206 14.986 36.242 ;
               RECT 14.932 36.435 14.986 36.471 ;
               RECT 14.932 36.729 14.986 36.765 ;
               RECT 14.932 36.958 14.986 36.994 ;
               RECT 14.932 37.406 14.986 37.442 ;
               RECT 14.932 37.635 14.986 37.671 ;
               RECT 14.932 37.929 14.986 37.965 ;
               RECT 14.932 38.158 14.986 38.194 ;
               RECT 14.932 38.606 14.986 38.642 ;
               RECT 14.932 38.835 14.986 38.871 ;
               RECT 14.932 39.129 14.986 39.165 ;
               RECT 14.932 39.358 14.986 39.394 ;
               RECT 14.932 39.806 14.986 39.842 ;
               RECT 14.932 40.035 14.986 40.071 ;
               RECT 14.932 40.329 14.986 40.365 ;
               RECT 14.932 40.558 14.986 40.594 ;
               RECT 14.932 41.006 14.986 41.042 ;
               RECT 14.932 41.235 14.986 41.271 ;
               RECT 14.932 41.529 14.986 41.565 ;
               RECT 14.932 41.758 14.986 41.794 ;
               RECT 14.932 42.206 14.986 42.242 ;
               RECT 14.932 42.435 14.986 42.471 ;
               RECT 14.932 42.729 14.986 42.765 ;
               RECT 14.932 42.958 14.986 42.994 ;
               RECT 14.932 43.406 14.986 43.442 ;
               RECT 14.932 43.635 14.986 43.671 ;
               RECT 14.932 43.929 14.986 43.965 ;
               RECT 14.932 44.158 14.986 44.194 ;
               RECT 14.932 44.606 14.986 44.642 ;
               RECT 14.932 44.835 14.986 44.871 ;
               RECT 14.932 45.129 14.986 45.165 ;
               RECT 14.932 45.358 14.986 45.394 ;
               RECT 14.932 45.806 14.986 45.842 ;
               RECT 14.932 46.035 14.986 46.071 ;
               RECT 14.932 46.329 14.986 46.365 ;
               RECT 14.932 46.558 14.986 46.594 ;
               RECT 14.932 47.006 14.986 47.042 ;
               RECT 14.932 47.235 14.986 47.271 ;
               RECT 14.932 47.529 14.986 47.565 ;
               RECT 14.932 47.758 14.986 47.794 ;
               RECT 14.932 48.206 14.986 48.242 ;
               RECT 14.932 48.435 14.986 48.471 ;
               RECT 14.932 49.062 14.986 49.098 ;
               RECT 14.932 49.182 14.986 49.218 ;
               RECT 14.932 49.542 14.986 49.578 ;
               RECT 14.932 49.662 14.986 49.698 ;
               RECT 14.932 49.782 14.986 49.818 ;
               RECT 14.932 50.262 14.986 50.298 ;
               RECT 14.932 50.622 14.986 50.658 ;
               RECT 14.932 51.102 14.986 51.138 ;
               RECT 14.932 51.582 14.986 51.618 ;
               RECT 14.932 52.062 14.986 52.098 ;
               RECT 14.932 52.182 14.986 52.218 ;
               RECT 14.932 52.542 14.986 52.578 ;
               RECT 14.932 52.902 14.986 52.938 ;
               RECT 14.932 53.022 14.986 53.058 ;
               RECT 14.932 53.502 14.986 53.538 ;
               RECT 14.932 53.982 14.986 54.018 ;
               RECT 14.932 54.462 14.986 54.498 ;
               RECT 14.932 54.822 14.986 54.858 ;
               RECT 14.932 54.942 14.986 54.978 ;
               RECT 14.932 55.302 14.986 55.338 ;
               RECT 14.932 55.422 14.986 55.458 ;
               RECT 14.932 55.542 14.986 55.578 ;
               RECT 14.932 55.902 14.986 55.938 ;
               RECT 14.932 56.649 14.986 56.685 ;
               RECT 14.932 56.878 14.986 56.914 ;
               RECT 14.932 57.326 14.986 57.362 ;
               RECT 14.932 57.555 14.986 57.591 ;
               RECT 14.932 57.849 14.986 57.885 ;
               RECT 14.932 58.078 14.986 58.114 ;
               RECT 14.932 58.526 14.986 58.562 ;
               RECT 14.932 58.755 14.986 58.791 ;
               RECT 14.932 59.049 14.986 59.085 ;
               RECT 14.932 59.278 14.986 59.314 ;
               RECT 14.932 59.726 14.986 59.762 ;
               RECT 14.932 59.955 14.986 59.991 ;
               RECT 14.932 60.249 14.986 60.285 ;
               RECT 14.932 60.478 14.986 60.514 ;
               RECT 14.932 60.926 14.986 60.962 ;
               RECT 14.932 61.155 14.986 61.191 ;
               RECT 14.932 61.449 14.986 61.485 ;
               RECT 14.932 61.678 14.986 61.714 ;
               RECT 14.932 62.126 14.986 62.162 ;
               RECT 14.932 62.355 14.986 62.391 ;
               RECT 14.932 62.649 14.986 62.685 ;
               RECT 14.932 62.878 14.986 62.914 ;
               RECT 14.932 63.326 14.986 63.362 ;
               RECT 14.932 63.555 14.986 63.591 ;
               RECT 14.932 63.849 14.986 63.885 ;
               RECT 14.932 64.078 14.986 64.114 ;
               RECT 14.932 64.526 14.986 64.562 ;
               RECT 14.932 64.755 14.986 64.791 ;
               RECT 14.932 65.049 14.986 65.085 ;
               RECT 14.932 65.278 14.986 65.314 ;
               RECT 14.932 65.726 14.986 65.762 ;
               RECT 14.932 65.955 14.986 65.991 ;
               RECT 14.932 66.249 14.986 66.285 ;
               RECT 14.932 66.478 14.986 66.514 ;
               RECT 14.932 66.926 14.986 66.962 ;
               RECT 14.932 67.155 14.986 67.191 ;
               RECT 14.932 67.449 14.986 67.485 ;
               RECT 14.932 67.678 14.986 67.714 ;
               RECT 14.932 68.126 14.986 68.162 ;
               RECT 14.932 68.355 14.986 68.391 ;
               RECT 14.932 68.649 14.986 68.685 ;
               RECT 14.932 68.878 14.986 68.914 ;
               RECT 14.932 69.326 14.986 69.362 ;
               RECT 14.932 69.555 14.986 69.591 ;
               RECT 14.932 69.849 14.986 69.885 ;
               RECT 14.932 70.078 14.986 70.114 ;
               RECT 14.932 70.526 14.986 70.562 ;
               RECT 14.932 70.755 14.986 70.791 ;
               RECT 14.932 71.049 14.986 71.085 ;
               RECT 14.932 71.278 14.986 71.314 ;
               RECT 14.932 71.726 14.986 71.762 ;
               RECT 14.932 71.955 14.986 71.991 ;
               RECT 14.932 72.249 14.986 72.285 ;
               RECT 14.932 72.478 14.986 72.514 ;
               RECT 14.932 72.926 14.986 72.962 ;
               RECT 14.932 73.155 14.986 73.191 ;
               RECT 14.932 73.449 14.986 73.485 ;
               RECT 14.932 73.678 14.986 73.714 ;
               RECT 14.932 74.126 14.986 74.162 ;
               RECT 14.932 74.355 14.986 74.391 ;
               RECT 14.932 74.649 14.986 74.685 ;
               RECT 14.932 74.878 14.986 74.914 ;
               RECT 14.932 75.326 14.986 75.362 ;
               RECT 14.932 75.555 14.986 75.591 ;
               RECT 14.932 75.849 14.986 75.885 ;
               RECT 14.932 76.078 14.986 76.114 ;
               RECT 14.932 76.526 14.986 76.562 ;
               RECT 14.932 76.755 14.986 76.791 ;
               RECT 14.932 77.049 14.986 77.085 ;
               RECT 14.932 77.278 14.986 77.314 ;
               RECT 14.932 77.726 14.986 77.762 ;
               RECT 14.932 77.955 14.986 77.991 ;
               RECT 14.932 78.249 14.986 78.285 ;
               RECT 14.932 78.478 14.986 78.514 ;
               RECT 14.932 78.926 14.986 78.962 ;
               RECT 14.932 79.155 14.986 79.191 ;
               RECT 14.932 79.449 14.986 79.485 ;
               RECT 14.932 79.678 14.986 79.714 ;
               RECT 14.932 80.126 14.986 80.162 ;
               RECT 14.932 80.355 14.986 80.391 ;
               RECT 14.932 80.649 14.986 80.685 ;
               RECT 14.932 80.878 14.986 80.914 ;
               RECT 14.932 81.326 14.986 81.362 ;
               RECT 14.932 81.555 14.986 81.591 ;
               RECT 14.932 81.849 14.986 81.885 ;
               RECT 14.932 82.078 14.986 82.114 ;
               RECT 14.932 82.526 14.986 82.562 ;
               RECT 14.932 82.755 14.986 82.791 ;
               RECT 14.932 83.049 14.986 83.085 ;
               RECT 14.932 83.278 14.986 83.314 ;
               RECT 14.932 83.726 14.986 83.762 ;
               RECT 14.932 83.955 14.986 83.991 ;
               RECT 14.932 84.249 14.986 84.285 ;
               RECT 14.932 84.478 14.986 84.514 ;
               RECT 14.932 84.926 14.986 84.962 ;
               RECT 14.932 85.155 14.986 85.191 ;
               RECT 14.932 85.449 14.986 85.485 ;
               RECT 14.932 85.678 14.986 85.714 ;
               RECT 14.932 86.126 14.986 86.162 ;
               RECT 14.932 86.355 14.986 86.391 ;
               RECT 14.932 86.649 14.986 86.685 ;
               RECT 14.932 86.878 14.986 86.914 ;
               RECT 14.932 87.326 14.986 87.362 ;
               RECT 14.932 87.555 14.986 87.591 ;
               RECT 14.932 87.849 14.986 87.885 ;
               RECT 14.932 88.078 14.986 88.114 ;
               RECT 14.932 88.526 14.986 88.562 ;
               RECT 14.932 88.755 14.986 88.791 ;
               RECT 14.932 89.049 14.986 89.085 ;
               RECT 14.932 89.278 14.986 89.314 ;
               RECT 14.932 89.726 14.986 89.762 ;
               RECT 14.932 89.955 14.986 89.991 ;
               RECT 14.932 90.249 14.986 90.285 ;
               RECT 14.932 90.478 14.986 90.514 ;
               RECT 14.932 90.926 14.986 90.962 ;
               RECT 14.932 91.155 14.986 91.191 ;
               RECT 14.932 91.449 14.986 91.485 ;
               RECT 14.932 91.678 14.986 91.714 ;
               RECT 14.932 92.126 14.986 92.162 ;
               RECT 14.932 92.355 14.986 92.391 ;
               RECT 14.932 92.649 14.986 92.685 ;
               RECT 14.932 92.878 14.986 92.914 ;
               RECT 14.932 93.326 14.986 93.362 ;
               RECT 14.932 93.555 14.986 93.591 ;
               RECT 14.932 93.849 14.986 93.885 ;
               RECT 14.932 94.078 14.986 94.114 ;
               RECT 14.932 94.526 14.986 94.562 ;
               RECT 14.932 94.755 14.986 94.791 ;
               RECT 14.932 95.049 14.986 95.085 ;
               RECT 14.932 95.278 14.986 95.314 ;
               RECT 14.932 95.726 14.986 95.762 ;
               RECT 14.932 95.955 14.986 95.991 ;
               RECT 14.932 96.249 14.986 96.285 ;
               RECT 14.932 96.478 14.986 96.514 ;
               RECT 14.932 96.926 14.986 96.962 ;
               RECT 14.932 97.155 14.986 97.191 ;
               RECT 14.932 97.449 14.986 97.485 ;
               RECT 14.932 97.678 14.986 97.714 ;
               RECT 14.932 98.126 14.986 98.162 ;
               RECT 14.932 98.355 14.986 98.391 ;
               RECT 14.932 98.649 14.986 98.685 ;
               RECT 14.932 98.878 14.986 98.914 ;
               RECT 14.932 99.326 14.986 99.362 ;
               RECT 14.932 99.555 14.986 99.591 ;
               RECT 14.932 99.849 14.986 99.885 ;
               RECT 14.932 100.078 14.986 100.114 ;
               RECT 14.932 100.526 14.986 100.562 ;
               RECT 14.932 100.755 14.986 100.791 ;
               RECT 14.932 101.049 14.986 101.085 ;
               RECT 14.932 101.278 14.986 101.314 ;
               RECT 14.932 101.726 14.986 101.762 ;
               RECT 14.932 101.955 14.986 101.991 ;
               RECT 14.932 102.249 14.986 102.285 ;
               RECT 14.932 102.478 14.986 102.514 ;
               RECT 14.932 102.926 14.986 102.962 ;
               RECT 14.932 103.155 14.986 103.191 ;
               RECT 14.932 103.449 14.986 103.485 ;
               RECT 14.932 103.678 14.986 103.714 ;
               RECT 14.932 104.126 14.986 104.162 ;
               RECT 14.932 104.355 14.986 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.318 0.5695 15.37 104.5505 ;
               LAYER v4 ;
               RECT 15.318 0.729 15.37 0.765 ;
               RECT 15.318 0.958 15.37 0.994 ;
               RECT 15.318 1.406 15.37 1.442 ;
               RECT 15.318 1.635 15.37 1.671 ;
               RECT 15.318 1.929 15.37 1.965 ;
               RECT 15.318 2.158 15.37 2.194 ;
               RECT 15.318 2.606 15.37 2.642 ;
               RECT 15.318 2.835 15.37 2.871 ;
               RECT 15.318 3.129 15.37 3.165 ;
               RECT 15.318 3.358 15.37 3.394 ;
               RECT 15.318 3.806 15.37 3.842 ;
               RECT 15.318 4.035 15.37 4.071 ;
               RECT 15.318 4.329 15.37 4.365 ;
               RECT 15.318 4.558 15.37 4.594 ;
               RECT 15.318 5.006 15.37 5.042 ;
               RECT 15.318 5.235 15.37 5.271 ;
               RECT 15.318 5.529 15.37 5.565 ;
               RECT 15.318 5.758 15.37 5.794 ;
               RECT 15.318 6.206 15.37 6.242 ;
               RECT 15.318 6.435 15.37 6.471 ;
               RECT 15.318 6.729 15.37 6.765 ;
               RECT 15.318 6.958 15.37 6.994 ;
               RECT 15.318 7.406 15.37 7.442 ;
               RECT 15.318 7.635 15.37 7.671 ;
               RECT 15.318 7.929 15.37 7.965 ;
               RECT 15.318 8.158 15.37 8.194 ;
               RECT 15.318 8.606 15.37 8.642 ;
               RECT 15.318 8.835 15.37 8.871 ;
               RECT 15.318 9.129 15.37 9.165 ;
               RECT 15.318 9.358 15.37 9.394 ;
               RECT 15.318 9.806 15.37 9.842 ;
               RECT 15.318 10.035 15.37 10.071 ;
               RECT 15.318 10.329 15.37 10.365 ;
               RECT 15.318 10.558 15.37 10.594 ;
               RECT 15.318 11.006 15.37 11.042 ;
               RECT 15.318 11.235 15.37 11.271 ;
               RECT 15.318 11.529 15.37 11.565 ;
               RECT 15.318 11.758 15.37 11.794 ;
               RECT 15.318 12.206 15.37 12.242 ;
               RECT 15.318 12.435 15.37 12.471 ;
               RECT 15.318 12.729 15.37 12.765 ;
               RECT 15.318 12.958 15.37 12.994 ;
               RECT 15.318 13.406 15.37 13.442 ;
               RECT 15.318 13.635 15.37 13.671 ;
               RECT 15.318 13.929 15.37 13.965 ;
               RECT 15.318 14.158 15.37 14.194 ;
               RECT 15.318 14.606 15.37 14.642 ;
               RECT 15.318 14.835 15.37 14.871 ;
               RECT 15.318 15.129 15.37 15.165 ;
               RECT 15.318 15.358 15.37 15.394 ;
               RECT 15.318 15.806 15.37 15.842 ;
               RECT 15.318 16.035 15.37 16.071 ;
               RECT 15.318 16.329 15.37 16.365 ;
               RECT 15.318 16.558 15.37 16.594 ;
               RECT 15.318 17.006 15.37 17.042 ;
               RECT 15.318 17.235 15.37 17.271 ;
               RECT 15.318 17.529 15.37 17.565 ;
               RECT 15.318 17.758 15.37 17.794 ;
               RECT 15.318 18.206 15.37 18.242 ;
               RECT 15.318 18.435 15.37 18.471 ;
               RECT 15.318 18.729 15.37 18.765 ;
               RECT 15.318 18.958 15.37 18.994 ;
               RECT 15.318 19.406 15.37 19.442 ;
               RECT 15.318 19.635 15.37 19.671 ;
               RECT 15.318 19.929 15.37 19.965 ;
               RECT 15.318 20.158 15.37 20.194 ;
               RECT 15.318 20.606 15.37 20.642 ;
               RECT 15.318 20.835 15.37 20.871 ;
               RECT 15.318 21.129 15.37 21.165 ;
               RECT 15.318 21.358 15.37 21.394 ;
               RECT 15.318 21.806 15.37 21.842 ;
               RECT 15.318 22.035 15.37 22.071 ;
               RECT 15.318 22.329 15.37 22.365 ;
               RECT 15.318 22.558 15.37 22.594 ;
               RECT 15.318 23.006 15.37 23.042 ;
               RECT 15.318 23.235 15.37 23.271 ;
               RECT 15.318 23.529 15.37 23.565 ;
               RECT 15.318 23.758 15.37 23.794 ;
               RECT 15.318 24.206 15.37 24.242 ;
               RECT 15.318 24.435 15.37 24.471 ;
               RECT 15.318 24.729 15.37 24.765 ;
               RECT 15.318 24.958 15.37 24.994 ;
               RECT 15.318 25.406 15.37 25.442 ;
               RECT 15.318 25.635 15.37 25.671 ;
               RECT 15.318 25.929 15.37 25.965 ;
               RECT 15.318 26.158 15.37 26.194 ;
               RECT 15.318 26.606 15.37 26.642 ;
               RECT 15.318 26.835 15.37 26.871 ;
               RECT 15.318 27.129 15.37 27.165 ;
               RECT 15.318 27.358 15.37 27.394 ;
               RECT 15.318 27.806 15.37 27.842 ;
               RECT 15.318 28.035 15.37 28.071 ;
               RECT 15.318 28.329 15.37 28.365 ;
               RECT 15.318 28.558 15.37 28.594 ;
               RECT 15.318 29.006 15.37 29.042 ;
               RECT 15.318 29.235 15.37 29.271 ;
               RECT 15.318 29.529 15.37 29.565 ;
               RECT 15.318 29.758 15.37 29.794 ;
               RECT 15.318 30.206 15.37 30.242 ;
               RECT 15.318 30.435 15.37 30.471 ;
               RECT 15.318 30.729 15.37 30.765 ;
               RECT 15.318 30.958 15.37 30.994 ;
               RECT 15.318 31.406 15.37 31.442 ;
               RECT 15.318 31.635 15.37 31.671 ;
               RECT 15.318 31.929 15.37 31.965 ;
               RECT 15.318 32.158 15.37 32.194 ;
               RECT 15.318 32.606 15.37 32.642 ;
               RECT 15.318 32.835 15.37 32.871 ;
               RECT 15.318 33.129 15.37 33.165 ;
               RECT 15.318 33.358 15.37 33.394 ;
               RECT 15.318 33.806 15.37 33.842 ;
               RECT 15.318 34.035 15.37 34.071 ;
               RECT 15.318 34.329 15.37 34.365 ;
               RECT 15.318 34.558 15.37 34.594 ;
               RECT 15.318 35.006 15.37 35.042 ;
               RECT 15.318 35.235 15.37 35.271 ;
               RECT 15.318 35.529 15.37 35.565 ;
               RECT 15.318 35.758 15.37 35.794 ;
               RECT 15.318 36.206 15.37 36.242 ;
               RECT 15.318 36.435 15.37 36.471 ;
               RECT 15.318 36.729 15.37 36.765 ;
               RECT 15.318 36.958 15.37 36.994 ;
               RECT 15.318 37.406 15.37 37.442 ;
               RECT 15.318 37.635 15.37 37.671 ;
               RECT 15.318 37.929 15.37 37.965 ;
               RECT 15.318 38.158 15.37 38.194 ;
               RECT 15.318 38.606 15.37 38.642 ;
               RECT 15.318 38.835 15.37 38.871 ;
               RECT 15.318 39.129 15.37 39.165 ;
               RECT 15.318 39.358 15.37 39.394 ;
               RECT 15.318 39.806 15.37 39.842 ;
               RECT 15.318 40.035 15.37 40.071 ;
               RECT 15.318 40.329 15.37 40.365 ;
               RECT 15.318 40.558 15.37 40.594 ;
               RECT 15.318 41.006 15.37 41.042 ;
               RECT 15.318 41.235 15.37 41.271 ;
               RECT 15.318 41.529 15.37 41.565 ;
               RECT 15.318 41.758 15.37 41.794 ;
               RECT 15.318 42.206 15.37 42.242 ;
               RECT 15.318 42.435 15.37 42.471 ;
               RECT 15.318 42.729 15.37 42.765 ;
               RECT 15.318 42.958 15.37 42.994 ;
               RECT 15.318 43.406 15.37 43.442 ;
               RECT 15.318 43.635 15.37 43.671 ;
               RECT 15.318 43.929 15.37 43.965 ;
               RECT 15.318 44.158 15.37 44.194 ;
               RECT 15.318 44.606 15.37 44.642 ;
               RECT 15.318 44.835 15.37 44.871 ;
               RECT 15.318 45.129 15.37 45.165 ;
               RECT 15.318 45.358 15.37 45.394 ;
               RECT 15.318 45.806 15.37 45.842 ;
               RECT 15.318 46.035 15.37 46.071 ;
               RECT 15.318 46.329 15.37 46.365 ;
               RECT 15.318 46.558 15.37 46.594 ;
               RECT 15.318 47.006 15.37 47.042 ;
               RECT 15.318 47.235 15.37 47.271 ;
               RECT 15.318 47.529 15.37 47.565 ;
               RECT 15.318 47.758 15.37 47.794 ;
               RECT 15.318 48.206 15.37 48.242 ;
               RECT 15.318 48.435 15.37 48.471 ;
               RECT 15.318 49.182 15.37 49.218 ;
               RECT 15.318 49.662 15.37 49.698 ;
               RECT 15.318 49.8435 15.37 49.8795 ;
               RECT 15.318 50.142 15.37 50.178 ;
               RECT 15.318 50.622 15.37 50.658 ;
               RECT 15.318 51.102 15.37 51.138 ;
               RECT 15.318 51.582 15.37 51.618 ;
               RECT 15.318 52.062 15.37 52.098 ;
               RECT 15.318 52.542 15.37 52.578 ;
               RECT 15.318 53.022 15.37 53.058 ;
               RECT 15.318 53.502 15.37 53.538 ;
               RECT 15.318 53.982 15.37 54.018 ;
               RECT 15.318 54.4675 15.37 54.4925 ;
               RECT 15.318 54.942 15.37 54.978 ;
               RECT 15.318 55.422 15.37 55.458 ;
               RECT 15.318 55.902 15.37 55.938 ;
               RECT 15.318 56.649 15.37 56.685 ;
               RECT 15.318 56.878 15.37 56.914 ;
               RECT 15.318 57.326 15.37 57.362 ;
               RECT 15.318 57.555 15.37 57.591 ;
               RECT 15.318 57.849 15.37 57.885 ;
               RECT 15.318 58.078 15.37 58.114 ;
               RECT 15.318 58.526 15.37 58.562 ;
               RECT 15.318 58.755 15.37 58.791 ;
               RECT 15.318 59.049 15.37 59.085 ;
               RECT 15.318 59.278 15.37 59.314 ;
               RECT 15.318 59.726 15.37 59.762 ;
               RECT 15.318 59.955 15.37 59.991 ;
               RECT 15.318 60.249 15.37 60.285 ;
               RECT 15.318 60.478 15.37 60.514 ;
               RECT 15.318 60.926 15.37 60.962 ;
               RECT 15.318 61.155 15.37 61.191 ;
               RECT 15.318 61.449 15.37 61.485 ;
               RECT 15.318 61.678 15.37 61.714 ;
               RECT 15.318 62.126 15.37 62.162 ;
               RECT 15.318 62.355 15.37 62.391 ;
               RECT 15.318 62.649 15.37 62.685 ;
               RECT 15.318 62.878 15.37 62.914 ;
               RECT 15.318 63.326 15.37 63.362 ;
               RECT 15.318 63.555 15.37 63.591 ;
               RECT 15.318 63.849 15.37 63.885 ;
               RECT 15.318 64.078 15.37 64.114 ;
               RECT 15.318 64.526 15.37 64.562 ;
               RECT 15.318 64.755 15.37 64.791 ;
               RECT 15.318 65.049 15.37 65.085 ;
               RECT 15.318 65.278 15.37 65.314 ;
               RECT 15.318 65.726 15.37 65.762 ;
               RECT 15.318 65.955 15.37 65.991 ;
               RECT 15.318 66.249 15.37 66.285 ;
               RECT 15.318 66.478 15.37 66.514 ;
               RECT 15.318 66.926 15.37 66.962 ;
               RECT 15.318 67.155 15.37 67.191 ;
               RECT 15.318 67.449 15.37 67.485 ;
               RECT 15.318 67.678 15.37 67.714 ;
               RECT 15.318 68.126 15.37 68.162 ;
               RECT 15.318 68.355 15.37 68.391 ;
               RECT 15.318 68.649 15.37 68.685 ;
               RECT 15.318 68.878 15.37 68.914 ;
               RECT 15.318 69.326 15.37 69.362 ;
               RECT 15.318 69.555 15.37 69.591 ;
               RECT 15.318 69.849 15.37 69.885 ;
               RECT 15.318 70.078 15.37 70.114 ;
               RECT 15.318 70.526 15.37 70.562 ;
               RECT 15.318 70.755 15.37 70.791 ;
               RECT 15.318 71.049 15.37 71.085 ;
               RECT 15.318 71.278 15.37 71.314 ;
               RECT 15.318 71.726 15.37 71.762 ;
               RECT 15.318 71.955 15.37 71.991 ;
               RECT 15.318 72.249 15.37 72.285 ;
               RECT 15.318 72.478 15.37 72.514 ;
               RECT 15.318 72.926 15.37 72.962 ;
               RECT 15.318 73.155 15.37 73.191 ;
               RECT 15.318 73.449 15.37 73.485 ;
               RECT 15.318 73.678 15.37 73.714 ;
               RECT 15.318 74.126 15.37 74.162 ;
               RECT 15.318 74.355 15.37 74.391 ;
               RECT 15.318 74.649 15.37 74.685 ;
               RECT 15.318 74.878 15.37 74.914 ;
               RECT 15.318 75.326 15.37 75.362 ;
               RECT 15.318 75.555 15.37 75.591 ;
               RECT 15.318 75.849 15.37 75.885 ;
               RECT 15.318 76.078 15.37 76.114 ;
               RECT 15.318 76.526 15.37 76.562 ;
               RECT 15.318 76.755 15.37 76.791 ;
               RECT 15.318 77.049 15.37 77.085 ;
               RECT 15.318 77.278 15.37 77.314 ;
               RECT 15.318 77.726 15.37 77.762 ;
               RECT 15.318 77.955 15.37 77.991 ;
               RECT 15.318 78.249 15.37 78.285 ;
               RECT 15.318 78.478 15.37 78.514 ;
               RECT 15.318 78.926 15.37 78.962 ;
               RECT 15.318 79.155 15.37 79.191 ;
               RECT 15.318 79.449 15.37 79.485 ;
               RECT 15.318 79.678 15.37 79.714 ;
               RECT 15.318 80.126 15.37 80.162 ;
               RECT 15.318 80.355 15.37 80.391 ;
               RECT 15.318 80.649 15.37 80.685 ;
               RECT 15.318 80.878 15.37 80.914 ;
               RECT 15.318 81.326 15.37 81.362 ;
               RECT 15.318 81.555 15.37 81.591 ;
               RECT 15.318 81.849 15.37 81.885 ;
               RECT 15.318 82.078 15.37 82.114 ;
               RECT 15.318 82.526 15.37 82.562 ;
               RECT 15.318 82.755 15.37 82.791 ;
               RECT 15.318 83.049 15.37 83.085 ;
               RECT 15.318 83.278 15.37 83.314 ;
               RECT 15.318 83.726 15.37 83.762 ;
               RECT 15.318 83.955 15.37 83.991 ;
               RECT 15.318 84.249 15.37 84.285 ;
               RECT 15.318 84.478 15.37 84.514 ;
               RECT 15.318 84.926 15.37 84.962 ;
               RECT 15.318 85.155 15.37 85.191 ;
               RECT 15.318 85.449 15.37 85.485 ;
               RECT 15.318 85.678 15.37 85.714 ;
               RECT 15.318 86.126 15.37 86.162 ;
               RECT 15.318 86.355 15.37 86.391 ;
               RECT 15.318 86.649 15.37 86.685 ;
               RECT 15.318 86.878 15.37 86.914 ;
               RECT 15.318 87.326 15.37 87.362 ;
               RECT 15.318 87.555 15.37 87.591 ;
               RECT 15.318 87.849 15.37 87.885 ;
               RECT 15.318 88.078 15.37 88.114 ;
               RECT 15.318 88.526 15.37 88.562 ;
               RECT 15.318 88.755 15.37 88.791 ;
               RECT 15.318 89.049 15.37 89.085 ;
               RECT 15.318 89.278 15.37 89.314 ;
               RECT 15.318 89.726 15.37 89.762 ;
               RECT 15.318 89.955 15.37 89.991 ;
               RECT 15.318 90.249 15.37 90.285 ;
               RECT 15.318 90.478 15.37 90.514 ;
               RECT 15.318 90.926 15.37 90.962 ;
               RECT 15.318 91.155 15.37 91.191 ;
               RECT 15.318 91.449 15.37 91.485 ;
               RECT 15.318 91.678 15.37 91.714 ;
               RECT 15.318 92.126 15.37 92.162 ;
               RECT 15.318 92.355 15.37 92.391 ;
               RECT 15.318 92.649 15.37 92.685 ;
               RECT 15.318 92.878 15.37 92.914 ;
               RECT 15.318 93.326 15.37 93.362 ;
               RECT 15.318 93.555 15.37 93.591 ;
               RECT 15.318 93.849 15.37 93.885 ;
               RECT 15.318 94.078 15.37 94.114 ;
               RECT 15.318 94.526 15.37 94.562 ;
               RECT 15.318 94.755 15.37 94.791 ;
               RECT 15.318 95.049 15.37 95.085 ;
               RECT 15.318 95.278 15.37 95.314 ;
               RECT 15.318 95.726 15.37 95.762 ;
               RECT 15.318 95.955 15.37 95.991 ;
               RECT 15.318 96.249 15.37 96.285 ;
               RECT 15.318 96.478 15.37 96.514 ;
               RECT 15.318 96.926 15.37 96.962 ;
               RECT 15.318 97.155 15.37 97.191 ;
               RECT 15.318 97.449 15.37 97.485 ;
               RECT 15.318 97.678 15.37 97.714 ;
               RECT 15.318 98.126 15.37 98.162 ;
               RECT 15.318 98.355 15.37 98.391 ;
               RECT 15.318 98.649 15.37 98.685 ;
               RECT 15.318 98.878 15.37 98.914 ;
               RECT 15.318 99.326 15.37 99.362 ;
               RECT 15.318 99.555 15.37 99.591 ;
               RECT 15.318 99.849 15.37 99.885 ;
               RECT 15.318 100.078 15.37 100.114 ;
               RECT 15.318 100.526 15.37 100.562 ;
               RECT 15.318 100.755 15.37 100.791 ;
               RECT 15.318 101.049 15.37 101.085 ;
               RECT 15.318 101.278 15.37 101.314 ;
               RECT 15.318 101.726 15.37 101.762 ;
               RECT 15.318 101.955 15.37 101.991 ;
               RECT 15.318 102.249 15.37 102.285 ;
               RECT 15.318 102.478 15.37 102.514 ;
               RECT 15.318 102.926 15.37 102.962 ;
               RECT 15.318 103.155 15.37 103.191 ;
               RECT 15.318 103.449 15.37 103.485 ;
               RECT 15.318 103.678 15.37 103.714 ;
               RECT 15.318 104.126 15.37 104.162 ;
               RECT 15.318 104.355 15.37 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.478 0.5695 15.53 49.6595 ;
               LAYER v4 ;
               RECT 15.478 0.729 15.53 0.765 ;
               RECT 15.478 0.958 15.53 0.994 ;
               RECT 15.478 1.635 15.53 1.671 ;
               RECT 15.478 1.929 15.53 1.965 ;
               RECT 15.478 2.158 15.53 2.194 ;
               RECT 15.478 2.835 15.53 2.871 ;
               RECT 15.478 3.129 15.53 3.165 ;
               RECT 15.478 3.358 15.53 3.394 ;
               RECT 15.478 4.035 15.53 4.071 ;
               RECT 15.478 4.329 15.53 4.365 ;
               RECT 15.478 4.558 15.53 4.594 ;
               RECT 15.478 5.235 15.53 5.271 ;
               RECT 15.478 5.529 15.53 5.565 ;
               RECT 15.478 5.758 15.53 5.794 ;
               RECT 15.478 6.435 15.53 6.471 ;
               RECT 15.478 6.729 15.53 6.765 ;
               RECT 15.478 6.958 15.53 6.994 ;
               RECT 15.478 7.635 15.53 7.671 ;
               RECT 15.478 7.929 15.53 7.965 ;
               RECT 15.478 8.158 15.53 8.194 ;
               RECT 15.478 8.835 15.53 8.871 ;
               RECT 15.478 9.129 15.53 9.165 ;
               RECT 15.478 9.358 15.53 9.394 ;
               RECT 15.478 10.035 15.53 10.071 ;
               RECT 15.478 10.329 15.53 10.365 ;
               RECT 15.478 10.558 15.53 10.594 ;
               RECT 15.478 11.235 15.53 11.271 ;
               RECT 15.478 11.529 15.53 11.565 ;
               RECT 15.478 11.758 15.53 11.794 ;
               RECT 15.478 12.435 15.53 12.471 ;
               RECT 15.478 12.729 15.53 12.765 ;
               RECT 15.478 12.958 15.53 12.994 ;
               RECT 15.478 13.635 15.53 13.671 ;
               RECT 15.478 13.929 15.53 13.965 ;
               RECT 15.478 14.158 15.53 14.194 ;
               RECT 15.478 14.835 15.53 14.871 ;
               RECT 15.478 15.129 15.53 15.165 ;
               RECT 15.478 15.358 15.53 15.394 ;
               RECT 15.478 16.035 15.53 16.071 ;
               RECT 15.478 16.329 15.53 16.365 ;
               RECT 15.478 16.558 15.53 16.594 ;
               RECT 15.478 17.235 15.53 17.271 ;
               RECT 15.478 17.529 15.53 17.565 ;
               RECT 15.478 17.758 15.53 17.794 ;
               RECT 15.478 18.435 15.53 18.471 ;
               RECT 15.478 18.729 15.53 18.765 ;
               RECT 15.478 18.958 15.53 18.994 ;
               RECT 15.478 19.635 15.53 19.671 ;
               RECT 15.478 19.929 15.53 19.965 ;
               RECT 15.478 20.158 15.53 20.194 ;
               RECT 15.478 20.835 15.53 20.871 ;
               RECT 15.478 21.129 15.53 21.165 ;
               RECT 15.478 21.358 15.53 21.394 ;
               RECT 15.478 22.035 15.53 22.071 ;
               RECT 15.478 22.329 15.53 22.365 ;
               RECT 15.478 22.558 15.53 22.594 ;
               RECT 15.478 23.235 15.53 23.271 ;
               RECT 15.478 23.529 15.53 23.565 ;
               RECT 15.478 23.758 15.53 23.794 ;
               RECT 15.478 24.435 15.53 24.471 ;
               RECT 15.478 24.729 15.53 24.765 ;
               RECT 15.478 24.958 15.53 24.994 ;
               RECT 15.478 25.635 15.53 25.671 ;
               RECT 15.478 25.929 15.53 25.965 ;
               RECT 15.478 26.158 15.53 26.194 ;
               RECT 15.478 26.835 15.53 26.871 ;
               RECT 15.478 27.129 15.53 27.165 ;
               RECT 15.478 27.358 15.53 27.394 ;
               RECT 15.478 28.035 15.53 28.071 ;
               RECT 15.478 28.329 15.53 28.365 ;
               RECT 15.478 28.558 15.53 28.594 ;
               RECT 15.478 29.235 15.53 29.271 ;
               RECT 15.478 29.529 15.53 29.565 ;
               RECT 15.478 29.758 15.53 29.794 ;
               RECT 15.478 30.435 15.53 30.471 ;
               RECT 15.478 30.729 15.53 30.765 ;
               RECT 15.478 30.958 15.53 30.994 ;
               RECT 15.478 31.635 15.53 31.671 ;
               RECT 15.478 31.929 15.53 31.965 ;
               RECT 15.478 32.158 15.53 32.194 ;
               RECT 15.478 32.835 15.53 32.871 ;
               RECT 15.478 33.129 15.53 33.165 ;
               RECT 15.478 33.358 15.53 33.394 ;
               RECT 15.478 34.035 15.53 34.071 ;
               RECT 15.478 34.329 15.53 34.365 ;
               RECT 15.478 34.558 15.53 34.594 ;
               RECT 15.478 35.235 15.53 35.271 ;
               RECT 15.478 35.529 15.53 35.565 ;
               RECT 15.478 35.758 15.53 35.794 ;
               RECT 15.478 36.435 15.53 36.471 ;
               RECT 15.478 36.729 15.53 36.765 ;
               RECT 15.478 36.958 15.53 36.994 ;
               RECT 15.478 37.635 15.53 37.671 ;
               RECT 15.478 37.929 15.53 37.965 ;
               RECT 15.478 38.158 15.53 38.194 ;
               RECT 15.478 38.835 15.53 38.871 ;
               RECT 15.478 39.129 15.53 39.165 ;
               RECT 15.478 39.358 15.53 39.394 ;
               RECT 15.478 40.035 15.53 40.071 ;
               RECT 15.478 40.329 15.53 40.365 ;
               RECT 15.478 40.558 15.53 40.594 ;
               RECT 15.478 41.235 15.53 41.271 ;
               RECT 15.478 41.529 15.53 41.565 ;
               RECT 15.478 41.758 15.53 41.794 ;
               RECT 15.478 42.435 15.53 42.471 ;
               RECT 15.478 42.729 15.53 42.765 ;
               RECT 15.478 42.958 15.53 42.994 ;
               RECT 15.478 43.635 15.53 43.671 ;
               RECT 15.478 43.929 15.53 43.965 ;
               RECT 15.478 44.158 15.53 44.194 ;
               RECT 15.478 44.835 15.53 44.871 ;
               RECT 15.478 45.129 15.53 45.165 ;
               RECT 15.478 45.358 15.53 45.394 ;
               RECT 15.478 46.035 15.53 46.071 ;
               RECT 15.478 46.329 15.53 46.365 ;
               RECT 15.478 46.558 15.53 46.594 ;
               RECT 15.478 47.235 15.53 47.271 ;
               RECT 15.478 47.529 15.53 47.565 ;
               RECT 15.478 47.758 15.53 47.794 ;
               RECT 15.478 48.435 15.53 48.471 ;
               RECT 15.478 49.182 15.53 49.218 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.478 54.999 15.53 104.5505 ;
               LAYER v4 ;
               RECT 15.478 55.422 15.53 55.458 ;
               RECT 15.478 55.902 15.53 55.938 ;
               RECT 15.478 56.649 15.53 56.685 ;
               RECT 15.478 56.878 15.53 56.914 ;
               RECT 15.478 57.555 15.53 57.591 ;
               RECT 15.478 57.849 15.53 57.885 ;
               RECT 15.478 58.078 15.53 58.114 ;
               RECT 15.478 58.755 15.53 58.791 ;
               RECT 15.478 59.049 15.53 59.085 ;
               RECT 15.478 59.278 15.53 59.314 ;
               RECT 15.478 59.955 15.53 59.991 ;
               RECT 15.478 60.249 15.53 60.285 ;
               RECT 15.478 60.478 15.53 60.514 ;
               RECT 15.478 61.155 15.53 61.191 ;
               RECT 15.478 61.449 15.53 61.485 ;
               RECT 15.478 61.678 15.53 61.714 ;
               RECT 15.478 62.355 15.53 62.391 ;
               RECT 15.478 62.649 15.53 62.685 ;
               RECT 15.478 62.878 15.53 62.914 ;
               RECT 15.478 63.555 15.53 63.591 ;
               RECT 15.478 63.849 15.53 63.885 ;
               RECT 15.478 64.078 15.53 64.114 ;
               RECT 15.478 64.755 15.53 64.791 ;
               RECT 15.478 65.049 15.53 65.085 ;
               RECT 15.478 65.278 15.53 65.314 ;
               RECT 15.478 65.955 15.53 65.991 ;
               RECT 15.478 66.249 15.53 66.285 ;
               RECT 15.478 66.478 15.53 66.514 ;
               RECT 15.478 67.155 15.53 67.191 ;
               RECT 15.478 67.449 15.53 67.485 ;
               RECT 15.478 67.678 15.53 67.714 ;
               RECT 15.478 68.355 15.53 68.391 ;
               RECT 15.478 68.649 15.53 68.685 ;
               RECT 15.478 68.878 15.53 68.914 ;
               RECT 15.478 69.555 15.53 69.591 ;
               RECT 15.478 69.849 15.53 69.885 ;
               RECT 15.478 70.078 15.53 70.114 ;
               RECT 15.478 70.755 15.53 70.791 ;
               RECT 15.478 71.049 15.53 71.085 ;
               RECT 15.478 71.278 15.53 71.314 ;
               RECT 15.478 71.955 15.53 71.991 ;
               RECT 15.478 72.249 15.53 72.285 ;
               RECT 15.478 72.478 15.53 72.514 ;
               RECT 15.478 73.155 15.53 73.191 ;
               RECT 15.478 73.449 15.53 73.485 ;
               RECT 15.478 73.678 15.53 73.714 ;
               RECT 15.478 74.355 15.53 74.391 ;
               RECT 15.478 74.649 15.53 74.685 ;
               RECT 15.478 74.878 15.53 74.914 ;
               RECT 15.478 75.555 15.53 75.591 ;
               RECT 15.478 75.849 15.53 75.885 ;
               RECT 15.478 76.078 15.53 76.114 ;
               RECT 15.478 76.755 15.53 76.791 ;
               RECT 15.478 77.049 15.53 77.085 ;
               RECT 15.478 77.278 15.53 77.314 ;
               RECT 15.478 77.955 15.53 77.991 ;
               RECT 15.478 78.249 15.53 78.285 ;
               RECT 15.478 78.478 15.53 78.514 ;
               RECT 15.478 79.155 15.53 79.191 ;
               RECT 15.478 79.449 15.53 79.485 ;
               RECT 15.478 79.678 15.53 79.714 ;
               RECT 15.478 80.355 15.53 80.391 ;
               RECT 15.478 80.649 15.53 80.685 ;
               RECT 15.478 80.878 15.53 80.914 ;
               RECT 15.478 81.555 15.53 81.591 ;
               RECT 15.478 81.849 15.53 81.885 ;
               RECT 15.478 82.078 15.53 82.114 ;
               RECT 15.478 82.755 15.53 82.791 ;
               RECT 15.478 83.049 15.53 83.085 ;
               RECT 15.478 83.278 15.53 83.314 ;
               RECT 15.478 83.955 15.53 83.991 ;
               RECT 15.478 84.249 15.53 84.285 ;
               RECT 15.478 84.478 15.53 84.514 ;
               RECT 15.478 85.155 15.53 85.191 ;
               RECT 15.478 85.449 15.53 85.485 ;
               RECT 15.478 85.678 15.53 85.714 ;
               RECT 15.478 86.355 15.53 86.391 ;
               RECT 15.478 86.649 15.53 86.685 ;
               RECT 15.478 86.878 15.53 86.914 ;
               RECT 15.478 87.555 15.53 87.591 ;
               RECT 15.478 87.849 15.53 87.885 ;
               RECT 15.478 88.078 15.53 88.114 ;
               RECT 15.478 88.755 15.53 88.791 ;
               RECT 15.478 89.049 15.53 89.085 ;
               RECT 15.478 89.278 15.53 89.314 ;
               RECT 15.478 89.955 15.53 89.991 ;
               RECT 15.478 90.249 15.53 90.285 ;
               RECT 15.478 90.478 15.53 90.514 ;
               RECT 15.478 91.155 15.53 91.191 ;
               RECT 15.478 91.449 15.53 91.485 ;
               RECT 15.478 91.678 15.53 91.714 ;
               RECT 15.478 92.355 15.53 92.391 ;
               RECT 15.478 92.649 15.53 92.685 ;
               RECT 15.478 92.878 15.53 92.914 ;
               RECT 15.478 93.555 15.53 93.591 ;
               RECT 15.478 93.849 15.53 93.885 ;
               RECT 15.478 94.078 15.53 94.114 ;
               RECT 15.478 94.755 15.53 94.791 ;
               RECT 15.478 95.049 15.53 95.085 ;
               RECT 15.478 95.278 15.53 95.314 ;
               RECT 15.478 95.955 15.53 95.991 ;
               RECT 15.478 96.249 15.53 96.285 ;
               RECT 15.478 96.478 15.53 96.514 ;
               RECT 15.478 97.155 15.53 97.191 ;
               RECT 15.478 97.449 15.53 97.485 ;
               RECT 15.478 97.678 15.53 97.714 ;
               RECT 15.478 98.355 15.53 98.391 ;
               RECT 15.478 98.649 15.53 98.685 ;
               RECT 15.478 98.878 15.53 98.914 ;
               RECT 15.478 99.555 15.53 99.591 ;
               RECT 15.478 99.849 15.53 99.885 ;
               RECT 15.478 100.078 15.53 100.114 ;
               RECT 15.478 100.755 15.53 100.791 ;
               RECT 15.478 101.049 15.53 101.085 ;
               RECT 15.478 101.278 15.53 101.314 ;
               RECT 15.478 101.955 15.53 101.991 ;
               RECT 15.478 102.249 15.53 102.285 ;
               RECT 15.478 102.478 15.53 102.514 ;
               RECT 15.478 103.155 15.53 103.191 ;
               RECT 15.478 103.449 15.53 103.485 ;
               RECT 15.478 103.678 15.53 103.714 ;
               RECT 15.478 104.355 15.53 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.874 0.6 15.926 104.52 ;
               LAYER v4 ;
               RECT 15.874 0.729 15.926 0.765 ;
               RECT 15.874 0.958 15.926 0.994 ;
               RECT 15.874 1.406 15.926 1.442 ;
               RECT 15.874 1.635 15.926 1.671 ;
               RECT 15.874 1.929 15.926 1.965 ;
               RECT 15.874 2.158 15.926 2.194 ;
               RECT 15.874 2.606 15.926 2.642 ;
               RECT 15.874 2.835 15.926 2.871 ;
               RECT 15.874 3.129 15.926 3.165 ;
               RECT 15.874 3.358 15.926 3.394 ;
               RECT 15.874 3.806 15.926 3.842 ;
               RECT 15.874 4.035 15.926 4.071 ;
               RECT 15.874 4.329 15.926 4.365 ;
               RECT 15.874 4.558 15.926 4.594 ;
               RECT 15.874 5.006 15.926 5.042 ;
               RECT 15.874 5.235 15.926 5.271 ;
               RECT 15.874 5.529 15.926 5.565 ;
               RECT 15.874 5.758 15.926 5.794 ;
               RECT 15.874 6.206 15.926 6.242 ;
               RECT 15.874 6.435 15.926 6.471 ;
               RECT 15.874 6.729 15.926 6.765 ;
               RECT 15.874 6.958 15.926 6.994 ;
               RECT 15.874 7.406 15.926 7.442 ;
               RECT 15.874 7.635 15.926 7.671 ;
               RECT 15.874 7.929 15.926 7.965 ;
               RECT 15.874 8.158 15.926 8.194 ;
               RECT 15.874 8.606 15.926 8.642 ;
               RECT 15.874 8.835 15.926 8.871 ;
               RECT 15.874 9.129 15.926 9.165 ;
               RECT 15.874 9.358 15.926 9.394 ;
               RECT 15.874 9.806 15.926 9.842 ;
               RECT 15.874 10.035 15.926 10.071 ;
               RECT 15.874 10.329 15.926 10.365 ;
               RECT 15.874 10.558 15.926 10.594 ;
               RECT 15.874 11.006 15.926 11.042 ;
               RECT 15.874 11.235 15.926 11.271 ;
               RECT 15.874 11.529 15.926 11.565 ;
               RECT 15.874 11.758 15.926 11.794 ;
               RECT 15.874 12.206 15.926 12.242 ;
               RECT 15.874 12.435 15.926 12.471 ;
               RECT 15.874 12.729 15.926 12.765 ;
               RECT 15.874 12.958 15.926 12.994 ;
               RECT 15.874 13.406 15.926 13.442 ;
               RECT 15.874 13.635 15.926 13.671 ;
               RECT 15.874 13.929 15.926 13.965 ;
               RECT 15.874 14.158 15.926 14.194 ;
               RECT 15.874 14.606 15.926 14.642 ;
               RECT 15.874 14.835 15.926 14.871 ;
               RECT 15.874 15.129 15.926 15.165 ;
               RECT 15.874 15.358 15.926 15.394 ;
               RECT 15.874 15.806 15.926 15.842 ;
               RECT 15.874 16.035 15.926 16.071 ;
               RECT 15.874 16.329 15.926 16.365 ;
               RECT 15.874 16.558 15.926 16.594 ;
               RECT 15.874 17.006 15.926 17.042 ;
               RECT 15.874 17.235 15.926 17.271 ;
               RECT 15.874 17.529 15.926 17.565 ;
               RECT 15.874 17.758 15.926 17.794 ;
               RECT 15.874 18.206 15.926 18.242 ;
               RECT 15.874 18.435 15.926 18.471 ;
               RECT 15.874 18.729 15.926 18.765 ;
               RECT 15.874 18.958 15.926 18.994 ;
               RECT 15.874 19.406 15.926 19.442 ;
               RECT 15.874 19.635 15.926 19.671 ;
               RECT 15.874 19.929 15.926 19.965 ;
               RECT 15.874 20.158 15.926 20.194 ;
               RECT 15.874 20.606 15.926 20.642 ;
               RECT 15.874 20.835 15.926 20.871 ;
               RECT 15.874 21.129 15.926 21.165 ;
               RECT 15.874 21.358 15.926 21.394 ;
               RECT 15.874 21.806 15.926 21.842 ;
               RECT 15.874 22.035 15.926 22.071 ;
               RECT 15.874 22.329 15.926 22.365 ;
               RECT 15.874 22.558 15.926 22.594 ;
               RECT 15.874 23.006 15.926 23.042 ;
               RECT 15.874 23.235 15.926 23.271 ;
               RECT 15.874 23.529 15.926 23.565 ;
               RECT 15.874 23.758 15.926 23.794 ;
               RECT 15.874 24.206 15.926 24.242 ;
               RECT 15.874 24.435 15.926 24.471 ;
               RECT 15.874 24.729 15.926 24.765 ;
               RECT 15.874 24.958 15.926 24.994 ;
               RECT 15.874 25.406 15.926 25.442 ;
               RECT 15.874 25.635 15.926 25.671 ;
               RECT 15.874 25.929 15.926 25.965 ;
               RECT 15.874 26.158 15.926 26.194 ;
               RECT 15.874 26.606 15.926 26.642 ;
               RECT 15.874 26.835 15.926 26.871 ;
               RECT 15.874 27.129 15.926 27.165 ;
               RECT 15.874 27.358 15.926 27.394 ;
               RECT 15.874 27.806 15.926 27.842 ;
               RECT 15.874 28.035 15.926 28.071 ;
               RECT 15.874 28.329 15.926 28.365 ;
               RECT 15.874 28.558 15.926 28.594 ;
               RECT 15.874 29.006 15.926 29.042 ;
               RECT 15.874 29.235 15.926 29.271 ;
               RECT 15.874 29.529 15.926 29.565 ;
               RECT 15.874 29.758 15.926 29.794 ;
               RECT 15.874 30.206 15.926 30.242 ;
               RECT 15.874 30.435 15.926 30.471 ;
               RECT 15.874 30.729 15.926 30.765 ;
               RECT 15.874 30.958 15.926 30.994 ;
               RECT 15.874 31.406 15.926 31.442 ;
               RECT 15.874 31.635 15.926 31.671 ;
               RECT 15.874 31.929 15.926 31.965 ;
               RECT 15.874 32.158 15.926 32.194 ;
               RECT 15.874 32.606 15.926 32.642 ;
               RECT 15.874 32.835 15.926 32.871 ;
               RECT 15.874 33.129 15.926 33.165 ;
               RECT 15.874 33.358 15.926 33.394 ;
               RECT 15.874 33.806 15.926 33.842 ;
               RECT 15.874 34.035 15.926 34.071 ;
               RECT 15.874 34.329 15.926 34.365 ;
               RECT 15.874 34.558 15.926 34.594 ;
               RECT 15.874 35.006 15.926 35.042 ;
               RECT 15.874 35.235 15.926 35.271 ;
               RECT 15.874 35.529 15.926 35.565 ;
               RECT 15.874 35.758 15.926 35.794 ;
               RECT 15.874 36.206 15.926 36.242 ;
               RECT 15.874 36.435 15.926 36.471 ;
               RECT 15.874 36.729 15.926 36.765 ;
               RECT 15.874 36.958 15.926 36.994 ;
               RECT 15.874 37.406 15.926 37.442 ;
               RECT 15.874 37.635 15.926 37.671 ;
               RECT 15.874 37.929 15.926 37.965 ;
               RECT 15.874 38.158 15.926 38.194 ;
               RECT 15.874 38.606 15.926 38.642 ;
               RECT 15.874 38.835 15.926 38.871 ;
               RECT 15.874 39.129 15.926 39.165 ;
               RECT 15.874 39.358 15.926 39.394 ;
               RECT 15.874 39.806 15.926 39.842 ;
               RECT 15.874 40.035 15.926 40.071 ;
               RECT 15.874 40.329 15.926 40.365 ;
               RECT 15.874 40.558 15.926 40.594 ;
               RECT 15.874 41.006 15.926 41.042 ;
               RECT 15.874 41.235 15.926 41.271 ;
               RECT 15.874 41.529 15.926 41.565 ;
               RECT 15.874 41.758 15.926 41.794 ;
               RECT 15.874 42.206 15.926 42.242 ;
               RECT 15.874 42.435 15.926 42.471 ;
               RECT 15.874 42.729 15.926 42.765 ;
               RECT 15.874 42.958 15.926 42.994 ;
               RECT 15.874 43.406 15.926 43.442 ;
               RECT 15.874 43.635 15.926 43.671 ;
               RECT 15.874 43.929 15.926 43.965 ;
               RECT 15.874 44.158 15.926 44.194 ;
               RECT 15.874 44.606 15.926 44.642 ;
               RECT 15.874 44.835 15.926 44.871 ;
               RECT 15.874 45.129 15.926 45.165 ;
               RECT 15.874 45.358 15.926 45.394 ;
               RECT 15.874 45.806 15.926 45.842 ;
               RECT 15.874 46.035 15.926 46.071 ;
               RECT 15.874 46.329 15.926 46.365 ;
               RECT 15.874 46.558 15.926 46.594 ;
               RECT 15.874 47.006 15.926 47.042 ;
               RECT 15.874 47.235 15.926 47.271 ;
               RECT 15.874 47.529 15.926 47.565 ;
               RECT 15.874 47.758 15.926 47.794 ;
               RECT 15.874 48.206 15.926 48.242 ;
               RECT 15.874 48.435 15.926 48.471 ;
               RECT 15.874 49.182 15.926 49.218 ;
               RECT 15.874 49.662 15.926 49.698 ;
               RECT 15.874 50.142 15.926 50.178 ;
               RECT 15.874 50.622 15.926 50.658 ;
               RECT 15.874 51.102 15.926 51.138 ;
               RECT 15.874 51.582 15.926 51.618 ;
               RECT 15.874 52.062 15.926 52.098 ;
               RECT 15.874 52.542 15.926 52.578 ;
               RECT 15.874 53.0275 15.926 53.0525 ;
               RECT 15.874 53.502 15.926 53.538 ;
               RECT 15.874 53.982 15.926 54.018 ;
               RECT 15.874 54.462 15.926 54.498 ;
               RECT 15.874 54.9475 15.926 54.9725 ;
               RECT 15.874 55.422 15.926 55.458 ;
               RECT 15.874 55.902 15.926 55.938 ;
               RECT 15.874 56.649 15.926 56.685 ;
               RECT 15.874 56.878 15.926 56.914 ;
               RECT 15.874 57.326 15.926 57.362 ;
               RECT 15.874 57.555 15.926 57.591 ;
               RECT 15.874 57.849 15.926 57.885 ;
               RECT 15.874 58.078 15.926 58.114 ;
               RECT 15.874 58.526 15.926 58.562 ;
               RECT 15.874 58.755 15.926 58.791 ;
               RECT 15.874 59.049 15.926 59.085 ;
               RECT 15.874 59.278 15.926 59.314 ;
               RECT 15.874 59.726 15.926 59.762 ;
               RECT 15.874 59.955 15.926 59.991 ;
               RECT 15.874 60.249 15.926 60.285 ;
               RECT 15.874 60.478 15.926 60.514 ;
               RECT 15.874 60.926 15.926 60.962 ;
               RECT 15.874 61.155 15.926 61.191 ;
               RECT 15.874 61.449 15.926 61.485 ;
               RECT 15.874 61.678 15.926 61.714 ;
               RECT 15.874 62.126 15.926 62.162 ;
               RECT 15.874 62.355 15.926 62.391 ;
               RECT 15.874 62.649 15.926 62.685 ;
               RECT 15.874 62.878 15.926 62.914 ;
               RECT 15.874 63.326 15.926 63.362 ;
               RECT 15.874 63.555 15.926 63.591 ;
               RECT 15.874 63.849 15.926 63.885 ;
               RECT 15.874 64.078 15.926 64.114 ;
               RECT 15.874 64.526 15.926 64.562 ;
               RECT 15.874 64.755 15.926 64.791 ;
               RECT 15.874 65.049 15.926 65.085 ;
               RECT 15.874 65.278 15.926 65.314 ;
               RECT 15.874 65.726 15.926 65.762 ;
               RECT 15.874 65.955 15.926 65.991 ;
               RECT 15.874 66.249 15.926 66.285 ;
               RECT 15.874 66.478 15.926 66.514 ;
               RECT 15.874 66.926 15.926 66.962 ;
               RECT 15.874 67.155 15.926 67.191 ;
               RECT 15.874 67.449 15.926 67.485 ;
               RECT 15.874 67.678 15.926 67.714 ;
               RECT 15.874 68.126 15.926 68.162 ;
               RECT 15.874 68.355 15.926 68.391 ;
               RECT 15.874 68.649 15.926 68.685 ;
               RECT 15.874 68.878 15.926 68.914 ;
               RECT 15.874 69.326 15.926 69.362 ;
               RECT 15.874 69.555 15.926 69.591 ;
               RECT 15.874 69.849 15.926 69.885 ;
               RECT 15.874 70.078 15.926 70.114 ;
               RECT 15.874 70.526 15.926 70.562 ;
               RECT 15.874 70.755 15.926 70.791 ;
               RECT 15.874 71.049 15.926 71.085 ;
               RECT 15.874 71.278 15.926 71.314 ;
               RECT 15.874 71.726 15.926 71.762 ;
               RECT 15.874 71.955 15.926 71.991 ;
               RECT 15.874 72.249 15.926 72.285 ;
               RECT 15.874 72.478 15.926 72.514 ;
               RECT 15.874 72.926 15.926 72.962 ;
               RECT 15.874 73.155 15.926 73.191 ;
               RECT 15.874 73.449 15.926 73.485 ;
               RECT 15.874 73.678 15.926 73.714 ;
               RECT 15.874 74.126 15.926 74.162 ;
               RECT 15.874 74.355 15.926 74.391 ;
               RECT 15.874 74.649 15.926 74.685 ;
               RECT 15.874 74.878 15.926 74.914 ;
               RECT 15.874 75.326 15.926 75.362 ;
               RECT 15.874 75.555 15.926 75.591 ;
               RECT 15.874 75.849 15.926 75.885 ;
               RECT 15.874 76.078 15.926 76.114 ;
               RECT 15.874 76.526 15.926 76.562 ;
               RECT 15.874 76.755 15.926 76.791 ;
               RECT 15.874 77.049 15.926 77.085 ;
               RECT 15.874 77.278 15.926 77.314 ;
               RECT 15.874 77.726 15.926 77.762 ;
               RECT 15.874 77.955 15.926 77.991 ;
               RECT 15.874 78.249 15.926 78.285 ;
               RECT 15.874 78.478 15.926 78.514 ;
               RECT 15.874 78.926 15.926 78.962 ;
               RECT 15.874 79.155 15.926 79.191 ;
               RECT 15.874 79.449 15.926 79.485 ;
               RECT 15.874 79.678 15.926 79.714 ;
               RECT 15.874 80.126 15.926 80.162 ;
               RECT 15.874 80.355 15.926 80.391 ;
               RECT 15.874 80.649 15.926 80.685 ;
               RECT 15.874 80.878 15.926 80.914 ;
               RECT 15.874 81.326 15.926 81.362 ;
               RECT 15.874 81.555 15.926 81.591 ;
               RECT 15.874 81.849 15.926 81.885 ;
               RECT 15.874 82.078 15.926 82.114 ;
               RECT 15.874 82.526 15.926 82.562 ;
               RECT 15.874 82.755 15.926 82.791 ;
               RECT 15.874 83.049 15.926 83.085 ;
               RECT 15.874 83.278 15.926 83.314 ;
               RECT 15.874 83.726 15.926 83.762 ;
               RECT 15.874 83.955 15.926 83.991 ;
               RECT 15.874 84.249 15.926 84.285 ;
               RECT 15.874 84.478 15.926 84.514 ;
               RECT 15.874 84.926 15.926 84.962 ;
               RECT 15.874 85.155 15.926 85.191 ;
               RECT 15.874 85.449 15.926 85.485 ;
               RECT 15.874 85.678 15.926 85.714 ;
               RECT 15.874 86.126 15.926 86.162 ;
               RECT 15.874 86.355 15.926 86.391 ;
               RECT 15.874 86.649 15.926 86.685 ;
               RECT 15.874 86.878 15.926 86.914 ;
               RECT 15.874 87.326 15.926 87.362 ;
               RECT 15.874 87.555 15.926 87.591 ;
               RECT 15.874 87.849 15.926 87.885 ;
               RECT 15.874 88.078 15.926 88.114 ;
               RECT 15.874 88.526 15.926 88.562 ;
               RECT 15.874 88.755 15.926 88.791 ;
               RECT 15.874 89.049 15.926 89.085 ;
               RECT 15.874 89.278 15.926 89.314 ;
               RECT 15.874 89.726 15.926 89.762 ;
               RECT 15.874 89.955 15.926 89.991 ;
               RECT 15.874 90.249 15.926 90.285 ;
               RECT 15.874 90.478 15.926 90.514 ;
               RECT 15.874 90.926 15.926 90.962 ;
               RECT 15.874 91.155 15.926 91.191 ;
               RECT 15.874 91.449 15.926 91.485 ;
               RECT 15.874 91.678 15.926 91.714 ;
               RECT 15.874 92.126 15.926 92.162 ;
               RECT 15.874 92.355 15.926 92.391 ;
               RECT 15.874 92.649 15.926 92.685 ;
               RECT 15.874 92.878 15.926 92.914 ;
               RECT 15.874 93.326 15.926 93.362 ;
               RECT 15.874 93.555 15.926 93.591 ;
               RECT 15.874 93.849 15.926 93.885 ;
               RECT 15.874 94.078 15.926 94.114 ;
               RECT 15.874 94.526 15.926 94.562 ;
               RECT 15.874 94.755 15.926 94.791 ;
               RECT 15.874 95.049 15.926 95.085 ;
               RECT 15.874 95.278 15.926 95.314 ;
               RECT 15.874 95.726 15.926 95.762 ;
               RECT 15.874 95.955 15.926 95.991 ;
               RECT 15.874 96.249 15.926 96.285 ;
               RECT 15.874 96.478 15.926 96.514 ;
               RECT 15.874 96.926 15.926 96.962 ;
               RECT 15.874 97.155 15.926 97.191 ;
               RECT 15.874 97.449 15.926 97.485 ;
               RECT 15.874 97.678 15.926 97.714 ;
               RECT 15.874 98.126 15.926 98.162 ;
               RECT 15.874 98.355 15.926 98.391 ;
               RECT 15.874 98.649 15.926 98.685 ;
               RECT 15.874 98.878 15.926 98.914 ;
               RECT 15.874 99.326 15.926 99.362 ;
               RECT 15.874 99.555 15.926 99.591 ;
               RECT 15.874 99.849 15.926 99.885 ;
               RECT 15.874 100.078 15.926 100.114 ;
               RECT 15.874 100.526 15.926 100.562 ;
               RECT 15.874 100.755 15.926 100.791 ;
               RECT 15.874 101.049 15.926 101.085 ;
               RECT 15.874 101.278 15.926 101.314 ;
               RECT 15.874 101.726 15.926 101.762 ;
               RECT 15.874 101.955 15.926 101.991 ;
               RECT 15.874 102.249 15.926 102.285 ;
               RECT 15.874 102.478 15.926 102.514 ;
               RECT 15.874 102.926 15.926 102.962 ;
               RECT 15.874 103.155 15.926 103.191 ;
               RECT 15.874 103.449 15.926 103.485 ;
               RECT 15.874 103.678 15.926 103.714 ;
               RECT 15.874 104.126 15.926 104.162 ;
               RECT 15.874 104.355 15.926 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.034 0.5695 16.086 104.5505 ;
               LAYER v4 ;
               RECT 16.034 0.729 16.086 0.765 ;
               RECT 16.034 0.958 16.086 0.994 ;
               RECT 16.034 1.406 16.086 1.442 ;
               RECT 16.034 1.929 16.086 1.965 ;
               RECT 16.034 2.158 16.086 2.194 ;
               RECT 16.034 2.606 16.086 2.642 ;
               RECT 16.034 3.129 16.086 3.165 ;
               RECT 16.034 3.358 16.086 3.394 ;
               RECT 16.034 3.806 16.086 3.842 ;
               RECT 16.034 4.329 16.086 4.365 ;
               RECT 16.034 4.558 16.086 4.594 ;
               RECT 16.034 5.006 16.086 5.042 ;
               RECT 16.034 5.529 16.086 5.565 ;
               RECT 16.034 5.758 16.086 5.794 ;
               RECT 16.034 6.206 16.086 6.242 ;
               RECT 16.034 6.729 16.086 6.765 ;
               RECT 16.034 6.958 16.086 6.994 ;
               RECT 16.034 7.406 16.086 7.442 ;
               RECT 16.034 7.929 16.086 7.965 ;
               RECT 16.034 8.158 16.086 8.194 ;
               RECT 16.034 8.606 16.086 8.642 ;
               RECT 16.034 9.129 16.086 9.165 ;
               RECT 16.034 9.358 16.086 9.394 ;
               RECT 16.034 9.806 16.086 9.842 ;
               RECT 16.034 10.329 16.086 10.365 ;
               RECT 16.034 10.558 16.086 10.594 ;
               RECT 16.034 11.006 16.086 11.042 ;
               RECT 16.034 11.529 16.086 11.565 ;
               RECT 16.034 11.758 16.086 11.794 ;
               RECT 16.034 12.206 16.086 12.242 ;
               RECT 16.034 12.729 16.086 12.765 ;
               RECT 16.034 12.958 16.086 12.994 ;
               RECT 16.034 13.406 16.086 13.442 ;
               RECT 16.034 13.929 16.086 13.965 ;
               RECT 16.034 14.158 16.086 14.194 ;
               RECT 16.034 14.606 16.086 14.642 ;
               RECT 16.034 15.129 16.086 15.165 ;
               RECT 16.034 15.358 16.086 15.394 ;
               RECT 16.034 15.806 16.086 15.842 ;
               RECT 16.034 16.329 16.086 16.365 ;
               RECT 16.034 16.558 16.086 16.594 ;
               RECT 16.034 17.006 16.086 17.042 ;
               RECT 16.034 17.529 16.086 17.565 ;
               RECT 16.034 17.758 16.086 17.794 ;
               RECT 16.034 18.206 16.086 18.242 ;
               RECT 16.034 18.729 16.086 18.765 ;
               RECT 16.034 18.958 16.086 18.994 ;
               RECT 16.034 19.406 16.086 19.442 ;
               RECT 16.034 19.929 16.086 19.965 ;
               RECT 16.034 20.158 16.086 20.194 ;
               RECT 16.034 20.606 16.086 20.642 ;
               RECT 16.034 21.129 16.086 21.165 ;
               RECT 16.034 21.358 16.086 21.394 ;
               RECT 16.034 21.806 16.086 21.842 ;
               RECT 16.034 22.329 16.086 22.365 ;
               RECT 16.034 22.558 16.086 22.594 ;
               RECT 16.034 23.006 16.086 23.042 ;
               RECT 16.034 23.529 16.086 23.565 ;
               RECT 16.034 23.758 16.086 23.794 ;
               RECT 16.034 24.206 16.086 24.242 ;
               RECT 16.034 24.729 16.086 24.765 ;
               RECT 16.034 24.958 16.086 24.994 ;
               RECT 16.034 25.406 16.086 25.442 ;
               RECT 16.034 25.929 16.086 25.965 ;
               RECT 16.034 26.158 16.086 26.194 ;
               RECT 16.034 26.606 16.086 26.642 ;
               RECT 16.034 27.129 16.086 27.165 ;
               RECT 16.034 27.358 16.086 27.394 ;
               RECT 16.034 27.806 16.086 27.842 ;
               RECT 16.034 28.329 16.086 28.365 ;
               RECT 16.034 28.558 16.086 28.594 ;
               RECT 16.034 29.006 16.086 29.042 ;
               RECT 16.034 29.529 16.086 29.565 ;
               RECT 16.034 29.758 16.086 29.794 ;
               RECT 16.034 30.206 16.086 30.242 ;
               RECT 16.034 30.729 16.086 30.765 ;
               RECT 16.034 30.958 16.086 30.994 ;
               RECT 16.034 31.406 16.086 31.442 ;
               RECT 16.034 31.929 16.086 31.965 ;
               RECT 16.034 32.158 16.086 32.194 ;
               RECT 16.034 32.606 16.086 32.642 ;
               RECT 16.034 33.129 16.086 33.165 ;
               RECT 16.034 33.358 16.086 33.394 ;
               RECT 16.034 33.806 16.086 33.842 ;
               RECT 16.034 34.329 16.086 34.365 ;
               RECT 16.034 34.558 16.086 34.594 ;
               RECT 16.034 35.006 16.086 35.042 ;
               RECT 16.034 35.529 16.086 35.565 ;
               RECT 16.034 35.758 16.086 35.794 ;
               RECT 16.034 36.206 16.086 36.242 ;
               RECT 16.034 36.729 16.086 36.765 ;
               RECT 16.034 36.958 16.086 36.994 ;
               RECT 16.034 37.406 16.086 37.442 ;
               RECT 16.034 37.929 16.086 37.965 ;
               RECT 16.034 38.158 16.086 38.194 ;
               RECT 16.034 38.606 16.086 38.642 ;
               RECT 16.034 39.129 16.086 39.165 ;
               RECT 16.034 39.358 16.086 39.394 ;
               RECT 16.034 39.806 16.086 39.842 ;
               RECT 16.034 40.329 16.086 40.365 ;
               RECT 16.034 40.558 16.086 40.594 ;
               RECT 16.034 41.006 16.086 41.042 ;
               RECT 16.034 41.529 16.086 41.565 ;
               RECT 16.034 41.758 16.086 41.794 ;
               RECT 16.034 42.206 16.086 42.242 ;
               RECT 16.034 42.729 16.086 42.765 ;
               RECT 16.034 42.958 16.086 42.994 ;
               RECT 16.034 43.406 16.086 43.442 ;
               RECT 16.034 43.929 16.086 43.965 ;
               RECT 16.034 44.158 16.086 44.194 ;
               RECT 16.034 44.606 16.086 44.642 ;
               RECT 16.034 45.129 16.086 45.165 ;
               RECT 16.034 45.358 16.086 45.394 ;
               RECT 16.034 45.806 16.086 45.842 ;
               RECT 16.034 46.329 16.086 46.365 ;
               RECT 16.034 46.558 16.086 46.594 ;
               RECT 16.034 47.006 16.086 47.042 ;
               RECT 16.034 47.529 16.086 47.565 ;
               RECT 16.034 47.758 16.086 47.794 ;
               RECT 16.034 48.206 16.086 48.242 ;
               RECT 16.034 49.182 16.086 49.218 ;
               RECT 16.034 49.662 16.086 49.698 ;
               RECT 16.034 50.142 16.086 50.178 ;
               RECT 16.034 50.622 16.086 50.658 ;
               RECT 16.034 51.1075 16.086 51.1325 ;
               RECT 16.034 51.582 16.086 51.618 ;
               RECT 16.034 52.062 16.086 52.098 ;
               RECT 16.034 52.542 16.086 52.578 ;
               RECT 16.034 53.022 16.086 53.058 ;
               RECT 16.034 53.502 16.086 53.538 ;
               RECT 16.034 53.982 16.086 54.018 ;
               RECT 16.034 54.462 16.086 54.498 ;
               RECT 16.034 54.942 16.086 54.978 ;
               RECT 16.034 55.422 16.086 55.458 ;
               RECT 16.034 55.902 16.086 55.938 ;
               RECT 16.034 56.649 16.086 56.685 ;
               RECT 16.034 56.878 16.086 56.914 ;
               RECT 16.034 57.326 16.086 57.362 ;
               RECT 16.034 57.849 16.086 57.885 ;
               RECT 16.034 58.078 16.086 58.114 ;
               RECT 16.034 58.526 16.086 58.562 ;
               RECT 16.034 59.049 16.086 59.085 ;
               RECT 16.034 59.278 16.086 59.314 ;
               RECT 16.034 59.726 16.086 59.762 ;
               RECT 16.034 60.249 16.086 60.285 ;
               RECT 16.034 60.478 16.086 60.514 ;
               RECT 16.034 60.926 16.086 60.962 ;
               RECT 16.034 61.449 16.086 61.485 ;
               RECT 16.034 61.678 16.086 61.714 ;
               RECT 16.034 62.126 16.086 62.162 ;
               RECT 16.034 62.649 16.086 62.685 ;
               RECT 16.034 62.878 16.086 62.914 ;
               RECT 16.034 63.326 16.086 63.362 ;
               RECT 16.034 63.849 16.086 63.885 ;
               RECT 16.034 64.078 16.086 64.114 ;
               RECT 16.034 64.526 16.086 64.562 ;
               RECT 16.034 65.049 16.086 65.085 ;
               RECT 16.034 65.278 16.086 65.314 ;
               RECT 16.034 65.726 16.086 65.762 ;
               RECT 16.034 66.249 16.086 66.285 ;
               RECT 16.034 66.478 16.086 66.514 ;
               RECT 16.034 66.926 16.086 66.962 ;
               RECT 16.034 67.449 16.086 67.485 ;
               RECT 16.034 67.678 16.086 67.714 ;
               RECT 16.034 68.126 16.086 68.162 ;
               RECT 16.034 68.649 16.086 68.685 ;
               RECT 16.034 68.878 16.086 68.914 ;
               RECT 16.034 69.326 16.086 69.362 ;
               RECT 16.034 69.849 16.086 69.885 ;
               RECT 16.034 70.078 16.086 70.114 ;
               RECT 16.034 70.526 16.086 70.562 ;
               RECT 16.034 71.049 16.086 71.085 ;
               RECT 16.034 71.278 16.086 71.314 ;
               RECT 16.034 71.726 16.086 71.762 ;
               RECT 16.034 72.249 16.086 72.285 ;
               RECT 16.034 72.478 16.086 72.514 ;
               RECT 16.034 72.926 16.086 72.962 ;
               RECT 16.034 73.449 16.086 73.485 ;
               RECT 16.034 73.678 16.086 73.714 ;
               RECT 16.034 74.126 16.086 74.162 ;
               RECT 16.034 74.649 16.086 74.685 ;
               RECT 16.034 74.878 16.086 74.914 ;
               RECT 16.034 75.326 16.086 75.362 ;
               RECT 16.034 75.849 16.086 75.885 ;
               RECT 16.034 76.078 16.086 76.114 ;
               RECT 16.034 76.526 16.086 76.562 ;
               RECT 16.034 77.049 16.086 77.085 ;
               RECT 16.034 77.278 16.086 77.314 ;
               RECT 16.034 77.726 16.086 77.762 ;
               RECT 16.034 78.249 16.086 78.285 ;
               RECT 16.034 78.478 16.086 78.514 ;
               RECT 16.034 78.926 16.086 78.962 ;
               RECT 16.034 79.449 16.086 79.485 ;
               RECT 16.034 79.678 16.086 79.714 ;
               RECT 16.034 80.126 16.086 80.162 ;
               RECT 16.034 80.649 16.086 80.685 ;
               RECT 16.034 80.878 16.086 80.914 ;
               RECT 16.034 81.326 16.086 81.362 ;
               RECT 16.034 81.849 16.086 81.885 ;
               RECT 16.034 82.078 16.086 82.114 ;
               RECT 16.034 82.526 16.086 82.562 ;
               RECT 16.034 83.049 16.086 83.085 ;
               RECT 16.034 83.278 16.086 83.314 ;
               RECT 16.034 83.726 16.086 83.762 ;
               RECT 16.034 84.249 16.086 84.285 ;
               RECT 16.034 84.478 16.086 84.514 ;
               RECT 16.034 84.926 16.086 84.962 ;
               RECT 16.034 85.449 16.086 85.485 ;
               RECT 16.034 85.678 16.086 85.714 ;
               RECT 16.034 86.126 16.086 86.162 ;
               RECT 16.034 86.649 16.086 86.685 ;
               RECT 16.034 86.878 16.086 86.914 ;
               RECT 16.034 87.326 16.086 87.362 ;
               RECT 16.034 87.849 16.086 87.885 ;
               RECT 16.034 88.078 16.086 88.114 ;
               RECT 16.034 88.526 16.086 88.562 ;
               RECT 16.034 89.049 16.086 89.085 ;
               RECT 16.034 89.278 16.086 89.314 ;
               RECT 16.034 89.726 16.086 89.762 ;
               RECT 16.034 90.249 16.086 90.285 ;
               RECT 16.034 90.478 16.086 90.514 ;
               RECT 16.034 90.926 16.086 90.962 ;
               RECT 16.034 91.449 16.086 91.485 ;
               RECT 16.034 91.678 16.086 91.714 ;
               RECT 16.034 92.126 16.086 92.162 ;
               RECT 16.034 92.649 16.086 92.685 ;
               RECT 16.034 92.878 16.086 92.914 ;
               RECT 16.034 93.326 16.086 93.362 ;
               RECT 16.034 93.849 16.086 93.885 ;
               RECT 16.034 94.078 16.086 94.114 ;
               RECT 16.034 94.526 16.086 94.562 ;
               RECT 16.034 95.049 16.086 95.085 ;
               RECT 16.034 95.278 16.086 95.314 ;
               RECT 16.034 95.726 16.086 95.762 ;
               RECT 16.034 96.249 16.086 96.285 ;
               RECT 16.034 96.478 16.086 96.514 ;
               RECT 16.034 96.926 16.086 96.962 ;
               RECT 16.034 97.449 16.086 97.485 ;
               RECT 16.034 97.678 16.086 97.714 ;
               RECT 16.034 98.126 16.086 98.162 ;
               RECT 16.034 98.649 16.086 98.685 ;
               RECT 16.034 98.878 16.086 98.914 ;
               RECT 16.034 99.326 16.086 99.362 ;
               RECT 16.034 99.849 16.086 99.885 ;
               RECT 16.034 100.078 16.086 100.114 ;
               RECT 16.034 100.526 16.086 100.562 ;
               RECT 16.034 101.049 16.086 101.085 ;
               RECT 16.034 101.278 16.086 101.314 ;
               RECT 16.034 101.726 16.086 101.762 ;
               RECT 16.034 102.249 16.086 102.285 ;
               RECT 16.034 102.478 16.086 102.514 ;
               RECT 16.034 102.926 16.086 102.962 ;
               RECT 16.034 103.449 16.086 103.485 ;
               RECT 16.034 103.678 16.086 103.714 ;
               RECT 16.034 104.126 16.086 104.162 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.8 0.5695 16.854 104.5505 ;
               LAYER v4 ;
               RECT 16.8 0.729 16.854 0.765 ;
               RECT 16.8 0.958 16.854 0.994 ;
               RECT 16.8 1.929 16.854 1.965 ;
               RECT 16.8 2.158 16.854 2.194 ;
               RECT 16.8 3.129 16.854 3.165 ;
               RECT 16.8 3.358 16.854 3.394 ;
               RECT 16.8 4.329 16.854 4.365 ;
               RECT 16.8 4.558 16.854 4.594 ;
               RECT 16.8 5.529 16.854 5.565 ;
               RECT 16.8 5.758 16.854 5.794 ;
               RECT 16.8 6.729 16.854 6.765 ;
               RECT 16.8 6.958 16.854 6.994 ;
               RECT 16.8 7.929 16.854 7.965 ;
               RECT 16.8 8.158 16.854 8.194 ;
               RECT 16.8 9.129 16.854 9.165 ;
               RECT 16.8 9.358 16.854 9.394 ;
               RECT 16.8 10.329 16.854 10.365 ;
               RECT 16.8 10.558 16.854 10.594 ;
               RECT 16.8 11.529 16.854 11.565 ;
               RECT 16.8 11.758 16.854 11.794 ;
               RECT 16.8 12.729 16.854 12.765 ;
               RECT 16.8 12.958 16.854 12.994 ;
               RECT 16.8 13.929 16.854 13.965 ;
               RECT 16.8 14.158 16.854 14.194 ;
               RECT 16.8 15.129 16.854 15.165 ;
               RECT 16.8 15.358 16.854 15.394 ;
               RECT 16.8 16.329 16.854 16.365 ;
               RECT 16.8 16.558 16.854 16.594 ;
               RECT 16.8 17.529 16.854 17.565 ;
               RECT 16.8 17.758 16.854 17.794 ;
               RECT 16.8 18.729 16.854 18.765 ;
               RECT 16.8 18.958 16.854 18.994 ;
               RECT 16.8 19.929 16.854 19.965 ;
               RECT 16.8 20.158 16.854 20.194 ;
               RECT 16.8 21.129 16.854 21.165 ;
               RECT 16.8 21.358 16.854 21.394 ;
               RECT 16.8 22.329 16.854 22.365 ;
               RECT 16.8 22.558 16.854 22.594 ;
               RECT 16.8 23.529 16.854 23.565 ;
               RECT 16.8 23.758 16.854 23.794 ;
               RECT 16.8 24.729 16.854 24.765 ;
               RECT 16.8 24.958 16.854 24.994 ;
               RECT 16.8 25.929 16.854 25.965 ;
               RECT 16.8 26.158 16.854 26.194 ;
               RECT 16.8 27.129 16.854 27.165 ;
               RECT 16.8 27.358 16.854 27.394 ;
               RECT 16.8 28.329 16.854 28.365 ;
               RECT 16.8 28.558 16.854 28.594 ;
               RECT 16.8 29.529 16.854 29.565 ;
               RECT 16.8 29.758 16.854 29.794 ;
               RECT 16.8 30.729 16.854 30.765 ;
               RECT 16.8 30.958 16.854 30.994 ;
               RECT 16.8 31.929 16.854 31.965 ;
               RECT 16.8 32.158 16.854 32.194 ;
               RECT 16.8 33.129 16.854 33.165 ;
               RECT 16.8 33.358 16.854 33.394 ;
               RECT 16.8 34.329 16.854 34.365 ;
               RECT 16.8 34.558 16.854 34.594 ;
               RECT 16.8 35.529 16.854 35.565 ;
               RECT 16.8 35.758 16.854 35.794 ;
               RECT 16.8 36.729 16.854 36.765 ;
               RECT 16.8 36.958 16.854 36.994 ;
               RECT 16.8 37.929 16.854 37.965 ;
               RECT 16.8 38.158 16.854 38.194 ;
               RECT 16.8 39.129 16.854 39.165 ;
               RECT 16.8 39.358 16.854 39.394 ;
               RECT 16.8 40.329 16.854 40.365 ;
               RECT 16.8 40.558 16.854 40.594 ;
               RECT 16.8 41.529 16.854 41.565 ;
               RECT 16.8 41.758 16.854 41.794 ;
               RECT 16.8 42.729 16.854 42.765 ;
               RECT 16.8 42.958 16.854 42.994 ;
               RECT 16.8 43.929 16.854 43.965 ;
               RECT 16.8 44.158 16.854 44.194 ;
               RECT 16.8 45.129 16.854 45.165 ;
               RECT 16.8 45.358 16.854 45.394 ;
               RECT 16.8 46.329 16.854 46.365 ;
               RECT 16.8 46.558 16.854 46.594 ;
               RECT 16.8 47.529 16.854 47.565 ;
               RECT 16.8 47.758 16.854 47.794 ;
               RECT 16.8 49.182 16.854 49.218 ;
               RECT 16.8 49.662 16.854 49.698 ;
               RECT 16.8 49.8435 16.854 49.8795 ;
               RECT 16.8 50.142 16.854 50.178 ;
               RECT 16.8 50.622 16.854 50.658 ;
               RECT 16.8 51.102 16.854 51.138 ;
               RECT 16.8 51.582 16.854 51.618 ;
               RECT 16.8 52.062 16.854 52.098 ;
               RECT 16.8 52.542 16.854 52.578 ;
               RECT 16.8 53.022 16.854 53.058 ;
               RECT 16.8 53.502 16.854 53.538 ;
               RECT 16.8 53.982 16.854 54.018 ;
               RECT 16.8 54.462 16.854 54.498 ;
               RECT 16.8 54.942 16.854 54.978 ;
               RECT 16.8 55.422 16.854 55.458 ;
               RECT 16.8 55.902 16.854 55.938 ;
               RECT 16.8 56.649 16.854 56.685 ;
               RECT 16.8 56.878 16.854 56.914 ;
               RECT 16.8 57.849 16.854 57.885 ;
               RECT 16.8 58.078 16.854 58.114 ;
               RECT 16.8 59.049 16.854 59.085 ;
               RECT 16.8 59.278 16.854 59.314 ;
               RECT 16.8 60.249 16.854 60.285 ;
               RECT 16.8 60.478 16.854 60.514 ;
               RECT 16.8 61.449 16.854 61.485 ;
               RECT 16.8 61.678 16.854 61.714 ;
               RECT 16.8 62.649 16.854 62.685 ;
               RECT 16.8 62.878 16.854 62.914 ;
               RECT 16.8 63.849 16.854 63.885 ;
               RECT 16.8 64.078 16.854 64.114 ;
               RECT 16.8 65.049 16.854 65.085 ;
               RECT 16.8 65.278 16.854 65.314 ;
               RECT 16.8 66.249 16.854 66.285 ;
               RECT 16.8 66.478 16.854 66.514 ;
               RECT 16.8 67.449 16.854 67.485 ;
               RECT 16.8 67.678 16.854 67.714 ;
               RECT 16.8 68.649 16.854 68.685 ;
               RECT 16.8 68.878 16.854 68.914 ;
               RECT 16.8 69.849 16.854 69.885 ;
               RECT 16.8 70.078 16.854 70.114 ;
               RECT 16.8 71.049 16.854 71.085 ;
               RECT 16.8 71.278 16.854 71.314 ;
               RECT 16.8 72.249 16.854 72.285 ;
               RECT 16.8 72.478 16.854 72.514 ;
               RECT 16.8 73.449 16.854 73.485 ;
               RECT 16.8 73.678 16.854 73.714 ;
               RECT 16.8 74.649 16.854 74.685 ;
               RECT 16.8 74.878 16.854 74.914 ;
               RECT 16.8 75.849 16.854 75.885 ;
               RECT 16.8 76.078 16.854 76.114 ;
               RECT 16.8 77.049 16.854 77.085 ;
               RECT 16.8 77.278 16.854 77.314 ;
               RECT 16.8 78.249 16.854 78.285 ;
               RECT 16.8 78.478 16.854 78.514 ;
               RECT 16.8 79.449 16.854 79.485 ;
               RECT 16.8 79.678 16.854 79.714 ;
               RECT 16.8 80.649 16.854 80.685 ;
               RECT 16.8 80.878 16.854 80.914 ;
               RECT 16.8 81.849 16.854 81.885 ;
               RECT 16.8 82.078 16.854 82.114 ;
               RECT 16.8 83.049 16.854 83.085 ;
               RECT 16.8 83.278 16.854 83.314 ;
               RECT 16.8 84.249 16.854 84.285 ;
               RECT 16.8 84.478 16.854 84.514 ;
               RECT 16.8 85.449 16.854 85.485 ;
               RECT 16.8 85.678 16.854 85.714 ;
               RECT 16.8 86.649 16.854 86.685 ;
               RECT 16.8 86.878 16.854 86.914 ;
               RECT 16.8 87.849 16.854 87.885 ;
               RECT 16.8 88.078 16.854 88.114 ;
               RECT 16.8 89.049 16.854 89.085 ;
               RECT 16.8 89.278 16.854 89.314 ;
               RECT 16.8 90.249 16.854 90.285 ;
               RECT 16.8 90.478 16.854 90.514 ;
               RECT 16.8 91.449 16.854 91.485 ;
               RECT 16.8 91.678 16.854 91.714 ;
               RECT 16.8 92.649 16.854 92.685 ;
               RECT 16.8 92.878 16.854 92.914 ;
               RECT 16.8 93.849 16.854 93.885 ;
               RECT 16.8 94.078 16.854 94.114 ;
               RECT 16.8 95.049 16.854 95.085 ;
               RECT 16.8 95.278 16.854 95.314 ;
               RECT 16.8 96.249 16.854 96.285 ;
               RECT 16.8 96.478 16.854 96.514 ;
               RECT 16.8 97.449 16.854 97.485 ;
               RECT 16.8 97.678 16.854 97.714 ;
               RECT 16.8 98.649 16.854 98.685 ;
               RECT 16.8 98.878 16.854 98.914 ;
               RECT 16.8 99.849 16.854 99.885 ;
               RECT 16.8 100.078 16.854 100.114 ;
               RECT 16.8 101.049 16.854 101.085 ;
               RECT 16.8 101.278 16.854 101.314 ;
               RECT 16.8 102.249 16.854 102.285 ;
               RECT 16.8 102.478 16.854 102.514 ;
               RECT 16.8 103.449 16.854 103.485 ;
               RECT 16.8 103.678 16.854 103.714 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.964 0.5695 17.036 104.5505 ;
               LAYER v4 ;
               RECT 16.964 0.7345 17.036 0.7595 ;
               RECT 16.964 1.4115 17.036 1.4365 ;
               RECT 16.964 1.9345 17.036 1.9595 ;
               RECT 16.964 2.6115 17.036 2.6365 ;
               RECT 16.964 3.1345 17.036 3.1595 ;
               RECT 16.964 3.8115 17.036 3.8365 ;
               RECT 16.964 4.3345 17.036 4.3595 ;
               RECT 16.964 5.0115 17.036 5.0365 ;
               RECT 16.964 5.5345 17.036 5.5595 ;
               RECT 16.964 6.2115 17.036 6.2365 ;
               RECT 16.964 6.7345 17.036 6.7595 ;
               RECT 16.964 7.4115 17.036 7.4365 ;
               RECT 16.964 7.9345 17.036 7.9595 ;
               RECT 16.964 8.6115 17.036 8.6365 ;
               RECT 16.964 9.1345 17.036 9.1595 ;
               RECT 16.964 9.8115 17.036 9.8365 ;
               RECT 16.964 10.3345 17.036 10.3595 ;
               RECT 16.964 11.0115 17.036 11.0365 ;
               RECT 16.964 11.5345 17.036 11.5595 ;
               RECT 16.964 12.2115 17.036 12.2365 ;
               RECT 16.964 12.7345 17.036 12.7595 ;
               RECT 16.964 13.4115 17.036 13.4365 ;
               RECT 16.964 13.9345 17.036 13.9595 ;
               RECT 16.964 14.6115 17.036 14.6365 ;
               RECT 16.964 15.1345 17.036 15.1595 ;
               RECT 16.964 15.8115 17.036 15.8365 ;
               RECT 16.964 16.3345 17.036 16.3595 ;
               RECT 16.964 17.0115 17.036 17.0365 ;
               RECT 16.964 17.5345 17.036 17.5595 ;
               RECT 16.964 18.2115 17.036 18.2365 ;
               RECT 16.964 18.7345 17.036 18.7595 ;
               RECT 16.964 19.4115 17.036 19.4365 ;
               RECT 16.964 19.9345 17.036 19.9595 ;
               RECT 16.964 20.6115 17.036 20.6365 ;
               RECT 16.964 21.1345 17.036 21.1595 ;
               RECT 16.964 21.8115 17.036 21.8365 ;
               RECT 16.964 22.3345 17.036 22.3595 ;
               RECT 16.964 23.0115 17.036 23.0365 ;
               RECT 16.964 23.5345 17.036 23.5595 ;
               RECT 16.964 24.2115 17.036 24.2365 ;
               RECT 16.964 24.7345 17.036 24.7595 ;
               RECT 16.964 25.4115 17.036 25.4365 ;
               RECT 16.964 25.9345 17.036 25.9595 ;
               RECT 16.964 26.6115 17.036 26.6365 ;
               RECT 16.964 27.1345 17.036 27.1595 ;
               RECT 16.964 27.8115 17.036 27.8365 ;
               RECT 16.964 28.3345 17.036 28.3595 ;
               RECT 16.964 29.0115 17.036 29.0365 ;
               RECT 16.964 29.5345 17.036 29.5595 ;
               RECT 16.964 30.2115 17.036 30.2365 ;
               RECT 16.964 30.7345 17.036 30.7595 ;
               RECT 16.964 31.4115 17.036 31.4365 ;
               RECT 16.964 31.9345 17.036 31.9595 ;
               RECT 16.964 32.6115 17.036 32.6365 ;
               RECT 16.964 33.1345 17.036 33.1595 ;
               RECT 16.964 33.8115 17.036 33.8365 ;
               RECT 16.964 34.3345 17.036 34.3595 ;
               RECT 16.964 35.0115 17.036 35.0365 ;
               RECT 16.964 35.5345 17.036 35.5595 ;
               RECT 16.964 36.2115 17.036 36.2365 ;
               RECT 16.964 36.7345 17.036 36.7595 ;
               RECT 16.964 37.4115 17.036 37.4365 ;
               RECT 16.964 37.9345 17.036 37.9595 ;
               RECT 16.964 38.6115 17.036 38.6365 ;
               RECT 16.964 39.1345 17.036 39.1595 ;
               RECT 16.964 39.8115 17.036 39.8365 ;
               RECT 16.964 40.3345 17.036 40.3595 ;
               RECT 16.964 41.0115 17.036 41.0365 ;
               RECT 16.964 41.5345 17.036 41.5595 ;
               RECT 16.964 42.2115 17.036 42.2365 ;
               RECT 16.964 42.7345 17.036 42.7595 ;
               RECT 16.964 43.4115 17.036 43.4365 ;
               RECT 16.964 43.9345 17.036 43.9595 ;
               RECT 16.964 44.6115 17.036 44.6365 ;
               RECT 16.964 45.1345 17.036 45.1595 ;
               RECT 16.964 45.8115 17.036 45.8365 ;
               RECT 16.964 46.3345 17.036 46.3595 ;
               RECT 16.964 47.0115 17.036 47.0365 ;
               RECT 16.964 47.5345 17.036 47.5595 ;
               RECT 16.964 48.2115 17.036 48.2365 ;
               RECT 16.964 49.1875 17.036 49.2125 ;
               RECT 16.964 49.6675 17.036 49.6925 ;
               RECT 16.964 49.849 17.036 49.874 ;
               RECT 16.964 50.1475 17.036 50.1725 ;
               RECT 16.964 50.6275 17.036 50.6525 ;
               RECT 16.964 51.1075 17.036 51.1325 ;
               RECT 16.964 51.5875 17.036 51.6125 ;
               RECT 16.964 52.0675 17.036 52.0925 ;
               RECT 16.964 52.5475 17.036 52.5725 ;
               RECT 16.964 53.0275 17.036 53.0525 ;
               RECT 16.964 53.5075 17.036 53.5325 ;
               RECT 16.964 53.9875 17.036 54.0125 ;
               RECT 16.964 54.4675 17.036 54.4925 ;
               RECT 16.964 54.9475 17.036 54.9725 ;
               RECT 16.964 55.4275 17.036 55.4525 ;
               RECT 16.964 55.9075 17.036 55.9325 ;
               RECT 16.964 56.6545 17.036 56.6795 ;
               RECT 16.964 57.3315 17.036 57.3565 ;
               RECT 16.964 57.8545 17.036 57.8795 ;
               RECT 16.964 58.5315 17.036 58.5565 ;
               RECT 16.964 59.0545 17.036 59.0795 ;
               RECT 16.964 59.7315 17.036 59.7565 ;
               RECT 16.964 60.2545 17.036 60.2795 ;
               RECT 16.964 60.9315 17.036 60.9565 ;
               RECT 16.964 61.4545 17.036 61.4795 ;
               RECT 16.964 62.1315 17.036 62.1565 ;
               RECT 16.964 62.6545 17.036 62.6795 ;
               RECT 16.964 63.3315 17.036 63.3565 ;
               RECT 16.964 63.8545 17.036 63.8795 ;
               RECT 16.964 64.5315 17.036 64.5565 ;
               RECT 16.964 65.0545 17.036 65.0795 ;
               RECT 16.964 65.7315 17.036 65.7565 ;
               RECT 16.964 66.2545 17.036 66.2795 ;
               RECT 16.964 66.9315 17.036 66.9565 ;
               RECT 16.964 67.4545 17.036 67.4795 ;
               RECT 16.964 68.1315 17.036 68.1565 ;
               RECT 16.964 68.6545 17.036 68.6795 ;
               RECT 16.964 69.3315 17.036 69.3565 ;
               RECT 16.964 69.8545 17.036 69.8795 ;
               RECT 16.964 70.5315 17.036 70.5565 ;
               RECT 16.964 71.0545 17.036 71.0795 ;
               RECT 16.964 71.7315 17.036 71.7565 ;
               RECT 16.964 72.2545 17.036 72.2795 ;
               RECT 16.964 72.9315 17.036 72.9565 ;
               RECT 16.964 73.4545 17.036 73.4795 ;
               RECT 16.964 74.1315 17.036 74.1565 ;
               RECT 16.964 74.6545 17.036 74.6795 ;
               RECT 16.964 75.3315 17.036 75.3565 ;
               RECT 16.964 75.8545 17.036 75.8795 ;
               RECT 16.964 76.5315 17.036 76.5565 ;
               RECT 16.964 77.0545 17.036 77.0795 ;
               RECT 16.964 77.7315 17.036 77.7565 ;
               RECT 16.964 78.2545 17.036 78.2795 ;
               RECT 16.964 78.9315 17.036 78.9565 ;
               RECT 16.964 79.4545 17.036 79.4795 ;
               RECT 16.964 80.1315 17.036 80.1565 ;
               RECT 16.964 80.6545 17.036 80.6795 ;
               RECT 16.964 81.3315 17.036 81.3565 ;
               RECT 16.964 81.8545 17.036 81.8795 ;
               RECT 16.964 82.5315 17.036 82.5565 ;
               RECT 16.964 83.0545 17.036 83.0795 ;
               RECT 16.964 83.7315 17.036 83.7565 ;
               RECT 16.964 84.2545 17.036 84.2795 ;
               RECT 16.964 84.9315 17.036 84.9565 ;
               RECT 16.964 85.4545 17.036 85.4795 ;
               RECT 16.964 86.1315 17.036 86.1565 ;
               RECT 16.964 86.6545 17.036 86.6795 ;
               RECT 16.964 87.3315 17.036 87.3565 ;
               RECT 16.964 87.8545 17.036 87.8795 ;
               RECT 16.964 88.5315 17.036 88.5565 ;
               RECT 16.964 89.0545 17.036 89.0795 ;
               RECT 16.964 89.7315 17.036 89.7565 ;
               RECT 16.964 90.2545 17.036 90.2795 ;
               RECT 16.964 90.9315 17.036 90.9565 ;
               RECT 16.964 91.4545 17.036 91.4795 ;
               RECT 16.964 92.1315 17.036 92.1565 ;
               RECT 16.964 92.6545 17.036 92.6795 ;
               RECT 16.964 93.3315 17.036 93.3565 ;
               RECT 16.964 93.8545 17.036 93.8795 ;
               RECT 16.964 94.5315 17.036 94.5565 ;
               RECT 16.964 95.0545 17.036 95.0795 ;
               RECT 16.964 95.7315 17.036 95.7565 ;
               RECT 16.964 96.2545 17.036 96.2795 ;
               RECT 16.964 96.9315 17.036 96.9565 ;
               RECT 16.964 97.4545 17.036 97.4795 ;
               RECT 16.964 98.1315 17.036 98.1565 ;
               RECT 16.964 98.6545 17.036 98.6795 ;
               RECT 16.964 99.3315 17.036 99.3565 ;
               RECT 16.964 99.8545 17.036 99.8795 ;
               RECT 16.964 100.5315 17.036 100.5565 ;
               RECT 16.964 101.0545 17.036 101.0795 ;
               RECT 16.964 101.7315 17.036 101.7565 ;
               RECT 16.964 102.2545 17.036 102.2795 ;
               RECT 16.964 102.9315 17.036 102.9565 ;
               RECT 16.964 103.4545 17.036 103.4795 ;
               RECT 16.964 104.1315 17.036 104.1565 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.412 48.98 17.452 56.14 ;
               LAYER v4 ;
               RECT 17.412 49.182 17.452 49.218 ;
               RECT 17.412 49.662 17.452 49.698 ;
               RECT 17.412 49.8435 17.452 49.8795 ;
               RECT 17.412 50.142 17.452 50.178 ;
               RECT 17.412 50.622 17.452 50.658 ;
               RECT 17.412 51.102 17.452 51.138 ;
               RECT 17.412 51.582 17.452 51.618 ;
               RECT 17.412 52.062 17.452 52.098 ;
               RECT 17.412 52.542 17.452 52.578 ;
               RECT 17.412 53.022 17.452 53.058 ;
               RECT 17.412 53.502 17.452 53.538 ;
               RECT 17.412 53.982 17.452 54.018 ;
               RECT 17.412 54.462 17.452 54.498 ;
               RECT 17.412 54.942 17.452 54.978 ;
               RECT 17.412 55.422 17.452 55.458 ;
               RECT 17.412 55.902 17.452 55.938 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.844 0.5695 17.916 104.5505 ;
               LAYER v4 ;
               RECT 17.844 1.0405 17.916 1.0655 ;
               RECT 17.844 1.5635 17.916 1.5885 ;
               RECT 17.844 2.2405 17.916 2.2655 ;
               RECT 17.844 2.7635 17.916 2.7885 ;
               RECT 17.844 3.4405 17.916 3.4655 ;
               RECT 17.844 3.9635 17.916 3.9885 ;
               RECT 17.844 4.6405 17.916 4.6655 ;
               RECT 17.844 5.1635 17.916 5.1885 ;
               RECT 17.844 5.8405 17.916 5.8655 ;
               RECT 17.844 6.3635 17.916 6.3885 ;
               RECT 17.844 7.0405 17.916 7.0655 ;
               RECT 17.844 7.5635 17.916 7.5885 ;
               RECT 17.844 8.2405 17.916 8.2655 ;
               RECT 17.844 8.7635 17.916 8.7885 ;
               RECT 17.844 9.4405 17.916 9.4655 ;
               RECT 17.844 9.9635 17.916 9.9885 ;
               RECT 17.844 10.6405 17.916 10.6655 ;
               RECT 17.844 11.1635 17.916 11.1885 ;
               RECT 17.844 11.8405 17.916 11.8655 ;
               RECT 17.844 12.3635 17.916 12.3885 ;
               RECT 17.844 13.0405 17.916 13.0655 ;
               RECT 17.844 13.5635 17.916 13.5885 ;
               RECT 17.844 14.2405 17.916 14.2655 ;
               RECT 17.844 14.7635 17.916 14.7885 ;
               RECT 17.844 15.4405 17.916 15.4655 ;
               RECT 17.844 15.9635 17.916 15.9885 ;
               RECT 17.844 16.6405 17.916 16.6655 ;
               RECT 17.844 17.1635 17.916 17.1885 ;
               RECT 17.844 17.8405 17.916 17.8655 ;
               RECT 17.844 18.3635 17.916 18.3885 ;
               RECT 17.844 19.0405 17.916 19.0655 ;
               RECT 17.844 19.5635 17.916 19.5885 ;
               RECT 17.844 20.2405 17.916 20.2655 ;
               RECT 17.844 20.7635 17.916 20.7885 ;
               RECT 17.844 21.4405 17.916 21.4655 ;
               RECT 17.844 21.9635 17.916 21.9885 ;
               RECT 17.844 22.6405 17.916 22.6655 ;
               RECT 17.844 23.1635 17.916 23.1885 ;
               RECT 17.844 23.8405 17.916 23.8655 ;
               RECT 17.844 24.3635 17.916 24.3885 ;
               RECT 17.844 25.0405 17.916 25.0655 ;
               RECT 17.844 25.5635 17.916 25.5885 ;
               RECT 17.844 26.2405 17.916 26.2655 ;
               RECT 17.844 26.7635 17.916 26.7885 ;
               RECT 17.844 27.4405 17.916 27.4655 ;
               RECT 17.844 27.9635 17.916 27.9885 ;
               RECT 17.844 28.6405 17.916 28.6655 ;
               RECT 17.844 29.1635 17.916 29.1885 ;
               RECT 17.844 29.8405 17.916 29.8655 ;
               RECT 17.844 30.3635 17.916 30.3885 ;
               RECT 17.844 31.0405 17.916 31.0655 ;
               RECT 17.844 31.5635 17.916 31.5885 ;
               RECT 17.844 32.2405 17.916 32.2655 ;
               RECT 17.844 32.7635 17.916 32.7885 ;
               RECT 17.844 33.4405 17.916 33.4655 ;
               RECT 17.844 33.9635 17.916 33.9885 ;
               RECT 17.844 34.6405 17.916 34.6655 ;
               RECT 17.844 35.1635 17.916 35.1885 ;
               RECT 17.844 35.8405 17.916 35.8655 ;
               RECT 17.844 36.3635 17.916 36.3885 ;
               RECT 17.844 37.0405 17.916 37.0655 ;
               RECT 17.844 37.5635 17.916 37.5885 ;
               RECT 17.844 38.2405 17.916 38.2655 ;
               RECT 17.844 38.7635 17.916 38.7885 ;
               RECT 17.844 39.4405 17.916 39.4655 ;
               RECT 17.844 39.9635 17.916 39.9885 ;
               RECT 17.844 40.6405 17.916 40.6655 ;
               RECT 17.844 41.1635 17.916 41.1885 ;
               RECT 17.844 41.8405 17.916 41.8655 ;
               RECT 17.844 42.3635 17.916 42.3885 ;
               RECT 17.844 43.0405 17.916 43.0655 ;
               RECT 17.844 43.5635 17.916 43.5885 ;
               RECT 17.844 44.2405 17.916 44.2655 ;
               RECT 17.844 44.7635 17.916 44.7885 ;
               RECT 17.844 45.4405 17.916 45.4655 ;
               RECT 17.844 45.9635 17.916 45.9885 ;
               RECT 17.844 46.6405 17.916 46.6655 ;
               RECT 17.844 47.1635 17.916 47.1885 ;
               RECT 17.844 47.8405 17.916 47.8655 ;
               RECT 17.844 48.3635 17.916 48.3885 ;
               RECT 17.844 49.1875 17.916 49.2125 ;
               RECT 17.844 49.849 17.916 49.874 ;
               RECT 17.844 50.1475 17.916 50.1725 ;
               RECT 17.844 50.6275 17.916 50.6525 ;
               RECT 17.844 51.1075 17.916 51.1325 ;
               RECT 17.844 51.5875 17.916 51.6125 ;
               RECT 17.844 52.0675 17.916 52.0925 ;
               RECT 17.844 52.5475 17.916 52.5725 ;
               RECT 17.844 53.0275 17.916 53.0525 ;
               RECT 17.844 53.5075 17.916 53.5325 ;
               RECT 17.844 54.4675 17.916 54.4925 ;
               RECT 17.844 54.9475 17.916 54.9725 ;
               RECT 17.844 55.4275 17.916 55.4525 ;
               RECT 17.844 55.9075 17.916 55.9325 ;
               RECT 17.844 56.9605 17.916 56.9855 ;
               RECT 17.844 57.4835 17.916 57.5085 ;
               RECT 17.844 58.1605 17.916 58.1855 ;
               RECT 17.844 58.6835 17.916 58.7085 ;
               RECT 17.844 59.3605 17.916 59.3855 ;
               RECT 17.844 59.8835 17.916 59.9085 ;
               RECT 17.844 60.5605 17.916 60.5855 ;
               RECT 17.844 61.0835 17.916 61.1085 ;
               RECT 17.844 61.7605 17.916 61.7855 ;
               RECT 17.844 62.2835 17.916 62.3085 ;
               RECT 17.844 62.9605 17.916 62.9855 ;
               RECT 17.844 63.4835 17.916 63.5085 ;
               RECT 17.844 64.1605 17.916 64.1855 ;
               RECT 17.844 64.6835 17.916 64.7085 ;
               RECT 17.844 65.3605 17.916 65.3855 ;
               RECT 17.844 65.8835 17.916 65.9085 ;
               RECT 17.844 66.5605 17.916 66.5855 ;
               RECT 17.844 67.0835 17.916 67.1085 ;
               RECT 17.844 67.7605 17.916 67.7855 ;
               RECT 17.844 68.2835 17.916 68.3085 ;
               RECT 17.844 68.9605 17.916 68.9855 ;
               RECT 17.844 69.4835 17.916 69.5085 ;
               RECT 17.844 70.1605 17.916 70.1855 ;
               RECT 17.844 70.6835 17.916 70.7085 ;
               RECT 17.844 71.3605 17.916 71.3855 ;
               RECT 17.844 71.8835 17.916 71.9085 ;
               RECT 17.844 72.5605 17.916 72.5855 ;
               RECT 17.844 73.0835 17.916 73.1085 ;
               RECT 17.844 73.7605 17.916 73.7855 ;
               RECT 17.844 74.2835 17.916 74.3085 ;
               RECT 17.844 74.9605 17.916 74.9855 ;
               RECT 17.844 75.4835 17.916 75.5085 ;
               RECT 17.844 76.1605 17.916 76.1855 ;
               RECT 17.844 76.6835 17.916 76.7085 ;
               RECT 17.844 77.3605 17.916 77.3855 ;
               RECT 17.844 77.8835 17.916 77.9085 ;
               RECT 17.844 78.5605 17.916 78.5855 ;
               RECT 17.844 79.0835 17.916 79.1085 ;
               RECT 17.844 79.7605 17.916 79.7855 ;
               RECT 17.844 80.2835 17.916 80.3085 ;
               RECT 17.844 80.9605 17.916 80.9855 ;
               RECT 17.844 81.4835 17.916 81.5085 ;
               RECT 17.844 82.1605 17.916 82.1855 ;
               RECT 17.844 82.6835 17.916 82.7085 ;
               RECT 17.844 83.3605 17.916 83.3855 ;
               RECT 17.844 83.8835 17.916 83.9085 ;
               RECT 17.844 84.5605 17.916 84.5855 ;
               RECT 17.844 85.0835 17.916 85.1085 ;
               RECT 17.844 85.7605 17.916 85.7855 ;
               RECT 17.844 86.2835 17.916 86.3085 ;
               RECT 17.844 86.9605 17.916 86.9855 ;
               RECT 17.844 87.4835 17.916 87.5085 ;
               RECT 17.844 88.1605 17.916 88.1855 ;
               RECT 17.844 88.6835 17.916 88.7085 ;
               RECT 17.844 89.3605 17.916 89.3855 ;
               RECT 17.844 89.8835 17.916 89.9085 ;
               RECT 17.844 90.5605 17.916 90.5855 ;
               RECT 17.844 91.0835 17.916 91.1085 ;
               RECT 17.844 91.7605 17.916 91.7855 ;
               RECT 17.844 92.2835 17.916 92.3085 ;
               RECT 17.844 92.9605 17.916 92.9855 ;
               RECT 17.844 93.4835 17.916 93.5085 ;
               RECT 17.844 94.1605 17.916 94.1855 ;
               RECT 17.844 94.6835 17.916 94.7085 ;
               RECT 17.844 95.3605 17.916 95.3855 ;
               RECT 17.844 95.8835 17.916 95.9085 ;
               RECT 17.844 96.5605 17.916 96.5855 ;
               RECT 17.844 97.0835 17.916 97.1085 ;
               RECT 17.844 97.7605 17.916 97.7855 ;
               RECT 17.844 98.2835 17.916 98.3085 ;
               RECT 17.844 98.9605 17.916 98.9855 ;
               RECT 17.844 99.4835 17.916 99.5085 ;
               RECT 17.844 100.1605 17.916 100.1855 ;
               RECT 17.844 100.6835 17.916 100.7085 ;
               RECT 17.844 101.3605 17.916 101.3855 ;
               RECT 17.844 101.8835 17.916 101.9085 ;
               RECT 17.844 102.5605 17.916 102.5855 ;
               RECT 17.844 103.0835 17.916 103.1085 ;
               RECT 17.844 103.7605 17.916 103.7855 ;
               RECT 17.844 104.2835 17.916 104.3085 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.148 0.6 18.188 104.52 ;
               LAYER v4 ;
               RECT 18.148 0.729 18.188 0.765 ;
               RECT 18.148 0.958 18.188 0.994 ;
               RECT 18.148 1.635 18.188 1.671 ;
               RECT 18.148 1.929 18.188 1.965 ;
               RECT 18.148 2.158 18.188 2.194 ;
               RECT 18.148 2.835 18.188 2.871 ;
               RECT 18.148 3.129 18.188 3.165 ;
               RECT 18.148 3.358 18.188 3.394 ;
               RECT 18.148 4.035 18.188 4.071 ;
               RECT 18.148 4.329 18.188 4.365 ;
               RECT 18.148 4.558 18.188 4.594 ;
               RECT 18.148 5.235 18.188 5.271 ;
               RECT 18.148 5.529 18.188 5.565 ;
               RECT 18.148 5.758 18.188 5.794 ;
               RECT 18.148 6.435 18.188 6.471 ;
               RECT 18.148 6.729 18.188 6.765 ;
               RECT 18.148 6.958 18.188 6.994 ;
               RECT 18.148 7.635 18.188 7.671 ;
               RECT 18.148 7.929 18.188 7.965 ;
               RECT 18.148 8.158 18.188 8.194 ;
               RECT 18.148 8.835 18.188 8.871 ;
               RECT 18.148 9.129 18.188 9.165 ;
               RECT 18.148 9.358 18.188 9.394 ;
               RECT 18.148 10.035 18.188 10.071 ;
               RECT 18.148 10.329 18.188 10.365 ;
               RECT 18.148 10.558 18.188 10.594 ;
               RECT 18.148 11.235 18.188 11.271 ;
               RECT 18.148 11.529 18.188 11.565 ;
               RECT 18.148 11.758 18.188 11.794 ;
               RECT 18.148 12.435 18.188 12.471 ;
               RECT 18.148 12.729 18.188 12.765 ;
               RECT 18.148 12.958 18.188 12.994 ;
               RECT 18.148 13.635 18.188 13.671 ;
               RECT 18.148 13.929 18.188 13.965 ;
               RECT 18.148 14.158 18.188 14.194 ;
               RECT 18.148 14.835 18.188 14.871 ;
               RECT 18.148 15.129 18.188 15.165 ;
               RECT 18.148 15.358 18.188 15.394 ;
               RECT 18.148 16.035 18.188 16.071 ;
               RECT 18.148 16.329 18.188 16.365 ;
               RECT 18.148 16.558 18.188 16.594 ;
               RECT 18.148 17.235 18.188 17.271 ;
               RECT 18.148 17.529 18.188 17.565 ;
               RECT 18.148 17.758 18.188 17.794 ;
               RECT 18.148 18.435 18.188 18.471 ;
               RECT 18.148 18.729 18.188 18.765 ;
               RECT 18.148 18.958 18.188 18.994 ;
               RECT 18.148 19.635 18.188 19.671 ;
               RECT 18.148 19.929 18.188 19.965 ;
               RECT 18.148 20.158 18.188 20.194 ;
               RECT 18.148 20.835 18.188 20.871 ;
               RECT 18.148 21.129 18.188 21.165 ;
               RECT 18.148 21.358 18.188 21.394 ;
               RECT 18.148 22.035 18.188 22.071 ;
               RECT 18.148 22.329 18.188 22.365 ;
               RECT 18.148 22.558 18.188 22.594 ;
               RECT 18.148 23.235 18.188 23.271 ;
               RECT 18.148 23.529 18.188 23.565 ;
               RECT 18.148 23.758 18.188 23.794 ;
               RECT 18.148 24.435 18.188 24.471 ;
               RECT 18.148 24.729 18.188 24.765 ;
               RECT 18.148 24.958 18.188 24.994 ;
               RECT 18.148 25.635 18.188 25.671 ;
               RECT 18.148 25.929 18.188 25.965 ;
               RECT 18.148 26.158 18.188 26.194 ;
               RECT 18.148 26.835 18.188 26.871 ;
               RECT 18.148 27.129 18.188 27.165 ;
               RECT 18.148 27.358 18.188 27.394 ;
               RECT 18.148 28.035 18.188 28.071 ;
               RECT 18.148 28.329 18.188 28.365 ;
               RECT 18.148 28.558 18.188 28.594 ;
               RECT 18.148 29.235 18.188 29.271 ;
               RECT 18.148 29.529 18.188 29.565 ;
               RECT 18.148 29.758 18.188 29.794 ;
               RECT 18.148 30.435 18.188 30.471 ;
               RECT 18.148 30.729 18.188 30.765 ;
               RECT 18.148 30.958 18.188 30.994 ;
               RECT 18.148 31.635 18.188 31.671 ;
               RECT 18.148 31.929 18.188 31.965 ;
               RECT 18.148 32.158 18.188 32.194 ;
               RECT 18.148 32.835 18.188 32.871 ;
               RECT 18.148 33.129 18.188 33.165 ;
               RECT 18.148 33.358 18.188 33.394 ;
               RECT 18.148 34.035 18.188 34.071 ;
               RECT 18.148 34.329 18.188 34.365 ;
               RECT 18.148 34.558 18.188 34.594 ;
               RECT 18.148 35.235 18.188 35.271 ;
               RECT 18.148 35.529 18.188 35.565 ;
               RECT 18.148 35.758 18.188 35.794 ;
               RECT 18.148 36.435 18.188 36.471 ;
               RECT 18.148 36.729 18.188 36.765 ;
               RECT 18.148 36.958 18.188 36.994 ;
               RECT 18.148 37.635 18.188 37.671 ;
               RECT 18.148 37.929 18.188 37.965 ;
               RECT 18.148 38.158 18.188 38.194 ;
               RECT 18.148 38.835 18.188 38.871 ;
               RECT 18.148 39.129 18.188 39.165 ;
               RECT 18.148 39.358 18.188 39.394 ;
               RECT 18.148 40.035 18.188 40.071 ;
               RECT 18.148 40.329 18.188 40.365 ;
               RECT 18.148 40.558 18.188 40.594 ;
               RECT 18.148 41.235 18.188 41.271 ;
               RECT 18.148 41.529 18.188 41.565 ;
               RECT 18.148 41.758 18.188 41.794 ;
               RECT 18.148 42.435 18.188 42.471 ;
               RECT 18.148 42.729 18.188 42.765 ;
               RECT 18.148 42.958 18.188 42.994 ;
               RECT 18.148 43.635 18.188 43.671 ;
               RECT 18.148 43.929 18.188 43.965 ;
               RECT 18.148 44.158 18.188 44.194 ;
               RECT 18.148 44.835 18.188 44.871 ;
               RECT 18.148 45.129 18.188 45.165 ;
               RECT 18.148 45.358 18.188 45.394 ;
               RECT 18.148 46.035 18.188 46.071 ;
               RECT 18.148 46.329 18.188 46.365 ;
               RECT 18.148 46.558 18.188 46.594 ;
               RECT 18.148 47.235 18.188 47.271 ;
               RECT 18.148 47.529 18.188 47.565 ;
               RECT 18.148 47.758 18.188 47.794 ;
               RECT 18.148 48.435 18.188 48.471 ;
               RECT 18.148 49.182 18.188 49.218 ;
               RECT 18.148 49.662 18.188 49.698 ;
               RECT 18.148 50.142 18.188 50.178 ;
               RECT 18.148 50.622 18.188 50.658 ;
               RECT 18.148 51.102 18.188 51.138 ;
               RECT 18.148 51.582 18.188 51.618 ;
               RECT 18.148 52.062 18.188 52.098 ;
               RECT 18.148 52.542 18.188 52.578 ;
               RECT 18.148 53.022 18.188 53.058 ;
               RECT 18.148 53.502 18.188 53.538 ;
               RECT 18.148 53.982 18.188 54.018 ;
               RECT 18.148 54.462 18.188 54.498 ;
               RECT 18.148 54.942 18.188 54.978 ;
               RECT 18.148 55.422 18.188 55.458 ;
               RECT 18.148 55.902 18.188 55.938 ;
               RECT 18.148 56.649 18.188 56.685 ;
               RECT 18.148 56.878 18.188 56.914 ;
               RECT 18.148 57.555 18.188 57.591 ;
               RECT 18.148 57.849 18.188 57.885 ;
               RECT 18.148 58.078 18.188 58.114 ;
               RECT 18.148 58.755 18.188 58.791 ;
               RECT 18.148 59.049 18.188 59.085 ;
               RECT 18.148 59.278 18.188 59.314 ;
               RECT 18.148 59.955 18.188 59.991 ;
               RECT 18.148 60.249 18.188 60.285 ;
               RECT 18.148 60.478 18.188 60.514 ;
               RECT 18.148 61.155 18.188 61.191 ;
               RECT 18.148 61.449 18.188 61.485 ;
               RECT 18.148 61.678 18.188 61.714 ;
               RECT 18.148 62.355 18.188 62.391 ;
               RECT 18.148 62.649 18.188 62.685 ;
               RECT 18.148 62.878 18.188 62.914 ;
               RECT 18.148 63.555 18.188 63.591 ;
               RECT 18.148 63.849 18.188 63.885 ;
               RECT 18.148 64.078 18.188 64.114 ;
               RECT 18.148 64.755 18.188 64.791 ;
               RECT 18.148 65.049 18.188 65.085 ;
               RECT 18.148 65.278 18.188 65.314 ;
               RECT 18.148 65.955 18.188 65.991 ;
               RECT 18.148 66.249 18.188 66.285 ;
               RECT 18.148 66.478 18.188 66.514 ;
               RECT 18.148 67.155 18.188 67.191 ;
               RECT 18.148 67.449 18.188 67.485 ;
               RECT 18.148 67.678 18.188 67.714 ;
               RECT 18.148 68.355 18.188 68.391 ;
               RECT 18.148 68.649 18.188 68.685 ;
               RECT 18.148 68.878 18.188 68.914 ;
               RECT 18.148 69.555 18.188 69.591 ;
               RECT 18.148 69.849 18.188 69.885 ;
               RECT 18.148 70.078 18.188 70.114 ;
               RECT 18.148 70.755 18.188 70.791 ;
               RECT 18.148 71.049 18.188 71.085 ;
               RECT 18.148 71.278 18.188 71.314 ;
               RECT 18.148 71.955 18.188 71.991 ;
               RECT 18.148 72.249 18.188 72.285 ;
               RECT 18.148 72.478 18.188 72.514 ;
               RECT 18.148 73.155 18.188 73.191 ;
               RECT 18.148 73.449 18.188 73.485 ;
               RECT 18.148 73.678 18.188 73.714 ;
               RECT 18.148 74.355 18.188 74.391 ;
               RECT 18.148 74.649 18.188 74.685 ;
               RECT 18.148 74.878 18.188 74.914 ;
               RECT 18.148 75.555 18.188 75.591 ;
               RECT 18.148 75.849 18.188 75.885 ;
               RECT 18.148 76.078 18.188 76.114 ;
               RECT 18.148 76.755 18.188 76.791 ;
               RECT 18.148 77.049 18.188 77.085 ;
               RECT 18.148 77.278 18.188 77.314 ;
               RECT 18.148 77.955 18.188 77.991 ;
               RECT 18.148 78.249 18.188 78.285 ;
               RECT 18.148 78.478 18.188 78.514 ;
               RECT 18.148 79.155 18.188 79.191 ;
               RECT 18.148 79.449 18.188 79.485 ;
               RECT 18.148 79.678 18.188 79.714 ;
               RECT 18.148 80.355 18.188 80.391 ;
               RECT 18.148 80.649 18.188 80.685 ;
               RECT 18.148 80.878 18.188 80.914 ;
               RECT 18.148 81.555 18.188 81.591 ;
               RECT 18.148 81.849 18.188 81.885 ;
               RECT 18.148 82.078 18.188 82.114 ;
               RECT 18.148 82.755 18.188 82.791 ;
               RECT 18.148 83.049 18.188 83.085 ;
               RECT 18.148 83.278 18.188 83.314 ;
               RECT 18.148 83.955 18.188 83.991 ;
               RECT 18.148 84.249 18.188 84.285 ;
               RECT 18.148 84.478 18.188 84.514 ;
               RECT 18.148 85.155 18.188 85.191 ;
               RECT 18.148 85.449 18.188 85.485 ;
               RECT 18.148 85.678 18.188 85.714 ;
               RECT 18.148 86.355 18.188 86.391 ;
               RECT 18.148 86.649 18.188 86.685 ;
               RECT 18.148 86.878 18.188 86.914 ;
               RECT 18.148 87.555 18.188 87.591 ;
               RECT 18.148 87.849 18.188 87.885 ;
               RECT 18.148 88.078 18.188 88.114 ;
               RECT 18.148 88.755 18.188 88.791 ;
               RECT 18.148 89.049 18.188 89.085 ;
               RECT 18.148 89.278 18.188 89.314 ;
               RECT 18.148 89.955 18.188 89.991 ;
               RECT 18.148 90.249 18.188 90.285 ;
               RECT 18.148 90.478 18.188 90.514 ;
               RECT 18.148 91.155 18.188 91.191 ;
               RECT 18.148 91.449 18.188 91.485 ;
               RECT 18.148 91.678 18.188 91.714 ;
               RECT 18.148 92.355 18.188 92.391 ;
               RECT 18.148 92.649 18.188 92.685 ;
               RECT 18.148 92.878 18.188 92.914 ;
               RECT 18.148 93.555 18.188 93.591 ;
               RECT 18.148 93.849 18.188 93.885 ;
               RECT 18.148 94.078 18.188 94.114 ;
               RECT 18.148 94.755 18.188 94.791 ;
               RECT 18.148 95.049 18.188 95.085 ;
               RECT 18.148 95.278 18.188 95.314 ;
               RECT 18.148 95.955 18.188 95.991 ;
               RECT 18.148 96.249 18.188 96.285 ;
               RECT 18.148 96.478 18.188 96.514 ;
               RECT 18.148 97.155 18.188 97.191 ;
               RECT 18.148 97.449 18.188 97.485 ;
               RECT 18.148 97.678 18.188 97.714 ;
               RECT 18.148 98.355 18.188 98.391 ;
               RECT 18.148 98.649 18.188 98.685 ;
               RECT 18.148 98.878 18.188 98.914 ;
               RECT 18.148 99.555 18.188 99.591 ;
               RECT 18.148 99.849 18.188 99.885 ;
               RECT 18.148 100.078 18.188 100.114 ;
               RECT 18.148 100.755 18.188 100.791 ;
               RECT 18.148 101.049 18.188 101.085 ;
               RECT 18.148 101.278 18.188 101.314 ;
               RECT 18.148 101.955 18.188 101.991 ;
               RECT 18.148 102.249 18.188 102.285 ;
               RECT 18.148 102.478 18.188 102.514 ;
               RECT 18.148 103.155 18.188 103.191 ;
               RECT 18.148 103.449 18.188 103.485 ;
               RECT 18.148 103.678 18.188 103.714 ;
               RECT 18.148 104.355 18.188 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.356 0.5695 18.396 104.5505 ;
               LAYER v4 ;
               RECT 18.356 1.035 18.396 1.071 ;
               RECT 18.356 1.558 18.396 1.594 ;
               RECT 18.356 2.235 18.396 2.271 ;
               RECT 18.356 2.758 18.396 2.794 ;
               RECT 18.356 3.435 18.396 3.471 ;
               RECT 18.356 3.958 18.396 3.994 ;
               RECT 18.356 4.635 18.396 4.671 ;
               RECT 18.356 5.158 18.396 5.194 ;
               RECT 18.356 5.835 18.396 5.871 ;
               RECT 18.356 6.358 18.396 6.394 ;
               RECT 18.356 7.035 18.396 7.071 ;
               RECT 18.356 7.558 18.396 7.594 ;
               RECT 18.356 8.235 18.396 8.271 ;
               RECT 18.356 8.758 18.396 8.794 ;
               RECT 18.356 9.435 18.396 9.471 ;
               RECT 18.356 9.958 18.396 9.994 ;
               RECT 18.356 10.635 18.396 10.671 ;
               RECT 18.356 11.158 18.396 11.194 ;
               RECT 18.356 11.835 18.396 11.871 ;
               RECT 18.356 12.358 18.396 12.394 ;
               RECT 18.356 13.035 18.396 13.071 ;
               RECT 18.356 13.558 18.396 13.594 ;
               RECT 18.356 14.235 18.396 14.271 ;
               RECT 18.356 14.758 18.396 14.794 ;
               RECT 18.356 15.435 18.396 15.471 ;
               RECT 18.356 15.958 18.396 15.994 ;
               RECT 18.356 16.635 18.396 16.671 ;
               RECT 18.356 17.158 18.396 17.194 ;
               RECT 18.356 17.835 18.396 17.871 ;
               RECT 18.356 18.358 18.396 18.394 ;
               RECT 18.356 19.035 18.396 19.071 ;
               RECT 18.356 19.558 18.396 19.594 ;
               RECT 18.356 20.235 18.396 20.271 ;
               RECT 18.356 20.758 18.396 20.794 ;
               RECT 18.356 21.435 18.396 21.471 ;
               RECT 18.356 21.958 18.396 21.994 ;
               RECT 18.356 22.635 18.396 22.671 ;
               RECT 18.356 23.158 18.396 23.194 ;
               RECT 18.356 23.835 18.396 23.871 ;
               RECT 18.356 24.358 18.396 24.394 ;
               RECT 18.356 25.035 18.396 25.071 ;
               RECT 18.356 25.558 18.396 25.594 ;
               RECT 18.356 26.235 18.396 26.271 ;
               RECT 18.356 26.758 18.396 26.794 ;
               RECT 18.356 27.435 18.396 27.471 ;
               RECT 18.356 27.958 18.396 27.994 ;
               RECT 18.356 28.635 18.396 28.671 ;
               RECT 18.356 29.158 18.396 29.194 ;
               RECT 18.356 29.835 18.396 29.871 ;
               RECT 18.356 30.358 18.396 30.394 ;
               RECT 18.356 31.035 18.396 31.071 ;
               RECT 18.356 31.558 18.396 31.594 ;
               RECT 18.356 32.235 18.396 32.271 ;
               RECT 18.356 32.758 18.396 32.794 ;
               RECT 18.356 33.435 18.396 33.471 ;
               RECT 18.356 33.958 18.396 33.994 ;
               RECT 18.356 34.635 18.396 34.671 ;
               RECT 18.356 35.158 18.396 35.194 ;
               RECT 18.356 35.835 18.396 35.871 ;
               RECT 18.356 36.358 18.396 36.394 ;
               RECT 18.356 37.035 18.396 37.071 ;
               RECT 18.356 37.558 18.396 37.594 ;
               RECT 18.356 38.235 18.396 38.271 ;
               RECT 18.356 38.758 18.396 38.794 ;
               RECT 18.356 39.435 18.396 39.471 ;
               RECT 18.356 39.958 18.396 39.994 ;
               RECT 18.356 40.635 18.396 40.671 ;
               RECT 18.356 41.158 18.396 41.194 ;
               RECT 18.356 41.835 18.396 41.871 ;
               RECT 18.356 42.358 18.396 42.394 ;
               RECT 18.356 43.035 18.396 43.071 ;
               RECT 18.356 43.558 18.396 43.594 ;
               RECT 18.356 44.235 18.396 44.271 ;
               RECT 18.356 44.758 18.396 44.794 ;
               RECT 18.356 45.435 18.396 45.471 ;
               RECT 18.356 45.958 18.396 45.994 ;
               RECT 18.356 46.635 18.396 46.671 ;
               RECT 18.356 47.158 18.396 47.194 ;
               RECT 18.356 47.835 18.396 47.871 ;
               RECT 18.356 48.358 18.396 48.394 ;
               RECT 18.356 49.182 18.396 49.218 ;
               RECT 18.356 49.6675 18.396 49.6925 ;
               RECT 18.356 49.8435 18.396 49.8795 ;
               RECT 18.356 50.142 18.396 50.178 ;
               RECT 18.356 50.622 18.396 50.658 ;
               RECT 18.356 51.102 18.396 51.138 ;
               RECT 18.356 51.582 18.396 51.618 ;
               RECT 18.356 52.062 18.396 52.098 ;
               RECT 18.356 52.542 18.396 52.578 ;
               RECT 18.356 53.022 18.396 53.058 ;
               RECT 18.356 53.502 18.396 53.538 ;
               RECT 18.356 53.982 18.396 54.018 ;
               RECT 18.356 54.942 18.396 54.978 ;
               RECT 18.356 55.422 18.396 55.458 ;
               RECT 18.356 55.902 18.396 55.938 ;
               RECT 18.356 56.955 18.396 56.991 ;
               RECT 18.356 57.478 18.396 57.514 ;
               RECT 18.356 58.155 18.396 58.191 ;
               RECT 18.356 58.678 18.396 58.714 ;
               RECT 18.356 59.355 18.396 59.391 ;
               RECT 18.356 59.878 18.396 59.914 ;
               RECT 18.356 60.555 18.396 60.591 ;
               RECT 18.356 61.078 18.396 61.114 ;
               RECT 18.356 61.755 18.396 61.791 ;
               RECT 18.356 62.278 18.396 62.314 ;
               RECT 18.356 62.955 18.396 62.991 ;
               RECT 18.356 63.478 18.396 63.514 ;
               RECT 18.356 64.155 18.396 64.191 ;
               RECT 18.356 64.678 18.396 64.714 ;
               RECT 18.356 65.355 18.396 65.391 ;
               RECT 18.356 65.878 18.396 65.914 ;
               RECT 18.356 66.555 18.396 66.591 ;
               RECT 18.356 67.078 18.396 67.114 ;
               RECT 18.356 67.755 18.396 67.791 ;
               RECT 18.356 68.278 18.396 68.314 ;
               RECT 18.356 68.955 18.396 68.991 ;
               RECT 18.356 69.478 18.396 69.514 ;
               RECT 18.356 70.155 18.396 70.191 ;
               RECT 18.356 70.678 18.396 70.714 ;
               RECT 18.356 71.355 18.396 71.391 ;
               RECT 18.356 71.878 18.396 71.914 ;
               RECT 18.356 72.555 18.396 72.591 ;
               RECT 18.356 73.078 18.396 73.114 ;
               RECT 18.356 73.755 18.396 73.791 ;
               RECT 18.356 74.278 18.396 74.314 ;
               RECT 18.356 74.955 18.396 74.991 ;
               RECT 18.356 75.478 18.396 75.514 ;
               RECT 18.356 76.155 18.396 76.191 ;
               RECT 18.356 76.678 18.396 76.714 ;
               RECT 18.356 77.355 18.396 77.391 ;
               RECT 18.356 77.878 18.396 77.914 ;
               RECT 18.356 78.555 18.396 78.591 ;
               RECT 18.356 79.078 18.396 79.114 ;
               RECT 18.356 79.755 18.396 79.791 ;
               RECT 18.356 80.278 18.396 80.314 ;
               RECT 18.356 80.955 18.396 80.991 ;
               RECT 18.356 81.478 18.396 81.514 ;
               RECT 18.356 82.155 18.396 82.191 ;
               RECT 18.356 82.678 18.396 82.714 ;
               RECT 18.356 83.355 18.396 83.391 ;
               RECT 18.356 83.878 18.396 83.914 ;
               RECT 18.356 84.555 18.396 84.591 ;
               RECT 18.356 85.078 18.396 85.114 ;
               RECT 18.356 85.755 18.396 85.791 ;
               RECT 18.356 86.278 18.396 86.314 ;
               RECT 18.356 86.955 18.396 86.991 ;
               RECT 18.356 87.478 18.396 87.514 ;
               RECT 18.356 88.155 18.396 88.191 ;
               RECT 18.356 88.678 18.396 88.714 ;
               RECT 18.356 89.355 18.396 89.391 ;
               RECT 18.356 89.878 18.396 89.914 ;
               RECT 18.356 90.555 18.396 90.591 ;
               RECT 18.356 91.078 18.396 91.114 ;
               RECT 18.356 91.755 18.396 91.791 ;
               RECT 18.356 92.278 18.396 92.314 ;
               RECT 18.356 92.955 18.396 92.991 ;
               RECT 18.356 93.478 18.396 93.514 ;
               RECT 18.356 94.155 18.396 94.191 ;
               RECT 18.356 94.678 18.396 94.714 ;
               RECT 18.356 95.355 18.396 95.391 ;
               RECT 18.356 95.878 18.396 95.914 ;
               RECT 18.356 96.555 18.396 96.591 ;
               RECT 18.356 97.078 18.396 97.114 ;
               RECT 18.356 97.755 18.396 97.791 ;
               RECT 18.356 98.278 18.396 98.314 ;
               RECT 18.356 98.955 18.396 98.991 ;
               RECT 18.356 99.478 18.396 99.514 ;
               RECT 18.356 100.155 18.396 100.191 ;
               RECT 18.356 100.678 18.396 100.714 ;
               RECT 18.356 101.355 18.396 101.391 ;
               RECT 18.356 101.878 18.396 101.914 ;
               RECT 18.356 102.555 18.396 102.591 ;
               RECT 18.356 103.078 18.396 103.114 ;
               RECT 18.356 103.755 18.396 103.791 ;
               RECT 18.356 104.278 18.396 104.314 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.664 0.5695 18.736 104.5505 ;
               LAYER v4 ;
               RECT 18.664 0.7345 18.736 0.7595 ;
               RECT 18.664 0.9635 18.736 0.9885 ;
               RECT 18.664 1.6405 18.736 1.6655 ;
               RECT 18.664 1.9345 18.736 1.9595 ;
               RECT 18.664 2.1635 18.736 2.1885 ;
               RECT 18.664 2.6115 18.736 2.6365 ;
               RECT 18.664 2.8405 18.736 2.8655 ;
               RECT 18.664 3.1345 18.736 3.1595 ;
               RECT 18.664 3.3635 18.736 3.3885 ;
               RECT 18.664 4.0405 18.736 4.0655 ;
               RECT 18.664 4.3345 18.736 4.3595 ;
               RECT 18.664 4.5635 18.736 4.5885 ;
               RECT 18.664 5.0115 18.736 5.0365 ;
               RECT 18.664 5.2405 18.736 5.2655 ;
               RECT 18.664 5.5345 18.736 5.5595 ;
               RECT 18.664 5.7635 18.736 5.7885 ;
               RECT 18.664 6.4405 18.736 6.4655 ;
               RECT 18.664 6.7345 18.736 6.7595 ;
               RECT 18.664 6.9635 18.736 6.9885 ;
               RECT 18.664 7.4115 18.736 7.4365 ;
               RECT 18.664 7.6405 18.736 7.6655 ;
               RECT 18.664 7.9345 18.736 7.9595 ;
               RECT 18.664 8.1635 18.736 8.1885 ;
               RECT 18.664 8.8405 18.736 8.8655 ;
               RECT 18.664 9.1345 18.736 9.1595 ;
               RECT 18.664 9.3635 18.736 9.3885 ;
               RECT 18.664 9.8115 18.736 9.8365 ;
               RECT 18.664 10.0405 18.736 10.0655 ;
               RECT 18.664 10.3345 18.736 10.3595 ;
               RECT 18.664 10.5635 18.736 10.5885 ;
               RECT 18.664 11.2405 18.736 11.2655 ;
               RECT 18.664 11.5345 18.736 11.5595 ;
               RECT 18.664 11.7635 18.736 11.7885 ;
               RECT 18.664 12.2115 18.736 12.2365 ;
               RECT 18.664 12.4405 18.736 12.4655 ;
               RECT 18.664 12.7345 18.736 12.7595 ;
               RECT 18.664 12.9635 18.736 12.9885 ;
               RECT 18.664 13.6405 18.736 13.6655 ;
               RECT 18.664 13.9345 18.736 13.9595 ;
               RECT 18.664 14.1635 18.736 14.1885 ;
               RECT 18.664 14.6115 18.736 14.6365 ;
               RECT 18.664 14.8405 18.736 14.8655 ;
               RECT 18.664 15.1345 18.736 15.1595 ;
               RECT 18.664 15.3635 18.736 15.3885 ;
               RECT 18.664 16.0405 18.736 16.0655 ;
               RECT 18.664 16.3345 18.736 16.3595 ;
               RECT 18.664 16.5635 18.736 16.5885 ;
               RECT 18.664 17.0115 18.736 17.0365 ;
               RECT 18.664 17.2405 18.736 17.2655 ;
               RECT 18.664 17.5345 18.736 17.5595 ;
               RECT 18.664 17.7635 18.736 17.7885 ;
               RECT 18.664 18.4405 18.736 18.4655 ;
               RECT 18.664 18.7345 18.736 18.7595 ;
               RECT 18.664 18.9635 18.736 18.9885 ;
               RECT 18.664 19.4115 18.736 19.4365 ;
               RECT 18.664 19.6405 18.736 19.6655 ;
               RECT 18.664 19.9345 18.736 19.9595 ;
               RECT 18.664 20.1635 18.736 20.1885 ;
               RECT 18.664 20.8405 18.736 20.8655 ;
               RECT 18.664 21.1345 18.736 21.1595 ;
               RECT 18.664 21.3635 18.736 21.3885 ;
               RECT 18.664 21.8115 18.736 21.8365 ;
               RECT 18.664 22.0405 18.736 22.0655 ;
               RECT 18.664 22.3345 18.736 22.3595 ;
               RECT 18.664 22.5635 18.736 22.5885 ;
               RECT 18.664 23.2405 18.736 23.2655 ;
               RECT 18.664 23.5345 18.736 23.5595 ;
               RECT 18.664 23.7635 18.736 23.7885 ;
               RECT 18.664 24.2115 18.736 24.2365 ;
               RECT 18.664 24.4405 18.736 24.4655 ;
               RECT 18.664 24.7345 18.736 24.7595 ;
               RECT 18.664 24.9635 18.736 24.9885 ;
               RECT 18.664 25.6405 18.736 25.6655 ;
               RECT 18.664 25.9345 18.736 25.9595 ;
               RECT 18.664 26.1635 18.736 26.1885 ;
               RECT 18.664 26.6115 18.736 26.6365 ;
               RECT 18.664 26.8405 18.736 26.8655 ;
               RECT 18.664 27.1345 18.736 27.1595 ;
               RECT 18.664 27.3635 18.736 27.3885 ;
               RECT 18.664 28.0405 18.736 28.0655 ;
               RECT 18.664 28.3345 18.736 28.3595 ;
               RECT 18.664 28.5635 18.736 28.5885 ;
               RECT 18.664 29.0115 18.736 29.0365 ;
               RECT 18.664 29.2405 18.736 29.2655 ;
               RECT 18.664 29.5345 18.736 29.5595 ;
               RECT 18.664 29.7635 18.736 29.7885 ;
               RECT 18.664 30.4405 18.736 30.4655 ;
               RECT 18.664 30.7345 18.736 30.7595 ;
               RECT 18.664 30.9635 18.736 30.9885 ;
               RECT 18.664 31.4115 18.736 31.4365 ;
               RECT 18.664 31.6405 18.736 31.6655 ;
               RECT 18.664 31.9345 18.736 31.9595 ;
               RECT 18.664 32.1635 18.736 32.1885 ;
               RECT 18.664 32.8405 18.736 32.8655 ;
               RECT 18.664 33.1345 18.736 33.1595 ;
               RECT 18.664 33.3635 18.736 33.3885 ;
               RECT 18.664 33.8115 18.736 33.8365 ;
               RECT 18.664 34.0405 18.736 34.0655 ;
               RECT 18.664 34.3345 18.736 34.3595 ;
               RECT 18.664 34.5635 18.736 34.5885 ;
               RECT 18.664 35.2405 18.736 35.2655 ;
               RECT 18.664 35.5345 18.736 35.5595 ;
               RECT 18.664 35.7635 18.736 35.7885 ;
               RECT 18.664 36.2115 18.736 36.2365 ;
               RECT 18.664 36.4405 18.736 36.4655 ;
               RECT 18.664 36.7345 18.736 36.7595 ;
               RECT 18.664 36.9635 18.736 36.9885 ;
               RECT 18.664 37.6405 18.736 37.6655 ;
               RECT 18.664 37.9345 18.736 37.9595 ;
               RECT 18.664 38.1635 18.736 38.1885 ;
               RECT 18.664 38.6115 18.736 38.6365 ;
               RECT 18.664 38.8405 18.736 38.8655 ;
               RECT 18.664 39.1345 18.736 39.1595 ;
               RECT 18.664 39.3635 18.736 39.3885 ;
               RECT 18.664 40.0405 18.736 40.0655 ;
               RECT 18.664 40.3345 18.736 40.3595 ;
               RECT 18.664 40.5635 18.736 40.5885 ;
               RECT 18.664 41.0115 18.736 41.0365 ;
               RECT 18.664 41.2405 18.736 41.2655 ;
               RECT 18.664 41.5345 18.736 41.5595 ;
               RECT 18.664 41.7635 18.736 41.7885 ;
               RECT 18.664 42.4405 18.736 42.4655 ;
               RECT 18.664 42.7345 18.736 42.7595 ;
               RECT 18.664 42.9635 18.736 42.9885 ;
               RECT 18.664 43.4115 18.736 43.4365 ;
               RECT 18.664 43.6405 18.736 43.6655 ;
               RECT 18.664 43.9345 18.736 43.9595 ;
               RECT 18.664 44.1635 18.736 44.1885 ;
               RECT 18.664 44.8405 18.736 44.8655 ;
               RECT 18.664 45.1345 18.736 45.1595 ;
               RECT 18.664 45.3635 18.736 45.3885 ;
               RECT 18.664 45.8115 18.736 45.8365 ;
               RECT 18.664 46.0405 18.736 46.0655 ;
               RECT 18.664 46.3345 18.736 46.3595 ;
               RECT 18.664 46.5635 18.736 46.5885 ;
               RECT 18.664 47.2405 18.736 47.2655 ;
               RECT 18.664 47.5345 18.736 47.5595 ;
               RECT 18.664 47.7635 18.736 47.7885 ;
               RECT 18.664 48.2115 18.736 48.2365 ;
               RECT 18.664 48.4405 18.736 48.4655 ;
               RECT 18.664 49.1875 18.736 49.2125 ;
               RECT 18.664 49.6675 18.736 49.6925 ;
               RECT 18.664 49.849 18.736 49.874 ;
               RECT 18.664 50.1475 18.736 50.1725 ;
               RECT 18.664 50.6275 18.736 50.6525 ;
               RECT 18.664 51.1075 18.736 51.1325 ;
               RECT 18.664 51.5875 18.736 51.6125 ;
               RECT 18.664 52.0675 18.736 52.0925 ;
               RECT 18.664 52.5475 18.736 52.5725 ;
               RECT 18.664 53.0275 18.736 53.0525 ;
               RECT 18.664 53.5075 18.736 53.5325 ;
               RECT 18.664 53.9875 18.736 54.0125 ;
               RECT 18.664 54.4675 18.736 54.4925 ;
               RECT 18.664 54.9475 18.736 54.9725 ;
               RECT 18.664 55.4275 18.736 55.4525 ;
               RECT 18.664 55.9075 18.736 55.9325 ;
               RECT 18.664 56.6545 18.736 56.6795 ;
               RECT 18.664 56.8835 18.736 56.9085 ;
               RECT 18.664 57.5605 18.736 57.5855 ;
               RECT 18.664 57.8545 18.736 57.8795 ;
               RECT 18.664 58.0835 18.736 58.1085 ;
               RECT 18.664 58.5315 18.736 58.5565 ;
               RECT 18.664 58.7605 18.736 58.7855 ;
               RECT 18.664 59.0545 18.736 59.0795 ;
               RECT 18.664 59.2835 18.736 59.3085 ;
               RECT 18.664 59.9605 18.736 59.9855 ;
               RECT 18.664 60.2545 18.736 60.2795 ;
               RECT 18.664 60.4835 18.736 60.5085 ;
               RECT 18.664 60.9315 18.736 60.9565 ;
               RECT 18.664 61.1605 18.736 61.1855 ;
               RECT 18.664 61.4545 18.736 61.4795 ;
               RECT 18.664 61.6835 18.736 61.7085 ;
               RECT 18.664 62.3605 18.736 62.3855 ;
               RECT 18.664 62.6545 18.736 62.6795 ;
               RECT 18.664 62.8835 18.736 62.9085 ;
               RECT 18.664 63.3315 18.736 63.3565 ;
               RECT 18.664 63.5605 18.736 63.5855 ;
               RECT 18.664 63.8545 18.736 63.8795 ;
               RECT 18.664 64.0835 18.736 64.1085 ;
               RECT 18.664 64.7605 18.736 64.7855 ;
               RECT 18.664 65.0545 18.736 65.0795 ;
               RECT 18.664 65.2835 18.736 65.3085 ;
               RECT 18.664 65.7315 18.736 65.7565 ;
               RECT 18.664 65.9605 18.736 65.9855 ;
               RECT 18.664 66.2545 18.736 66.2795 ;
               RECT 18.664 66.4835 18.736 66.5085 ;
               RECT 18.664 67.1605 18.736 67.1855 ;
               RECT 18.664 67.4545 18.736 67.4795 ;
               RECT 18.664 67.6835 18.736 67.7085 ;
               RECT 18.664 68.1315 18.736 68.1565 ;
               RECT 18.664 68.3605 18.736 68.3855 ;
               RECT 18.664 68.6545 18.736 68.6795 ;
               RECT 18.664 68.8835 18.736 68.9085 ;
               RECT 18.664 69.5605 18.736 69.5855 ;
               RECT 18.664 69.8545 18.736 69.8795 ;
               RECT 18.664 70.0835 18.736 70.1085 ;
               RECT 18.664 70.5315 18.736 70.5565 ;
               RECT 18.664 70.7605 18.736 70.7855 ;
               RECT 18.664 71.0545 18.736 71.0795 ;
               RECT 18.664 71.2835 18.736 71.3085 ;
               RECT 18.664 71.9605 18.736 71.9855 ;
               RECT 18.664 72.2545 18.736 72.2795 ;
               RECT 18.664 72.4835 18.736 72.5085 ;
               RECT 18.664 72.9315 18.736 72.9565 ;
               RECT 18.664 73.1605 18.736 73.1855 ;
               RECT 18.664 73.4545 18.736 73.4795 ;
               RECT 18.664 73.6835 18.736 73.7085 ;
               RECT 18.664 74.3605 18.736 74.3855 ;
               RECT 18.664 74.6545 18.736 74.6795 ;
               RECT 18.664 74.8835 18.736 74.9085 ;
               RECT 18.664 75.3315 18.736 75.3565 ;
               RECT 18.664 75.5605 18.736 75.5855 ;
               RECT 18.664 75.8545 18.736 75.8795 ;
               RECT 18.664 76.0835 18.736 76.1085 ;
               RECT 18.664 76.7605 18.736 76.7855 ;
               RECT 18.664 77.0545 18.736 77.0795 ;
               RECT 18.664 77.2835 18.736 77.3085 ;
               RECT 18.664 77.7315 18.736 77.7565 ;
               RECT 18.664 77.9605 18.736 77.9855 ;
               RECT 18.664 78.2545 18.736 78.2795 ;
               RECT 18.664 78.4835 18.736 78.5085 ;
               RECT 18.664 79.1605 18.736 79.1855 ;
               RECT 18.664 79.4545 18.736 79.4795 ;
               RECT 18.664 79.6835 18.736 79.7085 ;
               RECT 18.664 80.1315 18.736 80.1565 ;
               RECT 18.664 80.3605 18.736 80.3855 ;
               RECT 18.664 80.6545 18.736 80.6795 ;
               RECT 18.664 80.8835 18.736 80.9085 ;
               RECT 18.664 81.5605 18.736 81.5855 ;
               RECT 18.664 81.8545 18.736 81.8795 ;
               RECT 18.664 82.0835 18.736 82.1085 ;
               RECT 18.664 82.5315 18.736 82.5565 ;
               RECT 18.664 82.7605 18.736 82.7855 ;
               RECT 18.664 83.0545 18.736 83.0795 ;
               RECT 18.664 83.2835 18.736 83.3085 ;
               RECT 18.664 83.9605 18.736 83.9855 ;
               RECT 18.664 84.2545 18.736 84.2795 ;
               RECT 18.664 84.4835 18.736 84.5085 ;
               RECT 18.664 84.9315 18.736 84.9565 ;
               RECT 18.664 85.1605 18.736 85.1855 ;
               RECT 18.664 85.4545 18.736 85.4795 ;
               RECT 18.664 85.6835 18.736 85.7085 ;
               RECT 18.664 86.3605 18.736 86.3855 ;
               RECT 18.664 86.6545 18.736 86.6795 ;
               RECT 18.664 86.8835 18.736 86.9085 ;
               RECT 18.664 87.3315 18.736 87.3565 ;
               RECT 18.664 87.5605 18.736 87.5855 ;
               RECT 18.664 87.8545 18.736 87.8795 ;
               RECT 18.664 88.0835 18.736 88.1085 ;
               RECT 18.664 88.7605 18.736 88.7855 ;
               RECT 18.664 89.0545 18.736 89.0795 ;
               RECT 18.664 89.2835 18.736 89.3085 ;
               RECT 18.664 89.7315 18.736 89.7565 ;
               RECT 18.664 89.9605 18.736 89.9855 ;
               RECT 18.664 90.2545 18.736 90.2795 ;
               RECT 18.664 90.4835 18.736 90.5085 ;
               RECT 18.664 91.1605 18.736 91.1855 ;
               RECT 18.664 91.4545 18.736 91.4795 ;
               RECT 18.664 91.6835 18.736 91.7085 ;
               RECT 18.664 92.1315 18.736 92.1565 ;
               RECT 18.664 92.3605 18.736 92.3855 ;
               RECT 18.664 92.6545 18.736 92.6795 ;
               RECT 18.664 92.8835 18.736 92.9085 ;
               RECT 18.664 93.5605 18.736 93.5855 ;
               RECT 18.664 93.8545 18.736 93.8795 ;
               RECT 18.664 94.0835 18.736 94.1085 ;
               RECT 18.664 94.5315 18.736 94.5565 ;
               RECT 18.664 94.7605 18.736 94.7855 ;
               RECT 18.664 95.0545 18.736 95.0795 ;
               RECT 18.664 95.2835 18.736 95.3085 ;
               RECT 18.664 95.9605 18.736 95.9855 ;
               RECT 18.664 96.2545 18.736 96.2795 ;
               RECT 18.664 96.4835 18.736 96.5085 ;
               RECT 18.664 96.9315 18.736 96.9565 ;
               RECT 18.664 97.1605 18.736 97.1855 ;
               RECT 18.664 97.4545 18.736 97.4795 ;
               RECT 18.664 97.6835 18.736 97.7085 ;
               RECT 18.664 98.3605 18.736 98.3855 ;
               RECT 18.664 98.6545 18.736 98.6795 ;
               RECT 18.664 98.8835 18.736 98.9085 ;
               RECT 18.664 99.3315 18.736 99.3565 ;
               RECT 18.664 99.5605 18.736 99.5855 ;
               RECT 18.664 99.8545 18.736 99.8795 ;
               RECT 18.664 100.0835 18.736 100.1085 ;
               RECT 18.664 100.7605 18.736 100.7855 ;
               RECT 18.664 101.0545 18.736 101.0795 ;
               RECT 18.664 101.2835 18.736 101.3085 ;
               RECT 18.664 101.7315 18.736 101.7565 ;
               RECT 18.664 101.9605 18.736 101.9855 ;
               RECT 18.664 102.2545 18.736 102.2795 ;
               RECT 18.664 102.4835 18.736 102.5085 ;
               RECT 18.664 103.1605 18.736 103.1855 ;
               RECT 18.664 103.4545 18.736 103.4795 ;
               RECT 18.664 103.6835 18.736 103.7085 ;
               RECT 18.664 104.1315 18.736 104.1565 ;
               RECT 18.664 104.3605 18.736 104.3855 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.964 0.5695 19.036 104.5505 ;
               LAYER v4 ;
               RECT 18.964 0.7345 19.036 0.7595 ;
               RECT 18.964 0.9635 19.036 0.9885 ;
               RECT 18.964 1.4115 19.036 1.4365 ;
               RECT 18.964 1.6405 19.036 1.6655 ;
               RECT 18.964 1.9345 19.036 1.9595 ;
               RECT 18.964 2.1635 19.036 2.1885 ;
               RECT 18.964 2.6115 19.036 2.6365 ;
               RECT 18.964 2.8405 19.036 2.8655 ;
               RECT 18.964 3.1345 19.036 3.1595 ;
               RECT 18.964 3.3635 19.036 3.3885 ;
               RECT 18.964 3.8115 19.036 3.8365 ;
               RECT 18.964 4.0405 19.036 4.0655 ;
               RECT 18.964 4.3345 19.036 4.3595 ;
               RECT 18.964 4.5635 19.036 4.5885 ;
               RECT 18.964 5.0115 19.036 5.0365 ;
               RECT 18.964 5.2405 19.036 5.2655 ;
               RECT 18.964 5.5345 19.036 5.5595 ;
               RECT 18.964 5.7635 19.036 5.7885 ;
               RECT 18.964 6.2115 19.036 6.2365 ;
               RECT 18.964 6.4405 19.036 6.4655 ;
               RECT 18.964 6.7345 19.036 6.7595 ;
               RECT 18.964 6.9635 19.036 6.9885 ;
               RECT 18.964 7.4115 19.036 7.4365 ;
               RECT 18.964 7.6405 19.036 7.6655 ;
               RECT 18.964 7.9345 19.036 7.9595 ;
               RECT 18.964 8.1635 19.036 8.1885 ;
               RECT 18.964 8.6115 19.036 8.6365 ;
               RECT 18.964 8.8405 19.036 8.8655 ;
               RECT 18.964 9.1345 19.036 9.1595 ;
               RECT 18.964 9.3635 19.036 9.3885 ;
               RECT 18.964 9.8115 19.036 9.8365 ;
               RECT 18.964 10.0405 19.036 10.0655 ;
               RECT 18.964 10.3345 19.036 10.3595 ;
               RECT 18.964 10.5635 19.036 10.5885 ;
               RECT 18.964 11.0115 19.036 11.0365 ;
               RECT 18.964 11.2405 19.036 11.2655 ;
               RECT 18.964 11.5345 19.036 11.5595 ;
               RECT 18.964 11.7635 19.036 11.7885 ;
               RECT 18.964 12.2115 19.036 12.2365 ;
               RECT 18.964 12.4405 19.036 12.4655 ;
               RECT 18.964 12.7345 19.036 12.7595 ;
               RECT 18.964 12.9635 19.036 12.9885 ;
               RECT 18.964 13.4115 19.036 13.4365 ;
               RECT 18.964 13.6405 19.036 13.6655 ;
               RECT 18.964 13.9345 19.036 13.9595 ;
               RECT 18.964 14.1635 19.036 14.1885 ;
               RECT 18.964 14.6115 19.036 14.6365 ;
               RECT 18.964 14.8405 19.036 14.8655 ;
               RECT 18.964 15.1345 19.036 15.1595 ;
               RECT 18.964 15.3635 19.036 15.3885 ;
               RECT 18.964 15.8115 19.036 15.8365 ;
               RECT 18.964 16.0405 19.036 16.0655 ;
               RECT 18.964 16.3345 19.036 16.3595 ;
               RECT 18.964 16.5635 19.036 16.5885 ;
               RECT 18.964 17.0115 19.036 17.0365 ;
               RECT 18.964 17.2405 19.036 17.2655 ;
               RECT 18.964 17.5345 19.036 17.5595 ;
               RECT 18.964 17.7635 19.036 17.7885 ;
               RECT 18.964 18.2115 19.036 18.2365 ;
               RECT 18.964 18.4405 19.036 18.4655 ;
               RECT 18.964 18.7345 19.036 18.7595 ;
               RECT 18.964 18.9635 19.036 18.9885 ;
               RECT 18.964 19.4115 19.036 19.4365 ;
               RECT 18.964 19.6405 19.036 19.6655 ;
               RECT 18.964 19.9345 19.036 19.9595 ;
               RECT 18.964 20.1635 19.036 20.1885 ;
               RECT 18.964 20.6115 19.036 20.6365 ;
               RECT 18.964 20.8405 19.036 20.8655 ;
               RECT 18.964 21.1345 19.036 21.1595 ;
               RECT 18.964 21.3635 19.036 21.3885 ;
               RECT 18.964 21.8115 19.036 21.8365 ;
               RECT 18.964 22.0405 19.036 22.0655 ;
               RECT 18.964 22.3345 19.036 22.3595 ;
               RECT 18.964 22.5635 19.036 22.5885 ;
               RECT 18.964 23.0115 19.036 23.0365 ;
               RECT 18.964 23.2405 19.036 23.2655 ;
               RECT 18.964 23.5345 19.036 23.5595 ;
               RECT 18.964 23.7635 19.036 23.7885 ;
               RECT 18.964 24.2115 19.036 24.2365 ;
               RECT 18.964 24.4405 19.036 24.4655 ;
               RECT 18.964 24.7345 19.036 24.7595 ;
               RECT 18.964 24.9635 19.036 24.9885 ;
               RECT 18.964 25.4115 19.036 25.4365 ;
               RECT 18.964 25.6405 19.036 25.6655 ;
               RECT 18.964 25.9345 19.036 25.9595 ;
               RECT 18.964 26.1635 19.036 26.1885 ;
               RECT 18.964 26.6115 19.036 26.6365 ;
               RECT 18.964 26.8405 19.036 26.8655 ;
               RECT 18.964 27.1345 19.036 27.1595 ;
               RECT 18.964 27.3635 19.036 27.3885 ;
               RECT 18.964 27.8115 19.036 27.8365 ;
               RECT 18.964 28.0405 19.036 28.0655 ;
               RECT 18.964 28.3345 19.036 28.3595 ;
               RECT 18.964 28.5635 19.036 28.5885 ;
               RECT 18.964 29.0115 19.036 29.0365 ;
               RECT 18.964 29.2405 19.036 29.2655 ;
               RECT 18.964 29.5345 19.036 29.5595 ;
               RECT 18.964 29.7635 19.036 29.7885 ;
               RECT 18.964 30.2115 19.036 30.2365 ;
               RECT 18.964 30.4405 19.036 30.4655 ;
               RECT 18.964 30.7345 19.036 30.7595 ;
               RECT 18.964 30.9635 19.036 30.9885 ;
               RECT 18.964 31.4115 19.036 31.4365 ;
               RECT 18.964 31.6405 19.036 31.6655 ;
               RECT 18.964 31.9345 19.036 31.9595 ;
               RECT 18.964 32.1635 19.036 32.1885 ;
               RECT 18.964 32.6115 19.036 32.6365 ;
               RECT 18.964 32.8405 19.036 32.8655 ;
               RECT 18.964 33.1345 19.036 33.1595 ;
               RECT 18.964 33.3635 19.036 33.3885 ;
               RECT 18.964 33.8115 19.036 33.8365 ;
               RECT 18.964 34.0405 19.036 34.0655 ;
               RECT 18.964 34.3345 19.036 34.3595 ;
               RECT 18.964 34.5635 19.036 34.5885 ;
               RECT 18.964 35.0115 19.036 35.0365 ;
               RECT 18.964 35.2405 19.036 35.2655 ;
               RECT 18.964 35.5345 19.036 35.5595 ;
               RECT 18.964 35.7635 19.036 35.7885 ;
               RECT 18.964 36.2115 19.036 36.2365 ;
               RECT 18.964 36.4405 19.036 36.4655 ;
               RECT 18.964 36.7345 19.036 36.7595 ;
               RECT 18.964 36.9635 19.036 36.9885 ;
               RECT 18.964 37.4115 19.036 37.4365 ;
               RECT 18.964 37.6405 19.036 37.6655 ;
               RECT 18.964 37.9345 19.036 37.9595 ;
               RECT 18.964 38.1635 19.036 38.1885 ;
               RECT 18.964 38.6115 19.036 38.6365 ;
               RECT 18.964 38.8405 19.036 38.8655 ;
               RECT 18.964 39.1345 19.036 39.1595 ;
               RECT 18.964 39.3635 19.036 39.3885 ;
               RECT 18.964 39.8115 19.036 39.8365 ;
               RECT 18.964 40.0405 19.036 40.0655 ;
               RECT 18.964 40.3345 19.036 40.3595 ;
               RECT 18.964 40.5635 19.036 40.5885 ;
               RECT 18.964 41.0115 19.036 41.0365 ;
               RECT 18.964 41.2405 19.036 41.2655 ;
               RECT 18.964 41.5345 19.036 41.5595 ;
               RECT 18.964 41.7635 19.036 41.7885 ;
               RECT 18.964 42.2115 19.036 42.2365 ;
               RECT 18.964 42.4405 19.036 42.4655 ;
               RECT 18.964 42.7345 19.036 42.7595 ;
               RECT 18.964 42.9635 19.036 42.9885 ;
               RECT 18.964 43.4115 19.036 43.4365 ;
               RECT 18.964 43.6405 19.036 43.6655 ;
               RECT 18.964 43.9345 19.036 43.9595 ;
               RECT 18.964 44.1635 19.036 44.1885 ;
               RECT 18.964 44.6115 19.036 44.6365 ;
               RECT 18.964 44.8405 19.036 44.8655 ;
               RECT 18.964 45.1345 19.036 45.1595 ;
               RECT 18.964 45.3635 19.036 45.3885 ;
               RECT 18.964 45.8115 19.036 45.8365 ;
               RECT 18.964 46.0405 19.036 46.0655 ;
               RECT 18.964 46.3345 19.036 46.3595 ;
               RECT 18.964 46.5635 19.036 46.5885 ;
               RECT 18.964 47.0115 19.036 47.0365 ;
               RECT 18.964 47.2405 19.036 47.2655 ;
               RECT 18.964 47.5345 19.036 47.5595 ;
               RECT 18.964 47.7635 19.036 47.7885 ;
               RECT 18.964 48.2115 19.036 48.2365 ;
               RECT 18.964 48.4405 19.036 48.4655 ;
               RECT 18.964 49.1875 19.036 49.2125 ;
               RECT 18.964 49.6675 19.036 49.6925 ;
               RECT 18.964 50.1475 19.036 50.1725 ;
               RECT 18.964 50.6275 19.036 50.6525 ;
               RECT 18.964 51.1075 19.036 51.1325 ;
               RECT 18.964 51.5875 19.036 51.6125 ;
               RECT 18.964 52.0675 19.036 52.0925 ;
               RECT 18.964 52.5475 19.036 52.5725 ;
               RECT 18.964 53.0275 19.036 53.0525 ;
               RECT 18.964 53.5075 19.036 53.5325 ;
               RECT 18.964 53.9875 19.036 54.0125 ;
               RECT 18.964 54.4675 19.036 54.4925 ;
               RECT 18.964 54.9475 19.036 54.9725 ;
               RECT 18.964 55.4275 19.036 55.4525 ;
               RECT 18.964 55.9075 19.036 55.9325 ;
               RECT 18.964 56.6545 19.036 56.6795 ;
               RECT 18.964 56.8835 19.036 56.9085 ;
               RECT 18.964 57.3315 19.036 57.3565 ;
               RECT 18.964 57.5605 19.036 57.5855 ;
               RECT 18.964 57.8545 19.036 57.8795 ;
               RECT 18.964 58.0835 19.036 58.1085 ;
               RECT 18.964 58.5315 19.036 58.5565 ;
               RECT 18.964 58.7605 19.036 58.7855 ;
               RECT 18.964 59.0545 19.036 59.0795 ;
               RECT 18.964 59.2835 19.036 59.3085 ;
               RECT 18.964 59.7315 19.036 59.7565 ;
               RECT 18.964 59.9605 19.036 59.9855 ;
               RECT 18.964 60.2545 19.036 60.2795 ;
               RECT 18.964 60.4835 19.036 60.5085 ;
               RECT 18.964 60.9315 19.036 60.9565 ;
               RECT 18.964 61.1605 19.036 61.1855 ;
               RECT 18.964 61.4545 19.036 61.4795 ;
               RECT 18.964 61.6835 19.036 61.7085 ;
               RECT 18.964 62.1315 19.036 62.1565 ;
               RECT 18.964 62.3605 19.036 62.3855 ;
               RECT 18.964 62.6545 19.036 62.6795 ;
               RECT 18.964 62.8835 19.036 62.9085 ;
               RECT 18.964 63.3315 19.036 63.3565 ;
               RECT 18.964 63.5605 19.036 63.5855 ;
               RECT 18.964 63.8545 19.036 63.8795 ;
               RECT 18.964 64.0835 19.036 64.1085 ;
               RECT 18.964 64.5315 19.036 64.5565 ;
               RECT 18.964 64.7605 19.036 64.7855 ;
               RECT 18.964 65.0545 19.036 65.0795 ;
               RECT 18.964 65.2835 19.036 65.3085 ;
               RECT 18.964 65.7315 19.036 65.7565 ;
               RECT 18.964 65.9605 19.036 65.9855 ;
               RECT 18.964 66.2545 19.036 66.2795 ;
               RECT 18.964 66.4835 19.036 66.5085 ;
               RECT 18.964 66.9315 19.036 66.9565 ;
               RECT 18.964 67.1605 19.036 67.1855 ;
               RECT 18.964 67.4545 19.036 67.4795 ;
               RECT 18.964 67.6835 19.036 67.7085 ;
               RECT 18.964 68.1315 19.036 68.1565 ;
               RECT 18.964 68.3605 19.036 68.3855 ;
               RECT 18.964 68.6545 19.036 68.6795 ;
               RECT 18.964 68.8835 19.036 68.9085 ;
               RECT 18.964 69.3315 19.036 69.3565 ;
               RECT 18.964 69.5605 19.036 69.5855 ;
               RECT 18.964 69.8545 19.036 69.8795 ;
               RECT 18.964 70.0835 19.036 70.1085 ;
               RECT 18.964 70.5315 19.036 70.5565 ;
               RECT 18.964 70.7605 19.036 70.7855 ;
               RECT 18.964 71.0545 19.036 71.0795 ;
               RECT 18.964 71.2835 19.036 71.3085 ;
               RECT 18.964 71.7315 19.036 71.7565 ;
               RECT 18.964 71.9605 19.036 71.9855 ;
               RECT 18.964 72.2545 19.036 72.2795 ;
               RECT 18.964 72.4835 19.036 72.5085 ;
               RECT 18.964 72.9315 19.036 72.9565 ;
               RECT 18.964 73.1605 19.036 73.1855 ;
               RECT 18.964 73.4545 19.036 73.4795 ;
               RECT 18.964 73.6835 19.036 73.7085 ;
               RECT 18.964 74.1315 19.036 74.1565 ;
               RECT 18.964 74.3605 19.036 74.3855 ;
               RECT 18.964 74.6545 19.036 74.6795 ;
               RECT 18.964 74.8835 19.036 74.9085 ;
               RECT 18.964 75.3315 19.036 75.3565 ;
               RECT 18.964 75.5605 19.036 75.5855 ;
               RECT 18.964 75.8545 19.036 75.8795 ;
               RECT 18.964 76.0835 19.036 76.1085 ;
               RECT 18.964 76.5315 19.036 76.5565 ;
               RECT 18.964 76.7605 19.036 76.7855 ;
               RECT 18.964 77.0545 19.036 77.0795 ;
               RECT 18.964 77.2835 19.036 77.3085 ;
               RECT 18.964 77.7315 19.036 77.7565 ;
               RECT 18.964 77.9605 19.036 77.9855 ;
               RECT 18.964 78.2545 19.036 78.2795 ;
               RECT 18.964 78.4835 19.036 78.5085 ;
               RECT 18.964 78.9315 19.036 78.9565 ;
               RECT 18.964 79.1605 19.036 79.1855 ;
               RECT 18.964 79.4545 19.036 79.4795 ;
               RECT 18.964 79.6835 19.036 79.7085 ;
               RECT 18.964 80.1315 19.036 80.1565 ;
               RECT 18.964 80.3605 19.036 80.3855 ;
               RECT 18.964 80.6545 19.036 80.6795 ;
               RECT 18.964 80.8835 19.036 80.9085 ;
               RECT 18.964 81.3315 19.036 81.3565 ;
               RECT 18.964 81.5605 19.036 81.5855 ;
               RECT 18.964 81.8545 19.036 81.8795 ;
               RECT 18.964 82.0835 19.036 82.1085 ;
               RECT 18.964 82.5315 19.036 82.5565 ;
               RECT 18.964 82.7605 19.036 82.7855 ;
               RECT 18.964 83.0545 19.036 83.0795 ;
               RECT 18.964 83.2835 19.036 83.3085 ;
               RECT 18.964 83.7315 19.036 83.7565 ;
               RECT 18.964 83.9605 19.036 83.9855 ;
               RECT 18.964 84.2545 19.036 84.2795 ;
               RECT 18.964 84.4835 19.036 84.5085 ;
               RECT 18.964 84.9315 19.036 84.9565 ;
               RECT 18.964 85.1605 19.036 85.1855 ;
               RECT 18.964 85.4545 19.036 85.4795 ;
               RECT 18.964 85.6835 19.036 85.7085 ;
               RECT 18.964 86.1315 19.036 86.1565 ;
               RECT 18.964 86.3605 19.036 86.3855 ;
               RECT 18.964 86.6545 19.036 86.6795 ;
               RECT 18.964 86.8835 19.036 86.9085 ;
               RECT 18.964 87.3315 19.036 87.3565 ;
               RECT 18.964 87.5605 19.036 87.5855 ;
               RECT 18.964 87.8545 19.036 87.8795 ;
               RECT 18.964 88.0835 19.036 88.1085 ;
               RECT 18.964 88.5315 19.036 88.5565 ;
               RECT 18.964 88.7605 19.036 88.7855 ;
               RECT 18.964 89.0545 19.036 89.0795 ;
               RECT 18.964 89.2835 19.036 89.3085 ;
               RECT 18.964 89.7315 19.036 89.7565 ;
               RECT 18.964 89.9605 19.036 89.9855 ;
               RECT 18.964 90.2545 19.036 90.2795 ;
               RECT 18.964 90.4835 19.036 90.5085 ;
               RECT 18.964 90.9315 19.036 90.9565 ;
               RECT 18.964 91.1605 19.036 91.1855 ;
               RECT 18.964 91.4545 19.036 91.4795 ;
               RECT 18.964 91.6835 19.036 91.7085 ;
               RECT 18.964 92.1315 19.036 92.1565 ;
               RECT 18.964 92.3605 19.036 92.3855 ;
               RECT 18.964 92.6545 19.036 92.6795 ;
               RECT 18.964 92.8835 19.036 92.9085 ;
               RECT 18.964 93.3315 19.036 93.3565 ;
               RECT 18.964 93.5605 19.036 93.5855 ;
               RECT 18.964 93.8545 19.036 93.8795 ;
               RECT 18.964 94.0835 19.036 94.1085 ;
               RECT 18.964 94.5315 19.036 94.5565 ;
               RECT 18.964 94.7605 19.036 94.7855 ;
               RECT 18.964 95.0545 19.036 95.0795 ;
               RECT 18.964 95.2835 19.036 95.3085 ;
               RECT 18.964 95.7315 19.036 95.7565 ;
               RECT 18.964 95.9605 19.036 95.9855 ;
               RECT 18.964 96.2545 19.036 96.2795 ;
               RECT 18.964 96.4835 19.036 96.5085 ;
               RECT 18.964 96.9315 19.036 96.9565 ;
               RECT 18.964 97.1605 19.036 97.1855 ;
               RECT 18.964 97.4545 19.036 97.4795 ;
               RECT 18.964 97.6835 19.036 97.7085 ;
               RECT 18.964 98.1315 19.036 98.1565 ;
               RECT 18.964 98.3605 19.036 98.3855 ;
               RECT 18.964 98.6545 19.036 98.6795 ;
               RECT 18.964 98.8835 19.036 98.9085 ;
               RECT 18.964 99.3315 19.036 99.3565 ;
               RECT 18.964 99.5605 19.036 99.5855 ;
               RECT 18.964 99.8545 19.036 99.8795 ;
               RECT 18.964 100.0835 19.036 100.1085 ;
               RECT 18.964 100.5315 19.036 100.5565 ;
               RECT 18.964 100.7605 19.036 100.7855 ;
               RECT 18.964 101.0545 19.036 101.0795 ;
               RECT 18.964 101.2835 19.036 101.3085 ;
               RECT 18.964 101.7315 19.036 101.7565 ;
               RECT 18.964 101.9605 19.036 101.9855 ;
               RECT 18.964 102.2545 19.036 102.2795 ;
               RECT 18.964 102.4835 19.036 102.5085 ;
               RECT 18.964 102.9315 19.036 102.9565 ;
               RECT 18.964 103.1605 19.036 103.1855 ;
               RECT 18.964 103.4545 19.036 103.4795 ;
               RECT 18.964 103.6835 19.036 103.7085 ;
               RECT 18.964 104.1315 19.036 104.1565 ;
               RECT 18.964 104.3605 19.036 104.3855 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.31 48.6 19.35 56.52 ;
               LAYER v4 ;
               RECT 19.31 49.182 19.35 49.218 ;
               RECT 19.31 49.662 19.35 49.698 ;
               RECT 19.31 50.142 19.35 50.178 ;
               RECT 19.31 50.622 19.35 50.658 ;
               RECT 19.31 51.102 19.35 51.138 ;
               RECT 19.31 51.582 19.35 51.618 ;
               RECT 19.31 52.062 19.35 52.098 ;
               RECT 19.31 52.542 19.35 52.578 ;
               RECT 19.31 53.022 19.35 53.058 ;
               RECT 19.31 53.502 19.35 53.538 ;
               RECT 19.31 53.982 19.35 54.018 ;
               RECT 19.31 54.462 19.35 54.498 ;
               RECT 19.31 54.942 19.35 54.978 ;
               RECT 19.31 55.422 19.35 55.458 ;
               RECT 19.31 55.902 19.35 55.938 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.914 0.5695 19.966 104.5505 ;
               LAYER v4 ;
               RECT 19.914 0.729 19.966 0.765 ;
               RECT 19.914 0.958 19.966 0.994 ;
               RECT 19.914 1.406 19.966 1.442 ;
               RECT 19.914 1.929 19.966 1.965 ;
               RECT 19.914 2.158 19.966 2.194 ;
               RECT 19.914 2.606 19.966 2.642 ;
               RECT 19.914 3.129 19.966 3.165 ;
               RECT 19.914 3.358 19.966 3.394 ;
               RECT 19.914 3.806 19.966 3.842 ;
               RECT 19.914 4.329 19.966 4.365 ;
               RECT 19.914 4.558 19.966 4.594 ;
               RECT 19.914 5.006 19.966 5.042 ;
               RECT 19.914 5.529 19.966 5.565 ;
               RECT 19.914 5.758 19.966 5.794 ;
               RECT 19.914 6.206 19.966 6.242 ;
               RECT 19.914 6.729 19.966 6.765 ;
               RECT 19.914 6.958 19.966 6.994 ;
               RECT 19.914 7.406 19.966 7.442 ;
               RECT 19.914 7.929 19.966 7.965 ;
               RECT 19.914 8.158 19.966 8.194 ;
               RECT 19.914 8.606 19.966 8.642 ;
               RECT 19.914 9.129 19.966 9.165 ;
               RECT 19.914 9.358 19.966 9.394 ;
               RECT 19.914 9.806 19.966 9.842 ;
               RECT 19.914 10.329 19.966 10.365 ;
               RECT 19.914 10.558 19.966 10.594 ;
               RECT 19.914 11.006 19.966 11.042 ;
               RECT 19.914 11.529 19.966 11.565 ;
               RECT 19.914 11.758 19.966 11.794 ;
               RECT 19.914 12.206 19.966 12.242 ;
               RECT 19.914 12.729 19.966 12.765 ;
               RECT 19.914 12.958 19.966 12.994 ;
               RECT 19.914 13.406 19.966 13.442 ;
               RECT 19.914 13.929 19.966 13.965 ;
               RECT 19.914 14.158 19.966 14.194 ;
               RECT 19.914 14.606 19.966 14.642 ;
               RECT 19.914 15.129 19.966 15.165 ;
               RECT 19.914 15.358 19.966 15.394 ;
               RECT 19.914 15.806 19.966 15.842 ;
               RECT 19.914 16.329 19.966 16.365 ;
               RECT 19.914 16.558 19.966 16.594 ;
               RECT 19.914 17.006 19.966 17.042 ;
               RECT 19.914 17.529 19.966 17.565 ;
               RECT 19.914 17.758 19.966 17.794 ;
               RECT 19.914 18.206 19.966 18.242 ;
               RECT 19.914 18.729 19.966 18.765 ;
               RECT 19.914 18.958 19.966 18.994 ;
               RECT 19.914 19.406 19.966 19.442 ;
               RECT 19.914 19.929 19.966 19.965 ;
               RECT 19.914 20.158 19.966 20.194 ;
               RECT 19.914 20.606 19.966 20.642 ;
               RECT 19.914 21.129 19.966 21.165 ;
               RECT 19.914 21.358 19.966 21.394 ;
               RECT 19.914 21.806 19.966 21.842 ;
               RECT 19.914 22.329 19.966 22.365 ;
               RECT 19.914 22.558 19.966 22.594 ;
               RECT 19.914 23.006 19.966 23.042 ;
               RECT 19.914 23.529 19.966 23.565 ;
               RECT 19.914 23.758 19.966 23.794 ;
               RECT 19.914 24.206 19.966 24.242 ;
               RECT 19.914 24.729 19.966 24.765 ;
               RECT 19.914 24.958 19.966 24.994 ;
               RECT 19.914 25.406 19.966 25.442 ;
               RECT 19.914 25.929 19.966 25.965 ;
               RECT 19.914 26.158 19.966 26.194 ;
               RECT 19.914 26.606 19.966 26.642 ;
               RECT 19.914 27.129 19.966 27.165 ;
               RECT 19.914 27.358 19.966 27.394 ;
               RECT 19.914 27.806 19.966 27.842 ;
               RECT 19.914 28.329 19.966 28.365 ;
               RECT 19.914 28.558 19.966 28.594 ;
               RECT 19.914 29.006 19.966 29.042 ;
               RECT 19.914 29.529 19.966 29.565 ;
               RECT 19.914 29.758 19.966 29.794 ;
               RECT 19.914 30.206 19.966 30.242 ;
               RECT 19.914 30.729 19.966 30.765 ;
               RECT 19.914 30.958 19.966 30.994 ;
               RECT 19.914 31.406 19.966 31.442 ;
               RECT 19.914 31.929 19.966 31.965 ;
               RECT 19.914 32.158 19.966 32.194 ;
               RECT 19.914 32.606 19.966 32.642 ;
               RECT 19.914 33.129 19.966 33.165 ;
               RECT 19.914 33.358 19.966 33.394 ;
               RECT 19.914 33.806 19.966 33.842 ;
               RECT 19.914 34.329 19.966 34.365 ;
               RECT 19.914 34.558 19.966 34.594 ;
               RECT 19.914 35.006 19.966 35.042 ;
               RECT 19.914 35.529 19.966 35.565 ;
               RECT 19.914 35.758 19.966 35.794 ;
               RECT 19.914 36.206 19.966 36.242 ;
               RECT 19.914 36.729 19.966 36.765 ;
               RECT 19.914 36.958 19.966 36.994 ;
               RECT 19.914 37.406 19.966 37.442 ;
               RECT 19.914 37.929 19.966 37.965 ;
               RECT 19.914 38.158 19.966 38.194 ;
               RECT 19.914 38.606 19.966 38.642 ;
               RECT 19.914 39.129 19.966 39.165 ;
               RECT 19.914 39.358 19.966 39.394 ;
               RECT 19.914 39.806 19.966 39.842 ;
               RECT 19.914 40.329 19.966 40.365 ;
               RECT 19.914 40.558 19.966 40.594 ;
               RECT 19.914 41.006 19.966 41.042 ;
               RECT 19.914 41.529 19.966 41.565 ;
               RECT 19.914 41.758 19.966 41.794 ;
               RECT 19.914 42.206 19.966 42.242 ;
               RECT 19.914 42.729 19.966 42.765 ;
               RECT 19.914 42.958 19.966 42.994 ;
               RECT 19.914 43.406 19.966 43.442 ;
               RECT 19.914 43.929 19.966 43.965 ;
               RECT 19.914 44.158 19.966 44.194 ;
               RECT 19.914 44.606 19.966 44.642 ;
               RECT 19.914 45.129 19.966 45.165 ;
               RECT 19.914 45.358 19.966 45.394 ;
               RECT 19.914 45.806 19.966 45.842 ;
               RECT 19.914 46.329 19.966 46.365 ;
               RECT 19.914 46.558 19.966 46.594 ;
               RECT 19.914 47.006 19.966 47.042 ;
               RECT 19.914 47.529 19.966 47.565 ;
               RECT 19.914 47.758 19.966 47.794 ;
               RECT 19.914 48.206 19.966 48.242 ;
               RECT 19.914 49.182 19.966 49.218 ;
               RECT 19.914 49.662 19.966 49.698 ;
               RECT 19.914 50.142 19.966 50.178 ;
               RECT 19.914 50.622 19.966 50.658 ;
               RECT 19.914 51.1075 19.966 51.1325 ;
               RECT 19.914 51.582 19.966 51.618 ;
               RECT 19.914 52.062 19.966 52.098 ;
               RECT 19.914 52.542 19.966 52.578 ;
               RECT 19.914 53.022 19.966 53.058 ;
               RECT 19.914 53.502 19.966 53.538 ;
               RECT 19.914 53.982 19.966 54.018 ;
               RECT 19.914 54.462 19.966 54.498 ;
               RECT 19.914 54.942 19.966 54.978 ;
               RECT 19.914 55.422 19.966 55.458 ;
               RECT 19.914 55.902 19.966 55.938 ;
               RECT 19.914 56.649 19.966 56.685 ;
               RECT 19.914 56.878 19.966 56.914 ;
               RECT 19.914 57.326 19.966 57.362 ;
               RECT 19.914 57.849 19.966 57.885 ;
               RECT 19.914 58.078 19.966 58.114 ;
               RECT 19.914 58.526 19.966 58.562 ;
               RECT 19.914 59.049 19.966 59.085 ;
               RECT 19.914 59.278 19.966 59.314 ;
               RECT 19.914 59.726 19.966 59.762 ;
               RECT 19.914 60.249 19.966 60.285 ;
               RECT 19.914 60.478 19.966 60.514 ;
               RECT 19.914 60.926 19.966 60.962 ;
               RECT 19.914 61.449 19.966 61.485 ;
               RECT 19.914 61.678 19.966 61.714 ;
               RECT 19.914 62.126 19.966 62.162 ;
               RECT 19.914 62.649 19.966 62.685 ;
               RECT 19.914 62.878 19.966 62.914 ;
               RECT 19.914 63.326 19.966 63.362 ;
               RECT 19.914 63.849 19.966 63.885 ;
               RECT 19.914 64.078 19.966 64.114 ;
               RECT 19.914 64.526 19.966 64.562 ;
               RECT 19.914 65.049 19.966 65.085 ;
               RECT 19.914 65.278 19.966 65.314 ;
               RECT 19.914 65.726 19.966 65.762 ;
               RECT 19.914 66.249 19.966 66.285 ;
               RECT 19.914 66.478 19.966 66.514 ;
               RECT 19.914 66.926 19.966 66.962 ;
               RECT 19.914 67.449 19.966 67.485 ;
               RECT 19.914 67.678 19.966 67.714 ;
               RECT 19.914 68.126 19.966 68.162 ;
               RECT 19.914 68.649 19.966 68.685 ;
               RECT 19.914 68.878 19.966 68.914 ;
               RECT 19.914 69.326 19.966 69.362 ;
               RECT 19.914 69.849 19.966 69.885 ;
               RECT 19.914 70.078 19.966 70.114 ;
               RECT 19.914 70.526 19.966 70.562 ;
               RECT 19.914 71.049 19.966 71.085 ;
               RECT 19.914 71.278 19.966 71.314 ;
               RECT 19.914 71.726 19.966 71.762 ;
               RECT 19.914 72.249 19.966 72.285 ;
               RECT 19.914 72.478 19.966 72.514 ;
               RECT 19.914 72.926 19.966 72.962 ;
               RECT 19.914 73.449 19.966 73.485 ;
               RECT 19.914 73.678 19.966 73.714 ;
               RECT 19.914 74.126 19.966 74.162 ;
               RECT 19.914 74.649 19.966 74.685 ;
               RECT 19.914 74.878 19.966 74.914 ;
               RECT 19.914 75.326 19.966 75.362 ;
               RECT 19.914 75.849 19.966 75.885 ;
               RECT 19.914 76.078 19.966 76.114 ;
               RECT 19.914 76.526 19.966 76.562 ;
               RECT 19.914 77.049 19.966 77.085 ;
               RECT 19.914 77.278 19.966 77.314 ;
               RECT 19.914 77.726 19.966 77.762 ;
               RECT 19.914 78.249 19.966 78.285 ;
               RECT 19.914 78.478 19.966 78.514 ;
               RECT 19.914 78.926 19.966 78.962 ;
               RECT 19.914 79.449 19.966 79.485 ;
               RECT 19.914 79.678 19.966 79.714 ;
               RECT 19.914 80.126 19.966 80.162 ;
               RECT 19.914 80.649 19.966 80.685 ;
               RECT 19.914 80.878 19.966 80.914 ;
               RECT 19.914 81.326 19.966 81.362 ;
               RECT 19.914 81.849 19.966 81.885 ;
               RECT 19.914 82.078 19.966 82.114 ;
               RECT 19.914 82.526 19.966 82.562 ;
               RECT 19.914 83.049 19.966 83.085 ;
               RECT 19.914 83.278 19.966 83.314 ;
               RECT 19.914 83.726 19.966 83.762 ;
               RECT 19.914 84.249 19.966 84.285 ;
               RECT 19.914 84.478 19.966 84.514 ;
               RECT 19.914 84.926 19.966 84.962 ;
               RECT 19.914 85.449 19.966 85.485 ;
               RECT 19.914 85.678 19.966 85.714 ;
               RECT 19.914 86.126 19.966 86.162 ;
               RECT 19.914 86.649 19.966 86.685 ;
               RECT 19.914 86.878 19.966 86.914 ;
               RECT 19.914 87.326 19.966 87.362 ;
               RECT 19.914 87.849 19.966 87.885 ;
               RECT 19.914 88.078 19.966 88.114 ;
               RECT 19.914 88.526 19.966 88.562 ;
               RECT 19.914 89.049 19.966 89.085 ;
               RECT 19.914 89.278 19.966 89.314 ;
               RECT 19.914 89.726 19.966 89.762 ;
               RECT 19.914 90.249 19.966 90.285 ;
               RECT 19.914 90.478 19.966 90.514 ;
               RECT 19.914 90.926 19.966 90.962 ;
               RECT 19.914 91.449 19.966 91.485 ;
               RECT 19.914 91.678 19.966 91.714 ;
               RECT 19.914 92.126 19.966 92.162 ;
               RECT 19.914 92.649 19.966 92.685 ;
               RECT 19.914 92.878 19.966 92.914 ;
               RECT 19.914 93.326 19.966 93.362 ;
               RECT 19.914 93.849 19.966 93.885 ;
               RECT 19.914 94.078 19.966 94.114 ;
               RECT 19.914 94.526 19.966 94.562 ;
               RECT 19.914 95.049 19.966 95.085 ;
               RECT 19.914 95.278 19.966 95.314 ;
               RECT 19.914 95.726 19.966 95.762 ;
               RECT 19.914 96.249 19.966 96.285 ;
               RECT 19.914 96.478 19.966 96.514 ;
               RECT 19.914 96.926 19.966 96.962 ;
               RECT 19.914 97.449 19.966 97.485 ;
               RECT 19.914 97.678 19.966 97.714 ;
               RECT 19.914 98.126 19.966 98.162 ;
               RECT 19.914 98.649 19.966 98.685 ;
               RECT 19.914 98.878 19.966 98.914 ;
               RECT 19.914 99.326 19.966 99.362 ;
               RECT 19.914 99.849 19.966 99.885 ;
               RECT 19.914 100.078 19.966 100.114 ;
               RECT 19.914 100.526 19.966 100.562 ;
               RECT 19.914 101.049 19.966 101.085 ;
               RECT 19.914 101.278 19.966 101.314 ;
               RECT 19.914 101.726 19.966 101.762 ;
               RECT 19.914 102.249 19.966 102.285 ;
               RECT 19.914 102.478 19.966 102.514 ;
               RECT 19.914 102.926 19.966 102.962 ;
               RECT 19.914 103.449 19.966 103.485 ;
               RECT 19.914 103.678 19.966 103.714 ;
               RECT 19.914 104.126 19.966 104.162 ;
          END
          PORT
               LAYER m5 ;
               RECT 2.254 49.7505 2.306 55.3695 ;
               LAYER v4 ;
               RECT 2.254 49.782 2.306 49.818 ;
               RECT 2.254 50.262 2.306 50.298 ;
               RECT 2.254 50.502 2.306 50.538 ;
               RECT 2.254 50.982 2.306 51.018 ;
               RECT 2.254 51.102 2.306 51.138 ;
               RECT 2.254 51.582 2.306 51.618 ;
               RECT 2.254 52.062 2.306 52.098 ;
               RECT 2.254 52.182 2.306 52.218 ;
               RECT 2.254 52.542 2.306 52.578 ;
               RECT 2.254 52.662 2.306 52.698 ;
               RECT 2.254 52.902 2.306 52.938 ;
               RECT 2.254 53.022 2.306 53.058 ;
               RECT 2.254 53.502 2.306 53.538 ;
               RECT 2.254 53.982 2.306 54.018 ;
               RECT 2.254 54.102 2.306 54.138 ;
               RECT 2.254 54.582 2.306 54.618 ;
               RECT 2.254 54.822 2.306 54.858 ;
               RECT 2.254 55.302 2.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 2.574 0.6 2.626 104.52 ;
               LAYER v4 ;
               RECT 2.574 49.542 2.626 49.578 ;
               RECT 2.574 49.782 2.626 49.818 ;
               RECT 2.574 50.262 2.626 50.298 ;
               RECT 2.574 50.502 2.626 50.538 ;
               RECT 2.574 50.982 2.626 51.018 ;
               RECT 2.574 51.102 2.626 51.138 ;
               RECT 2.574 51.582 2.626 51.618 ;
               RECT 2.574 52.062 2.626 52.098 ;
               RECT 2.574 52.182 2.626 52.218 ;
               RECT 2.574 52.542 2.626 52.578 ;
               RECT 2.574 52.662 2.626 52.698 ;
               RECT 2.574 52.902 2.626 52.938 ;
               RECT 2.574 53.502 2.626 53.538 ;
               RECT 2.574 53.982 2.626 54.018 ;
               RECT 2.574 54.102 2.626 54.138 ;
               RECT 2.574 54.582 2.626 54.618 ;
               RECT 2.574 54.822 2.626 54.858 ;
               RECT 2.574 55.302 2.626 55.338 ;
               RECT 2.574 55.542 2.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 20.074 0.6 20.126 104.52 ;
               LAYER v4 ;
               RECT 20.074 0.729 20.126 0.765 ;
               RECT 20.074 0.958 20.126 0.994 ;
               RECT 20.074 1.406 20.126 1.442 ;
               RECT 20.074 1.635 20.126 1.671 ;
               RECT 20.074 1.929 20.126 1.965 ;
               RECT 20.074 2.158 20.126 2.194 ;
               RECT 20.074 2.606 20.126 2.642 ;
               RECT 20.074 2.835 20.126 2.871 ;
               RECT 20.074 3.129 20.126 3.165 ;
               RECT 20.074 3.358 20.126 3.394 ;
               RECT 20.074 3.806 20.126 3.842 ;
               RECT 20.074 4.035 20.126 4.071 ;
               RECT 20.074 4.329 20.126 4.365 ;
               RECT 20.074 4.558 20.126 4.594 ;
               RECT 20.074 5.006 20.126 5.042 ;
               RECT 20.074 5.235 20.126 5.271 ;
               RECT 20.074 5.529 20.126 5.565 ;
               RECT 20.074 5.758 20.126 5.794 ;
               RECT 20.074 6.206 20.126 6.242 ;
               RECT 20.074 6.435 20.126 6.471 ;
               RECT 20.074 6.729 20.126 6.765 ;
               RECT 20.074 6.958 20.126 6.994 ;
               RECT 20.074 7.406 20.126 7.442 ;
               RECT 20.074 7.635 20.126 7.671 ;
               RECT 20.074 7.929 20.126 7.965 ;
               RECT 20.074 8.158 20.126 8.194 ;
               RECT 20.074 8.606 20.126 8.642 ;
               RECT 20.074 8.835 20.126 8.871 ;
               RECT 20.074 9.129 20.126 9.165 ;
               RECT 20.074 9.358 20.126 9.394 ;
               RECT 20.074 9.806 20.126 9.842 ;
               RECT 20.074 10.035 20.126 10.071 ;
               RECT 20.074 10.329 20.126 10.365 ;
               RECT 20.074 10.558 20.126 10.594 ;
               RECT 20.074 11.006 20.126 11.042 ;
               RECT 20.074 11.235 20.126 11.271 ;
               RECT 20.074 11.529 20.126 11.565 ;
               RECT 20.074 11.758 20.126 11.794 ;
               RECT 20.074 12.206 20.126 12.242 ;
               RECT 20.074 12.435 20.126 12.471 ;
               RECT 20.074 12.729 20.126 12.765 ;
               RECT 20.074 12.958 20.126 12.994 ;
               RECT 20.074 13.406 20.126 13.442 ;
               RECT 20.074 13.635 20.126 13.671 ;
               RECT 20.074 13.929 20.126 13.965 ;
               RECT 20.074 14.158 20.126 14.194 ;
               RECT 20.074 14.606 20.126 14.642 ;
               RECT 20.074 14.835 20.126 14.871 ;
               RECT 20.074 15.129 20.126 15.165 ;
               RECT 20.074 15.358 20.126 15.394 ;
               RECT 20.074 15.806 20.126 15.842 ;
               RECT 20.074 16.035 20.126 16.071 ;
               RECT 20.074 16.329 20.126 16.365 ;
               RECT 20.074 16.558 20.126 16.594 ;
               RECT 20.074 17.006 20.126 17.042 ;
               RECT 20.074 17.235 20.126 17.271 ;
               RECT 20.074 17.529 20.126 17.565 ;
               RECT 20.074 17.758 20.126 17.794 ;
               RECT 20.074 18.206 20.126 18.242 ;
               RECT 20.074 18.435 20.126 18.471 ;
               RECT 20.074 18.729 20.126 18.765 ;
               RECT 20.074 18.958 20.126 18.994 ;
               RECT 20.074 19.406 20.126 19.442 ;
               RECT 20.074 19.635 20.126 19.671 ;
               RECT 20.074 19.929 20.126 19.965 ;
               RECT 20.074 20.158 20.126 20.194 ;
               RECT 20.074 20.606 20.126 20.642 ;
               RECT 20.074 20.835 20.126 20.871 ;
               RECT 20.074 21.129 20.126 21.165 ;
               RECT 20.074 21.358 20.126 21.394 ;
               RECT 20.074 21.806 20.126 21.842 ;
               RECT 20.074 22.035 20.126 22.071 ;
               RECT 20.074 22.329 20.126 22.365 ;
               RECT 20.074 22.558 20.126 22.594 ;
               RECT 20.074 23.006 20.126 23.042 ;
               RECT 20.074 23.235 20.126 23.271 ;
               RECT 20.074 23.529 20.126 23.565 ;
               RECT 20.074 23.758 20.126 23.794 ;
               RECT 20.074 24.206 20.126 24.242 ;
               RECT 20.074 24.435 20.126 24.471 ;
               RECT 20.074 24.729 20.126 24.765 ;
               RECT 20.074 24.958 20.126 24.994 ;
               RECT 20.074 25.406 20.126 25.442 ;
               RECT 20.074 25.635 20.126 25.671 ;
               RECT 20.074 25.929 20.126 25.965 ;
               RECT 20.074 26.158 20.126 26.194 ;
               RECT 20.074 26.606 20.126 26.642 ;
               RECT 20.074 26.835 20.126 26.871 ;
               RECT 20.074 27.129 20.126 27.165 ;
               RECT 20.074 27.358 20.126 27.394 ;
               RECT 20.074 27.806 20.126 27.842 ;
               RECT 20.074 28.035 20.126 28.071 ;
               RECT 20.074 28.329 20.126 28.365 ;
               RECT 20.074 28.558 20.126 28.594 ;
               RECT 20.074 29.006 20.126 29.042 ;
               RECT 20.074 29.235 20.126 29.271 ;
               RECT 20.074 29.529 20.126 29.565 ;
               RECT 20.074 29.758 20.126 29.794 ;
               RECT 20.074 30.206 20.126 30.242 ;
               RECT 20.074 30.435 20.126 30.471 ;
               RECT 20.074 30.729 20.126 30.765 ;
               RECT 20.074 30.958 20.126 30.994 ;
               RECT 20.074 31.406 20.126 31.442 ;
               RECT 20.074 31.635 20.126 31.671 ;
               RECT 20.074 31.929 20.126 31.965 ;
               RECT 20.074 32.158 20.126 32.194 ;
               RECT 20.074 32.606 20.126 32.642 ;
               RECT 20.074 32.835 20.126 32.871 ;
               RECT 20.074 33.129 20.126 33.165 ;
               RECT 20.074 33.358 20.126 33.394 ;
               RECT 20.074 33.806 20.126 33.842 ;
               RECT 20.074 34.035 20.126 34.071 ;
               RECT 20.074 34.329 20.126 34.365 ;
               RECT 20.074 34.558 20.126 34.594 ;
               RECT 20.074 35.006 20.126 35.042 ;
               RECT 20.074 35.235 20.126 35.271 ;
               RECT 20.074 35.529 20.126 35.565 ;
               RECT 20.074 35.758 20.126 35.794 ;
               RECT 20.074 36.206 20.126 36.242 ;
               RECT 20.074 36.435 20.126 36.471 ;
               RECT 20.074 36.729 20.126 36.765 ;
               RECT 20.074 36.958 20.126 36.994 ;
               RECT 20.074 37.406 20.126 37.442 ;
               RECT 20.074 37.635 20.126 37.671 ;
               RECT 20.074 37.929 20.126 37.965 ;
               RECT 20.074 38.158 20.126 38.194 ;
               RECT 20.074 38.606 20.126 38.642 ;
               RECT 20.074 38.835 20.126 38.871 ;
               RECT 20.074 39.129 20.126 39.165 ;
               RECT 20.074 39.358 20.126 39.394 ;
               RECT 20.074 39.806 20.126 39.842 ;
               RECT 20.074 40.035 20.126 40.071 ;
               RECT 20.074 40.329 20.126 40.365 ;
               RECT 20.074 40.558 20.126 40.594 ;
               RECT 20.074 41.006 20.126 41.042 ;
               RECT 20.074 41.235 20.126 41.271 ;
               RECT 20.074 41.529 20.126 41.565 ;
               RECT 20.074 41.758 20.126 41.794 ;
               RECT 20.074 42.206 20.126 42.242 ;
               RECT 20.074 42.435 20.126 42.471 ;
               RECT 20.074 42.729 20.126 42.765 ;
               RECT 20.074 42.958 20.126 42.994 ;
               RECT 20.074 43.406 20.126 43.442 ;
               RECT 20.074 43.635 20.126 43.671 ;
               RECT 20.074 43.929 20.126 43.965 ;
               RECT 20.074 44.158 20.126 44.194 ;
               RECT 20.074 44.606 20.126 44.642 ;
               RECT 20.074 44.835 20.126 44.871 ;
               RECT 20.074 45.129 20.126 45.165 ;
               RECT 20.074 45.358 20.126 45.394 ;
               RECT 20.074 45.806 20.126 45.842 ;
               RECT 20.074 46.035 20.126 46.071 ;
               RECT 20.074 46.329 20.126 46.365 ;
               RECT 20.074 46.558 20.126 46.594 ;
               RECT 20.074 47.006 20.126 47.042 ;
               RECT 20.074 47.235 20.126 47.271 ;
               RECT 20.074 47.529 20.126 47.565 ;
               RECT 20.074 47.758 20.126 47.794 ;
               RECT 20.074 48.206 20.126 48.242 ;
               RECT 20.074 48.435 20.126 48.471 ;
               RECT 20.074 49.182 20.126 49.218 ;
               RECT 20.074 49.662 20.126 49.698 ;
               RECT 20.074 50.142 20.126 50.178 ;
               RECT 20.074 50.622 20.126 50.658 ;
               RECT 20.074 51.102 20.126 51.138 ;
               RECT 20.074 51.582 20.126 51.618 ;
               RECT 20.074 52.062 20.126 52.098 ;
               RECT 20.074 52.542 20.126 52.578 ;
               RECT 20.074 53.0275 20.126 53.0525 ;
               RECT 20.074 53.502 20.126 53.538 ;
               RECT 20.074 53.982 20.126 54.018 ;
               RECT 20.074 54.462 20.126 54.498 ;
               RECT 20.074 54.9475 20.126 54.9725 ;
               RECT 20.074 55.422 20.126 55.458 ;
               RECT 20.074 55.902 20.126 55.938 ;
               RECT 20.074 56.649 20.126 56.685 ;
               RECT 20.074 56.878 20.126 56.914 ;
               RECT 20.074 57.326 20.126 57.362 ;
               RECT 20.074 57.555 20.126 57.591 ;
               RECT 20.074 57.849 20.126 57.885 ;
               RECT 20.074 58.078 20.126 58.114 ;
               RECT 20.074 58.526 20.126 58.562 ;
               RECT 20.074 58.755 20.126 58.791 ;
               RECT 20.074 59.049 20.126 59.085 ;
               RECT 20.074 59.278 20.126 59.314 ;
               RECT 20.074 59.726 20.126 59.762 ;
               RECT 20.074 59.955 20.126 59.991 ;
               RECT 20.074 60.249 20.126 60.285 ;
               RECT 20.074 60.478 20.126 60.514 ;
               RECT 20.074 60.926 20.126 60.962 ;
               RECT 20.074 61.155 20.126 61.191 ;
               RECT 20.074 61.449 20.126 61.485 ;
               RECT 20.074 61.678 20.126 61.714 ;
               RECT 20.074 62.126 20.126 62.162 ;
               RECT 20.074 62.355 20.126 62.391 ;
               RECT 20.074 62.649 20.126 62.685 ;
               RECT 20.074 62.878 20.126 62.914 ;
               RECT 20.074 63.326 20.126 63.362 ;
               RECT 20.074 63.555 20.126 63.591 ;
               RECT 20.074 63.849 20.126 63.885 ;
               RECT 20.074 64.078 20.126 64.114 ;
               RECT 20.074 64.526 20.126 64.562 ;
               RECT 20.074 64.755 20.126 64.791 ;
               RECT 20.074 65.049 20.126 65.085 ;
               RECT 20.074 65.278 20.126 65.314 ;
               RECT 20.074 65.726 20.126 65.762 ;
               RECT 20.074 65.955 20.126 65.991 ;
               RECT 20.074 66.249 20.126 66.285 ;
               RECT 20.074 66.478 20.126 66.514 ;
               RECT 20.074 66.926 20.126 66.962 ;
               RECT 20.074 67.155 20.126 67.191 ;
               RECT 20.074 67.449 20.126 67.485 ;
               RECT 20.074 67.678 20.126 67.714 ;
               RECT 20.074 68.126 20.126 68.162 ;
               RECT 20.074 68.355 20.126 68.391 ;
               RECT 20.074 68.649 20.126 68.685 ;
               RECT 20.074 68.878 20.126 68.914 ;
               RECT 20.074 69.326 20.126 69.362 ;
               RECT 20.074 69.555 20.126 69.591 ;
               RECT 20.074 69.849 20.126 69.885 ;
               RECT 20.074 70.078 20.126 70.114 ;
               RECT 20.074 70.526 20.126 70.562 ;
               RECT 20.074 70.755 20.126 70.791 ;
               RECT 20.074 71.049 20.126 71.085 ;
               RECT 20.074 71.278 20.126 71.314 ;
               RECT 20.074 71.726 20.126 71.762 ;
               RECT 20.074 71.955 20.126 71.991 ;
               RECT 20.074 72.249 20.126 72.285 ;
               RECT 20.074 72.478 20.126 72.514 ;
               RECT 20.074 72.926 20.126 72.962 ;
               RECT 20.074 73.155 20.126 73.191 ;
               RECT 20.074 73.449 20.126 73.485 ;
               RECT 20.074 73.678 20.126 73.714 ;
               RECT 20.074 74.126 20.126 74.162 ;
               RECT 20.074 74.355 20.126 74.391 ;
               RECT 20.074 74.649 20.126 74.685 ;
               RECT 20.074 74.878 20.126 74.914 ;
               RECT 20.074 75.326 20.126 75.362 ;
               RECT 20.074 75.555 20.126 75.591 ;
               RECT 20.074 75.849 20.126 75.885 ;
               RECT 20.074 76.078 20.126 76.114 ;
               RECT 20.074 76.526 20.126 76.562 ;
               RECT 20.074 76.755 20.126 76.791 ;
               RECT 20.074 77.049 20.126 77.085 ;
               RECT 20.074 77.278 20.126 77.314 ;
               RECT 20.074 77.726 20.126 77.762 ;
               RECT 20.074 77.955 20.126 77.991 ;
               RECT 20.074 78.249 20.126 78.285 ;
               RECT 20.074 78.478 20.126 78.514 ;
               RECT 20.074 78.926 20.126 78.962 ;
               RECT 20.074 79.155 20.126 79.191 ;
               RECT 20.074 79.449 20.126 79.485 ;
               RECT 20.074 79.678 20.126 79.714 ;
               RECT 20.074 80.126 20.126 80.162 ;
               RECT 20.074 80.355 20.126 80.391 ;
               RECT 20.074 80.649 20.126 80.685 ;
               RECT 20.074 80.878 20.126 80.914 ;
               RECT 20.074 81.326 20.126 81.362 ;
               RECT 20.074 81.555 20.126 81.591 ;
               RECT 20.074 81.849 20.126 81.885 ;
               RECT 20.074 82.078 20.126 82.114 ;
               RECT 20.074 82.526 20.126 82.562 ;
               RECT 20.074 82.755 20.126 82.791 ;
               RECT 20.074 83.049 20.126 83.085 ;
               RECT 20.074 83.278 20.126 83.314 ;
               RECT 20.074 83.726 20.126 83.762 ;
               RECT 20.074 83.955 20.126 83.991 ;
               RECT 20.074 84.249 20.126 84.285 ;
               RECT 20.074 84.478 20.126 84.514 ;
               RECT 20.074 84.926 20.126 84.962 ;
               RECT 20.074 85.155 20.126 85.191 ;
               RECT 20.074 85.449 20.126 85.485 ;
               RECT 20.074 85.678 20.126 85.714 ;
               RECT 20.074 86.126 20.126 86.162 ;
               RECT 20.074 86.355 20.126 86.391 ;
               RECT 20.074 86.649 20.126 86.685 ;
               RECT 20.074 86.878 20.126 86.914 ;
               RECT 20.074 87.326 20.126 87.362 ;
               RECT 20.074 87.555 20.126 87.591 ;
               RECT 20.074 87.849 20.126 87.885 ;
               RECT 20.074 88.078 20.126 88.114 ;
               RECT 20.074 88.526 20.126 88.562 ;
               RECT 20.074 88.755 20.126 88.791 ;
               RECT 20.074 89.049 20.126 89.085 ;
               RECT 20.074 89.278 20.126 89.314 ;
               RECT 20.074 89.726 20.126 89.762 ;
               RECT 20.074 89.955 20.126 89.991 ;
               RECT 20.074 90.249 20.126 90.285 ;
               RECT 20.074 90.478 20.126 90.514 ;
               RECT 20.074 90.926 20.126 90.962 ;
               RECT 20.074 91.155 20.126 91.191 ;
               RECT 20.074 91.449 20.126 91.485 ;
               RECT 20.074 91.678 20.126 91.714 ;
               RECT 20.074 92.126 20.126 92.162 ;
               RECT 20.074 92.355 20.126 92.391 ;
               RECT 20.074 92.649 20.126 92.685 ;
               RECT 20.074 92.878 20.126 92.914 ;
               RECT 20.074 93.326 20.126 93.362 ;
               RECT 20.074 93.555 20.126 93.591 ;
               RECT 20.074 93.849 20.126 93.885 ;
               RECT 20.074 94.078 20.126 94.114 ;
               RECT 20.074 94.526 20.126 94.562 ;
               RECT 20.074 94.755 20.126 94.791 ;
               RECT 20.074 95.049 20.126 95.085 ;
               RECT 20.074 95.278 20.126 95.314 ;
               RECT 20.074 95.726 20.126 95.762 ;
               RECT 20.074 95.955 20.126 95.991 ;
               RECT 20.074 96.249 20.126 96.285 ;
               RECT 20.074 96.478 20.126 96.514 ;
               RECT 20.074 96.926 20.126 96.962 ;
               RECT 20.074 97.155 20.126 97.191 ;
               RECT 20.074 97.449 20.126 97.485 ;
               RECT 20.074 97.678 20.126 97.714 ;
               RECT 20.074 98.126 20.126 98.162 ;
               RECT 20.074 98.355 20.126 98.391 ;
               RECT 20.074 98.649 20.126 98.685 ;
               RECT 20.074 98.878 20.126 98.914 ;
               RECT 20.074 99.326 20.126 99.362 ;
               RECT 20.074 99.555 20.126 99.591 ;
               RECT 20.074 99.849 20.126 99.885 ;
               RECT 20.074 100.078 20.126 100.114 ;
               RECT 20.074 100.526 20.126 100.562 ;
               RECT 20.074 100.755 20.126 100.791 ;
               RECT 20.074 101.049 20.126 101.085 ;
               RECT 20.074 101.278 20.126 101.314 ;
               RECT 20.074 101.726 20.126 101.762 ;
               RECT 20.074 101.955 20.126 101.991 ;
               RECT 20.074 102.249 20.126 102.285 ;
               RECT 20.074 102.478 20.126 102.514 ;
               RECT 20.074 102.926 20.126 102.962 ;
               RECT 20.074 103.155 20.126 103.191 ;
               RECT 20.074 103.449 20.126 103.485 ;
               RECT 20.074 103.678 20.126 103.714 ;
               RECT 20.074 104.126 20.126 104.162 ;
               RECT 20.074 104.355 20.126 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 20.47 0.5695 20.522 49.6595 ;
               LAYER v4 ;
               RECT 20.47 0.729 20.522 0.765 ;
               RECT 20.47 0.958 20.522 0.994 ;
               RECT 20.47 1.635 20.522 1.671 ;
               RECT 20.47 1.929 20.522 1.965 ;
               RECT 20.47 2.158 20.522 2.194 ;
               RECT 20.47 2.835 20.522 2.871 ;
               RECT 20.47 3.129 20.522 3.165 ;
               RECT 20.47 3.358 20.522 3.394 ;
               RECT 20.47 4.035 20.522 4.071 ;
               RECT 20.47 4.329 20.522 4.365 ;
               RECT 20.47 4.558 20.522 4.594 ;
               RECT 20.47 5.235 20.522 5.271 ;
               RECT 20.47 5.529 20.522 5.565 ;
               RECT 20.47 5.758 20.522 5.794 ;
               RECT 20.47 6.435 20.522 6.471 ;
               RECT 20.47 6.729 20.522 6.765 ;
               RECT 20.47 6.958 20.522 6.994 ;
               RECT 20.47 7.635 20.522 7.671 ;
               RECT 20.47 7.929 20.522 7.965 ;
               RECT 20.47 8.158 20.522 8.194 ;
               RECT 20.47 8.835 20.522 8.871 ;
               RECT 20.47 9.129 20.522 9.165 ;
               RECT 20.47 9.358 20.522 9.394 ;
               RECT 20.47 10.035 20.522 10.071 ;
               RECT 20.47 10.329 20.522 10.365 ;
               RECT 20.47 10.558 20.522 10.594 ;
               RECT 20.47 11.235 20.522 11.271 ;
               RECT 20.47 11.529 20.522 11.565 ;
               RECT 20.47 11.758 20.522 11.794 ;
               RECT 20.47 12.435 20.522 12.471 ;
               RECT 20.47 12.729 20.522 12.765 ;
               RECT 20.47 12.958 20.522 12.994 ;
               RECT 20.47 13.635 20.522 13.671 ;
               RECT 20.47 13.929 20.522 13.965 ;
               RECT 20.47 14.158 20.522 14.194 ;
               RECT 20.47 14.835 20.522 14.871 ;
               RECT 20.47 15.129 20.522 15.165 ;
               RECT 20.47 15.358 20.522 15.394 ;
               RECT 20.47 16.035 20.522 16.071 ;
               RECT 20.47 16.329 20.522 16.365 ;
               RECT 20.47 16.558 20.522 16.594 ;
               RECT 20.47 17.235 20.522 17.271 ;
               RECT 20.47 17.529 20.522 17.565 ;
               RECT 20.47 17.758 20.522 17.794 ;
               RECT 20.47 18.435 20.522 18.471 ;
               RECT 20.47 18.729 20.522 18.765 ;
               RECT 20.47 18.958 20.522 18.994 ;
               RECT 20.47 19.635 20.522 19.671 ;
               RECT 20.47 19.929 20.522 19.965 ;
               RECT 20.47 20.158 20.522 20.194 ;
               RECT 20.47 20.835 20.522 20.871 ;
               RECT 20.47 21.129 20.522 21.165 ;
               RECT 20.47 21.358 20.522 21.394 ;
               RECT 20.47 22.035 20.522 22.071 ;
               RECT 20.47 22.329 20.522 22.365 ;
               RECT 20.47 22.558 20.522 22.594 ;
               RECT 20.47 23.235 20.522 23.271 ;
               RECT 20.47 23.529 20.522 23.565 ;
               RECT 20.47 23.758 20.522 23.794 ;
               RECT 20.47 24.435 20.522 24.471 ;
               RECT 20.47 24.729 20.522 24.765 ;
               RECT 20.47 24.958 20.522 24.994 ;
               RECT 20.47 25.635 20.522 25.671 ;
               RECT 20.47 25.929 20.522 25.965 ;
               RECT 20.47 26.158 20.522 26.194 ;
               RECT 20.47 26.835 20.522 26.871 ;
               RECT 20.47 27.129 20.522 27.165 ;
               RECT 20.47 27.358 20.522 27.394 ;
               RECT 20.47 28.035 20.522 28.071 ;
               RECT 20.47 28.329 20.522 28.365 ;
               RECT 20.47 28.558 20.522 28.594 ;
               RECT 20.47 29.235 20.522 29.271 ;
               RECT 20.47 29.529 20.522 29.565 ;
               RECT 20.47 29.758 20.522 29.794 ;
               RECT 20.47 30.435 20.522 30.471 ;
               RECT 20.47 30.729 20.522 30.765 ;
               RECT 20.47 30.958 20.522 30.994 ;
               RECT 20.47 31.635 20.522 31.671 ;
               RECT 20.47 31.929 20.522 31.965 ;
               RECT 20.47 32.158 20.522 32.194 ;
               RECT 20.47 32.835 20.522 32.871 ;
               RECT 20.47 33.129 20.522 33.165 ;
               RECT 20.47 33.358 20.522 33.394 ;
               RECT 20.47 34.035 20.522 34.071 ;
               RECT 20.47 34.329 20.522 34.365 ;
               RECT 20.47 34.558 20.522 34.594 ;
               RECT 20.47 35.235 20.522 35.271 ;
               RECT 20.47 35.529 20.522 35.565 ;
               RECT 20.47 35.758 20.522 35.794 ;
               RECT 20.47 36.435 20.522 36.471 ;
               RECT 20.47 36.729 20.522 36.765 ;
               RECT 20.47 36.958 20.522 36.994 ;
               RECT 20.47 37.635 20.522 37.671 ;
               RECT 20.47 37.929 20.522 37.965 ;
               RECT 20.47 38.158 20.522 38.194 ;
               RECT 20.47 38.835 20.522 38.871 ;
               RECT 20.47 39.129 20.522 39.165 ;
               RECT 20.47 39.358 20.522 39.394 ;
               RECT 20.47 40.035 20.522 40.071 ;
               RECT 20.47 40.329 20.522 40.365 ;
               RECT 20.47 40.558 20.522 40.594 ;
               RECT 20.47 41.235 20.522 41.271 ;
               RECT 20.47 41.529 20.522 41.565 ;
               RECT 20.47 41.758 20.522 41.794 ;
               RECT 20.47 42.435 20.522 42.471 ;
               RECT 20.47 42.729 20.522 42.765 ;
               RECT 20.47 42.958 20.522 42.994 ;
               RECT 20.47 43.635 20.522 43.671 ;
               RECT 20.47 43.929 20.522 43.965 ;
               RECT 20.47 44.158 20.522 44.194 ;
               RECT 20.47 44.835 20.522 44.871 ;
               RECT 20.47 45.129 20.522 45.165 ;
               RECT 20.47 45.358 20.522 45.394 ;
               RECT 20.47 46.035 20.522 46.071 ;
               RECT 20.47 46.329 20.522 46.365 ;
               RECT 20.47 46.558 20.522 46.594 ;
               RECT 20.47 47.235 20.522 47.271 ;
               RECT 20.47 47.529 20.522 47.565 ;
               RECT 20.47 47.758 20.522 47.794 ;
               RECT 20.47 48.435 20.522 48.471 ;
               RECT 20.47 49.182 20.522 49.218 ;
          END
          PORT
               LAYER m5 ;
               RECT 20.47 54.999 20.522 104.5505 ;
               LAYER v4 ;
               RECT 20.47 55.422 20.522 55.458 ;
               RECT 20.47 55.902 20.522 55.938 ;
               RECT 20.47 56.649 20.522 56.685 ;
               RECT 20.47 56.878 20.522 56.914 ;
               RECT 20.47 57.555 20.522 57.591 ;
               RECT 20.47 57.849 20.522 57.885 ;
               RECT 20.47 58.078 20.522 58.114 ;
               RECT 20.47 58.755 20.522 58.791 ;
               RECT 20.47 59.049 20.522 59.085 ;
               RECT 20.47 59.278 20.522 59.314 ;
               RECT 20.47 59.955 20.522 59.991 ;
               RECT 20.47 60.249 20.522 60.285 ;
               RECT 20.47 60.478 20.522 60.514 ;
               RECT 20.47 61.155 20.522 61.191 ;
               RECT 20.47 61.449 20.522 61.485 ;
               RECT 20.47 61.678 20.522 61.714 ;
               RECT 20.47 62.355 20.522 62.391 ;
               RECT 20.47 62.649 20.522 62.685 ;
               RECT 20.47 62.878 20.522 62.914 ;
               RECT 20.47 63.555 20.522 63.591 ;
               RECT 20.47 63.849 20.522 63.885 ;
               RECT 20.47 64.078 20.522 64.114 ;
               RECT 20.47 64.755 20.522 64.791 ;
               RECT 20.47 65.049 20.522 65.085 ;
               RECT 20.47 65.278 20.522 65.314 ;
               RECT 20.47 65.955 20.522 65.991 ;
               RECT 20.47 66.249 20.522 66.285 ;
               RECT 20.47 66.478 20.522 66.514 ;
               RECT 20.47 67.155 20.522 67.191 ;
               RECT 20.47 67.449 20.522 67.485 ;
               RECT 20.47 67.678 20.522 67.714 ;
               RECT 20.47 68.355 20.522 68.391 ;
               RECT 20.47 68.649 20.522 68.685 ;
               RECT 20.47 68.878 20.522 68.914 ;
               RECT 20.47 69.555 20.522 69.591 ;
               RECT 20.47 69.849 20.522 69.885 ;
               RECT 20.47 70.078 20.522 70.114 ;
               RECT 20.47 70.755 20.522 70.791 ;
               RECT 20.47 71.049 20.522 71.085 ;
               RECT 20.47 71.278 20.522 71.314 ;
               RECT 20.47 71.955 20.522 71.991 ;
               RECT 20.47 72.249 20.522 72.285 ;
               RECT 20.47 72.478 20.522 72.514 ;
               RECT 20.47 73.155 20.522 73.191 ;
               RECT 20.47 73.449 20.522 73.485 ;
               RECT 20.47 73.678 20.522 73.714 ;
               RECT 20.47 74.355 20.522 74.391 ;
               RECT 20.47 74.649 20.522 74.685 ;
               RECT 20.47 74.878 20.522 74.914 ;
               RECT 20.47 75.555 20.522 75.591 ;
               RECT 20.47 75.849 20.522 75.885 ;
               RECT 20.47 76.078 20.522 76.114 ;
               RECT 20.47 76.755 20.522 76.791 ;
               RECT 20.47 77.049 20.522 77.085 ;
               RECT 20.47 77.278 20.522 77.314 ;
               RECT 20.47 77.955 20.522 77.991 ;
               RECT 20.47 78.249 20.522 78.285 ;
               RECT 20.47 78.478 20.522 78.514 ;
               RECT 20.47 79.155 20.522 79.191 ;
               RECT 20.47 79.449 20.522 79.485 ;
               RECT 20.47 79.678 20.522 79.714 ;
               RECT 20.47 80.355 20.522 80.391 ;
               RECT 20.47 80.649 20.522 80.685 ;
               RECT 20.47 80.878 20.522 80.914 ;
               RECT 20.47 81.555 20.522 81.591 ;
               RECT 20.47 81.849 20.522 81.885 ;
               RECT 20.47 82.078 20.522 82.114 ;
               RECT 20.47 82.755 20.522 82.791 ;
               RECT 20.47 83.049 20.522 83.085 ;
               RECT 20.47 83.278 20.522 83.314 ;
               RECT 20.47 83.955 20.522 83.991 ;
               RECT 20.47 84.249 20.522 84.285 ;
               RECT 20.47 84.478 20.522 84.514 ;
               RECT 20.47 85.155 20.522 85.191 ;
               RECT 20.47 85.449 20.522 85.485 ;
               RECT 20.47 85.678 20.522 85.714 ;
               RECT 20.47 86.355 20.522 86.391 ;
               RECT 20.47 86.649 20.522 86.685 ;
               RECT 20.47 86.878 20.522 86.914 ;
               RECT 20.47 87.555 20.522 87.591 ;
               RECT 20.47 87.849 20.522 87.885 ;
               RECT 20.47 88.078 20.522 88.114 ;
               RECT 20.47 88.755 20.522 88.791 ;
               RECT 20.47 89.049 20.522 89.085 ;
               RECT 20.47 89.278 20.522 89.314 ;
               RECT 20.47 89.955 20.522 89.991 ;
               RECT 20.47 90.249 20.522 90.285 ;
               RECT 20.47 90.478 20.522 90.514 ;
               RECT 20.47 91.155 20.522 91.191 ;
               RECT 20.47 91.449 20.522 91.485 ;
               RECT 20.47 91.678 20.522 91.714 ;
               RECT 20.47 92.355 20.522 92.391 ;
               RECT 20.47 92.649 20.522 92.685 ;
               RECT 20.47 92.878 20.522 92.914 ;
               RECT 20.47 93.555 20.522 93.591 ;
               RECT 20.47 93.849 20.522 93.885 ;
               RECT 20.47 94.078 20.522 94.114 ;
               RECT 20.47 94.755 20.522 94.791 ;
               RECT 20.47 95.049 20.522 95.085 ;
               RECT 20.47 95.278 20.522 95.314 ;
               RECT 20.47 95.955 20.522 95.991 ;
               RECT 20.47 96.249 20.522 96.285 ;
               RECT 20.47 96.478 20.522 96.514 ;
               RECT 20.47 97.155 20.522 97.191 ;
               RECT 20.47 97.449 20.522 97.485 ;
               RECT 20.47 97.678 20.522 97.714 ;
               RECT 20.47 98.355 20.522 98.391 ;
               RECT 20.47 98.649 20.522 98.685 ;
               RECT 20.47 98.878 20.522 98.914 ;
               RECT 20.47 99.555 20.522 99.591 ;
               RECT 20.47 99.849 20.522 99.885 ;
               RECT 20.47 100.078 20.522 100.114 ;
               RECT 20.47 100.755 20.522 100.791 ;
               RECT 20.47 101.049 20.522 101.085 ;
               RECT 20.47 101.278 20.522 101.314 ;
               RECT 20.47 101.955 20.522 101.991 ;
               RECT 20.47 102.249 20.522 102.285 ;
               RECT 20.47 102.478 20.522 102.514 ;
               RECT 20.47 103.155 20.522 103.191 ;
               RECT 20.47 103.449 20.522 103.485 ;
               RECT 20.47 103.678 20.522 103.714 ;
               RECT 20.47 104.355 20.522 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 20.63 0.5695 20.682 104.5505 ;
               LAYER v4 ;
               RECT 20.63 0.729 20.682 0.765 ;
               RECT 20.63 0.958 20.682 0.994 ;
               RECT 20.63 1.406 20.682 1.442 ;
               RECT 20.63 1.635 20.682 1.671 ;
               RECT 20.63 1.929 20.682 1.965 ;
               RECT 20.63 2.158 20.682 2.194 ;
               RECT 20.63 2.606 20.682 2.642 ;
               RECT 20.63 2.835 20.682 2.871 ;
               RECT 20.63 3.129 20.682 3.165 ;
               RECT 20.63 3.358 20.682 3.394 ;
               RECT 20.63 3.806 20.682 3.842 ;
               RECT 20.63 4.035 20.682 4.071 ;
               RECT 20.63 4.329 20.682 4.365 ;
               RECT 20.63 4.558 20.682 4.594 ;
               RECT 20.63 5.006 20.682 5.042 ;
               RECT 20.63 5.235 20.682 5.271 ;
               RECT 20.63 5.529 20.682 5.565 ;
               RECT 20.63 5.758 20.682 5.794 ;
               RECT 20.63 6.206 20.682 6.242 ;
               RECT 20.63 6.435 20.682 6.471 ;
               RECT 20.63 6.729 20.682 6.765 ;
               RECT 20.63 6.958 20.682 6.994 ;
               RECT 20.63 7.406 20.682 7.442 ;
               RECT 20.63 7.635 20.682 7.671 ;
               RECT 20.63 7.929 20.682 7.965 ;
               RECT 20.63 8.158 20.682 8.194 ;
               RECT 20.63 8.606 20.682 8.642 ;
               RECT 20.63 8.835 20.682 8.871 ;
               RECT 20.63 9.129 20.682 9.165 ;
               RECT 20.63 9.358 20.682 9.394 ;
               RECT 20.63 9.806 20.682 9.842 ;
               RECT 20.63 10.035 20.682 10.071 ;
               RECT 20.63 10.329 20.682 10.365 ;
               RECT 20.63 10.558 20.682 10.594 ;
               RECT 20.63 11.006 20.682 11.042 ;
               RECT 20.63 11.235 20.682 11.271 ;
               RECT 20.63 11.529 20.682 11.565 ;
               RECT 20.63 11.758 20.682 11.794 ;
               RECT 20.63 12.206 20.682 12.242 ;
               RECT 20.63 12.435 20.682 12.471 ;
               RECT 20.63 12.729 20.682 12.765 ;
               RECT 20.63 12.958 20.682 12.994 ;
               RECT 20.63 13.406 20.682 13.442 ;
               RECT 20.63 13.635 20.682 13.671 ;
               RECT 20.63 13.929 20.682 13.965 ;
               RECT 20.63 14.158 20.682 14.194 ;
               RECT 20.63 14.606 20.682 14.642 ;
               RECT 20.63 14.835 20.682 14.871 ;
               RECT 20.63 15.129 20.682 15.165 ;
               RECT 20.63 15.358 20.682 15.394 ;
               RECT 20.63 15.806 20.682 15.842 ;
               RECT 20.63 16.035 20.682 16.071 ;
               RECT 20.63 16.329 20.682 16.365 ;
               RECT 20.63 16.558 20.682 16.594 ;
               RECT 20.63 17.006 20.682 17.042 ;
               RECT 20.63 17.235 20.682 17.271 ;
               RECT 20.63 17.529 20.682 17.565 ;
               RECT 20.63 17.758 20.682 17.794 ;
               RECT 20.63 18.206 20.682 18.242 ;
               RECT 20.63 18.435 20.682 18.471 ;
               RECT 20.63 18.729 20.682 18.765 ;
               RECT 20.63 18.958 20.682 18.994 ;
               RECT 20.63 19.406 20.682 19.442 ;
               RECT 20.63 19.635 20.682 19.671 ;
               RECT 20.63 19.929 20.682 19.965 ;
               RECT 20.63 20.158 20.682 20.194 ;
               RECT 20.63 20.606 20.682 20.642 ;
               RECT 20.63 20.835 20.682 20.871 ;
               RECT 20.63 21.129 20.682 21.165 ;
               RECT 20.63 21.358 20.682 21.394 ;
               RECT 20.63 21.806 20.682 21.842 ;
               RECT 20.63 22.035 20.682 22.071 ;
               RECT 20.63 22.329 20.682 22.365 ;
               RECT 20.63 22.558 20.682 22.594 ;
               RECT 20.63 23.006 20.682 23.042 ;
               RECT 20.63 23.235 20.682 23.271 ;
               RECT 20.63 23.529 20.682 23.565 ;
               RECT 20.63 23.758 20.682 23.794 ;
               RECT 20.63 24.206 20.682 24.242 ;
               RECT 20.63 24.435 20.682 24.471 ;
               RECT 20.63 24.729 20.682 24.765 ;
               RECT 20.63 24.958 20.682 24.994 ;
               RECT 20.63 25.406 20.682 25.442 ;
               RECT 20.63 25.635 20.682 25.671 ;
               RECT 20.63 25.929 20.682 25.965 ;
               RECT 20.63 26.158 20.682 26.194 ;
               RECT 20.63 26.606 20.682 26.642 ;
               RECT 20.63 26.835 20.682 26.871 ;
               RECT 20.63 27.129 20.682 27.165 ;
               RECT 20.63 27.358 20.682 27.394 ;
               RECT 20.63 27.806 20.682 27.842 ;
               RECT 20.63 28.035 20.682 28.071 ;
               RECT 20.63 28.329 20.682 28.365 ;
               RECT 20.63 28.558 20.682 28.594 ;
               RECT 20.63 29.006 20.682 29.042 ;
               RECT 20.63 29.235 20.682 29.271 ;
               RECT 20.63 29.529 20.682 29.565 ;
               RECT 20.63 29.758 20.682 29.794 ;
               RECT 20.63 30.206 20.682 30.242 ;
               RECT 20.63 30.435 20.682 30.471 ;
               RECT 20.63 30.729 20.682 30.765 ;
               RECT 20.63 30.958 20.682 30.994 ;
               RECT 20.63 31.406 20.682 31.442 ;
               RECT 20.63 31.635 20.682 31.671 ;
               RECT 20.63 31.929 20.682 31.965 ;
               RECT 20.63 32.158 20.682 32.194 ;
               RECT 20.63 32.606 20.682 32.642 ;
               RECT 20.63 32.835 20.682 32.871 ;
               RECT 20.63 33.129 20.682 33.165 ;
               RECT 20.63 33.358 20.682 33.394 ;
               RECT 20.63 33.806 20.682 33.842 ;
               RECT 20.63 34.035 20.682 34.071 ;
               RECT 20.63 34.329 20.682 34.365 ;
               RECT 20.63 34.558 20.682 34.594 ;
               RECT 20.63 35.006 20.682 35.042 ;
               RECT 20.63 35.235 20.682 35.271 ;
               RECT 20.63 35.529 20.682 35.565 ;
               RECT 20.63 35.758 20.682 35.794 ;
               RECT 20.63 36.206 20.682 36.242 ;
               RECT 20.63 36.435 20.682 36.471 ;
               RECT 20.63 36.729 20.682 36.765 ;
               RECT 20.63 36.958 20.682 36.994 ;
               RECT 20.63 37.406 20.682 37.442 ;
               RECT 20.63 37.635 20.682 37.671 ;
               RECT 20.63 37.929 20.682 37.965 ;
               RECT 20.63 38.158 20.682 38.194 ;
               RECT 20.63 38.606 20.682 38.642 ;
               RECT 20.63 38.835 20.682 38.871 ;
               RECT 20.63 39.129 20.682 39.165 ;
               RECT 20.63 39.358 20.682 39.394 ;
               RECT 20.63 39.806 20.682 39.842 ;
               RECT 20.63 40.035 20.682 40.071 ;
               RECT 20.63 40.329 20.682 40.365 ;
               RECT 20.63 40.558 20.682 40.594 ;
               RECT 20.63 41.006 20.682 41.042 ;
               RECT 20.63 41.235 20.682 41.271 ;
               RECT 20.63 41.529 20.682 41.565 ;
               RECT 20.63 41.758 20.682 41.794 ;
               RECT 20.63 42.206 20.682 42.242 ;
               RECT 20.63 42.435 20.682 42.471 ;
               RECT 20.63 42.729 20.682 42.765 ;
               RECT 20.63 42.958 20.682 42.994 ;
               RECT 20.63 43.406 20.682 43.442 ;
               RECT 20.63 43.635 20.682 43.671 ;
               RECT 20.63 43.929 20.682 43.965 ;
               RECT 20.63 44.158 20.682 44.194 ;
               RECT 20.63 44.606 20.682 44.642 ;
               RECT 20.63 44.835 20.682 44.871 ;
               RECT 20.63 45.129 20.682 45.165 ;
               RECT 20.63 45.358 20.682 45.394 ;
               RECT 20.63 45.806 20.682 45.842 ;
               RECT 20.63 46.035 20.682 46.071 ;
               RECT 20.63 46.329 20.682 46.365 ;
               RECT 20.63 46.558 20.682 46.594 ;
               RECT 20.63 47.006 20.682 47.042 ;
               RECT 20.63 47.235 20.682 47.271 ;
               RECT 20.63 47.529 20.682 47.565 ;
               RECT 20.63 47.758 20.682 47.794 ;
               RECT 20.63 48.206 20.682 48.242 ;
               RECT 20.63 48.435 20.682 48.471 ;
               RECT 20.63 49.182 20.682 49.218 ;
               RECT 20.63 49.662 20.682 49.698 ;
               RECT 20.63 49.8435 20.682 49.8795 ;
               RECT 20.63 50.142 20.682 50.178 ;
               RECT 20.63 50.622 20.682 50.658 ;
               RECT 20.63 51.102 20.682 51.138 ;
               RECT 20.63 51.582 20.682 51.618 ;
               RECT 20.63 52.062 20.682 52.098 ;
               RECT 20.63 52.542 20.682 52.578 ;
               RECT 20.63 53.022 20.682 53.058 ;
               RECT 20.63 53.502 20.682 53.538 ;
               RECT 20.63 53.982 20.682 54.018 ;
               RECT 20.63 54.4675 20.682 54.4925 ;
               RECT 20.63 54.942 20.682 54.978 ;
               RECT 20.63 55.422 20.682 55.458 ;
               RECT 20.63 55.902 20.682 55.938 ;
               RECT 20.63 56.649 20.682 56.685 ;
               RECT 20.63 56.878 20.682 56.914 ;
               RECT 20.63 57.326 20.682 57.362 ;
               RECT 20.63 57.555 20.682 57.591 ;
               RECT 20.63 57.849 20.682 57.885 ;
               RECT 20.63 58.078 20.682 58.114 ;
               RECT 20.63 58.526 20.682 58.562 ;
               RECT 20.63 58.755 20.682 58.791 ;
               RECT 20.63 59.049 20.682 59.085 ;
               RECT 20.63 59.278 20.682 59.314 ;
               RECT 20.63 59.726 20.682 59.762 ;
               RECT 20.63 59.955 20.682 59.991 ;
               RECT 20.63 60.249 20.682 60.285 ;
               RECT 20.63 60.478 20.682 60.514 ;
               RECT 20.63 60.926 20.682 60.962 ;
               RECT 20.63 61.155 20.682 61.191 ;
               RECT 20.63 61.449 20.682 61.485 ;
               RECT 20.63 61.678 20.682 61.714 ;
               RECT 20.63 62.126 20.682 62.162 ;
               RECT 20.63 62.355 20.682 62.391 ;
               RECT 20.63 62.649 20.682 62.685 ;
               RECT 20.63 62.878 20.682 62.914 ;
               RECT 20.63 63.326 20.682 63.362 ;
               RECT 20.63 63.555 20.682 63.591 ;
               RECT 20.63 63.849 20.682 63.885 ;
               RECT 20.63 64.078 20.682 64.114 ;
               RECT 20.63 64.526 20.682 64.562 ;
               RECT 20.63 64.755 20.682 64.791 ;
               RECT 20.63 65.049 20.682 65.085 ;
               RECT 20.63 65.278 20.682 65.314 ;
               RECT 20.63 65.726 20.682 65.762 ;
               RECT 20.63 65.955 20.682 65.991 ;
               RECT 20.63 66.249 20.682 66.285 ;
               RECT 20.63 66.478 20.682 66.514 ;
               RECT 20.63 66.926 20.682 66.962 ;
               RECT 20.63 67.155 20.682 67.191 ;
               RECT 20.63 67.449 20.682 67.485 ;
               RECT 20.63 67.678 20.682 67.714 ;
               RECT 20.63 68.126 20.682 68.162 ;
               RECT 20.63 68.355 20.682 68.391 ;
               RECT 20.63 68.649 20.682 68.685 ;
               RECT 20.63 68.878 20.682 68.914 ;
               RECT 20.63 69.326 20.682 69.362 ;
               RECT 20.63 69.555 20.682 69.591 ;
               RECT 20.63 69.849 20.682 69.885 ;
               RECT 20.63 70.078 20.682 70.114 ;
               RECT 20.63 70.526 20.682 70.562 ;
               RECT 20.63 70.755 20.682 70.791 ;
               RECT 20.63 71.049 20.682 71.085 ;
               RECT 20.63 71.278 20.682 71.314 ;
               RECT 20.63 71.726 20.682 71.762 ;
               RECT 20.63 71.955 20.682 71.991 ;
               RECT 20.63 72.249 20.682 72.285 ;
               RECT 20.63 72.478 20.682 72.514 ;
               RECT 20.63 72.926 20.682 72.962 ;
               RECT 20.63 73.155 20.682 73.191 ;
               RECT 20.63 73.449 20.682 73.485 ;
               RECT 20.63 73.678 20.682 73.714 ;
               RECT 20.63 74.126 20.682 74.162 ;
               RECT 20.63 74.355 20.682 74.391 ;
               RECT 20.63 74.649 20.682 74.685 ;
               RECT 20.63 74.878 20.682 74.914 ;
               RECT 20.63 75.326 20.682 75.362 ;
               RECT 20.63 75.555 20.682 75.591 ;
               RECT 20.63 75.849 20.682 75.885 ;
               RECT 20.63 76.078 20.682 76.114 ;
               RECT 20.63 76.526 20.682 76.562 ;
               RECT 20.63 76.755 20.682 76.791 ;
               RECT 20.63 77.049 20.682 77.085 ;
               RECT 20.63 77.278 20.682 77.314 ;
               RECT 20.63 77.726 20.682 77.762 ;
               RECT 20.63 77.955 20.682 77.991 ;
               RECT 20.63 78.249 20.682 78.285 ;
               RECT 20.63 78.478 20.682 78.514 ;
               RECT 20.63 78.926 20.682 78.962 ;
               RECT 20.63 79.155 20.682 79.191 ;
               RECT 20.63 79.449 20.682 79.485 ;
               RECT 20.63 79.678 20.682 79.714 ;
               RECT 20.63 80.126 20.682 80.162 ;
               RECT 20.63 80.355 20.682 80.391 ;
               RECT 20.63 80.649 20.682 80.685 ;
               RECT 20.63 80.878 20.682 80.914 ;
               RECT 20.63 81.326 20.682 81.362 ;
               RECT 20.63 81.555 20.682 81.591 ;
               RECT 20.63 81.849 20.682 81.885 ;
               RECT 20.63 82.078 20.682 82.114 ;
               RECT 20.63 82.526 20.682 82.562 ;
               RECT 20.63 82.755 20.682 82.791 ;
               RECT 20.63 83.049 20.682 83.085 ;
               RECT 20.63 83.278 20.682 83.314 ;
               RECT 20.63 83.726 20.682 83.762 ;
               RECT 20.63 83.955 20.682 83.991 ;
               RECT 20.63 84.249 20.682 84.285 ;
               RECT 20.63 84.478 20.682 84.514 ;
               RECT 20.63 84.926 20.682 84.962 ;
               RECT 20.63 85.155 20.682 85.191 ;
               RECT 20.63 85.449 20.682 85.485 ;
               RECT 20.63 85.678 20.682 85.714 ;
               RECT 20.63 86.126 20.682 86.162 ;
               RECT 20.63 86.355 20.682 86.391 ;
               RECT 20.63 86.649 20.682 86.685 ;
               RECT 20.63 86.878 20.682 86.914 ;
               RECT 20.63 87.326 20.682 87.362 ;
               RECT 20.63 87.555 20.682 87.591 ;
               RECT 20.63 87.849 20.682 87.885 ;
               RECT 20.63 88.078 20.682 88.114 ;
               RECT 20.63 88.526 20.682 88.562 ;
               RECT 20.63 88.755 20.682 88.791 ;
               RECT 20.63 89.049 20.682 89.085 ;
               RECT 20.63 89.278 20.682 89.314 ;
               RECT 20.63 89.726 20.682 89.762 ;
               RECT 20.63 89.955 20.682 89.991 ;
               RECT 20.63 90.249 20.682 90.285 ;
               RECT 20.63 90.478 20.682 90.514 ;
               RECT 20.63 90.926 20.682 90.962 ;
               RECT 20.63 91.155 20.682 91.191 ;
               RECT 20.63 91.449 20.682 91.485 ;
               RECT 20.63 91.678 20.682 91.714 ;
               RECT 20.63 92.126 20.682 92.162 ;
               RECT 20.63 92.355 20.682 92.391 ;
               RECT 20.63 92.649 20.682 92.685 ;
               RECT 20.63 92.878 20.682 92.914 ;
               RECT 20.63 93.326 20.682 93.362 ;
               RECT 20.63 93.555 20.682 93.591 ;
               RECT 20.63 93.849 20.682 93.885 ;
               RECT 20.63 94.078 20.682 94.114 ;
               RECT 20.63 94.526 20.682 94.562 ;
               RECT 20.63 94.755 20.682 94.791 ;
               RECT 20.63 95.049 20.682 95.085 ;
               RECT 20.63 95.278 20.682 95.314 ;
               RECT 20.63 95.726 20.682 95.762 ;
               RECT 20.63 95.955 20.682 95.991 ;
               RECT 20.63 96.249 20.682 96.285 ;
               RECT 20.63 96.478 20.682 96.514 ;
               RECT 20.63 96.926 20.682 96.962 ;
               RECT 20.63 97.155 20.682 97.191 ;
               RECT 20.63 97.449 20.682 97.485 ;
               RECT 20.63 97.678 20.682 97.714 ;
               RECT 20.63 98.126 20.682 98.162 ;
               RECT 20.63 98.355 20.682 98.391 ;
               RECT 20.63 98.649 20.682 98.685 ;
               RECT 20.63 98.878 20.682 98.914 ;
               RECT 20.63 99.326 20.682 99.362 ;
               RECT 20.63 99.555 20.682 99.591 ;
               RECT 20.63 99.849 20.682 99.885 ;
               RECT 20.63 100.078 20.682 100.114 ;
               RECT 20.63 100.526 20.682 100.562 ;
               RECT 20.63 100.755 20.682 100.791 ;
               RECT 20.63 101.049 20.682 101.085 ;
               RECT 20.63 101.278 20.682 101.314 ;
               RECT 20.63 101.726 20.682 101.762 ;
               RECT 20.63 101.955 20.682 101.991 ;
               RECT 20.63 102.249 20.682 102.285 ;
               RECT 20.63 102.478 20.682 102.514 ;
               RECT 20.63 102.926 20.682 102.962 ;
               RECT 20.63 103.155 20.682 103.191 ;
               RECT 20.63 103.449 20.682 103.485 ;
               RECT 20.63 103.678 20.682 103.714 ;
               RECT 20.63 104.126 20.682 104.162 ;
               RECT 20.63 104.355 20.682 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 21.014 0.5695 21.068 104.5505 ;
               LAYER v4 ;
               RECT 21.014 0.729 21.068 0.765 ;
               RECT 21.014 0.958 21.068 0.994 ;
               RECT 21.014 1.406 21.068 1.442 ;
               RECT 21.014 1.635 21.068 1.671 ;
               RECT 21.014 1.929 21.068 1.965 ;
               RECT 21.014 2.158 21.068 2.194 ;
               RECT 21.014 2.606 21.068 2.642 ;
               RECT 21.014 2.835 21.068 2.871 ;
               RECT 21.014 3.129 21.068 3.165 ;
               RECT 21.014 3.358 21.068 3.394 ;
               RECT 21.014 3.806 21.068 3.842 ;
               RECT 21.014 4.035 21.068 4.071 ;
               RECT 21.014 4.329 21.068 4.365 ;
               RECT 21.014 4.558 21.068 4.594 ;
               RECT 21.014 5.006 21.068 5.042 ;
               RECT 21.014 5.235 21.068 5.271 ;
               RECT 21.014 5.529 21.068 5.565 ;
               RECT 21.014 5.758 21.068 5.794 ;
               RECT 21.014 6.206 21.068 6.242 ;
               RECT 21.014 6.435 21.068 6.471 ;
               RECT 21.014 6.729 21.068 6.765 ;
               RECT 21.014 6.958 21.068 6.994 ;
               RECT 21.014 7.406 21.068 7.442 ;
               RECT 21.014 7.635 21.068 7.671 ;
               RECT 21.014 7.929 21.068 7.965 ;
               RECT 21.014 8.158 21.068 8.194 ;
               RECT 21.014 8.606 21.068 8.642 ;
               RECT 21.014 8.835 21.068 8.871 ;
               RECT 21.014 9.129 21.068 9.165 ;
               RECT 21.014 9.358 21.068 9.394 ;
               RECT 21.014 9.806 21.068 9.842 ;
               RECT 21.014 10.035 21.068 10.071 ;
               RECT 21.014 10.329 21.068 10.365 ;
               RECT 21.014 10.558 21.068 10.594 ;
               RECT 21.014 11.006 21.068 11.042 ;
               RECT 21.014 11.235 21.068 11.271 ;
               RECT 21.014 11.529 21.068 11.565 ;
               RECT 21.014 11.758 21.068 11.794 ;
               RECT 21.014 12.206 21.068 12.242 ;
               RECT 21.014 12.435 21.068 12.471 ;
               RECT 21.014 12.729 21.068 12.765 ;
               RECT 21.014 12.958 21.068 12.994 ;
               RECT 21.014 13.406 21.068 13.442 ;
               RECT 21.014 13.635 21.068 13.671 ;
               RECT 21.014 13.929 21.068 13.965 ;
               RECT 21.014 14.158 21.068 14.194 ;
               RECT 21.014 14.606 21.068 14.642 ;
               RECT 21.014 14.835 21.068 14.871 ;
               RECT 21.014 15.129 21.068 15.165 ;
               RECT 21.014 15.358 21.068 15.394 ;
               RECT 21.014 15.806 21.068 15.842 ;
               RECT 21.014 16.035 21.068 16.071 ;
               RECT 21.014 16.329 21.068 16.365 ;
               RECT 21.014 16.558 21.068 16.594 ;
               RECT 21.014 17.006 21.068 17.042 ;
               RECT 21.014 17.235 21.068 17.271 ;
               RECT 21.014 17.529 21.068 17.565 ;
               RECT 21.014 17.758 21.068 17.794 ;
               RECT 21.014 18.206 21.068 18.242 ;
               RECT 21.014 18.435 21.068 18.471 ;
               RECT 21.014 18.729 21.068 18.765 ;
               RECT 21.014 18.958 21.068 18.994 ;
               RECT 21.014 19.406 21.068 19.442 ;
               RECT 21.014 19.635 21.068 19.671 ;
               RECT 21.014 19.929 21.068 19.965 ;
               RECT 21.014 20.158 21.068 20.194 ;
               RECT 21.014 20.606 21.068 20.642 ;
               RECT 21.014 20.835 21.068 20.871 ;
               RECT 21.014 21.129 21.068 21.165 ;
               RECT 21.014 21.358 21.068 21.394 ;
               RECT 21.014 21.806 21.068 21.842 ;
               RECT 21.014 22.035 21.068 22.071 ;
               RECT 21.014 22.329 21.068 22.365 ;
               RECT 21.014 22.558 21.068 22.594 ;
               RECT 21.014 23.006 21.068 23.042 ;
               RECT 21.014 23.235 21.068 23.271 ;
               RECT 21.014 23.529 21.068 23.565 ;
               RECT 21.014 23.758 21.068 23.794 ;
               RECT 21.014 24.206 21.068 24.242 ;
               RECT 21.014 24.435 21.068 24.471 ;
               RECT 21.014 24.729 21.068 24.765 ;
               RECT 21.014 24.958 21.068 24.994 ;
               RECT 21.014 25.406 21.068 25.442 ;
               RECT 21.014 25.635 21.068 25.671 ;
               RECT 21.014 25.929 21.068 25.965 ;
               RECT 21.014 26.158 21.068 26.194 ;
               RECT 21.014 26.606 21.068 26.642 ;
               RECT 21.014 26.835 21.068 26.871 ;
               RECT 21.014 27.129 21.068 27.165 ;
               RECT 21.014 27.358 21.068 27.394 ;
               RECT 21.014 27.806 21.068 27.842 ;
               RECT 21.014 28.035 21.068 28.071 ;
               RECT 21.014 28.329 21.068 28.365 ;
               RECT 21.014 28.558 21.068 28.594 ;
               RECT 21.014 29.006 21.068 29.042 ;
               RECT 21.014 29.235 21.068 29.271 ;
               RECT 21.014 29.529 21.068 29.565 ;
               RECT 21.014 29.758 21.068 29.794 ;
               RECT 21.014 30.206 21.068 30.242 ;
               RECT 21.014 30.435 21.068 30.471 ;
               RECT 21.014 30.729 21.068 30.765 ;
               RECT 21.014 30.958 21.068 30.994 ;
               RECT 21.014 31.406 21.068 31.442 ;
               RECT 21.014 31.635 21.068 31.671 ;
               RECT 21.014 31.929 21.068 31.965 ;
               RECT 21.014 32.158 21.068 32.194 ;
               RECT 21.014 32.606 21.068 32.642 ;
               RECT 21.014 32.835 21.068 32.871 ;
               RECT 21.014 33.129 21.068 33.165 ;
               RECT 21.014 33.358 21.068 33.394 ;
               RECT 21.014 33.806 21.068 33.842 ;
               RECT 21.014 34.035 21.068 34.071 ;
               RECT 21.014 34.329 21.068 34.365 ;
               RECT 21.014 34.558 21.068 34.594 ;
               RECT 21.014 35.006 21.068 35.042 ;
               RECT 21.014 35.235 21.068 35.271 ;
               RECT 21.014 35.529 21.068 35.565 ;
               RECT 21.014 35.758 21.068 35.794 ;
               RECT 21.014 36.206 21.068 36.242 ;
               RECT 21.014 36.435 21.068 36.471 ;
               RECT 21.014 36.729 21.068 36.765 ;
               RECT 21.014 36.958 21.068 36.994 ;
               RECT 21.014 37.406 21.068 37.442 ;
               RECT 21.014 37.635 21.068 37.671 ;
               RECT 21.014 37.929 21.068 37.965 ;
               RECT 21.014 38.158 21.068 38.194 ;
               RECT 21.014 38.606 21.068 38.642 ;
               RECT 21.014 38.835 21.068 38.871 ;
               RECT 21.014 39.129 21.068 39.165 ;
               RECT 21.014 39.358 21.068 39.394 ;
               RECT 21.014 39.806 21.068 39.842 ;
               RECT 21.014 40.035 21.068 40.071 ;
               RECT 21.014 40.329 21.068 40.365 ;
               RECT 21.014 40.558 21.068 40.594 ;
               RECT 21.014 41.006 21.068 41.042 ;
               RECT 21.014 41.235 21.068 41.271 ;
               RECT 21.014 41.529 21.068 41.565 ;
               RECT 21.014 41.758 21.068 41.794 ;
               RECT 21.014 42.206 21.068 42.242 ;
               RECT 21.014 42.435 21.068 42.471 ;
               RECT 21.014 42.729 21.068 42.765 ;
               RECT 21.014 42.958 21.068 42.994 ;
               RECT 21.014 43.406 21.068 43.442 ;
               RECT 21.014 43.635 21.068 43.671 ;
               RECT 21.014 43.929 21.068 43.965 ;
               RECT 21.014 44.158 21.068 44.194 ;
               RECT 21.014 44.606 21.068 44.642 ;
               RECT 21.014 44.835 21.068 44.871 ;
               RECT 21.014 45.129 21.068 45.165 ;
               RECT 21.014 45.358 21.068 45.394 ;
               RECT 21.014 45.806 21.068 45.842 ;
               RECT 21.014 46.035 21.068 46.071 ;
               RECT 21.014 46.329 21.068 46.365 ;
               RECT 21.014 46.558 21.068 46.594 ;
               RECT 21.014 47.006 21.068 47.042 ;
               RECT 21.014 47.235 21.068 47.271 ;
               RECT 21.014 47.529 21.068 47.565 ;
               RECT 21.014 47.758 21.068 47.794 ;
               RECT 21.014 48.206 21.068 48.242 ;
               RECT 21.014 48.435 21.068 48.471 ;
               RECT 21.014 49.062 21.068 49.098 ;
               RECT 21.014 49.182 21.068 49.218 ;
               RECT 21.014 49.542 21.068 49.578 ;
               RECT 21.014 49.662 21.068 49.698 ;
               RECT 21.014 49.782 21.068 49.818 ;
               RECT 21.014 50.262 21.068 50.298 ;
               RECT 21.014 50.622 21.068 50.658 ;
               RECT 21.014 51.102 21.068 51.138 ;
               RECT 21.014 51.582 21.068 51.618 ;
               RECT 21.014 52.062 21.068 52.098 ;
               RECT 21.014 52.182 21.068 52.218 ;
               RECT 21.014 52.542 21.068 52.578 ;
               RECT 21.014 52.902 21.068 52.938 ;
               RECT 21.014 53.022 21.068 53.058 ;
               RECT 21.014 53.502 21.068 53.538 ;
               RECT 21.014 53.982 21.068 54.018 ;
               RECT 21.014 54.462 21.068 54.498 ;
               RECT 21.014 54.822 21.068 54.858 ;
               RECT 21.014 54.942 21.068 54.978 ;
               RECT 21.014 55.302 21.068 55.338 ;
               RECT 21.014 55.422 21.068 55.458 ;
               RECT 21.014 55.542 21.068 55.578 ;
               RECT 21.014 55.902 21.068 55.938 ;
               RECT 21.014 56.649 21.068 56.685 ;
               RECT 21.014 56.878 21.068 56.914 ;
               RECT 21.014 57.326 21.068 57.362 ;
               RECT 21.014 57.555 21.068 57.591 ;
               RECT 21.014 57.849 21.068 57.885 ;
               RECT 21.014 58.078 21.068 58.114 ;
               RECT 21.014 58.526 21.068 58.562 ;
               RECT 21.014 58.755 21.068 58.791 ;
               RECT 21.014 59.049 21.068 59.085 ;
               RECT 21.014 59.278 21.068 59.314 ;
               RECT 21.014 59.726 21.068 59.762 ;
               RECT 21.014 59.955 21.068 59.991 ;
               RECT 21.014 60.249 21.068 60.285 ;
               RECT 21.014 60.478 21.068 60.514 ;
               RECT 21.014 60.926 21.068 60.962 ;
               RECT 21.014 61.155 21.068 61.191 ;
               RECT 21.014 61.449 21.068 61.485 ;
               RECT 21.014 61.678 21.068 61.714 ;
               RECT 21.014 62.126 21.068 62.162 ;
               RECT 21.014 62.355 21.068 62.391 ;
               RECT 21.014 62.649 21.068 62.685 ;
               RECT 21.014 62.878 21.068 62.914 ;
               RECT 21.014 63.326 21.068 63.362 ;
               RECT 21.014 63.555 21.068 63.591 ;
               RECT 21.014 63.849 21.068 63.885 ;
               RECT 21.014 64.078 21.068 64.114 ;
               RECT 21.014 64.526 21.068 64.562 ;
               RECT 21.014 64.755 21.068 64.791 ;
               RECT 21.014 65.049 21.068 65.085 ;
               RECT 21.014 65.278 21.068 65.314 ;
               RECT 21.014 65.726 21.068 65.762 ;
               RECT 21.014 65.955 21.068 65.991 ;
               RECT 21.014 66.249 21.068 66.285 ;
               RECT 21.014 66.478 21.068 66.514 ;
               RECT 21.014 66.926 21.068 66.962 ;
               RECT 21.014 67.155 21.068 67.191 ;
               RECT 21.014 67.449 21.068 67.485 ;
               RECT 21.014 67.678 21.068 67.714 ;
               RECT 21.014 68.126 21.068 68.162 ;
               RECT 21.014 68.355 21.068 68.391 ;
               RECT 21.014 68.649 21.068 68.685 ;
               RECT 21.014 68.878 21.068 68.914 ;
               RECT 21.014 69.326 21.068 69.362 ;
               RECT 21.014 69.555 21.068 69.591 ;
               RECT 21.014 69.849 21.068 69.885 ;
               RECT 21.014 70.078 21.068 70.114 ;
               RECT 21.014 70.526 21.068 70.562 ;
               RECT 21.014 70.755 21.068 70.791 ;
               RECT 21.014 71.049 21.068 71.085 ;
               RECT 21.014 71.278 21.068 71.314 ;
               RECT 21.014 71.726 21.068 71.762 ;
               RECT 21.014 71.955 21.068 71.991 ;
               RECT 21.014 72.249 21.068 72.285 ;
               RECT 21.014 72.478 21.068 72.514 ;
               RECT 21.014 72.926 21.068 72.962 ;
               RECT 21.014 73.155 21.068 73.191 ;
               RECT 21.014 73.449 21.068 73.485 ;
               RECT 21.014 73.678 21.068 73.714 ;
               RECT 21.014 74.126 21.068 74.162 ;
               RECT 21.014 74.355 21.068 74.391 ;
               RECT 21.014 74.649 21.068 74.685 ;
               RECT 21.014 74.878 21.068 74.914 ;
               RECT 21.014 75.326 21.068 75.362 ;
               RECT 21.014 75.555 21.068 75.591 ;
               RECT 21.014 75.849 21.068 75.885 ;
               RECT 21.014 76.078 21.068 76.114 ;
               RECT 21.014 76.526 21.068 76.562 ;
               RECT 21.014 76.755 21.068 76.791 ;
               RECT 21.014 77.049 21.068 77.085 ;
               RECT 21.014 77.278 21.068 77.314 ;
               RECT 21.014 77.726 21.068 77.762 ;
               RECT 21.014 77.955 21.068 77.991 ;
               RECT 21.014 78.249 21.068 78.285 ;
               RECT 21.014 78.478 21.068 78.514 ;
               RECT 21.014 78.926 21.068 78.962 ;
               RECT 21.014 79.155 21.068 79.191 ;
               RECT 21.014 79.449 21.068 79.485 ;
               RECT 21.014 79.678 21.068 79.714 ;
               RECT 21.014 80.126 21.068 80.162 ;
               RECT 21.014 80.355 21.068 80.391 ;
               RECT 21.014 80.649 21.068 80.685 ;
               RECT 21.014 80.878 21.068 80.914 ;
               RECT 21.014 81.326 21.068 81.362 ;
               RECT 21.014 81.555 21.068 81.591 ;
               RECT 21.014 81.849 21.068 81.885 ;
               RECT 21.014 82.078 21.068 82.114 ;
               RECT 21.014 82.526 21.068 82.562 ;
               RECT 21.014 82.755 21.068 82.791 ;
               RECT 21.014 83.049 21.068 83.085 ;
               RECT 21.014 83.278 21.068 83.314 ;
               RECT 21.014 83.726 21.068 83.762 ;
               RECT 21.014 83.955 21.068 83.991 ;
               RECT 21.014 84.249 21.068 84.285 ;
               RECT 21.014 84.478 21.068 84.514 ;
               RECT 21.014 84.926 21.068 84.962 ;
               RECT 21.014 85.155 21.068 85.191 ;
               RECT 21.014 85.449 21.068 85.485 ;
               RECT 21.014 85.678 21.068 85.714 ;
               RECT 21.014 86.126 21.068 86.162 ;
               RECT 21.014 86.355 21.068 86.391 ;
               RECT 21.014 86.649 21.068 86.685 ;
               RECT 21.014 86.878 21.068 86.914 ;
               RECT 21.014 87.326 21.068 87.362 ;
               RECT 21.014 87.555 21.068 87.591 ;
               RECT 21.014 87.849 21.068 87.885 ;
               RECT 21.014 88.078 21.068 88.114 ;
               RECT 21.014 88.526 21.068 88.562 ;
               RECT 21.014 88.755 21.068 88.791 ;
               RECT 21.014 89.049 21.068 89.085 ;
               RECT 21.014 89.278 21.068 89.314 ;
               RECT 21.014 89.726 21.068 89.762 ;
               RECT 21.014 89.955 21.068 89.991 ;
               RECT 21.014 90.249 21.068 90.285 ;
               RECT 21.014 90.478 21.068 90.514 ;
               RECT 21.014 90.926 21.068 90.962 ;
               RECT 21.014 91.155 21.068 91.191 ;
               RECT 21.014 91.449 21.068 91.485 ;
               RECT 21.014 91.678 21.068 91.714 ;
               RECT 21.014 92.126 21.068 92.162 ;
               RECT 21.014 92.355 21.068 92.391 ;
               RECT 21.014 92.649 21.068 92.685 ;
               RECT 21.014 92.878 21.068 92.914 ;
               RECT 21.014 93.326 21.068 93.362 ;
               RECT 21.014 93.555 21.068 93.591 ;
               RECT 21.014 93.849 21.068 93.885 ;
               RECT 21.014 94.078 21.068 94.114 ;
               RECT 21.014 94.526 21.068 94.562 ;
               RECT 21.014 94.755 21.068 94.791 ;
               RECT 21.014 95.049 21.068 95.085 ;
               RECT 21.014 95.278 21.068 95.314 ;
               RECT 21.014 95.726 21.068 95.762 ;
               RECT 21.014 95.955 21.068 95.991 ;
               RECT 21.014 96.249 21.068 96.285 ;
               RECT 21.014 96.478 21.068 96.514 ;
               RECT 21.014 96.926 21.068 96.962 ;
               RECT 21.014 97.155 21.068 97.191 ;
               RECT 21.014 97.449 21.068 97.485 ;
               RECT 21.014 97.678 21.068 97.714 ;
               RECT 21.014 98.126 21.068 98.162 ;
               RECT 21.014 98.355 21.068 98.391 ;
               RECT 21.014 98.649 21.068 98.685 ;
               RECT 21.014 98.878 21.068 98.914 ;
               RECT 21.014 99.326 21.068 99.362 ;
               RECT 21.014 99.555 21.068 99.591 ;
               RECT 21.014 99.849 21.068 99.885 ;
               RECT 21.014 100.078 21.068 100.114 ;
               RECT 21.014 100.526 21.068 100.562 ;
               RECT 21.014 100.755 21.068 100.791 ;
               RECT 21.014 101.049 21.068 101.085 ;
               RECT 21.014 101.278 21.068 101.314 ;
               RECT 21.014 101.726 21.068 101.762 ;
               RECT 21.014 101.955 21.068 101.991 ;
               RECT 21.014 102.249 21.068 102.285 ;
               RECT 21.014 102.478 21.068 102.514 ;
               RECT 21.014 102.926 21.068 102.962 ;
               RECT 21.014 103.155 21.068 103.191 ;
               RECT 21.014 103.449 21.068 103.485 ;
               RECT 21.014 103.678 21.068 103.714 ;
               RECT 21.014 104.126 21.068 104.162 ;
               RECT 21.014 104.355 21.068 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 21.65 0.5695 21.704 104.5505 ;
               LAYER v4 ;
               RECT 21.65 0.958 21.704 0.994 ;
               RECT 21.65 1.406 21.704 1.442 ;
               RECT 21.65 1.635 21.704 1.671 ;
               RECT 21.65 2.158 21.704 2.194 ;
               RECT 21.65 2.606 21.704 2.642 ;
               RECT 21.65 2.835 21.704 2.871 ;
               RECT 21.65 3.358 21.704 3.394 ;
               RECT 21.65 3.806 21.704 3.842 ;
               RECT 21.65 4.035 21.704 4.071 ;
               RECT 21.65 4.558 21.704 4.594 ;
               RECT 21.65 5.006 21.704 5.042 ;
               RECT 21.65 5.235 21.704 5.271 ;
               RECT 21.65 5.758 21.704 5.794 ;
               RECT 21.65 6.206 21.704 6.242 ;
               RECT 21.65 6.435 21.704 6.471 ;
               RECT 21.65 6.958 21.704 6.994 ;
               RECT 21.65 7.406 21.704 7.442 ;
               RECT 21.65 7.635 21.704 7.671 ;
               RECT 21.65 8.158 21.704 8.194 ;
               RECT 21.65 8.606 21.704 8.642 ;
               RECT 21.65 8.835 21.704 8.871 ;
               RECT 21.65 9.358 21.704 9.394 ;
               RECT 21.65 9.806 21.704 9.842 ;
               RECT 21.65 10.035 21.704 10.071 ;
               RECT 21.65 10.558 21.704 10.594 ;
               RECT 21.65 11.006 21.704 11.042 ;
               RECT 21.65 11.235 21.704 11.271 ;
               RECT 21.65 11.758 21.704 11.794 ;
               RECT 21.65 12.206 21.704 12.242 ;
               RECT 21.65 12.435 21.704 12.471 ;
               RECT 21.65 12.958 21.704 12.994 ;
               RECT 21.65 13.406 21.704 13.442 ;
               RECT 21.65 13.635 21.704 13.671 ;
               RECT 21.65 14.158 21.704 14.194 ;
               RECT 21.65 14.606 21.704 14.642 ;
               RECT 21.65 14.835 21.704 14.871 ;
               RECT 21.65 15.358 21.704 15.394 ;
               RECT 21.65 15.806 21.704 15.842 ;
               RECT 21.65 16.035 21.704 16.071 ;
               RECT 21.65 16.558 21.704 16.594 ;
               RECT 21.65 17.006 21.704 17.042 ;
               RECT 21.65 17.235 21.704 17.271 ;
               RECT 21.65 17.758 21.704 17.794 ;
               RECT 21.65 18.206 21.704 18.242 ;
               RECT 21.65 18.435 21.704 18.471 ;
               RECT 21.65 18.958 21.704 18.994 ;
               RECT 21.65 19.406 21.704 19.442 ;
               RECT 21.65 19.635 21.704 19.671 ;
               RECT 21.65 20.158 21.704 20.194 ;
               RECT 21.65 20.606 21.704 20.642 ;
               RECT 21.65 20.835 21.704 20.871 ;
               RECT 21.65 21.358 21.704 21.394 ;
               RECT 21.65 21.806 21.704 21.842 ;
               RECT 21.65 22.035 21.704 22.071 ;
               RECT 21.65 22.558 21.704 22.594 ;
               RECT 21.65 23.006 21.704 23.042 ;
               RECT 21.65 23.235 21.704 23.271 ;
               RECT 21.65 23.758 21.704 23.794 ;
               RECT 21.65 24.206 21.704 24.242 ;
               RECT 21.65 24.435 21.704 24.471 ;
               RECT 21.65 24.958 21.704 24.994 ;
               RECT 21.65 25.406 21.704 25.442 ;
               RECT 21.65 25.635 21.704 25.671 ;
               RECT 21.65 26.158 21.704 26.194 ;
               RECT 21.65 26.606 21.704 26.642 ;
               RECT 21.65 26.835 21.704 26.871 ;
               RECT 21.65 27.358 21.704 27.394 ;
               RECT 21.65 27.806 21.704 27.842 ;
               RECT 21.65 28.035 21.704 28.071 ;
               RECT 21.65 28.558 21.704 28.594 ;
               RECT 21.65 29.006 21.704 29.042 ;
               RECT 21.65 29.235 21.704 29.271 ;
               RECT 21.65 29.758 21.704 29.794 ;
               RECT 21.65 30.206 21.704 30.242 ;
               RECT 21.65 30.435 21.704 30.471 ;
               RECT 21.65 30.958 21.704 30.994 ;
               RECT 21.65 31.406 21.704 31.442 ;
               RECT 21.65 31.635 21.704 31.671 ;
               RECT 21.65 32.158 21.704 32.194 ;
               RECT 21.65 32.606 21.704 32.642 ;
               RECT 21.65 32.835 21.704 32.871 ;
               RECT 21.65 33.358 21.704 33.394 ;
               RECT 21.65 33.806 21.704 33.842 ;
               RECT 21.65 34.035 21.704 34.071 ;
               RECT 21.65 34.558 21.704 34.594 ;
               RECT 21.65 35.006 21.704 35.042 ;
               RECT 21.65 35.235 21.704 35.271 ;
               RECT 21.65 35.758 21.704 35.794 ;
               RECT 21.65 36.206 21.704 36.242 ;
               RECT 21.65 36.435 21.704 36.471 ;
               RECT 21.65 36.958 21.704 36.994 ;
               RECT 21.65 37.406 21.704 37.442 ;
               RECT 21.65 37.635 21.704 37.671 ;
               RECT 21.65 38.158 21.704 38.194 ;
               RECT 21.65 38.606 21.704 38.642 ;
               RECT 21.65 38.835 21.704 38.871 ;
               RECT 21.65 39.358 21.704 39.394 ;
               RECT 21.65 39.806 21.704 39.842 ;
               RECT 21.65 40.035 21.704 40.071 ;
               RECT 21.65 40.558 21.704 40.594 ;
               RECT 21.65 41.006 21.704 41.042 ;
               RECT 21.65 41.235 21.704 41.271 ;
               RECT 21.65 41.758 21.704 41.794 ;
               RECT 21.65 42.206 21.704 42.242 ;
               RECT 21.65 42.435 21.704 42.471 ;
               RECT 21.65 42.958 21.704 42.994 ;
               RECT 21.65 43.406 21.704 43.442 ;
               RECT 21.65 43.635 21.704 43.671 ;
               RECT 21.65 44.158 21.704 44.194 ;
               RECT 21.65 44.606 21.704 44.642 ;
               RECT 21.65 44.835 21.704 44.871 ;
               RECT 21.65 45.358 21.704 45.394 ;
               RECT 21.65 45.806 21.704 45.842 ;
               RECT 21.65 46.035 21.704 46.071 ;
               RECT 21.65 46.558 21.704 46.594 ;
               RECT 21.65 47.006 21.704 47.042 ;
               RECT 21.65 47.235 21.704 47.271 ;
               RECT 21.65 47.758 21.704 47.794 ;
               RECT 21.65 48.206 21.704 48.242 ;
               RECT 21.65 48.435 21.704 48.471 ;
               RECT 21.65 49.062 21.704 49.098 ;
               RECT 21.65 49.1875 21.704 49.2125 ;
               RECT 21.65 49.542 21.704 49.578 ;
               RECT 21.65 49.662 21.704 49.698 ;
               RECT 21.65 49.782 21.704 49.818 ;
               RECT 21.65 50.142 21.704 50.178 ;
               RECT 21.65 50.262 21.704 50.298 ;
               RECT 21.65 50.622 21.704 50.658 ;
               RECT 21.65 51.102 21.704 51.138 ;
               RECT 21.65 51.582 21.704 51.618 ;
               RECT 21.65 52.062 21.704 52.098 ;
               RECT 21.65 52.182 21.704 52.218 ;
               RECT 21.65 52.542 21.704 52.578 ;
               RECT 21.65 52.902 21.704 52.938 ;
               RECT 21.65 53.022 21.704 53.058 ;
               RECT 21.65 53.5075 21.704 53.5325 ;
               RECT 21.65 53.9875 21.704 54.0125 ;
               RECT 21.65 54.462 21.704 54.498 ;
               RECT 21.65 54.822 21.704 54.858 ;
               RECT 21.65 54.942 21.704 54.978 ;
               RECT 21.65 55.302 21.704 55.338 ;
               RECT 21.65 55.4275 21.704 55.4525 ;
               RECT 21.65 55.542 21.704 55.578 ;
               RECT 21.65 55.902 21.704 55.938 ;
               RECT 21.65 56.878 21.704 56.914 ;
               RECT 21.65 57.326 21.704 57.362 ;
               RECT 21.65 57.555 21.704 57.591 ;
               RECT 21.65 58.078 21.704 58.114 ;
               RECT 21.65 58.526 21.704 58.562 ;
               RECT 21.65 58.755 21.704 58.791 ;
               RECT 21.65 59.278 21.704 59.314 ;
               RECT 21.65 59.726 21.704 59.762 ;
               RECT 21.65 59.955 21.704 59.991 ;
               RECT 21.65 60.478 21.704 60.514 ;
               RECT 21.65 60.926 21.704 60.962 ;
               RECT 21.65 61.155 21.704 61.191 ;
               RECT 21.65 61.678 21.704 61.714 ;
               RECT 21.65 62.126 21.704 62.162 ;
               RECT 21.65 62.355 21.704 62.391 ;
               RECT 21.65 62.878 21.704 62.914 ;
               RECT 21.65 63.326 21.704 63.362 ;
               RECT 21.65 63.555 21.704 63.591 ;
               RECT 21.65 64.078 21.704 64.114 ;
               RECT 21.65 64.526 21.704 64.562 ;
               RECT 21.65 64.755 21.704 64.791 ;
               RECT 21.65 65.278 21.704 65.314 ;
               RECT 21.65 65.726 21.704 65.762 ;
               RECT 21.65 65.955 21.704 65.991 ;
               RECT 21.65 66.478 21.704 66.514 ;
               RECT 21.65 66.926 21.704 66.962 ;
               RECT 21.65 67.155 21.704 67.191 ;
               RECT 21.65 67.678 21.704 67.714 ;
               RECT 21.65 68.126 21.704 68.162 ;
               RECT 21.65 68.355 21.704 68.391 ;
               RECT 21.65 68.878 21.704 68.914 ;
               RECT 21.65 69.326 21.704 69.362 ;
               RECT 21.65 69.555 21.704 69.591 ;
               RECT 21.65 70.078 21.704 70.114 ;
               RECT 21.65 70.526 21.704 70.562 ;
               RECT 21.65 70.755 21.704 70.791 ;
               RECT 21.65 71.278 21.704 71.314 ;
               RECT 21.65 71.726 21.704 71.762 ;
               RECT 21.65 71.955 21.704 71.991 ;
               RECT 21.65 72.478 21.704 72.514 ;
               RECT 21.65 72.926 21.704 72.962 ;
               RECT 21.65 73.155 21.704 73.191 ;
               RECT 21.65 73.678 21.704 73.714 ;
               RECT 21.65 74.126 21.704 74.162 ;
               RECT 21.65 74.355 21.704 74.391 ;
               RECT 21.65 74.878 21.704 74.914 ;
               RECT 21.65 75.326 21.704 75.362 ;
               RECT 21.65 75.555 21.704 75.591 ;
               RECT 21.65 76.078 21.704 76.114 ;
               RECT 21.65 76.526 21.704 76.562 ;
               RECT 21.65 76.755 21.704 76.791 ;
               RECT 21.65 77.278 21.704 77.314 ;
               RECT 21.65 77.726 21.704 77.762 ;
               RECT 21.65 77.955 21.704 77.991 ;
               RECT 21.65 78.478 21.704 78.514 ;
               RECT 21.65 78.926 21.704 78.962 ;
               RECT 21.65 79.155 21.704 79.191 ;
               RECT 21.65 79.678 21.704 79.714 ;
               RECT 21.65 80.126 21.704 80.162 ;
               RECT 21.65 80.355 21.704 80.391 ;
               RECT 21.65 80.878 21.704 80.914 ;
               RECT 21.65 81.326 21.704 81.362 ;
               RECT 21.65 81.555 21.704 81.591 ;
               RECT 21.65 82.078 21.704 82.114 ;
               RECT 21.65 82.526 21.704 82.562 ;
               RECT 21.65 82.755 21.704 82.791 ;
               RECT 21.65 83.278 21.704 83.314 ;
               RECT 21.65 83.726 21.704 83.762 ;
               RECT 21.65 83.955 21.704 83.991 ;
               RECT 21.65 84.478 21.704 84.514 ;
               RECT 21.65 84.926 21.704 84.962 ;
               RECT 21.65 85.155 21.704 85.191 ;
               RECT 21.65 85.678 21.704 85.714 ;
               RECT 21.65 86.126 21.704 86.162 ;
               RECT 21.65 86.355 21.704 86.391 ;
               RECT 21.65 86.878 21.704 86.914 ;
               RECT 21.65 87.326 21.704 87.362 ;
               RECT 21.65 87.555 21.704 87.591 ;
               RECT 21.65 88.078 21.704 88.114 ;
               RECT 21.65 88.526 21.704 88.562 ;
               RECT 21.65 88.755 21.704 88.791 ;
               RECT 21.65 89.278 21.704 89.314 ;
               RECT 21.65 89.726 21.704 89.762 ;
               RECT 21.65 89.955 21.704 89.991 ;
               RECT 21.65 90.478 21.704 90.514 ;
               RECT 21.65 90.926 21.704 90.962 ;
               RECT 21.65 91.155 21.704 91.191 ;
               RECT 21.65 91.678 21.704 91.714 ;
               RECT 21.65 92.126 21.704 92.162 ;
               RECT 21.65 92.355 21.704 92.391 ;
               RECT 21.65 92.878 21.704 92.914 ;
               RECT 21.65 93.326 21.704 93.362 ;
               RECT 21.65 93.555 21.704 93.591 ;
               RECT 21.65 94.078 21.704 94.114 ;
               RECT 21.65 94.526 21.704 94.562 ;
               RECT 21.65 94.755 21.704 94.791 ;
               RECT 21.65 95.278 21.704 95.314 ;
               RECT 21.65 95.726 21.704 95.762 ;
               RECT 21.65 95.955 21.704 95.991 ;
               RECT 21.65 96.478 21.704 96.514 ;
               RECT 21.65 96.926 21.704 96.962 ;
               RECT 21.65 97.155 21.704 97.191 ;
               RECT 21.65 97.678 21.704 97.714 ;
               RECT 21.65 98.126 21.704 98.162 ;
               RECT 21.65 98.355 21.704 98.391 ;
               RECT 21.65 98.878 21.704 98.914 ;
               RECT 21.65 99.326 21.704 99.362 ;
               RECT 21.65 99.555 21.704 99.591 ;
               RECT 21.65 100.078 21.704 100.114 ;
               RECT 21.65 100.526 21.704 100.562 ;
               RECT 21.65 100.755 21.704 100.791 ;
               RECT 21.65 101.278 21.704 101.314 ;
               RECT 21.65 101.726 21.704 101.762 ;
               RECT 21.65 101.955 21.704 101.991 ;
               RECT 21.65 102.478 21.704 102.514 ;
               RECT 21.65 102.926 21.704 102.962 ;
               RECT 21.65 103.155 21.704 103.191 ;
               RECT 21.65 103.678 21.704 103.714 ;
               RECT 21.65 104.126 21.704 104.162 ;
               RECT 21.65 104.355 21.704 104.391 ;
          END
          PORT
               LAYER m5 ;
               RECT 21.896 0.5695 21.95 104.5505 ;
               LAYER v4 ;
               RECT 21.896 0.729 21.95 0.765 ;
               RECT 21.896 0.958 21.95 0.994 ;
               RECT 21.896 1.406 21.95 1.442 ;
               RECT 21.896 1.929 21.95 1.965 ;
               RECT 21.896 2.158 21.95 2.194 ;
               RECT 21.896 2.606 21.95 2.642 ;
               RECT 21.896 3.129 21.95 3.165 ;
               RECT 21.896 3.358 21.95 3.394 ;
               RECT 21.896 3.806 21.95 3.842 ;
               RECT 21.896 4.329 21.95 4.365 ;
               RECT 21.896 4.558 21.95 4.594 ;
               RECT 21.896 5.006 21.95 5.042 ;
               RECT 21.896 5.529 21.95 5.565 ;
               RECT 21.896 5.758 21.95 5.794 ;
               RECT 21.896 6.206 21.95 6.242 ;
               RECT 21.896 6.729 21.95 6.765 ;
               RECT 21.896 6.958 21.95 6.994 ;
               RECT 21.896 7.406 21.95 7.442 ;
               RECT 21.896 7.929 21.95 7.965 ;
               RECT 21.896 8.158 21.95 8.194 ;
               RECT 21.896 8.606 21.95 8.642 ;
               RECT 21.896 9.129 21.95 9.165 ;
               RECT 21.896 9.358 21.95 9.394 ;
               RECT 21.896 9.806 21.95 9.842 ;
               RECT 21.896 10.329 21.95 10.365 ;
               RECT 21.896 10.558 21.95 10.594 ;
               RECT 21.896 11.006 21.95 11.042 ;
               RECT 21.896 11.529 21.95 11.565 ;
               RECT 21.896 11.758 21.95 11.794 ;
               RECT 21.896 12.206 21.95 12.242 ;
               RECT 21.896 12.729 21.95 12.765 ;
               RECT 21.896 12.958 21.95 12.994 ;
               RECT 21.896 13.406 21.95 13.442 ;
               RECT 21.896 13.929 21.95 13.965 ;
               RECT 21.896 14.158 21.95 14.194 ;
               RECT 21.896 14.606 21.95 14.642 ;
               RECT 21.896 15.129 21.95 15.165 ;
               RECT 21.896 15.358 21.95 15.394 ;
               RECT 21.896 15.806 21.95 15.842 ;
               RECT 21.896 16.329 21.95 16.365 ;
               RECT 21.896 16.558 21.95 16.594 ;
               RECT 21.896 17.006 21.95 17.042 ;
               RECT 21.896 17.529 21.95 17.565 ;
               RECT 21.896 17.758 21.95 17.794 ;
               RECT 21.896 18.206 21.95 18.242 ;
               RECT 21.896 18.729 21.95 18.765 ;
               RECT 21.896 18.958 21.95 18.994 ;
               RECT 21.896 19.406 21.95 19.442 ;
               RECT 21.896 19.929 21.95 19.965 ;
               RECT 21.896 20.158 21.95 20.194 ;
               RECT 21.896 20.606 21.95 20.642 ;
               RECT 21.896 21.129 21.95 21.165 ;
               RECT 21.896 21.358 21.95 21.394 ;
               RECT 21.896 21.806 21.95 21.842 ;
               RECT 21.896 22.329 21.95 22.365 ;
               RECT 21.896 22.558 21.95 22.594 ;
               RECT 21.896 23.006 21.95 23.042 ;
               RECT 21.896 23.529 21.95 23.565 ;
               RECT 21.896 23.758 21.95 23.794 ;
               RECT 21.896 24.206 21.95 24.242 ;
               RECT 21.896 24.729 21.95 24.765 ;
               RECT 21.896 24.958 21.95 24.994 ;
               RECT 21.896 25.406 21.95 25.442 ;
               RECT 21.896 25.929 21.95 25.965 ;
               RECT 21.896 26.158 21.95 26.194 ;
               RECT 21.896 26.606 21.95 26.642 ;
               RECT 21.896 27.129 21.95 27.165 ;
               RECT 21.896 27.358 21.95 27.394 ;
               RECT 21.896 27.806 21.95 27.842 ;
               RECT 21.896 28.329 21.95 28.365 ;
               RECT 21.896 28.558 21.95 28.594 ;
               RECT 21.896 29.006 21.95 29.042 ;
               RECT 21.896 29.529 21.95 29.565 ;
               RECT 21.896 29.758 21.95 29.794 ;
               RECT 21.896 30.206 21.95 30.242 ;
               RECT 21.896 30.729 21.95 30.765 ;
               RECT 21.896 30.958 21.95 30.994 ;
               RECT 21.896 31.406 21.95 31.442 ;
               RECT 21.896 31.929 21.95 31.965 ;
               RECT 21.896 32.158 21.95 32.194 ;
               RECT 21.896 32.606 21.95 32.642 ;
               RECT 21.896 33.129 21.95 33.165 ;
               RECT 21.896 33.358 21.95 33.394 ;
               RECT 21.896 33.806 21.95 33.842 ;
               RECT 21.896 34.329 21.95 34.365 ;
               RECT 21.896 34.558 21.95 34.594 ;
               RECT 21.896 35.006 21.95 35.042 ;
               RECT 21.896 35.529 21.95 35.565 ;
               RECT 21.896 35.758 21.95 35.794 ;
               RECT 21.896 36.206 21.95 36.242 ;
               RECT 21.896 36.729 21.95 36.765 ;
               RECT 21.896 36.958 21.95 36.994 ;
               RECT 21.896 37.406 21.95 37.442 ;
               RECT 21.896 37.929 21.95 37.965 ;
               RECT 21.896 38.158 21.95 38.194 ;
               RECT 21.896 38.606 21.95 38.642 ;
               RECT 21.896 39.129 21.95 39.165 ;
               RECT 21.896 39.358 21.95 39.394 ;
               RECT 21.896 39.806 21.95 39.842 ;
               RECT 21.896 40.329 21.95 40.365 ;
               RECT 21.896 40.558 21.95 40.594 ;
               RECT 21.896 41.006 21.95 41.042 ;
               RECT 21.896 41.529 21.95 41.565 ;
               RECT 21.896 41.758 21.95 41.794 ;
               RECT 21.896 42.206 21.95 42.242 ;
               RECT 21.896 42.729 21.95 42.765 ;
               RECT 21.896 42.958 21.95 42.994 ;
               RECT 21.896 43.406 21.95 43.442 ;
               RECT 21.896 43.929 21.95 43.965 ;
               RECT 21.896 44.158 21.95 44.194 ;
               RECT 21.896 44.606 21.95 44.642 ;
               RECT 21.896 45.129 21.95 45.165 ;
               RECT 21.896 45.358 21.95 45.394 ;
               RECT 21.896 45.806 21.95 45.842 ;
               RECT 21.896 46.329 21.95 46.365 ;
               RECT 21.896 46.558 21.95 46.594 ;
               RECT 21.896 47.006 21.95 47.042 ;
               RECT 21.896 47.529 21.95 47.565 ;
               RECT 21.896 47.758 21.95 47.794 ;
               RECT 21.896 48.206 21.95 48.242 ;
               RECT 21.896 49.062 21.95 49.098 ;
               RECT 21.896 49.182 21.95 49.218 ;
               RECT 21.896 49.542 21.95 49.578 ;
               RECT 21.896 49.662 21.95 49.698 ;
               RECT 21.896 49.782 21.95 49.818 ;
               RECT 21.896 50.142 21.95 50.178 ;
               RECT 21.896 50.262 21.95 50.298 ;
               RECT 21.896 50.622 21.95 50.658 ;
               RECT 21.896 51.5875 21.95 51.6125 ;
               RECT 21.896 52.062 21.95 52.098 ;
               RECT 21.896 52.182 21.95 52.218 ;
               RECT 21.896 52.542 21.95 52.578 ;
               RECT 21.896 52.902 21.95 52.938 ;
               RECT 21.896 53.022 21.95 53.058 ;
               RECT 21.896 53.502 21.95 53.538 ;
               RECT 21.896 53.9875 21.95 54.0125 ;
               RECT 21.896 54.462 21.95 54.498 ;
               RECT 21.896 54.822 21.95 54.858 ;
               RECT 21.896 54.942 21.95 54.978 ;
               RECT 21.896 55.302 21.95 55.338 ;
               RECT 21.896 55.422 21.95 55.458 ;
               RECT 21.896 55.542 21.95 55.578 ;
               RECT 21.896 55.902 21.95 55.938 ;
               RECT 21.896 56.649 21.95 56.685 ;
               RECT 21.896 56.878 21.95 56.914 ;
               RECT 21.896 57.326 21.95 57.362 ;
               RECT 21.896 57.849 21.95 57.885 ;
               RECT 21.896 58.078 21.95 58.114 ;
               RECT 21.896 58.526 21.95 58.562 ;
               RECT 21.896 59.049 21.95 59.085 ;
               RECT 21.896 59.278 21.95 59.314 ;
               RECT 21.896 59.726 21.95 59.762 ;
               RECT 21.896 60.249 21.95 60.285 ;
               RECT 21.896 60.478 21.95 60.514 ;
               RECT 21.896 60.926 21.95 60.962 ;
               RECT 21.896 61.449 21.95 61.485 ;
               RECT 21.896 61.678 21.95 61.714 ;
               RECT 21.896 62.126 21.95 62.162 ;
               RECT 21.896 62.649 21.95 62.685 ;
               RECT 21.896 62.878 21.95 62.914 ;
               RECT 21.896 63.326 21.95 63.362 ;
               RECT 21.896 63.849 21.95 63.885 ;
               RECT 21.896 64.078 21.95 64.114 ;
               RECT 21.896 64.526 21.95 64.562 ;
               RECT 21.896 65.049 21.95 65.085 ;
               RECT 21.896 65.278 21.95 65.314 ;
               RECT 21.896 65.726 21.95 65.762 ;
               RECT 21.896 66.249 21.95 66.285 ;
               RECT 21.896 66.478 21.95 66.514 ;
               RECT 21.896 66.926 21.95 66.962 ;
               RECT 21.896 67.449 21.95 67.485 ;
               RECT 21.896 67.678 21.95 67.714 ;
               RECT 21.896 68.126 21.95 68.162 ;
               RECT 21.896 68.649 21.95 68.685 ;
               RECT 21.896 68.878 21.95 68.914 ;
               RECT 21.896 69.326 21.95 69.362 ;
               RECT 21.896 69.849 21.95 69.885 ;
               RECT 21.896 70.078 21.95 70.114 ;
               RECT 21.896 70.526 21.95 70.562 ;
               RECT 21.896 71.049 21.95 71.085 ;
               RECT 21.896 71.278 21.95 71.314 ;
               RECT 21.896 71.726 21.95 71.762 ;
               RECT 21.896 72.249 21.95 72.285 ;
               RECT 21.896 72.478 21.95 72.514 ;
               RECT 21.896 72.926 21.95 72.962 ;
               RECT 21.896 73.449 21.95 73.485 ;
               RECT 21.896 73.678 21.95 73.714 ;
               RECT 21.896 74.126 21.95 74.162 ;
               RECT 21.896 74.649 21.95 74.685 ;
               RECT 21.896 74.878 21.95 74.914 ;
               RECT 21.896 75.326 21.95 75.362 ;
               RECT 21.896 75.849 21.95 75.885 ;
               RECT 21.896 76.078 21.95 76.114 ;
               RECT 21.896 76.526 21.95 76.562 ;
               RECT 21.896 77.049 21.95 77.085 ;
               RECT 21.896 77.278 21.95 77.314 ;
               RECT 21.896 77.726 21.95 77.762 ;
               RECT 21.896 78.249 21.95 78.285 ;
               RECT 21.896 78.478 21.95 78.514 ;
               RECT 21.896 78.926 21.95 78.962 ;
               RECT 21.896 79.449 21.95 79.485 ;
               RECT 21.896 79.678 21.95 79.714 ;
               RECT 21.896 80.126 21.95 80.162 ;
               RECT 21.896 80.649 21.95 80.685 ;
               RECT 21.896 80.878 21.95 80.914 ;
               RECT 21.896 81.326 21.95 81.362 ;
               RECT 21.896 81.849 21.95 81.885 ;
               RECT 21.896 82.078 21.95 82.114 ;
               RECT 21.896 82.526 21.95 82.562 ;
               RECT 21.896 83.049 21.95 83.085 ;
               RECT 21.896 83.278 21.95 83.314 ;
               RECT 21.896 83.726 21.95 83.762 ;
               RECT 21.896 84.249 21.95 84.285 ;
               RECT 21.896 84.478 21.95 84.514 ;
               RECT 21.896 84.926 21.95 84.962 ;
               RECT 21.896 85.449 21.95 85.485 ;
               RECT 21.896 85.678 21.95 85.714 ;
               RECT 21.896 86.126 21.95 86.162 ;
               RECT 21.896 86.649 21.95 86.685 ;
               RECT 21.896 86.878 21.95 86.914 ;
               RECT 21.896 87.326 21.95 87.362 ;
               RECT 21.896 87.849 21.95 87.885 ;
               RECT 21.896 88.078 21.95 88.114 ;
               RECT 21.896 88.526 21.95 88.562 ;
               RECT 21.896 89.049 21.95 89.085 ;
               RECT 21.896 89.278 21.95 89.314 ;
               RECT 21.896 89.726 21.95 89.762 ;
               RECT 21.896 90.249 21.95 90.285 ;
               RECT 21.896 90.478 21.95 90.514 ;
               RECT 21.896 90.926 21.95 90.962 ;
               RECT 21.896 91.449 21.95 91.485 ;
               RECT 21.896 91.678 21.95 91.714 ;
               RECT 21.896 92.126 21.95 92.162 ;
               RECT 21.896 92.649 21.95 92.685 ;
               RECT 21.896 92.878 21.95 92.914 ;
               RECT 21.896 93.326 21.95 93.362 ;
               RECT 21.896 93.849 21.95 93.885 ;
               RECT 21.896 94.078 21.95 94.114 ;
               RECT 21.896 94.526 21.95 94.562 ;
               RECT 21.896 95.049 21.95 95.085 ;
               RECT 21.896 95.278 21.95 95.314 ;
               RECT 21.896 95.726 21.95 95.762 ;
               RECT 21.896 96.249 21.95 96.285 ;
               RECT 21.896 96.478 21.95 96.514 ;
               RECT 21.896 96.926 21.95 96.962 ;
               RECT 21.896 97.449 21.95 97.485 ;
               RECT 21.896 97.678 21.95 97.714 ;
               RECT 21.896 98.126 21.95 98.162 ;
               RECT 21.896 98.649 21.95 98.685 ;
               RECT 21.896 98.878 21.95 98.914 ;
               RECT 21.896 99.326 21.95 99.362 ;
               RECT 21.896 99.849 21.95 99.885 ;
               RECT 21.896 100.078 21.95 100.114 ;
               RECT 21.896 100.526 21.95 100.562 ;
               RECT 21.896 101.049 21.95 101.085 ;
               RECT 21.896 101.278 21.95 101.314 ;
               RECT 21.896 101.726 21.95 101.762 ;
               RECT 21.896 102.249 21.95 102.285 ;
               RECT 21.896 102.478 21.95 102.514 ;
               RECT 21.896 102.926 21.95 102.962 ;
               RECT 21.896 103.449 21.95 103.485 ;
               RECT 21.896 103.678 21.95 103.714 ;
               RECT 21.896 104.126 21.95 104.162 ;
          END
          PORT
               LAYER m5 ;
               RECT 22.854 49.7505 22.906 55.3695 ;
               LAYER v4 ;
               RECT 22.854 49.782 22.906 49.818 ;
               RECT 22.854 50.262 22.906 50.298 ;
               RECT 22.854 50.502 22.906 50.538 ;
               RECT 22.854 50.982 22.906 51.018 ;
               RECT 22.854 51.102 22.906 51.138 ;
               RECT 22.854 51.582 22.906 51.618 ;
               RECT 22.854 52.062 22.906 52.098 ;
               RECT 22.854 52.182 22.906 52.218 ;
               RECT 22.854 52.542 22.906 52.578 ;
               RECT 22.854 52.662 22.906 52.698 ;
               RECT 22.854 52.902 22.906 52.938 ;
               RECT 22.854 53.022 22.906 53.058 ;
               RECT 22.854 53.502 22.906 53.538 ;
               RECT 22.854 53.982 22.906 54.018 ;
               RECT 22.854 54.102 22.906 54.138 ;
               RECT 22.854 54.582 22.906 54.618 ;
               RECT 22.854 54.822 22.906 54.858 ;
               RECT 22.854 55.302 22.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 23.174 0.6 23.226 104.52 ;
               LAYER v4 ;
               RECT 23.174 49.542 23.226 49.578 ;
               RECT 23.174 49.782 23.226 49.818 ;
               RECT 23.174 50.262 23.226 50.298 ;
               RECT 23.174 50.502 23.226 50.538 ;
               RECT 23.174 50.982 23.226 51.018 ;
               RECT 23.174 51.102 23.226 51.138 ;
               RECT 23.174 51.582 23.226 51.618 ;
               RECT 23.174 52.062 23.226 52.098 ;
               RECT 23.174 52.182 23.226 52.218 ;
               RECT 23.174 52.542 23.226 52.578 ;
               RECT 23.174 52.662 23.226 52.698 ;
               RECT 23.174 52.902 23.226 52.938 ;
               RECT 23.174 53.502 23.226 53.538 ;
               RECT 23.174 53.982 23.226 54.018 ;
               RECT 23.174 54.102 23.226 54.138 ;
               RECT 23.174 54.582 23.226 54.618 ;
               RECT 23.174 54.822 23.226 54.858 ;
               RECT 23.174 55.302 23.226 55.338 ;
               RECT 23.174 55.542 23.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 23.654 49.7505 23.706 55.3695 ;
               LAYER v4 ;
               RECT 23.654 49.782 23.706 49.818 ;
               RECT 23.654 50.262 23.706 50.298 ;
               RECT 23.654 50.502 23.706 50.538 ;
               RECT 23.654 50.982 23.706 51.018 ;
               RECT 23.654 51.102 23.706 51.138 ;
               RECT 23.654 51.582 23.706 51.618 ;
               RECT 23.654 52.062 23.706 52.098 ;
               RECT 23.654 52.182 23.706 52.218 ;
               RECT 23.654 52.542 23.706 52.578 ;
               RECT 23.654 52.662 23.706 52.698 ;
               RECT 23.654 52.902 23.706 52.938 ;
               RECT 23.654 53.022 23.706 53.058 ;
               RECT 23.654 53.502 23.706 53.538 ;
               RECT 23.654 53.982 23.706 54.018 ;
               RECT 23.654 54.102 23.706 54.138 ;
               RECT 23.654 54.582 23.706 54.618 ;
               RECT 23.654 54.822 23.706 54.858 ;
               RECT 23.654 55.302 23.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 23.974 0.6 24.026 104.52 ;
               LAYER v4 ;
               RECT 23.974 49.542 24.026 49.578 ;
               RECT 23.974 49.782 24.026 49.818 ;
               RECT 23.974 50.262 24.026 50.298 ;
               RECT 23.974 50.502 24.026 50.538 ;
               RECT 23.974 50.982 24.026 51.018 ;
               RECT 23.974 51.102 24.026 51.138 ;
               RECT 23.974 51.582 24.026 51.618 ;
               RECT 23.974 52.062 24.026 52.098 ;
               RECT 23.974 52.182 24.026 52.218 ;
               RECT 23.974 52.542 24.026 52.578 ;
               RECT 23.974 52.662 24.026 52.698 ;
               RECT 23.974 52.902 24.026 52.938 ;
               RECT 23.974 53.502 24.026 53.538 ;
               RECT 23.974 53.982 24.026 54.018 ;
               RECT 23.974 54.102 24.026 54.138 ;
               RECT 23.974 54.582 24.026 54.618 ;
               RECT 23.974 54.822 24.026 54.858 ;
               RECT 23.974 55.302 24.026 55.338 ;
               RECT 23.974 55.542 24.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 24.454 49.7505 24.506 55.3695 ;
               LAYER v4 ;
               RECT 24.454 49.782 24.506 49.818 ;
               RECT 24.454 50.262 24.506 50.298 ;
               RECT 24.454 50.502 24.506 50.538 ;
               RECT 24.454 50.982 24.506 51.018 ;
               RECT 24.454 51.102 24.506 51.138 ;
               RECT 24.454 51.582 24.506 51.618 ;
               RECT 24.454 52.062 24.506 52.098 ;
               RECT 24.454 52.182 24.506 52.218 ;
               RECT 24.454 52.542 24.506 52.578 ;
               RECT 24.454 52.662 24.506 52.698 ;
               RECT 24.454 52.902 24.506 52.938 ;
               RECT 24.454 53.022 24.506 53.058 ;
               RECT 24.454 53.502 24.506 53.538 ;
               RECT 24.454 53.982 24.506 54.018 ;
               RECT 24.454 54.102 24.506 54.138 ;
               RECT 24.454 54.582 24.506 54.618 ;
               RECT 24.454 54.822 24.506 54.858 ;
               RECT 24.454 55.302 24.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 24.774 0.6 24.826 104.52 ;
               LAYER v4 ;
               RECT 24.774 49.542 24.826 49.578 ;
               RECT 24.774 49.782 24.826 49.818 ;
               RECT 24.774 50.262 24.826 50.298 ;
               RECT 24.774 50.502 24.826 50.538 ;
               RECT 24.774 50.982 24.826 51.018 ;
               RECT 24.774 51.102 24.826 51.138 ;
               RECT 24.774 51.582 24.826 51.618 ;
               RECT 24.774 52.062 24.826 52.098 ;
               RECT 24.774 52.182 24.826 52.218 ;
               RECT 24.774 52.542 24.826 52.578 ;
               RECT 24.774 52.662 24.826 52.698 ;
               RECT 24.774 52.902 24.826 52.938 ;
               RECT 24.774 53.502 24.826 53.538 ;
               RECT 24.774 53.982 24.826 54.018 ;
               RECT 24.774 54.102 24.826 54.138 ;
               RECT 24.774 54.582 24.826 54.618 ;
               RECT 24.774 54.822 24.826 54.858 ;
               RECT 24.774 55.302 24.826 55.338 ;
               RECT 24.774 55.542 24.826 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 25.254 49.7505 25.306 55.3695 ;
               LAYER v4 ;
               RECT 25.254 49.782 25.306 49.818 ;
               RECT 25.254 50.262 25.306 50.298 ;
               RECT 25.254 50.502 25.306 50.538 ;
               RECT 25.254 50.982 25.306 51.018 ;
               RECT 25.254 51.102 25.306 51.138 ;
               RECT 25.254 51.582 25.306 51.618 ;
               RECT 25.254 52.062 25.306 52.098 ;
               RECT 25.254 52.182 25.306 52.218 ;
               RECT 25.254 52.542 25.306 52.578 ;
               RECT 25.254 52.662 25.306 52.698 ;
               RECT 25.254 52.902 25.306 52.938 ;
               RECT 25.254 53.022 25.306 53.058 ;
               RECT 25.254 53.502 25.306 53.538 ;
               RECT 25.254 53.982 25.306 54.018 ;
               RECT 25.254 54.102 25.306 54.138 ;
               RECT 25.254 54.582 25.306 54.618 ;
               RECT 25.254 54.822 25.306 54.858 ;
               RECT 25.254 55.302 25.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 25.574 0.6 25.626 104.52 ;
               LAYER v4 ;
               RECT 25.574 49.542 25.626 49.578 ;
               RECT 25.574 49.782 25.626 49.818 ;
               RECT 25.574 50.262 25.626 50.298 ;
               RECT 25.574 50.502 25.626 50.538 ;
               RECT 25.574 50.982 25.626 51.018 ;
               RECT 25.574 51.102 25.626 51.138 ;
               RECT 25.574 51.582 25.626 51.618 ;
               RECT 25.574 52.062 25.626 52.098 ;
               RECT 25.574 52.182 25.626 52.218 ;
               RECT 25.574 52.542 25.626 52.578 ;
               RECT 25.574 52.662 25.626 52.698 ;
               RECT 25.574 52.902 25.626 52.938 ;
               RECT 25.574 53.502 25.626 53.538 ;
               RECT 25.574 53.982 25.626 54.018 ;
               RECT 25.574 54.102 25.626 54.138 ;
               RECT 25.574 54.582 25.626 54.618 ;
               RECT 25.574 54.822 25.626 54.858 ;
               RECT 25.574 55.302 25.626 55.338 ;
               RECT 25.574 55.542 25.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 26.054 49.7505 26.106 55.3695 ;
               LAYER v4 ;
               RECT 26.054 49.782 26.106 49.818 ;
               RECT 26.054 50.262 26.106 50.298 ;
               RECT 26.054 50.502 26.106 50.538 ;
               RECT 26.054 50.982 26.106 51.018 ;
               RECT 26.054 51.102 26.106 51.138 ;
               RECT 26.054 51.582 26.106 51.618 ;
               RECT 26.054 52.062 26.106 52.098 ;
               RECT 26.054 52.182 26.106 52.218 ;
               RECT 26.054 52.542 26.106 52.578 ;
               RECT 26.054 52.662 26.106 52.698 ;
               RECT 26.054 52.902 26.106 52.938 ;
               RECT 26.054 53.022 26.106 53.058 ;
               RECT 26.054 53.502 26.106 53.538 ;
               RECT 26.054 53.982 26.106 54.018 ;
               RECT 26.054 54.102 26.106 54.138 ;
               RECT 26.054 54.582 26.106 54.618 ;
               RECT 26.054 54.822 26.106 54.858 ;
               RECT 26.054 55.302 26.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 26.374 0.6 26.426 104.52 ;
               LAYER v4 ;
               RECT 26.374 49.542 26.426 49.578 ;
               RECT 26.374 49.782 26.426 49.818 ;
               RECT 26.374 50.262 26.426 50.298 ;
               RECT 26.374 50.502 26.426 50.538 ;
               RECT 26.374 50.982 26.426 51.018 ;
               RECT 26.374 51.102 26.426 51.138 ;
               RECT 26.374 51.582 26.426 51.618 ;
               RECT 26.374 52.062 26.426 52.098 ;
               RECT 26.374 52.182 26.426 52.218 ;
               RECT 26.374 52.542 26.426 52.578 ;
               RECT 26.374 52.662 26.426 52.698 ;
               RECT 26.374 52.902 26.426 52.938 ;
               RECT 26.374 53.502 26.426 53.538 ;
               RECT 26.374 53.982 26.426 54.018 ;
               RECT 26.374 54.102 26.426 54.138 ;
               RECT 26.374 54.582 26.426 54.618 ;
               RECT 26.374 54.822 26.426 54.858 ;
               RECT 26.374 55.302 26.426 55.338 ;
               RECT 26.374 55.542 26.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 26.854 49.7505 26.906 55.3695 ;
               LAYER v4 ;
               RECT 26.854 49.782 26.906 49.818 ;
               RECT 26.854 50.262 26.906 50.298 ;
               RECT 26.854 50.502 26.906 50.538 ;
               RECT 26.854 50.982 26.906 51.018 ;
               RECT 26.854 51.102 26.906 51.138 ;
               RECT 26.854 51.582 26.906 51.618 ;
               RECT 26.854 52.062 26.906 52.098 ;
               RECT 26.854 52.182 26.906 52.218 ;
               RECT 26.854 52.542 26.906 52.578 ;
               RECT 26.854 52.662 26.906 52.698 ;
               RECT 26.854 52.902 26.906 52.938 ;
               RECT 26.854 53.022 26.906 53.058 ;
               RECT 26.854 53.502 26.906 53.538 ;
               RECT 26.854 53.982 26.906 54.018 ;
               RECT 26.854 54.102 26.906 54.138 ;
               RECT 26.854 54.582 26.906 54.618 ;
               RECT 26.854 54.822 26.906 54.858 ;
               RECT 26.854 55.302 26.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 27.174 0.6 27.226 104.52 ;
               LAYER v4 ;
               RECT 27.174 49.542 27.226 49.578 ;
               RECT 27.174 49.782 27.226 49.818 ;
               RECT 27.174 50.262 27.226 50.298 ;
               RECT 27.174 50.502 27.226 50.538 ;
               RECT 27.174 50.982 27.226 51.018 ;
               RECT 27.174 51.102 27.226 51.138 ;
               RECT 27.174 51.582 27.226 51.618 ;
               RECT 27.174 52.062 27.226 52.098 ;
               RECT 27.174 52.182 27.226 52.218 ;
               RECT 27.174 52.542 27.226 52.578 ;
               RECT 27.174 52.662 27.226 52.698 ;
               RECT 27.174 52.902 27.226 52.938 ;
               RECT 27.174 53.502 27.226 53.538 ;
               RECT 27.174 53.982 27.226 54.018 ;
               RECT 27.174 54.102 27.226 54.138 ;
               RECT 27.174 54.582 27.226 54.618 ;
               RECT 27.174 54.822 27.226 54.858 ;
               RECT 27.174 55.302 27.226 55.338 ;
               RECT 27.174 55.542 27.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 27.654 49.7505 27.706 55.3695 ;
               LAYER v4 ;
               RECT 27.654 49.782 27.706 49.818 ;
               RECT 27.654 50.262 27.706 50.298 ;
               RECT 27.654 50.502 27.706 50.538 ;
               RECT 27.654 50.982 27.706 51.018 ;
               RECT 27.654 51.102 27.706 51.138 ;
               RECT 27.654 51.582 27.706 51.618 ;
               RECT 27.654 52.062 27.706 52.098 ;
               RECT 27.654 52.182 27.706 52.218 ;
               RECT 27.654 52.542 27.706 52.578 ;
               RECT 27.654 52.662 27.706 52.698 ;
               RECT 27.654 52.902 27.706 52.938 ;
               RECT 27.654 53.022 27.706 53.058 ;
               RECT 27.654 53.502 27.706 53.538 ;
               RECT 27.654 53.982 27.706 54.018 ;
               RECT 27.654 54.102 27.706 54.138 ;
               RECT 27.654 54.582 27.706 54.618 ;
               RECT 27.654 54.822 27.706 54.858 ;
               RECT 27.654 55.302 27.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 27.974 0.6 28.026 104.52 ;
               LAYER v4 ;
               RECT 27.974 49.542 28.026 49.578 ;
               RECT 27.974 49.782 28.026 49.818 ;
               RECT 27.974 50.262 28.026 50.298 ;
               RECT 27.974 50.502 28.026 50.538 ;
               RECT 27.974 50.982 28.026 51.018 ;
               RECT 27.974 51.102 28.026 51.138 ;
               RECT 27.974 51.582 28.026 51.618 ;
               RECT 27.974 52.062 28.026 52.098 ;
               RECT 27.974 52.182 28.026 52.218 ;
               RECT 27.974 52.542 28.026 52.578 ;
               RECT 27.974 52.662 28.026 52.698 ;
               RECT 27.974 52.902 28.026 52.938 ;
               RECT 27.974 53.502 28.026 53.538 ;
               RECT 27.974 53.982 28.026 54.018 ;
               RECT 27.974 54.102 28.026 54.138 ;
               RECT 27.974 54.582 28.026 54.618 ;
               RECT 27.974 54.822 28.026 54.858 ;
               RECT 27.974 55.302 28.026 55.338 ;
               RECT 27.974 55.542 28.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 28.454 49.7505 28.506 55.3695 ;
               LAYER v4 ;
               RECT 28.454 49.782 28.506 49.818 ;
               RECT 28.454 50.262 28.506 50.298 ;
               RECT 28.454 50.502 28.506 50.538 ;
               RECT 28.454 50.982 28.506 51.018 ;
               RECT 28.454 51.102 28.506 51.138 ;
               RECT 28.454 51.582 28.506 51.618 ;
               RECT 28.454 52.062 28.506 52.098 ;
               RECT 28.454 52.182 28.506 52.218 ;
               RECT 28.454 52.542 28.506 52.578 ;
               RECT 28.454 52.662 28.506 52.698 ;
               RECT 28.454 52.902 28.506 52.938 ;
               RECT 28.454 53.022 28.506 53.058 ;
               RECT 28.454 53.502 28.506 53.538 ;
               RECT 28.454 53.982 28.506 54.018 ;
               RECT 28.454 54.102 28.506 54.138 ;
               RECT 28.454 54.582 28.506 54.618 ;
               RECT 28.454 54.822 28.506 54.858 ;
               RECT 28.454 55.302 28.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 28.774 0.6 28.826 104.52 ;
               LAYER v4 ;
               RECT 28.774 49.542 28.826 49.578 ;
               RECT 28.774 49.782 28.826 49.818 ;
               RECT 28.774 50.262 28.826 50.298 ;
               RECT 28.774 50.502 28.826 50.538 ;
               RECT 28.774 50.982 28.826 51.018 ;
               RECT 28.774 51.102 28.826 51.138 ;
               RECT 28.774 51.582 28.826 51.618 ;
               RECT 28.774 52.062 28.826 52.098 ;
               RECT 28.774 52.182 28.826 52.218 ;
               RECT 28.774 52.542 28.826 52.578 ;
               RECT 28.774 52.662 28.826 52.698 ;
               RECT 28.774 52.902 28.826 52.938 ;
               RECT 28.774 53.502 28.826 53.538 ;
               RECT 28.774 53.982 28.826 54.018 ;
               RECT 28.774 54.102 28.826 54.138 ;
               RECT 28.774 54.582 28.826 54.618 ;
               RECT 28.774 54.822 28.826 54.858 ;
               RECT 28.774 55.302 28.826 55.338 ;
               RECT 28.774 55.542 28.826 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 29.254 49.7505 29.306 55.3695 ;
               LAYER v4 ;
               RECT 29.254 49.782 29.306 49.818 ;
               RECT 29.254 50.262 29.306 50.298 ;
               RECT 29.254 50.502 29.306 50.538 ;
               RECT 29.254 50.982 29.306 51.018 ;
               RECT 29.254 51.102 29.306 51.138 ;
               RECT 29.254 51.582 29.306 51.618 ;
               RECT 29.254 52.062 29.306 52.098 ;
               RECT 29.254 52.182 29.306 52.218 ;
               RECT 29.254 52.542 29.306 52.578 ;
               RECT 29.254 52.662 29.306 52.698 ;
               RECT 29.254 52.902 29.306 52.938 ;
               RECT 29.254 53.022 29.306 53.058 ;
               RECT 29.254 53.502 29.306 53.538 ;
               RECT 29.254 53.982 29.306 54.018 ;
               RECT 29.254 54.102 29.306 54.138 ;
               RECT 29.254 54.582 29.306 54.618 ;
               RECT 29.254 54.822 29.306 54.858 ;
               RECT 29.254 55.302 29.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 29.574 0.6 29.626 104.52 ;
               LAYER v4 ;
               RECT 29.574 49.542 29.626 49.578 ;
               RECT 29.574 49.782 29.626 49.818 ;
               RECT 29.574 50.262 29.626 50.298 ;
               RECT 29.574 50.502 29.626 50.538 ;
               RECT 29.574 50.982 29.626 51.018 ;
               RECT 29.574 51.102 29.626 51.138 ;
               RECT 29.574 51.582 29.626 51.618 ;
               RECT 29.574 52.062 29.626 52.098 ;
               RECT 29.574 52.182 29.626 52.218 ;
               RECT 29.574 52.542 29.626 52.578 ;
               RECT 29.574 52.662 29.626 52.698 ;
               RECT 29.574 52.902 29.626 52.938 ;
               RECT 29.574 53.502 29.626 53.538 ;
               RECT 29.574 53.982 29.626 54.018 ;
               RECT 29.574 54.102 29.626 54.138 ;
               RECT 29.574 54.582 29.626 54.618 ;
               RECT 29.574 54.822 29.626 54.858 ;
               RECT 29.574 55.302 29.626 55.338 ;
               RECT 29.574 55.542 29.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 3.054 49.7505 3.106 55.3695 ;
               LAYER v4 ;
               RECT 3.054 49.782 3.106 49.818 ;
               RECT 3.054 50.262 3.106 50.298 ;
               RECT 3.054 50.502 3.106 50.538 ;
               RECT 3.054 50.982 3.106 51.018 ;
               RECT 3.054 51.102 3.106 51.138 ;
               RECT 3.054 51.582 3.106 51.618 ;
               RECT 3.054 52.062 3.106 52.098 ;
               RECT 3.054 52.182 3.106 52.218 ;
               RECT 3.054 52.542 3.106 52.578 ;
               RECT 3.054 52.662 3.106 52.698 ;
               RECT 3.054 52.902 3.106 52.938 ;
               RECT 3.054 53.022 3.106 53.058 ;
               RECT 3.054 53.502 3.106 53.538 ;
               RECT 3.054 53.982 3.106 54.018 ;
               RECT 3.054 54.102 3.106 54.138 ;
               RECT 3.054 54.582 3.106 54.618 ;
               RECT 3.054 54.822 3.106 54.858 ;
               RECT 3.054 55.302 3.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 3.374 0.6 3.426 104.52 ;
               LAYER v4 ;
               RECT 3.374 49.542 3.426 49.578 ;
               RECT 3.374 49.782 3.426 49.818 ;
               RECT 3.374 50.262 3.426 50.298 ;
               RECT 3.374 50.502 3.426 50.538 ;
               RECT 3.374 50.982 3.426 51.018 ;
               RECT 3.374 51.102 3.426 51.138 ;
               RECT 3.374 51.582 3.426 51.618 ;
               RECT 3.374 52.062 3.426 52.098 ;
               RECT 3.374 52.182 3.426 52.218 ;
               RECT 3.374 52.542 3.426 52.578 ;
               RECT 3.374 52.662 3.426 52.698 ;
               RECT 3.374 52.902 3.426 52.938 ;
               RECT 3.374 53.502 3.426 53.538 ;
               RECT 3.374 53.982 3.426 54.018 ;
               RECT 3.374 54.102 3.426 54.138 ;
               RECT 3.374 54.582 3.426 54.618 ;
               RECT 3.374 54.822 3.426 54.858 ;
               RECT 3.374 55.302 3.426 55.338 ;
               RECT 3.374 55.542 3.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 3.854 49.7505 3.906 55.3695 ;
               LAYER v4 ;
               RECT 3.854 49.782 3.906 49.818 ;
               RECT 3.854 50.262 3.906 50.298 ;
               RECT 3.854 50.502 3.906 50.538 ;
               RECT 3.854 50.982 3.906 51.018 ;
               RECT 3.854 51.102 3.906 51.138 ;
               RECT 3.854 51.582 3.906 51.618 ;
               RECT 3.854 52.062 3.906 52.098 ;
               RECT 3.854 52.182 3.906 52.218 ;
               RECT 3.854 52.542 3.906 52.578 ;
               RECT 3.854 52.662 3.906 52.698 ;
               RECT 3.854 52.902 3.906 52.938 ;
               RECT 3.854 53.022 3.906 53.058 ;
               RECT 3.854 53.502 3.906 53.538 ;
               RECT 3.854 53.982 3.906 54.018 ;
               RECT 3.854 54.102 3.906 54.138 ;
               RECT 3.854 54.582 3.906 54.618 ;
               RECT 3.854 54.822 3.906 54.858 ;
               RECT 3.854 55.302 3.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 30.054 49.7505 30.106 55.3695 ;
               LAYER v4 ;
               RECT 30.054 49.782 30.106 49.818 ;
               RECT 30.054 50.262 30.106 50.298 ;
               RECT 30.054 50.502 30.106 50.538 ;
               RECT 30.054 50.982 30.106 51.018 ;
               RECT 30.054 51.102 30.106 51.138 ;
               RECT 30.054 51.582 30.106 51.618 ;
               RECT 30.054 52.062 30.106 52.098 ;
               RECT 30.054 52.182 30.106 52.218 ;
               RECT 30.054 52.542 30.106 52.578 ;
               RECT 30.054 52.662 30.106 52.698 ;
               RECT 30.054 52.902 30.106 52.938 ;
               RECT 30.054 53.022 30.106 53.058 ;
               RECT 30.054 53.502 30.106 53.538 ;
               RECT 30.054 53.982 30.106 54.018 ;
               RECT 30.054 54.102 30.106 54.138 ;
               RECT 30.054 54.582 30.106 54.618 ;
               RECT 30.054 54.822 30.106 54.858 ;
               RECT 30.054 55.302 30.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 30.374 0.6 30.426 104.52 ;
               LAYER v4 ;
               RECT 30.374 49.542 30.426 49.578 ;
               RECT 30.374 49.782 30.426 49.818 ;
               RECT 30.374 50.262 30.426 50.298 ;
               RECT 30.374 50.502 30.426 50.538 ;
               RECT 30.374 50.982 30.426 51.018 ;
               RECT 30.374 51.102 30.426 51.138 ;
               RECT 30.374 51.582 30.426 51.618 ;
               RECT 30.374 52.062 30.426 52.098 ;
               RECT 30.374 52.182 30.426 52.218 ;
               RECT 30.374 52.542 30.426 52.578 ;
               RECT 30.374 52.662 30.426 52.698 ;
               RECT 30.374 52.902 30.426 52.938 ;
               RECT 30.374 53.502 30.426 53.538 ;
               RECT 30.374 53.982 30.426 54.018 ;
               RECT 30.374 54.102 30.426 54.138 ;
               RECT 30.374 54.582 30.426 54.618 ;
               RECT 30.374 54.822 30.426 54.858 ;
               RECT 30.374 55.302 30.426 55.338 ;
               RECT 30.374 55.542 30.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 30.854 49.7505 30.906 55.3695 ;
               LAYER v4 ;
               RECT 30.854 49.782 30.906 49.818 ;
               RECT 30.854 50.262 30.906 50.298 ;
               RECT 30.854 50.502 30.906 50.538 ;
               RECT 30.854 50.982 30.906 51.018 ;
               RECT 30.854 51.102 30.906 51.138 ;
               RECT 30.854 51.582 30.906 51.618 ;
               RECT 30.854 52.062 30.906 52.098 ;
               RECT 30.854 52.182 30.906 52.218 ;
               RECT 30.854 52.542 30.906 52.578 ;
               RECT 30.854 52.662 30.906 52.698 ;
               RECT 30.854 52.902 30.906 52.938 ;
               RECT 30.854 53.022 30.906 53.058 ;
               RECT 30.854 53.502 30.906 53.538 ;
               RECT 30.854 53.982 30.906 54.018 ;
               RECT 30.854 54.102 30.906 54.138 ;
               RECT 30.854 54.582 30.906 54.618 ;
               RECT 30.854 54.822 30.906 54.858 ;
               RECT 30.854 55.302 30.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 31.174 0.6 31.226 104.52 ;
               LAYER v4 ;
               RECT 31.174 49.542 31.226 49.578 ;
               RECT 31.174 49.782 31.226 49.818 ;
               RECT 31.174 50.262 31.226 50.298 ;
               RECT 31.174 50.502 31.226 50.538 ;
               RECT 31.174 50.982 31.226 51.018 ;
               RECT 31.174 51.102 31.226 51.138 ;
               RECT 31.174 51.582 31.226 51.618 ;
               RECT 31.174 52.062 31.226 52.098 ;
               RECT 31.174 52.182 31.226 52.218 ;
               RECT 31.174 52.542 31.226 52.578 ;
               RECT 31.174 52.662 31.226 52.698 ;
               RECT 31.174 52.902 31.226 52.938 ;
               RECT 31.174 53.502 31.226 53.538 ;
               RECT 31.174 53.982 31.226 54.018 ;
               RECT 31.174 54.102 31.226 54.138 ;
               RECT 31.174 54.582 31.226 54.618 ;
               RECT 31.174 54.822 31.226 54.858 ;
               RECT 31.174 55.302 31.226 55.338 ;
               RECT 31.174 55.542 31.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 31.654 49.7505 31.706 55.3695 ;
               LAYER v4 ;
               RECT 31.654 49.782 31.706 49.818 ;
               RECT 31.654 50.262 31.706 50.298 ;
               RECT 31.654 50.502 31.706 50.538 ;
               RECT 31.654 50.982 31.706 51.018 ;
               RECT 31.654 51.102 31.706 51.138 ;
               RECT 31.654 51.582 31.706 51.618 ;
               RECT 31.654 52.062 31.706 52.098 ;
               RECT 31.654 52.182 31.706 52.218 ;
               RECT 31.654 52.542 31.706 52.578 ;
               RECT 31.654 52.662 31.706 52.698 ;
               RECT 31.654 52.902 31.706 52.938 ;
               RECT 31.654 53.022 31.706 53.058 ;
               RECT 31.654 53.502 31.706 53.538 ;
               RECT 31.654 53.982 31.706 54.018 ;
               RECT 31.654 54.102 31.706 54.138 ;
               RECT 31.654 54.582 31.706 54.618 ;
               RECT 31.654 54.822 31.706 54.858 ;
               RECT 31.654 55.302 31.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 31.974 0.6 32.026 104.52 ;
               LAYER v4 ;
               RECT 31.974 49.542 32.026 49.578 ;
               RECT 31.974 49.782 32.026 49.818 ;
               RECT 31.974 50.262 32.026 50.298 ;
               RECT 31.974 50.502 32.026 50.538 ;
               RECT 31.974 50.982 32.026 51.018 ;
               RECT 31.974 51.102 32.026 51.138 ;
               RECT 31.974 51.582 32.026 51.618 ;
               RECT 31.974 52.062 32.026 52.098 ;
               RECT 31.974 52.182 32.026 52.218 ;
               RECT 31.974 52.542 32.026 52.578 ;
               RECT 31.974 52.662 32.026 52.698 ;
               RECT 31.974 52.902 32.026 52.938 ;
               RECT 31.974 53.502 32.026 53.538 ;
               RECT 31.974 53.982 32.026 54.018 ;
               RECT 31.974 54.102 32.026 54.138 ;
               RECT 31.974 54.582 32.026 54.618 ;
               RECT 31.974 54.822 32.026 54.858 ;
               RECT 31.974 55.302 32.026 55.338 ;
               RECT 31.974 55.542 32.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 32.454 49.7505 32.506 55.3695 ;
               LAYER v4 ;
               RECT 32.454 49.782 32.506 49.818 ;
               RECT 32.454 50.262 32.506 50.298 ;
               RECT 32.454 50.502 32.506 50.538 ;
               RECT 32.454 50.982 32.506 51.018 ;
               RECT 32.454 51.102 32.506 51.138 ;
               RECT 32.454 51.582 32.506 51.618 ;
               RECT 32.454 52.062 32.506 52.098 ;
               RECT 32.454 52.182 32.506 52.218 ;
               RECT 32.454 52.542 32.506 52.578 ;
               RECT 32.454 52.662 32.506 52.698 ;
               RECT 32.454 52.902 32.506 52.938 ;
               RECT 32.454 53.022 32.506 53.058 ;
               RECT 32.454 53.502 32.506 53.538 ;
               RECT 32.454 53.982 32.506 54.018 ;
               RECT 32.454 54.102 32.506 54.138 ;
               RECT 32.454 54.582 32.506 54.618 ;
               RECT 32.454 54.822 32.506 54.858 ;
               RECT 32.454 55.302 32.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 32.774 0.6 32.826 104.52 ;
               LAYER v4 ;
               RECT 32.774 49.542 32.826 49.578 ;
               RECT 32.774 49.782 32.826 49.818 ;
               RECT 32.774 50.262 32.826 50.298 ;
               RECT 32.774 50.502 32.826 50.538 ;
               RECT 32.774 50.982 32.826 51.018 ;
               RECT 32.774 51.102 32.826 51.138 ;
               RECT 32.774 51.582 32.826 51.618 ;
               RECT 32.774 52.062 32.826 52.098 ;
               RECT 32.774 52.182 32.826 52.218 ;
               RECT 32.774 52.542 32.826 52.578 ;
               RECT 32.774 52.662 32.826 52.698 ;
               RECT 32.774 52.902 32.826 52.938 ;
               RECT 32.774 53.502 32.826 53.538 ;
               RECT 32.774 53.982 32.826 54.018 ;
               RECT 32.774 54.102 32.826 54.138 ;
               RECT 32.774 54.582 32.826 54.618 ;
               RECT 32.774 54.822 32.826 54.858 ;
               RECT 32.774 55.302 32.826 55.338 ;
               RECT 32.774 55.542 32.826 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 33.254 49.7505 33.306 55.3695 ;
               LAYER v4 ;
               RECT 33.254 49.782 33.306 49.818 ;
               RECT 33.254 50.262 33.306 50.298 ;
               RECT 33.254 50.502 33.306 50.538 ;
               RECT 33.254 50.982 33.306 51.018 ;
               RECT 33.254 51.102 33.306 51.138 ;
               RECT 33.254 51.582 33.306 51.618 ;
               RECT 33.254 52.062 33.306 52.098 ;
               RECT 33.254 52.182 33.306 52.218 ;
               RECT 33.254 52.542 33.306 52.578 ;
               RECT 33.254 52.662 33.306 52.698 ;
               RECT 33.254 52.902 33.306 52.938 ;
               RECT 33.254 53.022 33.306 53.058 ;
               RECT 33.254 53.502 33.306 53.538 ;
               RECT 33.254 53.982 33.306 54.018 ;
               RECT 33.254 54.102 33.306 54.138 ;
               RECT 33.254 54.582 33.306 54.618 ;
               RECT 33.254 54.822 33.306 54.858 ;
               RECT 33.254 55.302 33.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 33.574 0.6 33.626 104.52 ;
               LAYER v4 ;
               RECT 33.574 49.542 33.626 49.578 ;
               RECT 33.574 49.782 33.626 49.818 ;
               RECT 33.574 50.262 33.626 50.298 ;
               RECT 33.574 50.502 33.626 50.538 ;
               RECT 33.574 50.982 33.626 51.018 ;
               RECT 33.574 51.102 33.626 51.138 ;
               RECT 33.574 51.582 33.626 51.618 ;
               RECT 33.574 52.062 33.626 52.098 ;
               RECT 33.574 52.182 33.626 52.218 ;
               RECT 33.574 52.542 33.626 52.578 ;
               RECT 33.574 52.662 33.626 52.698 ;
               RECT 33.574 52.902 33.626 52.938 ;
               RECT 33.574 53.502 33.626 53.538 ;
               RECT 33.574 53.982 33.626 54.018 ;
               RECT 33.574 54.102 33.626 54.138 ;
               RECT 33.574 54.582 33.626 54.618 ;
               RECT 33.574 54.822 33.626 54.858 ;
               RECT 33.574 55.302 33.626 55.338 ;
               RECT 33.574 55.542 33.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 34.054 49.7505 34.106 55.3695 ;
               LAYER v4 ;
               RECT 34.054 49.782 34.106 49.818 ;
               RECT 34.054 50.262 34.106 50.298 ;
               RECT 34.054 50.502 34.106 50.538 ;
               RECT 34.054 50.982 34.106 51.018 ;
               RECT 34.054 51.102 34.106 51.138 ;
               RECT 34.054 51.582 34.106 51.618 ;
               RECT 34.054 52.062 34.106 52.098 ;
               RECT 34.054 52.182 34.106 52.218 ;
               RECT 34.054 52.542 34.106 52.578 ;
               RECT 34.054 52.662 34.106 52.698 ;
               RECT 34.054 52.902 34.106 52.938 ;
               RECT 34.054 53.022 34.106 53.058 ;
               RECT 34.054 53.502 34.106 53.538 ;
               RECT 34.054 53.982 34.106 54.018 ;
               RECT 34.054 54.102 34.106 54.138 ;
               RECT 34.054 54.582 34.106 54.618 ;
               RECT 34.054 54.822 34.106 54.858 ;
               RECT 34.054 55.302 34.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 34.374 0.6 34.426 104.52 ;
               LAYER v4 ;
               RECT 34.374 49.542 34.426 49.578 ;
               RECT 34.374 49.782 34.426 49.818 ;
               RECT 34.374 50.262 34.426 50.298 ;
               RECT 34.374 50.502 34.426 50.538 ;
               RECT 34.374 50.982 34.426 51.018 ;
               RECT 34.374 51.102 34.426 51.138 ;
               RECT 34.374 51.582 34.426 51.618 ;
               RECT 34.374 52.062 34.426 52.098 ;
               RECT 34.374 52.182 34.426 52.218 ;
               RECT 34.374 52.542 34.426 52.578 ;
               RECT 34.374 52.662 34.426 52.698 ;
               RECT 34.374 52.902 34.426 52.938 ;
               RECT 34.374 53.502 34.426 53.538 ;
               RECT 34.374 53.982 34.426 54.018 ;
               RECT 34.374 54.102 34.426 54.138 ;
               RECT 34.374 54.582 34.426 54.618 ;
               RECT 34.374 54.822 34.426 54.858 ;
               RECT 34.374 55.302 34.426 55.338 ;
               RECT 34.374 55.542 34.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 34.854 49.7505 34.906 55.3695 ;
               LAYER v4 ;
               RECT 34.854 49.782 34.906 49.818 ;
               RECT 34.854 50.262 34.906 50.298 ;
               RECT 34.854 50.502 34.906 50.538 ;
               RECT 34.854 50.982 34.906 51.018 ;
               RECT 34.854 51.102 34.906 51.138 ;
               RECT 34.854 51.582 34.906 51.618 ;
               RECT 34.854 52.062 34.906 52.098 ;
               RECT 34.854 52.182 34.906 52.218 ;
               RECT 34.854 52.542 34.906 52.578 ;
               RECT 34.854 52.662 34.906 52.698 ;
               RECT 34.854 52.902 34.906 52.938 ;
               RECT 34.854 53.022 34.906 53.058 ;
               RECT 34.854 53.502 34.906 53.538 ;
               RECT 34.854 53.982 34.906 54.018 ;
               RECT 34.854 54.102 34.906 54.138 ;
               RECT 34.854 54.582 34.906 54.618 ;
               RECT 34.854 54.822 34.906 54.858 ;
               RECT 34.854 55.302 34.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 35.174 0.6 35.226 104.52 ;
               LAYER v4 ;
               RECT 35.174 49.542 35.226 49.578 ;
               RECT 35.174 49.782 35.226 49.818 ;
               RECT 35.174 50.262 35.226 50.298 ;
               RECT 35.174 50.502 35.226 50.538 ;
               RECT 35.174 50.982 35.226 51.018 ;
               RECT 35.174 51.102 35.226 51.138 ;
               RECT 35.174 51.582 35.226 51.618 ;
               RECT 35.174 52.062 35.226 52.098 ;
               RECT 35.174 52.182 35.226 52.218 ;
               RECT 35.174 52.542 35.226 52.578 ;
               RECT 35.174 52.662 35.226 52.698 ;
               RECT 35.174 52.902 35.226 52.938 ;
               RECT 35.174 53.502 35.226 53.538 ;
               RECT 35.174 53.982 35.226 54.018 ;
               RECT 35.174 54.102 35.226 54.138 ;
               RECT 35.174 54.582 35.226 54.618 ;
               RECT 35.174 54.822 35.226 54.858 ;
               RECT 35.174 55.302 35.226 55.338 ;
               RECT 35.174 55.542 35.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 4.174 0.6 4.226 104.52 ;
               LAYER v4 ;
               RECT 4.174 49.542 4.226 49.578 ;
               RECT 4.174 49.782 4.226 49.818 ;
               RECT 4.174 50.262 4.226 50.298 ;
               RECT 4.174 50.502 4.226 50.538 ;
               RECT 4.174 50.982 4.226 51.018 ;
               RECT 4.174 51.102 4.226 51.138 ;
               RECT 4.174 51.582 4.226 51.618 ;
               RECT 4.174 52.062 4.226 52.098 ;
               RECT 4.174 52.182 4.226 52.218 ;
               RECT 4.174 52.542 4.226 52.578 ;
               RECT 4.174 52.662 4.226 52.698 ;
               RECT 4.174 52.902 4.226 52.938 ;
               RECT 4.174 53.502 4.226 53.538 ;
               RECT 4.174 53.982 4.226 54.018 ;
               RECT 4.174 54.102 4.226 54.138 ;
               RECT 4.174 54.582 4.226 54.618 ;
               RECT 4.174 54.822 4.226 54.858 ;
               RECT 4.174 55.302 4.226 55.338 ;
               RECT 4.174 55.542 4.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 4.654 49.7505 4.706 55.3695 ;
               LAYER v4 ;
               RECT 4.654 49.782 4.706 49.818 ;
               RECT 4.654 50.262 4.706 50.298 ;
               RECT 4.654 50.502 4.706 50.538 ;
               RECT 4.654 50.982 4.706 51.018 ;
               RECT 4.654 51.102 4.706 51.138 ;
               RECT 4.654 51.582 4.706 51.618 ;
               RECT 4.654 52.062 4.706 52.098 ;
               RECT 4.654 52.182 4.706 52.218 ;
               RECT 4.654 52.542 4.706 52.578 ;
               RECT 4.654 52.662 4.706 52.698 ;
               RECT 4.654 52.902 4.706 52.938 ;
               RECT 4.654 53.022 4.706 53.058 ;
               RECT 4.654 53.502 4.706 53.538 ;
               RECT 4.654 53.982 4.706 54.018 ;
               RECT 4.654 54.102 4.706 54.138 ;
               RECT 4.654 54.582 4.706 54.618 ;
               RECT 4.654 54.822 4.706 54.858 ;
               RECT 4.654 55.302 4.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 4.974 0.6 5.026 104.52 ;
               LAYER v4 ;
               RECT 4.974 49.542 5.026 49.578 ;
               RECT 4.974 49.782 5.026 49.818 ;
               RECT 4.974 50.262 5.026 50.298 ;
               RECT 4.974 50.502 5.026 50.538 ;
               RECT 4.974 50.982 5.026 51.018 ;
               RECT 4.974 51.102 5.026 51.138 ;
               RECT 4.974 51.582 5.026 51.618 ;
               RECT 4.974 52.062 5.026 52.098 ;
               RECT 4.974 52.182 5.026 52.218 ;
               RECT 4.974 52.542 5.026 52.578 ;
               RECT 4.974 52.662 5.026 52.698 ;
               RECT 4.974 52.902 5.026 52.938 ;
               RECT 4.974 53.502 5.026 53.538 ;
               RECT 4.974 53.982 5.026 54.018 ;
               RECT 4.974 54.102 5.026 54.138 ;
               RECT 4.974 54.582 5.026 54.618 ;
               RECT 4.974 54.822 5.026 54.858 ;
               RECT 4.974 55.302 5.026 55.338 ;
               RECT 4.974 55.542 5.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 5.454 49.7505 5.506 55.3695 ;
               LAYER v4 ;
               RECT 5.454 49.782 5.506 49.818 ;
               RECT 5.454 50.262 5.506 50.298 ;
               RECT 5.454 50.502 5.506 50.538 ;
               RECT 5.454 50.982 5.506 51.018 ;
               RECT 5.454 51.102 5.506 51.138 ;
               RECT 5.454 51.582 5.506 51.618 ;
               RECT 5.454 52.062 5.506 52.098 ;
               RECT 5.454 52.182 5.506 52.218 ;
               RECT 5.454 52.542 5.506 52.578 ;
               RECT 5.454 52.662 5.506 52.698 ;
               RECT 5.454 52.902 5.506 52.938 ;
               RECT 5.454 53.022 5.506 53.058 ;
               RECT 5.454 53.502 5.506 53.538 ;
               RECT 5.454 53.982 5.506 54.018 ;
               RECT 5.454 54.102 5.506 54.138 ;
               RECT 5.454 54.582 5.506 54.618 ;
               RECT 5.454 54.822 5.506 54.858 ;
               RECT 5.454 55.302 5.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 5.774 0.6 5.826 104.52 ;
               LAYER v4 ;
               RECT 5.774 49.542 5.826 49.578 ;
               RECT 5.774 49.782 5.826 49.818 ;
               RECT 5.774 50.262 5.826 50.298 ;
               RECT 5.774 50.502 5.826 50.538 ;
               RECT 5.774 50.982 5.826 51.018 ;
               RECT 5.774 51.102 5.826 51.138 ;
               RECT 5.774 51.582 5.826 51.618 ;
               RECT 5.774 52.062 5.826 52.098 ;
               RECT 5.774 52.182 5.826 52.218 ;
               RECT 5.774 52.542 5.826 52.578 ;
               RECT 5.774 52.662 5.826 52.698 ;
               RECT 5.774 52.902 5.826 52.938 ;
               RECT 5.774 53.502 5.826 53.538 ;
               RECT 5.774 53.982 5.826 54.018 ;
               RECT 5.774 54.102 5.826 54.138 ;
               RECT 5.774 54.582 5.826 54.618 ;
               RECT 5.774 54.822 5.826 54.858 ;
               RECT 5.774 55.302 5.826 55.338 ;
               RECT 5.774 55.542 5.826 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 6.254 49.7505 6.306 55.3695 ;
               LAYER v4 ;
               RECT 6.254 49.782 6.306 49.818 ;
               RECT 6.254 50.262 6.306 50.298 ;
               RECT 6.254 50.502 6.306 50.538 ;
               RECT 6.254 50.982 6.306 51.018 ;
               RECT 6.254 51.102 6.306 51.138 ;
               RECT 6.254 51.582 6.306 51.618 ;
               RECT 6.254 52.062 6.306 52.098 ;
               RECT 6.254 52.182 6.306 52.218 ;
               RECT 6.254 52.542 6.306 52.578 ;
               RECT 6.254 52.662 6.306 52.698 ;
               RECT 6.254 52.902 6.306 52.938 ;
               RECT 6.254 53.022 6.306 53.058 ;
               RECT 6.254 53.502 6.306 53.538 ;
               RECT 6.254 53.982 6.306 54.018 ;
               RECT 6.254 54.102 6.306 54.138 ;
               RECT 6.254 54.582 6.306 54.618 ;
               RECT 6.254 54.822 6.306 54.858 ;
               RECT 6.254 55.302 6.306 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 6.574 0.6 6.626 104.52 ;
               LAYER v4 ;
               RECT 6.574 49.542 6.626 49.578 ;
               RECT 6.574 49.782 6.626 49.818 ;
               RECT 6.574 50.262 6.626 50.298 ;
               RECT 6.574 50.502 6.626 50.538 ;
               RECT 6.574 50.982 6.626 51.018 ;
               RECT 6.574 51.102 6.626 51.138 ;
               RECT 6.574 51.582 6.626 51.618 ;
               RECT 6.574 52.062 6.626 52.098 ;
               RECT 6.574 52.182 6.626 52.218 ;
               RECT 6.574 52.542 6.626 52.578 ;
               RECT 6.574 52.662 6.626 52.698 ;
               RECT 6.574 52.902 6.626 52.938 ;
               RECT 6.574 53.502 6.626 53.538 ;
               RECT 6.574 53.982 6.626 54.018 ;
               RECT 6.574 54.102 6.626 54.138 ;
               RECT 6.574 54.582 6.626 54.618 ;
               RECT 6.574 54.822 6.626 54.858 ;
               RECT 6.574 55.302 6.626 55.338 ;
               RECT 6.574 55.542 6.626 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 7.054 49.7505 7.106 55.3695 ;
               LAYER v4 ;
               RECT 7.054 49.782 7.106 49.818 ;
               RECT 7.054 50.262 7.106 50.298 ;
               RECT 7.054 50.502 7.106 50.538 ;
               RECT 7.054 50.982 7.106 51.018 ;
               RECT 7.054 51.102 7.106 51.138 ;
               RECT 7.054 51.582 7.106 51.618 ;
               RECT 7.054 52.062 7.106 52.098 ;
               RECT 7.054 52.182 7.106 52.218 ;
               RECT 7.054 52.542 7.106 52.578 ;
               RECT 7.054 52.662 7.106 52.698 ;
               RECT 7.054 52.902 7.106 52.938 ;
               RECT 7.054 53.022 7.106 53.058 ;
               RECT 7.054 53.502 7.106 53.538 ;
               RECT 7.054 53.982 7.106 54.018 ;
               RECT 7.054 54.102 7.106 54.138 ;
               RECT 7.054 54.582 7.106 54.618 ;
               RECT 7.054 54.822 7.106 54.858 ;
               RECT 7.054 55.302 7.106 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 7.374 0.6 7.426 104.52 ;
               LAYER v4 ;
               RECT 7.374 49.542 7.426 49.578 ;
               RECT 7.374 49.782 7.426 49.818 ;
               RECT 7.374 50.262 7.426 50.298 ;
               RECT 7.374 50.502 7.426 50.538 ;
               RECT 7.374 50.982 7.426 51.018 ;
               RECT 7.374 51.102 7.426 51.138 ;
               RECT 7.374 51.582 7.426 51.618 ;
               RECT 7.374 52.062 7.426 52.098 ;
               RECT 7.374 52.182 7.426 52.218 ;
               RECT 7.374 52.542 7.426 52.578 ;
               RECT 7.374 52.662 7.426 52.698 ;
               RECT 7.374 52.902 7.426 52.938 ;
               RECT 7.374 53.502 7.426 53.538 ;
               RECT 7.374 53.982 7.426 54.018 ;
               RECT 7.374 54.102 7.426 54.138 ;
               RECT 7.374 54.582 7.426 54.618 ;
               RECT 7.374 54.822 7.426 54.858 ;
               RECT 7.374 55.302 7.426 55.338 ;
               RECT 7.374 55.542 7.426 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 7.854 49.7505 7.906 55.3695 ;
               LAYER v4 ;
               RECT 7.854 49.782 7.906 49.818 ;
               RECT 7.854 50.262 7.906 50.298 ;
               RECT 7.854 50.502 7.906 50.538 ;
               RECT 7.854 50.982 7.906 51.018 ;
               RECT 7.854 51.102 7.906 51.138 ;
               RECT 7.854 51.582 7.906 51.618 ;
               RECT 7.854 52.062 7.906 52.098 ;
               RECT 7.854 52.182 7.906 52.218 ;
               RECT 7.854 52.542 7.906 52.578 ;
               RECT 7.854 52.662 7.906 52.698 ;
               RECT 7.854 52.902 7.906 52.938 ;
               RECT 7.854 53.022 7.906 53.058 ;
               RECT 7.854 53.502 7.906 53.538 ;
               RECT 7.854 53.982 7.906 54.018 ;
               RECT 7.854 54.102 7.906 54.138 ;
               RECT 7.854 54.582 7.906 54.618 ;
               RECT 7.854 54.822 7.906 54.858 ;
               RECT 7.854 55.302 7.906 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 8.174 0.6 8.226 104.52 ;
               LAYER v4 ;
               RECT 8.174 49.542 8.226 49.578 ;
               RECT 8.174 49.782 8.226 49.818 ;
               RECT 8.174 50.262 8.226 50.298 ;
               RECT 8.174 50.502 8.226 50.538 ;
               RECT 8.174 50.982 8.226 51.018 ;
               RECT 8.174 51.102 8.226 51.138 ;
               RECT 8.174 51.582 8.226 51.618 ;
               RECT 8.174 52.062 8.226 52.098 ;
               RECT 8.174 52.182 8.226 52.218 ;
               RECT 8.174 52.542 8.226 52.578 ;
               RECT 8.174 52.662 8.226 52.698 ;
               RECT 8.174 52.902 8.226 52.938 ;
               RECT 8.174 53.502 8.226 53.538 ;
               RECT 8.174 53.982 8.226 54.018 ;
               RECT 8.174 54.102 8.226 54.138 ;
               RECT 8.174 54.582 8.226 54.618 ;
               RECT 8.174 54.822 8.226 54.858 ;
               RECT 8.174 55.302 8.226 55.338 ;
               RECT 8.174 55.542 8.226 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 8.654 49.7505 8.706 55.3695 ;
               LAYER v4 ;
               RECT 8.654 49.782 8.706 49.818 ;
               RECT 8.654 50.262 8.706 50.298 ;
               RECT 8.654 50.502 8.706 50.538 ;
               RECT 8.654 50.982 8.706 51.018 ;
               RECT 8.654 51.102 8.706 51.138 ;
               RECT 8.654 51.582 8.706 51.618 ;
               RECT 8.654 52.062 8.706 52.098 ;
               RECT 8.654 52.182 8.706 52.218 ;
               RECT 8.654 52.542 8.706 52.578 ;
               RECT 8.654 52.662 8.706 52.698 ;
               RECT 8.654 52.902 8.706 52.938 ;
               RECT 8.654 53.022 8.706 53.058 ;
               RECT 8.654 53.502 8.706 53.538 ;
               RECT 8.654 53.982 8.706 54.018 ;
               RECT 8.654 54.102 8.706 54.138 ;
               RECT 8.654 54.582 8.706 54.618 ;
               RECT 8.654 54.822 8.706 54.858 ;
               RECT 8.654 55.302 8.706 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 8.974 0.6 9.026 104.52 ;
               LAYER v4 ;
               RECT 8.974 49.542 9.026 49.578 ;
               RECT 8.974 49.782 9.026 49.818 ;
               RECT 8.974 50.262 9.026 50.298 ;
               RECT 8.974 50.502 9.026 50.538 ;
               RECT 8.974 50.982 9.026 51.018 ;
               RECT 8.974 51.102 9.026 51.138 ;
               RECT 8.974 51.582 9.026 51.618 ;
               RECT 8.974 52.062 9.026 52.098 ;
               RECT 8.974 52.182 9.026 52.218 ;
               RECT 8.974 52.542 9.026 52.578 ;
               RECT 8.974 52.662 9.026 52.698 ;
               RECT 8.974 52.902 9.026 52.938 ;
               RECT 8.974 53.502 9.026 53.538 ;
               RECT 8.974 53.982 9.026 54.018 ;
               RECT 8.974 54.102 9.026 54.138 ;
               RECT 8.974 54.582 9.026 54.618 ;
               RECT 8.974 54.822 9.026 54.858 ;
               RECT 8.974 55.302 9.026 55.338 ;
               RECT 8.974 55.542 9.026 55.578 ;
          END
          PORT
               LAYER m5 ;
               RECT 9.454 49.7505 9.506 55.3695 ;
               LAYER v4 ;
               RECT 9.454 49.782 9.506 49.818 ;
               RECT 9.454 50.262 9.506 50.298 ;
               RECT 9.454 50.502 9.506 50.538 ;
               RECT 9.454 50.982 9.506 51.018 ;
               RECT 9.454 51.102 9.506 51.138 ;
               RECT 9.454 51.582 9.506 51.618 ;
               RECT 9.454 52.062 9.506 52.098 ;
               RECT 9.454 52.182 9.506 52.218 ;
               RECT 9.454 52.542 9.506 52.578 ;
               RECT 9.454 52.662 9.506 52.698 ;
               RECT 9.454 52.902 9.506 52.938 ;
               RECT 9.454 53.022 9.506 53.058 ;
               RECT 9.454 53.502 9.506 53.538 ;
               RECT 9.454 53.982 9.506 54.018 ;
               RECT 9.454 54.102 9.506 54.138 ;
               RECT 9.454 54.582 9.506 54.618 ;
               RECT 9.454 54.822 9.506 54.858 ;
               RECT 9.454 55.302 9.506 55.338 ;
          END
          PORT
               LAYER m5 ;
               RECT 9.774 0.6 9.826 104.52 ;
               LAYER v4 ;
               RECT 9.774 49.542 9.826 49.578 ;
               RECT 9.774 49.782 9.826 49.818 ;
               RECT 9.774 50.262 9.826 50.298 ;
               RECT 9.774 50.502 9.826 50.538 ;
               RECT 9.774 50.982 9.826 51.018 ;
               RECT 9.774 51.102 9.826 51.138 ;
               RECT 9.774 51.582 9.826 51.618 ;
               RECT 9.774 52.062 9.826 52.098 ;
               RECT 9.774 52.182 9.826 52.218 ;
               RECT 9.774 52.542 9.826 52.578 ;
               RECT 9.774 52.662 9.826 52.698 ;
               RECT 9.774 52.902 9.826 52.938 ;
               RECT 9.774 53.502 9.826 53.538 ;
               RECT 9.774 53.982 9.826 54.018 ;
               RECT 9.774 54.102 9.826 54.138 ;
               RECT 9.774 54.582 9.826 54.618 ;
               RECT 9.774 54.822 9.826 54.858 ;
               RECT 9.774 55.302 9.826 55.338 ;
               RECT 9.774 55.542 9.826 55.578 ;
          END
     END vddp
     PIN vss
     SHAPE ABUTMENT ;
     DIRECTION inout ;
          USE GROUND ;
          PORT
               LAYER m5 ;
               RECT 0.574 0.5695 0.626 104.5505 ;
               LAYER v4 ;
               RECT 0.574 0.582 0.626 0.618 ;
               RECT 0.574 1.182 0.626 1.218 ;
               RECT 0.574 1.782 0.626 1.818 ;
               RECT 0.574 2.382 0.626 2.418 ;
               RECT 0.574 2.982 0.626 3.018 ;
               RECT 0.574 3.582 0.626 3.618 ;
               RECT 0.574 4.182 0.626 4.218 ;
               RECT 0.574 4.782 0.626 4.818 ;
               RECT 0.574 5.382 0.626 5.418 ;
               RECT 0.574 5.982 0.626 6.018 ;
               RECT 0.574 6.582 0.626 6.618 ;
               RECT 0.574 7.182 0.626 7.218 ;
               RECT 0.574 7.782 0.626 7.818 ;
               RECT 0.574 8.382 0.626 8.418 ;
               RECT 0.574 8.982 0.626 9.018 ;
               RECT 0.574 9.582 0.626 9.618 ;
               RECT 0.574 10.182 0.626 10.218 ;
               RECT 0.574 10.782 0.626 10.818 ;
               RECT 0.574 11.382 0.626 11.418 ;
               RECT 0.574 11.982 0.626 12.018 ;
               RECT 0.574 12.582 0.626 12.618 ;
               RECT 0.574 13.182 0.626 13.218 ;
               RECT 0.574 13.782 0.626 13.818 ;
               RECT 0.574 14.382 0.626 14.418 ;
               RECT 0.574 14.982 0.626 15.018 ;
               RECT 0.574 15.582 0.626 15.618 ;
               RECT 0.574 16.182 0.626 16.218 ;
               RECT 0.574 16.782 0.626 16.818 ;
               RECT 0.574 17.382 0.626 17.418 ;
               RECT 0.574 17.982 0.626 18.018 ;
               RECT 0.574 18.582 0.626 18.618 ;
               RECT 0.574 19.182 0.626 19.218 ;
               RECT 0.574 19.782 0.626 19.818 ;
               RECT 0.574 20.382 0.626 20.418 ;
               RECT 0.574 20.982 0.626 21.018 ;
               RECT 0.574 21.582 0.626 21.618 ;
               RECT 0.574 22.182 0.626 22.218 ;
               RECT 0.574 22.782 0.626 22.818 ;
               RECT 0.574 23.382 0.626 23.418 ;
               RECT 0.574 23.982 0.626 24.018 ;
               RECT 0.574 24.582 0.626 24.618 ;
               RECT 0.574 25.182 0.626 25.218 ;
               RECT 0.574 25.782 0.626 25.818 ;
               RECT 0.574 26.382 0.626 26.418 ;
               RECT 0.574 26.982 0.626 27.018 ;
               RECT 0.574 27.582 0.626 27.618 ;
               RECT 0.574 28.182 0.626 28.218 ;
               RECT 0.574 28.782 0.626 28.818 ;
               RECT 0.574 29.382 0.626 29.418 ;
               RECT 0.574 29.982 0.626 30.018 ;
               RECT 0.574 30.582 0.626 30.618 ;
               RECT 0.574 31.182 0.626 31.218 ;
               RECT 0.574 31.782 0.626 31.818 ;
               RECT 0.574 32.382 0.626 32.418 ;
               RECT 0.574 32.982 0.626 33.018 ;
               RECT 0.574 33.582 0.626 33.618 ;
               RECT 0.574 34.182 0.626 34.218 ;
               RECT 0.574 34.782 0.626 34.818 ;
               RECT 0.574 35.382 0.626 35.418 ;
               RECT 0.574 35.982 0.626 36.018 ;
               RECT 0.574 36.582 0.626 36.618 ;
               RECT 0.574 37.182 0.626 37.218 ;
               RECT 0.574 37.782 0.626 37.818 ;
               RECT 0.574 38.382 0.626 38.418 ;
               RECT 0.574 38.982 0.626 39.018 ;
               RECT 0.574 39.582 0.626 39.618 ;
               RECT 0.574 40.182 0.626 40.218 ;
               RECT 0.574 40.782 0.626 40.818 ;
               RECT 0.574 41.382 0.626 41.418 ;
               RECT 0.574 41.982 0.626 42.018 ;
               RECT 0.574 42.582 0.626 42.618 ;
               RECT 0.574 43.182 0.626 43.218 ;
               RECT 0.574 43.782 0.626 43.818 ;
               RECT 0.574 44.382 0.626 44.418 ;
               RECT 0.574 44.982 0.626 45.018 ;
               RECT 0.574 45.582 0.626 45.618 ;
               RECT 0.574 46.182 0.626 46.218 ;
               RECT 0.574 46.782 0.626 46.818 ;
               RECT 0.574 47.382 0.626 47.418 ;
               RECT 0.574 47.982 0.626 48.018 ;
               RECT 0.574 48.582 0.626 48.618 ;
               RECT 0.574 48.942 0.626 48.978 ;
               RECT 0.574 49.182 0.626 49.218 ;
               RECT 0.574 49.902 0.626 49.938 ;
               RECT 0.574 50.622 0.626 50.658 ;
               RECT 0.574 50.862 0.626 50.898 ;
               RECT 0.574 51.342 0.626 51.378 ;
               RECT 0.574 51.822 0.626 51.858 ;
               RECT 0.574 52.302 0.626 52.338 ;
               RECT 0.574 52.782 0.626 52.818 ;
               RECT 0.574 53.262 0.626 53.298 ;
               RECT 0.574 53.742 0.626 53.778 ;
               RECT 0.574 54.222 0.626 54.258 ;
               RECT 0.574 54.462 0.626 54.498 ;
               RECT 0.574 55.182 0.626 55.218 ;
               RECT 0.574 55.902 0.626 55.938 ;
               RECT 0.574 56.142 0.626 56.178 ;
               RECT 0.574 56.502 0.626 56.538 ;
               RECT 0.574 57.102 0.626 57.138 ;
               RECT 0.574 57.702 0.626 57.738 ;
               RECT 0.574 58.302 0.626 58.338 ;
               RECT 0.574 58.902 0.626 58.938 ;
               RECT 0.574 59.502 0.626 59.538 ;
               RECT 0.574 60.102 0.626 60.138 ;
               RECT 0.574 60.702 0.626 60.738 ;
               RECT 0.574 61.302 0.626 61.338 ;
               RECT 0.574 61.902 0.626 61.938 ;
               RECT 0.574 62.502 0.626 62.538 ;
               RECT 0.574 63.102 0.626 63.138 ;
               RECT 0.574 63.702 0.626 63.738 ;
               RECT 0.574 64.302 0.626 64.338 ;
               RECT 0.574 64.902 0.626 64.938 ;
               RECT 0.574 65.502 0.626 65.538 ;
               RECT 0.574 66.102 0.626 66.138 ;
               RECT 0.574 66.702 0.626 66.738 ;
               RECT 0.574 67.302 0.626 67.338 ;
               RECT 0.574 67.902 0.626 67.938 ;
               RECT 0.574 68.502 0.626 68.538 ;
               RECT 0.574 69.102 0.626 69.138 ;
               RECT 0.574 69.702 0.626 69.738 ;
               RECT 0.574 70.302 0.626 70.338 ;
               RECT 0.574 70.902 0.626 70.938 ;
               RECT 0.574 71.502 0.626 71.538 ;
               RECT 0.574 72.102 0.626 72.138 ;
               RECT 0.574 72.702 0.626 72.738 ;
               RECT 0.574 73.302 0.626 73.338 ;
               RECT 0.574 73.902 0.626 73.938 ;
               RECT 0.574 74.502 0.626 74.538 ;
               RECT 0.574 75.102 0.626 75.138 ;
               RECT 0.574 75.702 0.626 75.738 ;
               RECT 0.574 76.302 0.626 76.338 ;
               RECT 0.574 76.902 0.626 76.938 ;
               RECT 0.574 77.502 0.626 77.538 ;
               RECT 0.574 78.102 0.626 78.138 ;
               RECT 0.574 78.702 0.626 78.738 ;
               RECT 0.574 79.302 0.626 79.338 ;
               RECT 0.574 79.902 0.626 79.938 ;
               RECT 0.574 80.502 0.626 80.538 ;
               RECT 0.574 81.102 0.626 81.138 ;
               RECT 0.574 81.702 0.626 81.738 ;
               RECT 0.574 82.302 0.626 82.338 ;
               RECT 0.574 82.902 0.626 82.938 ;
               RECT 0.574 83.502 0.626 83.538 ;
               RECT 0.574 84.102 0.626 84.138 ;
               RECT 0.574 84.702 0.626 84.738 ;
               RECT 0.574 85.302 0.626 85.338 ;
               RECT 0.574 85.902 0.626 85.938 ;
               RECT 0.574 86.502 0.626 86.538 ;
               RECT 0.574 87.102 0.626 87.138 ;
               RECT 0.574 87.702 0.626 87.738 ;
               RECT 0.574 88.302 0.626 88.338 ;
               RECT 0.574 88.902 0.626 88.938 ;
               RECT 0.574 89.502 0.626 89.538 ;
               RECT 0.574 90.102 0.626 90.138 ;
               RECT 0.574 90.702 0.626 90.738 ;
               RECT 0.574 91.302 0.626 91.338 ;
               RECT 0.574 91.902 0.626 91.938 ;
               RECT 0.574 92.502 0.626 92.538 ;
               RECT 0.574 93.102 0.626 93.138 ;
               RECT 0.574 93.702 0.626 93.738 ;
               RECT 0.574 94.302 0.626 94.338 ;
               RECT 0.574 94.902 0.626 94.938 ;
               RECT 0.574 95.502 0.626 95.538 ;
               RECT 0.574 96.102 0.626 96.138 ;
               RECT 0.574 96.702 0.626 96.738 ;
               RECT 0.574 97.302 0.626 97.338 ;
               RECT 0.574 97.902 0.626 97.938 ;
               RECT 0.574 98.502 0.626 98.538 ;
               RECT 0.574 99.102 0.626 99.138 ;
               RECT 0.574 99.702 0.626 99.738 ;
               RECT 0.574 100.302 0.626 100.338 ;
               RECT 0.574 100.902 0.626 100.938 ;
               RECT 0.574 101.502 0.626 101.538 ;
               RECT 0.574 102.102 0.626 102.138 ;
               RECT 0.574 102.702 0.626 102.738 ;
               RECT 0.574 103.302 0.626 103.338 ;
               RECT 0.574 103.902 0.626 103.938 ;
               RECT 0.574 104.502 0.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 1.374 0.5695 1.426 104.5505 ;
               LAYER v4 ;
               RECT 1.374 0.582 1.426 0.618 ;
               RECT 1.374 1.182 1.426 1.218 ;
               RECT 1.374 1.782 1.426 1.818 ;
               RECT 1.374 2.382 1.426 2.418 ;
               RECT 1.374 2.982 1.426 3.018 ;
               RECT 1.374 3.582 1.426 3.618 ;
               RECT 1.374 4.182 1.426 4.218 ;
               RECT 1.374 4.782 1.426 4.818 ;
               RECT 1.374 5.382 1.426 5.418 ;
               RECT 1.374 5.982 1.426 6.018 ;
               RECT 1.374 6.582 1.426 6.618 ;
               RECT 1.374 7.182 1.426 7.218 ;
               RECT 1.374 7.782 1.426 7.818 ;
               RECT 1.374 8.382 1.426 8.418 ;
               RECT 1.374 8.982 1.426 9.018 ;
               RECT 1.374 9.582 1.426 9.618 ;
               RECT 1.374 10.182 1.426 10.218 ;
               RECT 1.374 10.782 1.426 10.818 ;
               RECT 1.374 11.382 1.426 11.418 ;
               RECT 1.374 11.982 1.426 12.018 ;
               RECT 1.374 12.582 1.426 12.618 ;
               RECT 1.374 13.182 1.426 13.218 ;
               RECT 1.374 13.782 1.426 13.818 ;
               RECT 1.374 14.382 1.426 14.418 ;
               RECT 1.374 14.982 1.426 15.018 ;
               RECT 1.374 15.582 1.426 15.618 ;
               RECT 1.374 16.182 1.426 16.218 ;
               RECT 1.374 16.782 1.426 16.818 ;
               RECT 1.374 17.382 1.426 17.418 ;
               RECT 1.374 17.982 1.426 18.018 ;
               RECT 1.374 18.582 1.426 18.618 ;
               RECT 1.374 19.182 1.426 19.218 ;
               RECT 1.374 19.782 1.426 19.818 ;
               RECT 1.374 20.382 1.426 20.418 ;
               RECT 1.374 20.982 1.426 21.018 ;
               RECT 1.374 21.582 1.426 21.618 ;
               RECT 1.374 22.182 1.426 22.218 ;
               RECT 1.374 22.782 1.426 22.818 ;
               RECT 1.374 23.382 1.426 23.418 ;
               RECT 1.374 23.982 1.426 24.018 ;
               RECT 1.374 24.582 1.426 24.618 ;
               RECT 1.374 25.182 1.426 25.218 ;
               RECT 1.374 25.782 1.426 25.818 ;
               RECT 1.374 26.382 1.426 26.418 ;
               RECT 1.374 26.982 1.426 27.018 ;
               RECT 1.374 27.582 1.426 27.618 ;
               RECT 1.374 28.182 1.426 28.218 ;
               RECT 1.374 28.782 1.426 28.818 ;
               RECT 1.374 29.382 1.426 29.418 ;
               RECT 1.374 29.982 1.426 30.018 ;
               RECT 1.374 30.582 1.426 30.618 ;
               RECT 1.374 31.182 1.426 31.218 ;
               RECT 1.374 31.782 1.426 31.818 ;
               RECT 1.374 32.382 1.426 32.418 ;
               RECT 1.374 32.982 1.426 33.018 ;
               RECT 1.374 33.582 1.426 33.618 ;
               RECT 1.374 34.182 1.426 34.218 ;
               RECT 1.374 34.782 1.426 34.818 ;
               RECT 1.374 35.382 1.426 35.418 ;
               RECT 1.374 35.982 1.426 36.018 ;
               RECT 1.374 36.582 1.426 36.618 ;
               RECT 1.374 37.182 1.426 37.218 ;
               RECT 1.374 37.782 1.426 37.818 ;
               RECT 1.374 38.382 1.426 38.418 ;
               RECT 1.374 38.982 1.426 39.018 ;
               RECT 1.374 39.582 1.426 39.618 ;
               RECT 1.374 40.182 1.426 40.218 ;
               RECT 1.374 40.782 1.426 40.818 ;
               RECT 1.374 41.382 1.426 41.418 ;
               RECT 1.374 41.982 1.426 42.018 ;
               RECT 1.374 42.582 1.426 42.618 ;
               RECT 1.374 43.182 1.426 43.218 ;
               RECT 1.374 43.782 1.426 43.818 ;
               RECT 1.374 44.382 1.426 44.418 ;
               RECT 1.374 44.982 1.426 45.018 ;
               RECT 1.374 45.582 1.426 45.618 ;
               RECT 1.374 46.182 1.426 46.218 ;
               RECT 1.374 46.782 1.426 46.818 ;
               RECT 1.374 47.382 1.426 47.418 ;
               RECT 1.374 47.982 1.426 48.018 ;
               RECT 1.374 48.582 1.426 48.618 ;
               RECT 1.374 48.942 1.426 48.978 ;
               RECT 1.374 49.182 1.426 49.218 ;
               RECT 1.374 49.902 1.426 49.938 ;
               RECT 1.374 50.622 1.426 50.658 ;
               RECT 1.374 50.862 1.426 50.898 ;
               RECT 1.374 51.342 1.426 51.378 ;
               RECT 1.374 51.822 1.426 51.858 ;
               RECT 1.374 52.302 1.426 52.338 ;
               RECT 1.374 52.782 1.426 52.818 ;
               RECT 1.374 53.262 1.426 53.298 ;
               RECT 1.374 53.742 1.426 53.778 ;
               RECT 1.374 54.222 1.426 54.258 ;
               RECT 1.374 54.462 1.426 54.498 ;
               RECT 1.374 55.182 1.426 55.218 ;
               RECT 1.374 55.902 1.426 55.938 ;
               RECT 1.374 56.142 1.426 56.178 ;
               RECT 1.374 56.502 1.426 56.538 ;
               RECT 1.374 57.102 1.426 57.138 ;
               RECT 1.374 57.702 1.426 57.738 ;
               RECT 1.374 58.302 1.426 58.338 ;
               RECT 1.374 58.902 1.426 58.938 ;
               RECT 1.374 59.502 1.426 59.538 ;
               RECT 1.374 60.102 1.426 60.138 ;
               RECT 1.374 60.702 1.426 60.738 ;
               RECT 1.374 61.302 1.426 61.338 ;
               RECT 1.374 61.902 1.426 61.938 ;
               RECT 1.374 62.502 1.426 62.538 ;
               RECT 1.374 63.102 1.426 63.138 ;
               RECT 1.374 63.702 1.426 63.738 ;
               RECT 1.374 64.302 1.426 64.338 ;
               RECT 1.374 64.902 1.426 64.938 ;
               RECT 1.374 65.502 1.426 65.538 ;
               RECT 1.374 66.102 1.426 66.138 ;
               RECT 1.374 66.702 1.426 66.738 ;
               RECT 1.374 67.302 1.426 67.338 ;
               RECT 1.374 67.902 1.426 67.938 ;
               RECT 1.374 68.502 1.426 68.538 ;
               RECT 1.374 69.102 1.426 69.138 ;
               RECT 1.374 69.702 1.426 69.738 ;
               RECT 1.374 70.302 1.426 70.338 ;
               RECT 1.374 70.902 1.426 70.938 ;
               RECT 1.374 71.502 1.426 71.538 ;
               RECT 1.374 72.102 1.426 72.138 ;
               RECT 1.374 72.702 1.426 72.738 ;
               RECT 1.374 73.302 1.426 73.338 ;
               RECT 1.374 73.902 1.426 73.938 ;
               RECT 1.374 74.502 1.426 74.538 ;
               RECT 1.374 75.102 1.426 75.138 ;
               RECT 1.374 75.702 1.426 75.738 ;
               RECT 1.374 76.302 1.426 76.338 ;
               RECT 1.374 76.902 1.426 76.938 ;
               RECT 1.374 77.502 1.426 77.538 ;
               RECT 1.374 78.102 1.426 78.138 ;
               RECT 1.374 78.702 1.426 78.738 ;
               RECT 1.374 79.302 1.426 79.338 ;
               RECT 1.374 79.902 1.426 79.938 ;
               RECT 1.374 80.502 1.426 80.538 ;
               RECT 1.374 81.102 1.426 81.138 ;
               RECT 1.374 81.702 1.426 81.738 ;
               RECT 1.374 82.302 1.426 82.338 ;
               RECT 1.374 82.902 1.426 82.938 ;
               RECT 1.374 83.502 1.426 83.538 ;
               RECT 1.374 84.102 1.426 84.138 ;
               RECT 1.374 84.702 1.426 84.738 ;
               RECT 1.374 85.302 1.426 85.338 ;
               RECT 1.374 85.902 1.426 85.938 ;
               RECT 1.374 86.502 1.426 86.538 ;
               RECT 1.374 87.102 1.426 87.138 ;
               RECT 1.374 87.702 1.426 87.738 ;
               RECT 1.374 88.302 1.426 88.338 ;
               RECT 1.374 88.902 1.426 88.938 ;
               RECT 1.374 89.502 1.426 89.538 ;
               RECT 1.374 90.102 1.426 90.138 ;
               RECT 1.374 90.702 1.426 90.738 ;
               RECT 1.374 91.302 1.426 91.338 ;
               RECT 1.374 91.902 1.426 91.938 ;
               RECT 1.374 92.502 1.426 92.538 ;
               RECT 1.374 93.102 1.426 93.138 ;
               RECT 1.374 93.702 1.426 93.738 ;
               RECT 1.374 94.302 1.426 94.338 ;
               RECT 1.374 94.902 1.426 94.938 ;
               RECT 1.374 95.502 1.426 95.538 ;
               RECT 1.374 96.102 1.426 96.138 ;
               RECT 1.374 96.702 1.426 96.738 ;
               RECT 1.374 97.302 1.426 97.338 ;
               RECT 1.374 97.902 1.426 97.938 ;
               RECT 1.374 98.502 1.426 98.538 ;
               RECT 1.374 99.102 1.426 99.138 ;
               RECT 1.374 99.702 1.426 99.738 ;
               RECT 1.374 100.302 1.426 100.338 ;
               RECT 1.374 100.902 1.426 100.938 ;
               RECT 1.374 101.502 1.426 101.538 ;
               RECT 1.374 102.102 1.426 102.138 ;
               RECT 1.374 102.702 1.426 102.738 ;
               RECT 1.374 103.302 1.426 103.338 ;
               RECT 1.374 103.902 1.426 103.938 ;
               RECT 1.374 104.502 1.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 10.174 0.5695 10.226 104.5505 ;
               LAYER v4 ;
               RECT 10.174 0.582 10.226 0.618 ;
               RECT 10.174 1.182 10.226 1.218 ;
               RECT 10.174 1.782 10.226 1.818 ;
               RECT 10.174 2.382 10.226 2.418 ;
               RECT 10.174 2.982 10.226 3.018 ;
               RECT 10.174 3.582 10.226 3.618 ;
               RECT 10.174 4.182 10.226 4.218 ;
               RECT 10.174 4.782 10.226 4.818 ;
               RECT 10.174 5.382 10.226 5.418 ;
               RECT 10.174 5.982 10.226 6.018 ;
               RECT 10.174 6.582 10.226 6.618 ;
               RECT 10.174 7.182 10.226 7.218 ;
               RECT 10.174 7.782 10.226 7.818 ;
               RECT 10.174 8.382 10.226 8.418 ;
               RECT 10.174 8.982 10.226 9.018 ;
               RECT 10.174 9.582 10.226 9.618 ;
               RECT 10.174 10.182 10.226 10.218 ;
               RECT 10.174 10.782 10.226 10.818 ;
               RECT 10.174 11.382 10.226 11.418 ;
               RECT 10.174 11.982 10.226 12.018 ;
               RECT 10.174 12.582 10.226 12.618 ;
               RECT 10.174 13.182 10.226 13.218 ;
               RECT 10.174 13.782 10.226 13.818 ;
               RECT 10.174 14.382 10.226 14.418 ;
               RECT 10.174 14.982 10.226 15.018 ;
               RECT 10.174 15.582 10.226 15.618 ;
               RECT 10.174 16.182 10.226 16.218 ;
               RECT 10.174 16.782 10.226 16.818 ;
               RECT 10.174 17.382 10.226 17.418 ;
               RECT 10.174 17.982 10.226 18.018 ;
               RECT 10.174 18.582 10.226 18.618 ;
               RECT 10.174 19.182 10.226 19.218 ;
               RECT 10.174 19.782 10.226 19.818 ;
               RECT 10.174 20.382 10.226 20.418 ;
               RECT 10.174 20.982 10.226 21.018 ;
               RECT 10.174 21.582 10.226 21.618 ;
               RECT 10.174 22.182 10.226 22.218 ;
               RECT 10.174 22.782 10.226 22.818 ;
               RECT 10.174 23.382 10.226 23.418 ;
               RECT 10.174 23.982 10.226 24.018 ;
               RECT 10.174 24.582 10.226 24.618 ;
               RECT 10.174 25.182 10.226 25.218 ;
               RECT 10.174 25.782 10.226 25.818 ;
               RECT 10.174 26.382 10.226 26.418 ;
               RECT 10.174 26.982 10.226 27.018 ;
               RECT 10.174 27.582 10.226 27.618 ;
               RECT 10.174 28.182 10.226 28.218 ;
               RECT 10.174 28.782 10.226 28.818 ;
               RECT 10.174 29.382 10.226 29.418 ;
               RECT 10.174 29.982 10.226 30.018 ;
               RECT 10.174 30.582 10.226 30.618 ;
               RECT 10.174 31.182 10.226 31.218 ;
               RECT 10.174 31.782 10.226 31.818 ;
               RECT 10.174 32.382 10.226 32.418 ;
               RECT 10.174 32.982 10.226 33.018 ;
               RECT 10.174 33.582 10.226 33.618 ;
               RECT 10.174 34.182 10.226 34.218 ;
               RECT 10.174 34.782 10.226 34.818 ;
               RECT 10.174 35.382 10.226 35.418 ;
               RECT 10.174 35.982 10.226 36.018 ;
               RECT 10.174 36.582 10.226 36.618 ;
               RECT 10.174 37.182 10.226 37.218 ;
               RECT 10.174 37.782 10.226 37.818 ;
               RECT 10.174 38.382 10.226 38.418 ;
               RECT 10.174 38.982 10.226 39.018 ;
               RECT 10.174 39.582 10.226 39.618 ;
               RECT 10.174 40.182 10.226 40.218 ;
               RECT 10.174 40.782 10.226 40.818 ;
               RECT 10.174 41.382 10.226 41.418 ;
               RECT 10.174 41.982 10.226 42.018 ;
               RECT 10.174 42.582 10.226 42.618 ;
               RECT 10.174 43.182 10.226 43.218 ;
               RECT 10.174 43.782 10.226 43.818 ;
               RECT 10.174 44.382 10.226 44.418 ;
               RECT 10.174 44.982 10.226 45.018 ;
               RECT 10.174 45.582 10.226 45.618 ;
               RECT 10.174 46.182 10.226 46.218 ;
               RECT 10.174 46.782 10.226 46.818 ;
               RECT 10.174 47.382 10.226 47.418 ;
               RECT 10.174 47.982 10.226 48.018 ;
               RECT 10.174 48.582 10.226 48.618 ;
               RECT 10.174 48.942 10.226 48.978 ;
               RECT 10.174 48.9475 10.226 48.9725 ;
               RECT 10.174 49.182 10.226 49.218 ;
               RECT 10.174 49.902 10.226 49.938 ;
               RECT 10.174 50.622 10.226 50.658 ;
               RECT 10.174 50.862 10.226 50.898 ;
               RECT 10.174 51.342 10.226 51.378 ;
               RECT 10.174 51.822 10.226 51.858 ;
               RECT 10.174 52.302 10.226 52.338 ;
               RECT 10.174 52.782 10.226 52.818 ;
               RECT 10.174 53.262 10.226 53.298 ;
               RECT 10.174 53.742 10.226 53.778 ;
               RECT 10.174 54.222 10.226 54.258 ;
               RECT 10.174 54.462 10.226 54.498 ;
               RECT 10.174 55.182 10.226 55.218 ;
               RECT 10.174 55.902 10.226 55.938 ;
               RECT 10.174 56.142 10.226 56.178 ;
               RECT 10.174 56.1475 10.226 56.1725 ;
               RECT 10.174 56.502 10.226 56.538 ;
               RECT 10.174 57.102 10.226 57.138 ;
               RECT 10.174 57.702 10.226 57.738 ;
               RECT 10.174 58.302 10.226 58.338 ;
               RECT 10.174 58.902 10.226 58.938 ;
               RECT 10.174 59.502 10.226 59.538 ;
               RECT 10.174 60.102 10.226 60.138 ;
               RECT 10.174 60.702 10.226 60.738 ;
               RECT 10.174 61.302 10.226 61.338 ;
               RECT 10.174 61.902 10.226 61.938 ;
               RECT 10.174 62.502 10.226 62.538 ;
               RECT 10.174 63.102 10.226 63.138 ;
               RECT 10.174 63.702 10.226 63.738 ;
               RECT 10.174 64.302 10.226 64.338 ;
               RECT 10.174 64.902 10.226 64.938 ;
               RECT 10.174 65.502 10.226 65.538 ;
               RECT 10.174 66.102 10.226 66.138 ;
               RECT 10.174 66.702 10.226 66.738 ;
               RECT 10.174 67.302 10.226 67.338 ;
               RECT 10.174 67.902 10.226 67.938 ;
               RECT 10.174 68.502 10.226 68.538 ;
               RECT 10.174 69.102 10.226 69.138 ;
               RECT 10.174 69.702 10.226 69.738 ;
               RECT 10.174 70.302 10.226 70.338 ;
               RECT 10.174 70.902 10.226 70.938 ;
               RECT 10.174 71.502 10.226 71.538 ;
               RECT 10.174 72.102 10.226 72.138 ;
               RECT 10.174 72.702 10.226 72.738 ;
               RECT 10.174 73.302 10.226 73.338 ;
               RECT 10.174 73.902 10.226 73.938 ;
               RECT 10.174 74.502 10.226 74.538 ;
               RECT 10.174 75.102 10.226 75.138 ;
               RECT 10.174 75.702 10.226 75.738 ;
               RECT 10.174 76.302 10.226 76.338 ;
               RECT 10.174 76.902 10.226 76.938 ;
               RECT 10.174 77.502 10.226 77.538 ;
               RECT 10.174 78.102 10.226 78.138 ;
               RECT 10.174 78.702 10.226 78.738 ;
               RECT 10.174 79.302 10.226 79.338 ;
               RECT 10.174 79.902 10.226 79.938 ;
               RECT 10.174 80.502 10.226 80.538 ;
               RECT 10.174 81.102 10.226 81.138 ;
               RECT 10.174 81.702 10.226 81.738 ;
               RECT 10.174 82.302 10.226 82.338 ;
               RECT 10.174 82.902 10.226 82.938 ;
               RECT 10.174 83.502 10.226 83.538 ;
               RECT 10.174 84.102 10.226 84.138 ;
               RECT 10.174 84.702 10.226 84.738 ;
               RECT 10.174 85.302 10.226 85.338 ;
               RECT 10.174 85.902 10.226 85.938 ;
               RECT 10.174 86.502 10.226 86.538 ;
               RECT 10.174 87.102 10.226 87.138 ;
               RECT 10.174 87.702 10.226 87.738 ;
               RECT 10.174 88.302 10.226 88.338 ;
               RECT 10.174 88.902 10.226 88.938 ;
               RECT 10.174 89.502 10.226 89.538 ;
               RECT 10.174 90.102 10.226 90.138 ;
               RECT 10.174 90.702 10.226 90.738 ;
               RECT 10.174 91.302 10.226 91.338 ;
               RECT 10.174 91.902 10.226 91.938 ;
               RECT 10.174 92.502 10.226 92.538 ;
               RECT 10.174 93.102 10.226 93.138 ;
               RECT 10.174 93.702 10.226 93.738 ;
               RECT 10.174 94.302 10.226 94.338 ;
               RECT 10.174 94.902 10.226 94.938 ;
               RECT 10.174 95.502 10.226 95.538 ;
               RECT 10.174 96.102 10.226 96.138 ;
               RECT 10.174 96.702 10.226 96.738 ;
               RECT 10.174 97.302 10.226 97.338 ;
               RECT 10.174 97.902 10.226 97.938 ;
               RECT 10.174 98.502 10.226 98.538 ;
               RECT 10.174 99.102 10.226 99.138 ;
               RECT 10.174 99.702 10.226 99.738 ;
               RECT 10.174 100.302 10.226 100.338 ;
               RECT 10.174 100.902 10.226 100.938 ;
               RECT 10.174 101.502 10.226 101.538 ;
               RECT 10.174 102.102 10.226 102.138 ;
               RECT 10.174 102.702 10.226 102.738 ;
               RECT 10.174 103.302 10.226 103.338 ;
               RECT 10.174 103.902 10.226 103.938 ;
               RECT 10.174 104.502 10.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 10.974 0.5695 11.026 104.5505 ;
               LAYER v4 ;
               RECT 10.974 0.582 11.026 0.618 ;
               RECT 10.974 1.182 11.026 1.218 ;
               RECT 10.974 1.782 11.026 1.818 ;
               RECT 10.974 2.382 11.026 2.418 ;
               RECT 10.974 2.982 11.026 3.018 ;
               RECT 10.974 3.582 11.026 3.618 ;
               RECT 10.974 4.182 11.026 4.218 ;
               RECT 10.974 4.782 11.026 4.818 ;
               RECT 10.974 5.382 11.026 5.418 ;
               RECT 10.974 5.982 11.026 6.018 ;
               RECT 10.974 6.582 11.026 6.618 ;
               RECT 10.974 7.182 11.026 7.218 ;
               RECT 10.974 7.782 11.026 7.818 ;
               RECT 10.974 8.382 11.026 8.418 ;
               RECT 10.974 8.982 11.026 9.018 ;
               RECT 10.974 9.582 11.026 9.618 ;
               RECT 10.974 10.182 11.026 10.218 ;
               RECT 10.974 10.782 11.026 10.818 ;
               RECT 10.974 11.382 11.026 11.418 ;
               RECT 10.974 11.982 11.026 12.018 ;
               RECT 10.974 12.582 11.026 12.618 ;
               RECT 10.974 13.182 11.026 13.218 ;
               RECT 10.974 13.782 11.026 13.818 ;
               RECT 10.974 14.382 11.026 14.418 ;
               RECT 10.974 14.982 11.026 15.018 ;
               RECT 10.974 15.582 11.026 15.618 ;
               RECT 10.974 16.182 11.026 16.218 ;
               RECT 10.974 16.782 11.026 16.818 ;
               RECT 10.974 17.382 11.026 17.418 ;
               RECT 10.974 17.982 11.026 18.018 ;
               RECT 10.974 18.582 11.026 18.618 ;
               RECT 10.974 19.182 11.026 19.218 ;
               RECT 10.974 19.782 11.026 19.818 ;
               RECT 10.974 20.382 11.026 20.418 ;
               RECT 10.974 20.982 11.026 21.018 ;
               RECT 10.974 21.582 11.026 21.618 ;
               RECT 10.974 22.182 11.026 22.218 ;
               RECT 10.974 22.782 11.026 22.818 ;
               RECT 10.974 23.382 11.026 23.418 ;
               RECT 10.974 23.982 11.026 24.018 ;
               RECT 10.974 24.582 11.026 24.618 ;
               RECT 10.974 25.182 11.026 25.218 ;
               RECT 10.974 25.782 11.026 25.818 ;
               RECT 10.974 26.382 11.026 26.418 ;
               RECT 10.974 26.982 11.026 27.018 ;
               RECT 10.974 27.582 11.026 27.618 ;
               RECT 10.974 28.182 11.026 28.218 ;
               RECT 10.974 28.782 11.026 28.818 ;
               RECT 10.974 29.382 11.026 29.418 ;
               RECT 10.974 29.982 11.026 30.018 ;
               RECT 10.974 30.582 11.026 30.618 ;
               RECT 10.974 31.182 11.026 31.218 ;
               RECT 10.974 31.782 11.026 31.818 ;
               RECT 10.974 32.382 11.026 32.418 ;
               RECT 10.974 32.982 11.026 33.018 ;
               RECT 10.974 33.582 11.026 33.618 ;
               RECT 10.974 34.182 11.026 34.218 ;
               RECT 10.974 34.782 11.026 34.818 ;
               RECT 10.974 35.382 11.026 35.418 ;
               RECT 10.974 35.982 11.026 36.018 ;
               RECT 10.974 36.582 11.026 36.618 ;
               RECT 10.974 37.182 11.026 37.218 ;
               RECT 10.974 37.782 11.026 37.818 ;
               RECT 10.974 38.382 11.026 38.418 ;
               RECT 10.974 38.982 11.026 39.018 ;
               RECT 10.974 39.582 11.026 39.618 ;
               RECT 10.974 40.182 11.026 40.218 ;
               RECT 10.974 40.782 11.026 40.818 ;
               RECT 10.974 41.382 11.026 41.418 ;
               RECT 10.974 41.982 11.026 42.018 ;
               RECT 10.974 42.582 11.026 42.618 ;
               RECT 10.974 43.182 11.026 43.218 ;
               RECT 10.974 43.782 11.026 43.818 ;
               RECT 10.974 44.382 11.026 44.418 ;
               RECT 10.974 44.982 11.026 45.018 ;
               RECT 10.974 45.582 11.026 45.618 ;
               RECT 10.974 46.182 11.026 46.218 ;
               RECT 10.974 46.782 11.026 46.818 ;
               RECT 10.974 47.382 11.026 47.418 ;
               RECT 10.974 47.982 11.026 48.018 ;
               RECT 10.974 48.582 11.026 48.618 ;
               RECT 10.974 48.942 11.026 48.978 ;
               RECT 10.974 49.182 11.026 49.218 ;
               RECT 10.974 49.902 11.026 49.938 ;
               RECT 10.974 50.622 11.026 50.658 ;
               RECT 10.974 50.862 11.026 50.898 ;
               RECT 10.974 51.342 11.026 51.378 ;
               RECT 10.974 51.822 11.026 51.858 ;
               RECT 10.974 52.302 11.026 52.338 ;
               RECT 10.974 52.782 11.026 52.818 ;
               RECT 10.974 53.262 11.026 53.298 ;
               RECT 10.974 53.742 11.026 53.778 ;
               RECT 10.974 54.222 11.026 54.258 ;
               RECT 10.974 54.462 11.026 54.498 ;
               RECT 10.974 55.182 11.026 55.218 ;
               RECT 10.974 55.902 11.026 55.938 ;
               RECT 10.974 56.142 11.026 56.178 ;
               RECT 10.974 56.502 11.026 56.538 ;
               RECT 10.974 57.102 11.026 57.138 ;
               RECT 10.974 57.702 11.026 57.738 ;
               RECT 10.974 58.302 11.026 58.338 ;
               RECT 10.974 58.902 11.026 58.938 ;
               RECT 10.974 59.502 11.026 59.538 ;
               RECT 10.974 60.102 11.026 60.138 ;
               RECT 10.974 60.702 11.026 60.738 ;
               RECT 10.974 61.302 11.026 61.338 ;
               RECT 10.974 61.902 11.026 61.938 ;
               RECT 10.974 62.502 11.026 62.538 ;
               RECT 10.974 63.102 11.026 63.138 ;
               RECT 10.974 63.702 11.026 63.738 ;
               RECT 10.974 64.302 11.026 64.338 ;
               RECT 10.974 64.902 11.026 64.938 ;
               RECT 10.974 65.502 11.026 65.538 ;
               RECT 10.974 66.102 11.026 66.138 ;
               RECT 10.974 66.702 11.026 66.738 ;
               RECT 10.974 67.302 11.026 67.338 ;
               RECT 10.974 67.902 11.026 67.938 ;
               RECT 10.974 68.502 11.026 68.538 ;
               RECT 10.974 69.102 11.026 69.138 ;
               RECT 10.974 69.702 11.026 69.738 ;
               RECT 10.974 70.302 11.026 70.338 ;
               RECT 10.974 70.902 11.026 70.938 ;
               RECT 10.974 71.502 11.026 71.538 ;
               RECT 10.974 72.102 11.026 72.138 ;
               RECT 10.974 72.702 11.026 72.738 ;
               RECT 10.974 73.302 11.026 73.338 ;
               RECT 10.974 73.902 11.026 73.938 ;
               RECT 10.974 74.502 11.026 74.538 ;
               RECT 10.974 75.102 11.026 75.138 ;
               RECT 10.974 75.702 11.026 75.738 ;
               RECT 10.974 76.302 11.026 76.338 ;
               RECT 10.974 76.902 11.026 76.938 ;
               RECT 10.974 77.502 11.026 77.538 ;
               RECT 10.974 78.102 11.026 78.138 ;
               RECT 10.974 78.702 11.026 78.738 ;
               RECT 10.974 79.302 11.026 79.338 ;
               RECT 10.974 79.902 11.026 79.938 ;
               RECT 10.974 80.502 11.026 80.538 ;
               RECT 10.974 81.102 11.026 81.138 ;
               RECT 10.974 81.702 11.026 81.738 ;
               RECT 10.974 82.302 11.026 82.338 ;
               RECT 10.974 82.902 11.026 82.938 ;
               RECT 10.974 83.502 11.026 83.538 ;
               RECT 10.974 84.102 11.026 84.138 ;
               RECT 10.974 84.702 11.026 84.738 ;
               RECT 10.974 85.302 11.026 85.338 ;
               RECT 10.974 85.902 11.026 85.938 ;
               RECT 10.974 86.502 11.026 86.538 ;
               RECT 10.974 87.102 11.026 87.138 ;
               RECT 10.974 87.702 11.026 87.738 ;
               RECT 10.974 88.302 11.026 88.338 ;
               RECT 10.974 88.902 11.026 88.938 ;
               RECT 10.974 89.502 11.026 89.538 ;
               RECT 10.974 90.102 11.026 90.138 ;
               RECT 10.974 90.702 11.026 90.738 ;
               RECT 10.974 91.302 11.026 91.338 ;
               RECT 10.974 91.902 11.026 91.938 ;
               RECT 10.974 92.502 11.026 92.538 ;
               RECT 10.974 93.102 11.026 93.138 ;
               RECT 10.974 93.702 11.026 93.738 ;
               RECT 10.974 94.302 11.026 94.338 ;
               RECT 10.974 94.902 11.026 94.938 ;
               RECT 10.974 95.502 11.026 95.538 ;
               RECT 10.974 96.102 11.026 96.138 ;
               RECT 10.974 96.702 11.026 96.738 ;
               RECT 10.974 97.302 11.026 97.338 ;
               RECT 10.974 97.902 11.026 97.938 ;
               RECT 10.974 98.502 11.026 98.538 ;
               RECT 10.974 99.102 11.026 99.138 ;
               RECT 10.974 99.702 11.026 99.738 ;
               RECT 10.974 100.302 11.026 100.338 ;
               RECT 10.974 100.902 11.026 100.938 ;
               RECT 10.974 101.502 11.026 101.538 ;
               RECT 10.974 102.102 11.026 102.138 ;
               RECT 10.974 102.702 11.026 102.738 ;
               RECT 10.974 103.302 11.026 103.338 ;
               RECT 10.974 103.902 11.026 103.938 ;
               RECT 10.974 104.502 11.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 11.774 0.5695 11.826 104.5505 ;
               LAYER v4 ;
               RECT 11.774 0.582 11.826 0.618 ;
               RECT 11.774 1.182 11.826 1.218 ;
               RECT 11.774 1.782 11.826 1.818 ;
               RECT 11.774 2.382 11.826 2.418 ;
               RECT 11.774 2.982 11.826 3.018 ;
               RECT 11.774 3.582 11.826 3.618 ;
               RECT 11.774 4.182 11.826 4.218 ;
               RECT 11.774 4.782 11.826 4.818 ;
               RECT 11.774 5.382 11.826 5.418 ;
               RECT 11.774 5.982 11.826 6.018 ;
               RECT 11.774 6.582 11.826 6.618 ;
               RECT 11.774 7.182 11.826 7.218 ;
               RECT 11.774 7.782 11.826 7.818 ;
               RECT 11.774 8.382 11.826 8.418 ;
               RECT 11.774 8.982 11.826 9.018 ;
               RECT 11.774 9.582 11.826 9.618 ;
               RECT 11.774 10.182 11.826 10.218 ;
               RECT 11.774 10.782 11.826 10.818 ;
               RECT 11.774 11.382 11.826 11.418 ;
               RECT 11.774 11.982 11.826 12.018 ;
               RECT 11.774 12.582 11.826 12.618 ;
               RECT 11.774 13.182 11.826 13.218 ;
               RECT 11.774 13.782 11.826 13.818 ;
               RECT 11.774 14.382 11.826 14.418 ;
               RECT 11.774 14.982 11.826 15.018 ;
               RECT 11.774 15.582 11.826 15.618 ;
               RECT 11.774 16.182 11.826 16.218 ;
               RECT 11.774 16.782 11.826 16.818 ;
               RECT 11.774 17.382 11.826 17.418 ;
               RECT 11.774 17.982 11.826 18.018 ;
               RECT 11.774 18.582 11.826 18.618 ;
               RECT 11.774 19.182 11.826 19.218 ;
               RECT 11.774 19.782 11.826 19.818 ;
               RECT 11.774 20.382 11.826 20.418 ;
               RECT 11.774 20.982 11.826 21.018 ;
               RECT 11.774 21.582 11.826 21.618 ;
               RECT 11.774 22.182 11.826 22.218 ;
               RECT 11.774 22.782 11.826 22.818 ;
               RECT 11.774 23.382 11.826 23.418 ;
               RECT 11.774 23.982 11.826 24.018 ;
               RECT 11.774 24.582 11.826 24.618 ;
               RECT 11.774 25.182 11.826 25.218 ;
               RECT 11.774 25.782 11.826 25.818 ;
               RECT 11.774 26.382 11.826 26.418 ;
               RECT 11.774 26.982 11.826 27.018 ;
               RECT 11.774 27.582 11.826 27.618 ;
               RECT 11.774 28.182 11.826 28.218 ;
               RECT 11.774 28.782 11.826 28.818 ;
               RECT 11.774 29.382 11.826 29.418 ;
               RECT 11.774 29.982 11.826 30.018 ;
               RECT 11.774 30.582 11.826 30.618 ;
               RECT 11.774 31.182 11.826 31.218 ;
               RECT 11.774 31.782 11.826 31.818 ;
               RECT 11.774 32.382 11.826 32.418 ;
               RECT 11.774 32.982 11.826 33.018 ;
               RECT 11.774 33.582 11.826 33.618 ;
               RECT 11.774 34.182 11.826 34.218 ;
               RECT 11.774 34.782 11.826 34.818 ;
               RECT 11.774 35.382 11.826 35.418 ;
               RECT 11.774 35.982 11.826 36.018 ;
               RECT 11.774 36.582 11.826 36.618 ;
               RECT 11.774 37.182 11.826 37.218 ;
               RECT 11.774 37.782 11.826 37.818 ;
               RECT 11.774 38.382 11.826 38.418 ;
               RECT 11.774 38.982 11.826 39.018 ;
               RECT 11.774 39.582 11.826 39.618 ;
               RECT 11.774 40.182 11.826 40.218 ;
               RECT 11.774 40.782 11.826 40.818 ;
               RECT 11.774 41.382 11.826 41.418 ;
               RECT 11.774 41.982 11.826 42.018 ;
               RECT 11.774 42.582 11.826 42.618 ;
               RECT 11.774 43.182 11.826 43.218 ;
               RECT 11.774 43.782 11.826 43.818 ;
               RECT 11.774 44.382 11.826 44.418 ;
               RECT 11.774 44.982 11.826 45.018 ;
               RECT 11.774 45.582 11.826 45.618 ;
               RECT 11.774 46.182 11.826 46.218 ;
               RECT 11.774 46.782 11.826 46.818 ;
               RECT 11.774 47.382 11.826 47.418 ;
               RECT 11.774 47.982 11.826 48.018 ;
               RECT 11.774 48.582 11.826 48.618 ;
               RECT 11.774 48.942 11.826 48.978 ;
               RECT 11.774 48.9475 11.826 48.9725 ;
               RECT 11.774 49.182 11.826 49.218 ;
               RECT 11.774 49.902 11.826 49.938 ;
               RECT 11.774 50.622 11.826 50.658 ;
               RECT 11.774 50.862 11.826 50.898 ;
               RECT 11.774 51.342 11.826 51.378 ;
               RECT 11.774 51.822 11.826 51.858 ;
               RECT 11.774 52.302 11.826 52.338 ;
               RECT 11.774 52.782 11.826 52.818 ;
               RECT 11.774 53.262 11.826 53.298 ;
               RECT 11.774 53.742 11.826 53.778 ;
               RECT 11.774 54.222 11.826 54.258 ;
               RECT 11.774 54.462 11.826 54.498 ;
               RECT 11.774 55.182 11.826 55.218 ;
               RECT 11.774 55.902 11.826 55.938 ;
               RECT 11.774 56.142 11.826 56.178 ;
               RECT 11.774 56.1475 11.826 56.1725 ;
               RECT 11.774 56.502 11.826 56.538 ;
               RECT 11.774 57.102 11.826 57.138 ;
               RECT 11.774 57.702 11.826 57.738 ;
               RECT 11.774 58.302 11.826 58.338 ;
               RECT 11.774 58.902 11.826 58.938 ;
               RECT 11.774 59.502 11.826 59.538 ;
               RECT 11.774 60.102 11.826 60.138 ;
               RECT 11.774 60.702 11.826 60.738 ;
               RECT 11.774 61.302 11.826 61.338 ;
               RECT 11.774 61.902 11.826 61.938 ;
               RECT 11.774 62.502 11.826 62.538 ;
               RECT 11.774 63.102 11.826 63.138 ;
               RECT 11.774 63.702 11.826 63.738 ;
               RECT 11.774 64.302 11.826 64.338 ;
               RECT 11.774 64.902 11.826 64.938 ;
               RECT 11.774 65.502 11.826 65.538 ;
               RECT 11.774 66.102 11.826 66.138 ;
               RECT 11.774 66.702 11.826 66.738 ;
               RECT 11.774 67.302 11.826 67.338 ;
               RECT 11.774 67.902 11.826 67.938 ;
               RECT 11.774 68.502 11.826 68.538 ;
               RECT 11.774 69.102 11.826 69.138 ;
               RECT 11.774 69.702 11.826 69.738 ;
               RECT 11.774 70.302 11.826 70.338 ;
               RECT 11.774 70.902 11.826 70.938 ;
               RECT 11.774 71.502 11.826 71.538 ;
               RECT 11.774 72.102 11.826 72.138 ;
               RECT 11.774 72.702 11.826 72.738 ;
               RECT 11.774 73.302 11.826 73.338 ;
               RECT 11.774 73.902 11.826 73.938 ;
               RECT 11.774 74.502 11.826 74.538 ;
               RECT 11.774 75.102 11.826 75.138 ;
               RECT 11.774 75.702 11.826 75.738 ;
               RECT 11.774 76.302 11.826 76.338 ;
               RECT 11.774 76.902 11.826 76.938 ;
               RECT 11.774 77.502 11.826 77.538 ;
               RECT 11.774 78.102 11.826 78.138 ;
               RECT 11.774 78.702 11.826 78.738 ;
               RECT 11.774 79.302 11.826 79.338 ;
               RECT 11.774 79.902 11.826 79.938 ;
               RECT 11.774 80.502 11.826 80.538 ;
               RECT 11.774 81.102 11.826 81.138 ;
               RECT 11.774 81.702 11.826 81.738 ;
               RECT 11.774 82.302 11.826 82.338 ;
               RECT 11.774 82.902 11.826 82.938 ;
               RECT 11.774 83.502 11.826 83.538 ;
               RECT 11.774 84.102 11.826 84.138 ;
               RECT 11.774 84.702 11.826 84.738 ;
               RECT 11.774 85.302 11.826 85.338 ;
               RECT 11.774 85.902 11.826 85.938 ;
               RECT 11.774 86.502 11.826 86.538 ;
               RECT 11.774 87.102 11.826 87.138 ;
               RECT 11.774 87.702 11.826 87.738 ;
               RECT 11.774 88.302 11.826 88.338 ;
               RECT 11.774 88.902 11.826 88.938 ;
               RECT 11.774 89.502 11.826 89.538 ;
               RECT 11.774 90.102 11.826 90.138 ;
               RECT 11.774 90.702 11.826 90.738 ;
               RECT 11.774 91.302 11.826 91.338 ;
               RECT 11.774 91.902 11.826 91.938 ;
               RECT 11.774 92.502 11.826 92.538 ;
               RECT 11.774 93.102 11.826 93.138 ;
               RECT 11.774 93.702 11.826 93.738 ;
               RECT 11.774 94.302 11.826 94.338 ;
               RECT 11.774 94.902 11.826 94.938 ;
               RECT 11.774 95.502 11.826 95.538 ;
               RECT 11.774 96.102 11.826 96.138 ;
               RECT 11.774 96.702 11.826 96.738 ;
               RECT 11.774 97.302 11.826 97.338 ;
               RECT 11.774 97.902 11.826 97.938 ;
               RECT 11.774 98.502 11.826 98.538 ;
               RECT 11.774 99.102 11.826 99.138 ;
               RECT 11.774 99.702 11.826 99.738 ;
               RECT 11.774 100.302 11.826 100.338 ;
               RECT 11.774 100.902 11.826 100.938 ;
               RECT 11.774 101.502 11.826 101.538 ;
               RECT 11.774 102.102 11.826 102.138 ;
               RECT 11.774 102.702 11.826 102.738 ;
               RECT 11.774 103.302 11.826 103.338 ;
               RECT 11.774 103.902 11.826 103.938 ;
               RECT 11.774 104.502 11.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 12.574 0.5695 12.626 104.5505 ;
               LAYER v4 ;
               RECT 12.574 0.582 12.626 0.618 ;
               RECT 12.574 1.182 12.626 1.218 ;
               RECT 12.574 1.782 12.626 1.818 ;
               RECT 12.574 2.382 12.626 2.418 ;
               RECT 12.574 2.982 12.626 3.018 ;
               RECT 12.574 3.582 12.626 3.618 ;
               RECT 12.574 4.182 12.626 4.218 ;
               RECT 12.574 4.782 12.626 4.818 ;
               RECT 12.574 5.382 12.626 5.418 ;
               RECT 12.574 5.982 12.626 6.018 ;
               RECT 12.574 6.582 12.626 6.618 ;
               RECT 12.574 7.182 12.626 7.218 ;
               RECT 12.574 7.782 12.626 7.818 ;
               RECT 12.574 8.382 12.626 8.418 ;
               RECT 12.574 8.982 12.626 9.018 ;
               RECT 12.574 9.582 12.626 9.618 ;
               RECT 12.574 10.182 12.626 10.218 ;
               RECT 12.574 10.782 12.626 10.818 ;
               RECT 12.574 11.382 12.626 11.418 ;
               RECT 12.574 11.982 12.626 12.018 ;
               RECT 12.574 12.582 12.626 12.618 ;
               RECT 12.574 13.182 12.626 13.218 ;
               RECT 12.574 13.782 12.626 13.818 ;
               RECT 12.574 14.382 12.626 14.418 ;
               RECT 12.574 14.982 12.626 15.018 ;
               RECT 12.574 15.582 12.626 15.618 ;
               RECT 12.574 16.182 12.626 16.218 ;
               RECT 12.574 16.782 12.626 16.818 ;
               RECT 12.574 17.382 12.626 17.418 ;
               RECT 12.574 17.982 12.626 18.018 ;
               RECT 12.574 18.582 12.626 18.618 ;
               RECT 12.574 19.182 12.626 19.218 ;
               RECT 12.574 19.782 12.626 19.818 ;
               RECT 12.574 20.382 12.626 20.418 ;
               RECT 12.574 20.982 12.626 21.018 ;
               RECT 12.574 21.582 12.626 21.618 ;
               RECT 12.574 22.182 12.626 22.218 ;
               RECT 12.574 22.782 12.626 22.818 ;
               RECT 12.574 23.382 12.626 23.418 ;
               RECT 12.574 23.982 12.626 24.018 ;
               RECT 12.574 24.582 12.626 24.618 ;
               RECT 12.574 25.182 12.626 25.218 ;
               RECT 12.574 25.782 12.626 25.818 ;
               RECT 12.574 26.382 12.626 26.418 ;
               RECT 12.574 26.982 12.626 27.018 ;
               RECT 12.574 27.582 12.626 27.618 ;
               RECT 12.574 28.182 12.626 28.218 ;
               RECT 12.574 28.782 12.626 28.818 ;
               RECT 12.574 29.382 12.626 29.418 ;
               RECT 12.574 29.982 12.626 30.018 ;
               RECT 12.574 30.582 12.626 30.618 ;
               RECT 12.574 31.182 12.626 31.218 ;
               RECT 12.574 31.782 12.626 31.818 ;
               RECT 12.574 32.382 12.626 32.418 ;
               RECT 12.574 32.982 12.626 33.018 ;
               RECT 12.574 33.582 12.626 33.618 ;
               RECT 12.574 34.182 12.626 34.218 ;
               RECT 12.574 34.782 12.626 34.818 ;
               RECT 12.574 35.382 12.626 35.418 ;
               RECT 12.574 35.982 12.626 36.018 ;
               RECT 12.574 36.582 12.626 36.618 ;
               RECT 12.574 37.182 12.626 37.218 ;
               RECT 12.574 37.782 12.626 37.818 ;
               RECT 12.574 38.382 12.626 38.418 ;
               RECT 12.574 38.982 12.626 39.018 ;
               RECT 12.574 39.582 12.626 39.618 ;
               RECT 12.574 40.182 12.626 40.218 ;
               RECT 12.574 40.782 12.626 40.818 ;
               RECT 12.574 41.382 12.626 41.418 ;
               RECT 12.574 41.982 12.626 42.018 ;
               RECT 12.574 42.582 12.626 42.618 ;
               RECT 12.574 43.182 12.626 43.218 ;
               RECT 12.574 43.782 12.626 43.818 ;
               RECT 12.574 44.382 12.626 44.418 ;
               RECT 12.574 44.982 12.626 45.018 ;
               RECT 12.574 45.582 12.626 45.618 ;
               RECT 12.574 46.182 12.626 46.218 ;
               RECT 12.574 46.782 12.626 46.818 ;
               RECT 12.574 47.382 12.626 47.418 ;
               RECT 12.574 47.982 12.626 48.018 ;
               RECT 12.574 48.582 12.626 48.618 ;
               RECT 12.574 48.942 12.626 48.978 ;
               RECT 12.574 49.182 12.626 49.218 ;
               RECT 12.574 49.902 12.626 49.938 ;
               RECT 12.574 50.622 12.626 50.658 ;
               RECT 12.574 50.862 12.626 50.898 ;
               RECT 12.574 51.342 12.626 51.378 ;
               RECT 12.574 51.822 12.626 51.858 ;
               RECT 12.574 52.302 12.626 52.338 ;
               RECT 12.574 52.782 12.626 52.818 ;
               RECT 12.574 53.262 12.626 53.298 ;
               RECT 12.574 53.742 12.626 53.778 ;
               RECT 12.574 54.222 12.626 54.258 ;
               RECT 12.574 54.462 12.626 54.498 ;
               RECT 12.574 55.182 12.626 55.218 ;
               RECT 12.574 55.902 12.626 55.938 ;
               RECT 12.574 56.142 12.626 56.178 ;
               RECT 12.574 56.502 12.626 56.538 ;
               RECT 12.574 57.102 12.626 57.138 ;
               RECT 12.574 57.702 12.626 57.738 ;
               RECT 12.574 58.302 12.626 58.338 ;
               RECT 12.574 58.902 12.626 58.938 ;
               RECT 12.574 59.502 12.626 59.538 ;
               RECT 12.574 60.102 12.626 60.138 ;
               RECT 12.574 60.702 12.626 60.738 ;
               RECT 12.574 61.302 12.626 61.338 ;
               RECT 12.574 61.902 12.626 61.938 ;
               RECT 12.574 62.502 12.626 62.538 ;
               RECT 12.574 63.102 12.626 63.138 ;
               RECT 12.574 63.702 12.626 63.738 ;
               RECT 12.574 64.302 12.626 64.338 ;
               RECT 12.574 64.902 12.626 64.938 ;
               RECT 12.574 65.502 12.626 65.538 ;
               RECT 12.574 66.102 12.626 66.138 ;
               RECT 12.574 66.702 12.626 66.738 ;
               RECT 12.574 67.302 12.626 67.338 ;
               RECT 12.574 67.902 12.626 67.938 ;
               RECT 12.574 68.502 12.626 68.538 ;
               RECT 12.574 69.102 12.626 69.138 ;
               RECT 12.574 69.702 12.626 69.738 ;
               RECT 12.574 70.302 12.626 70.338 ;
               RECT 12.574 70.902 12.626 70.938 ;
               RECT 12.574 71.502 12.626 71.538 ;
               RECT 12.574 72.102 12.626 72.138 ;
               RECT 12.574 72.702 12.626 72.738 ;
               RECT 12.574 73.302 12.626 73.338 ;
               RECT 12.574 73.902 12.626 73.938 ;
               RECT 12.574 74.502 12.626 74.538 ;
               RECT 12.574 75.102 12.626 75.138 ;
               RECT 12.574 75.702 12.626 75.738 ;
               RECT 12.574 76.302 12.626 76.338 ;
               RECT 12.574 76.902 12.626 76.938 ;
               RECT 12.574 77.502 12.626 77.538 ;
               RECT 12.574 78.102 12.626 78.138 ;
               RECT 12.574 78.702 12.626 78.738 ;
               RECT 12.574 79.302 12.626 79.338 ;
               RECT 12.574 79.902 12.626 79.938 ;
               RECT 12.574 80.502 12.626 80.538 ;
               RECT 12.574 81.102 12.626 81.138 ;
               RECT 12.574 81.702 12.626 81.738 ;
               RECT 12.574 82.302 12.626 82.338 ;
               RECT 12.574 82.902 12.626 82.938 ;
               RECT 12.574 83.502 12.626 83.538 ;
               RECT 12.574 84.102 12.626 84.138 ;
               RECT 12.574 84.702 12.626 84.738 ;
               RECT 12.574 85.302 12.626 85.338 ;
               RECT 12.574 85.902 12.626 85.938 ;
               RECT 12.574 86.502 12.626 86.538 ;
               RECT 12.574 87.102 12.626 87.138 ;
               RECT 12.574 87.702 12.626 87.738 ;
               RECT 12.574 88.302 12.626 88.338 ;
               RECT 12.574 88.902 12.626 88.938 ;
               RECT 12.574 89.502 12.626 89.538 ;
               RECT 12.574 90.102 12.626 90.138 ;
               RECT 12.574 90.702 12.626 90.738 ;
               RECT 12.574 91.302 12.626 91.338 ;
               RECT 12.574 91.902 12.626 91.938 ;
               RECT 12.574 92.502 12.626 92.538 ;
               RECT 12.574 93.102 12.626 93.138 ;
               RECT 12.574 93.702 12.626 93.738 ;
               RECT 12.574 94.302 12.626 94.338 ;
               RECT 12.574 94.902 12.626 94.938 ;
               RECT 12.574 95.502 12.626 95.538 ;
               RECT 12.574 96.102 12.626 96.138 ;
               RECT 12.574 96.702 12.626 96.738 ;
               RECT 12.574 97.302 12.626 97.338 ;
               RECT 12.574 97.902 12.626 97.938 ;
               RECT 12.574 98.502 12.626 98.538 ;
               RECT 12.574 99.102 12.626 99.138 ;
               RECT 12.574 99.702 12.626 99.738 ;
               RECT 12.574 100.302 12.626 100.338 ;
               RECT 12.574 100.902 12.626 100.938 ;
               RECT 12.574 101.502 12.626 101.538 ;
               RECT 12.574 102.102 12.626 102.138 ;
               RECT 12.574 102.702 12.626 102.738 ;
               RECT 12.574 103.302 12.626 103.338 ;
               RECT 12.574 103.902 12.626 103.938 ;
               RECT 12.574 104.502 12.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 13.374 0.5695 13.426 104.5505 ;
               LAYER v4 ;
               RECT 13.374 0.582 13.426 0.618 ;
               RECT 13.374 1.182 13.426 1.218 ;
               RECT 13.374 1.782 13.426 1.818 ;
               RECT 13.374 2.382 13.426 2.418 ;
               RECT 13.374 2.982 13.426 3.018 ;
               RECT 13.374 3.582 13.426 3.618 ;
               RECT 13.374 4.182 13.426 4.218 ;
               RECT 13.374 4.782 13.426 4.818 ;
               RECT 13.374 5.382 13.426 5.418 ;
               RECT 13.374 5.982 13.426 6.018 ;
               RECT 13.374 6.582 13.426 6.618 ;
               RECT 13.374 7.182 13.426 7.218 ;
               RECT 13.374 7.782 13.426 7.818 ;
               RECT 13.374 8.382 13.426 8.418 ;
               RECT 13.374 8.982 13.426 9.018 ;
               RECT 13.374 9.582 13.426 9.618 ;
               RECT 13.374 10.182 13.426 10.218 ;
               RECT 13.374 10.782 13.426 10.818 ;
               RECT 13.374 11.382 13.426 11.418 ;
               RECT 13.374 11.982 13.426 12.018 ;
               RECT 13.374 12.582 13.426 12.618 ;
               RECT 13.374 13.182 13.426 13.218 ;
               RECT 13.374 13.782 13.426 13.818 ;
               RECT 13.374 14.382 13.426 14.418 ;
               RECT 13.374 14.982 13.426 15.018 ;
               RECT 13.374 15.582 13.426 15.618 ;
               RECT 13.374 16.182 13.426 16.218 ;
               RECT 13.374 16.782 13.426 16.818 ;
               RECT 13.374 17.382 13.426 17.418 ;
               RECT 13.374 17.982 13.426 18.018 ;
               RECT 13.374 18.582 13.426 18.618 ;
               RECT 13.374 19.182 13.426 19.218 ;
               RECT 13.374 19.782 13.426 19.818 ;
               RECT 13.374 20.382 13.426 20.418 ;
               RECT 13.374 20.982 13.426 21.018 ;
               RECT 13.374 21.582 13.426 21.618 ;
               RECT 13.374 22.182 13.426 22.218 ;
               RECT 13.374 22.782 13.426 22.818 ;
               RECT 13.374 23.382 13.426 23.418 ;
               RECT 13.374 23.982 13.426 24.018 ;
               RECT 13.374 24.582 13.426 24.618 ;
               RECT 13.374 25.182 13.426 25.218 ;
               RECT 13.374 25.782 13.426 25.818 ;
               RECT 13.374 26.382 13.426 26.418 ;
               RECT 13.374 26.982 13.426 27.018 ;
               RECT 13.374 27.582 13.426 27.618 ;
               RECT 13.374 28.182 13.426 28.218 ;
               RECT 13.374 28.782 13.426 28.818 ;
               RECT 13.374 29.382 13.426 29.418 ;
               RECT 13.374 29.982 13.426 30.018 ;
               RECT 13.374 30.582 13.426 30.618 ;
               RECT 13.374 31.182 13.426 31.218 ;
               RECT 13.374 31.782 13.426 31.818 ;
               RECT 13.374 32.382 13.426 32.418 ;
               RECT 13.374 32.982 13.426 33.018 ;
               RECT 13.374 33.582 13.426 33.618 ;
               RECT 13.374 34.182 13.426 34.218 ;
               RECT 13.374 34.782 13.426 34.818 ;
               RECT 13.374 35.382 13.426 35.418 ;
               RECT 13.374 35.982 13.426 36.018 ;
               RECT 13.374 36.582 13.426 36.618 ;
               RECT 13.374 37.182 13.426 37.218 ;
               RECT 13.374 37.782 13.426 37.818 ;
               RECT 13.374 38.382 13.426 38.418 ;
               RECT 13.374 38.982 13.426 39.018 ;
               RECT 13.374 39.582 13.426 39.618 ;
               RECT 13.374 40.182 13.426 40.218 ;
               RECT 13.374 40.782 13.426 40.818 ;
               RECT 13.374 41.382 13.426 41.418 ;
               RECT 13.374 41.982 13.426 42.018 ;
               RECT 13.374 42.582 13.426 42.618 ;
               RECT 13.374 43.182 13.426 43.218 ;
               RECT 13.374 43.782 13.426 43.818 ;
               RECT 13.374 44.382 13.426 44.418 ;
               RECT 13.374 44.982 13.426 45.018 ;
               RECT 13.374 45.582 13.426 45.618 ;
               RECT 13.374 46.182 13.426 46.218 ;
               RECT 13.374 46.782 13.426 46.818 ;
               RECT 13.374 47.382 13.426 47.418 ;
               RECT 13.374 47.982 13.426 48.018 ;
               RECT 13.374 48.582 13.426 48.618 ;
               RECT 13.374 48.9475 13.426 48.9725 ;
               RECT 13.374 49.182 13.426 49.218 ;
               RECT 13.374 49.902 13.426 49.938 ;
               RECT 13.374 50.622 13.426 50.658 ;
               RECT 13.374 50.862 13.426 50.898 ;
               RECT 13.374 51.342 13.426 51.378 ;
               RECT 13.374 51.822 13.426 51.858 ;
               RECT 13.374 52.302 13.426 52.338 ;
               RECT 13.374 52.782 13.426 52.818 ;
               RECT 13.374 53.262 13.426 53.298 ;
               RECT 13.374 53.742 13.426 53.778 ;
               RECT 13.374 54.222 13.426 54.258 ;
               RECT 13.374 54.462 13.426 54.498 ;
               RECT 13.374 55.182 13.426 55.218 ;
               RECT 13.374 55.902 13.426 55.938 ;
               RECT 13.374 56.1475 13.426 56.1725 ;
               RECT 13.374 56.502 13.426 56.538 ;
               RECT 13.374 57.102 13.426 57.138 ;
               RECT 13.374 57.702 13.426 57.738 ;
               RECT 13.374 58.302 13.426 58.338 ;
               RECT 13.374 58.902 13.426 58.938 ;
               RECT 13.374 59.502 13.426 59.538 ;
               RECT 13.374 60.102 13.426 60.138 ;
               RECT 13.374 60.702 13.426 60.738 ;
               RECT 13.374 61.302 13.426 61.338 ;
               RECT 13.374 61.902 13.426 61.938 ;
               RECT 13.374 62.502 13.426 62.538 ;
               RECT 13.374 63.102 13.426 63.138 ;
               RECT 13.374 63.702 13.426 63.738 ;
               RECT 13.374 64.302 13.426 64.338 ;
               RECT 13.374 64.902 13.426 64.938 ;
               RECT 13.374 65.502 13.426 65.538 ;
               RECT 13.374 66.102 13.426 66.138 ;
               RECT 13.374 66.702 13.426 66.738 ;
               RECT 13.374 67.302 13.426 67.338 ;
               RECT 13.374 67.902 13.426 67.938 ;
               RECT 13.374 68.502 13.426 68.538 ;
               RECT 13.374 69.102 13.426 69.138 ;
               RECT 13.374 69.702 13.426 69.738 ;
               RECT 13.374 70.302 13.426 70.338 ;
               RECT 13.374 70.902 13.426 70.938 ;
               RECT 13.374 71.502 13.426 71.538 ;
               RECT 13.374 72.102 13.426 72.138 ;
               RECT 13.374 72.702 13.426 72.738 ;
               RECT 13.374 73.302 13.426 73.338 ;
               RECT 13.374 73.902 13.426 73.938 ;
               RECT 13.374 74.502 13.426 74.538 ;
               RECT 13.374 75.102 13.426 75.138 ;
               RECT 13.374 75.702 13.426 75.738 ;
               RECT 13.374 76.302 13.426 76.338 ;
               RECT 13.374 76.902 13.426 76.938 ;
               RECT 13.374 77.502 13.426 77.538 ;
               RECT 13.374 78.102 13.426 78.138 ;
               RECT 13.374 78.702 13.426 78.738 ;
               RECT 13.374 79.302 13.426 79.338 ;
               RECT 13.374 79.902 13.426 79.938 ;
               RECT 13.374 80.502 13.426 80.538 ;
               RECT 13.374 81.102 13.426 81.138 ;
               RECT 13.374 81.702 13.426 81.738 ;
               RECT 13.374 82.302 13.426 82.338 ;
               RECT 13.374 82.902 13.426 82.938 ;
               RECT 13.374 83.502 13.426 83.538 ;
               RECT 13.374 84.102 13.426 84.138 ;
               RECT 13.374 84.702 13.426 84.738 ;
               RECT 13.374 85.302 13.426 85.338 ;
               RECT 13.374 85.902 13.426 85.938 ;
               RECT 13.374 86.502 13.426 86.538 ;
               RECT 13.374 87.102 13.426 87.138 ;
               RECT 13.374 87.702 13.426 87.738 ;
               RECT 13.374 88.302 13.426 88.338 ;
               RECT 13.374 88.902 13.426 88.938 ;
               RECT 13.374 89.502 13.426 89.538 ;
               RECT 13.374 90.102 13.426 90.138 ;
               RECT 13.374 90.702 13.426 90.738 ;
               RECT 13.374 91.302 13.426 91.338 ;
               RECT 13.374 91.902 13.426 91.938 ;
               RECT 13.374 92.502 13.426 92.538 ;
               RECT 13.374 93.102 13.426 93.138 ;
               RECT 13.374 93.702 13.426 93.738 ;
               RECT 13.374 94.302 13.426 94.338 ;
               RECT 13.374 94.902 13.426 94.938 ;
               RECT 13.374 95.502 13.426 95.538 ;
               RECT 13.374 96.102 13.426 96.138 ;
               RECT 13.374 96.702 13.426 96.738 ;
               RECT 13.374 97.302 13.426 97.338 ;
               RECT 13.374 97.902 13.426 97.938 ;
               RECT 13.374 98.502 13.426 98.538 ;
               RECT 13.374 99.102 13.426 99.138 ;
               RECT 13.374 99.702 13.426 99.738 ;
               RECT 13.374 100.302 13.426 100.338 ;
               RECT 13.374 100.902 13.426 100.938 ;
               RECT 13.374 101.502 13.426 101.538 ;
               RECT 13.374 102.102 13.426 102.138 ;
               RECT 13.374 102.702 13.426 102.738 ;
               RECT 13.374 103.302 13.426 103.338 ;
               RECT 13.374 103.902 13.426 103.938 ;
               RECT 13.374 104.502 13.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 14.45 0.5695 14.504 104.5505 ;
               LAYER v4 ;
               RECT 14.45 0.582 14.504 0.618 ;
               RECT 14.45 1.182 14.504 1.218 ;
               RECT 14.45 1.782 14.504 1.818 ;
               RECT 14.45 2.382 14.504 2.418 ;
               RECT 14.45 2.982 14.504 3.018 ;
               RECT 14.45 3.582 14.504 3.618 ;
               RECT 14.45 4.182 14.504 4.218 ;
               RECT 14.45 4.782 14.504 4.818 ;
               RECT 14.45 5.382 14.504 5.418 ;
               RECT 14.45 5.982 14.504 6.018 ;
               RECT 14.45 6.582 14.504 6.618 ;
               RECT 14.45 7.182 14.504 7.218 ;
               RECT 14.45 7.782 14.504 7.818 ;
               RECT 14.45 8.382 14.504 8.418 ;
               RECT 14.45 8.982 14.504 9.018 ;
               RECT 14.45 9.582 14.504 9.618 ;
               RECT 14.45 10.182 14.504 10.218 ;
               RECT 14.45 10.782 14.504 10.818 ;
               RECT 14.45 11.382 14.504 11.418 ;
               RECT 14.45 11.982 14.504 12.018 ;
               RECT 14.45 12.582 14.504 12.618 ;
               RECT 14.45 13.182 14.504 13.218 ;
               RECT 14.45 13.782 14.504 13.818 ;
               RECT 14.45 14.382 14.504 14.418 ;
               RECT 14.45 14.982 14.504 15.018 ;
               RECT 14.45 15.582 14.504 15.618 ;
               RECT 14.45 16.182 14.504 16.218 ;
               RECT 14.45 16.782 14.504 16.818 ;
               RECT 14.45 17.382 14.504 17.418 ;
               RECT 14.45 17.982 14.504 18.018 ;
               RECT 14.45 18.582 14.504 18.618 ;
               RECT 14.45 19.182 14.504 19.218 ;
               RECT 14.45 19.782 14.504 19.818 ;
               RECT 14.45 20.382 14.504 20.418 ;
               RECT 14.45 20.982 14.504 21.018 ;
               RECT 14.45 21.582 14.504 21.618 ;
               RECT 14.45 22.182 14.504 22.218 ;
               RECT 14.45 22.782 14.504 22.818 ;
               RECT 14.45 23.382 14.504 23.418 ;
               RECT 14.45 23.982 14.504 24.018 ;
               RECT 14.45 24.582 14.504 24.618 ;
               RECT 14.45 25.182 14.504 25.218 ;
               RECT 14.45 25.782 14.504 25.818 ;
               RECT 14.45 26.382 14.504 26.418 ;
               RECT 14.45 26.982 14.504 27.018 ;
               RECT 14.45 27.582 14.504 27.618 ;
               RECT 14.45 28.182 14.504 28.218 ;
               RECT 14.45 28.782 14.504 28.818 ;
               RECT 14.45 29.382 14.504 29.418 ;
               RECT 14.45 29.982 14.504 30.018 ;
               RECT 14.45 30.582 14.504 30.618 ;
               RECT 14.45 31.182 14.504 31.218 ;
               RECT 14.45 31.782 14.504 31.818 ;
               RECT 14.45 32.382 14.504 32.418 ;
               RECT 14.45 32.982 14.504 33.018 ;
               RECT 14.45 33.582 14.504 33.618 ;
               RECT 14.45 34.182 14.504 34.218 ;
               RECT 14.45 34.782 14.504 34.818 ;
               RECT 14.45 35.382 14.504 35.418 ;
               RECT 14.45 35.982 14.504 36.018 ;
               RECT 14.45 36.582 14.504 36.618 ;
               RECT 14.45 37.182 14.504 37.218 ;
               RECT 14.45 37.782 14.504 37.818 ;
               RECT 14.45 38.382 14.504 38.418 ;
               RECT 14.45 38.982 14.504 39.018 ;
               RECT 14.45 39.582 14.504 39.618 ;
               RECT 14.45 40.182 14.504 40.218 ;
               RECT 14.45 40.782 14.504 40.818 ;
               RECT 14.45 41.382 14.504 41.418 ;
               RECT 14.45 41.982 14.504 42.018 ;
               RECT 14.45 42.582 14.504 42.618 ;
               RECT 14.45 43.182 14.504 43.218 ;
               RECT 14.45 43.782 14.504 43.818 ;
               RECT 14.45 44.382 14.504 44.418 ;
               RECT 14.45 44.982 14.504 45.018 ;
               RECT 14.45 45.582 14.504 45.618 ;
               RECT 14.45 46.182 14.504 46.218 ;
               RECT 14.45 46.782 14.504 46.818 ;
               RECT 14.45 47.382 14.504 47.418 ;
               RECT 14.45 47.982 14.504 48.018 ;
               RECT 14.45 48.582 14.504 48.618 ;
               RECT 14.45 48.942 14.504 48.978 ;
               RECT 14.45 49.422 14.504 49.458 ;
               RECT 14.45 49.902 14.504 49.938 ;
               RECT 14.45 50.0835 14.504 50.1195 ;
               RECT 14.45 50.382 14.504 50.418 ;
               RECT 14.45 50.862 14.504 50.898 ;
               RECT 14.45 51.342 14.504 51.378 ;
               RECT 14.45 51.822 14.504 51.858 ;
               RECT 14.45 52.302 14.504 52.338 ;
               RECT 14.45 52.662 14.504 52.698 ;
               RECT 14.45 52.782 14.504 52.818 ;
               RECT 14.45 53.262 14.504 53.298 ;
               RECT 14.45 53.742 14.504 53.778 ;
               RECT 14.45 54.222 14.504 54.258 ;
               RECT 14.45 54.702 14.504 54.738 ;
               RECT 14.45 55.182 14.504 55.218 ;
               RECT 14.45 55.662 14.504 55.698 ;
               RECT 14.45 56.142 14.504 56.178 ;
               RECT 14.45 56.502 14.504 56.538 ;
               RECT 14.45 57.102 14.504 57.138 ;
               RECT 14.45 57.702 14.504 57.738 ;
               RECT 14.45 58.302 14.504 58.338 ;
               RECT 14.45 58.902 14.504 58.938 ;
               RECT 14.45 59.502 14.504 59.538 ;
               RECT 14.45 60.102 14.504 60.138 ;
               RECT 14.45 60.702 14.504 60.738 ;
               RECT 14.45 61.302 14.504 61.338 ;
               RECT 14.45 61.902 14.504 61.938 ;
               RECT 14.45 62.502 14.504 62.538 ;
               RECT 14.45 63.102 14.504 63.138 ;
               RECT 14.45 63.702 14.504 63.738 ;
               RECT 14.45 64.302 14.504 64.338 ;
               RECT 14.45 64.902 14.504 64.938 ;
               RECT 14.45 65.502 14.504 65.538 ;
               RECT 14.45 66.102 14.504 66.138 ;
               RECT 14.45 66.702 14.504 66.738 ;
               RECT 14.45 67.302 14.504 67.338 ;
               RECT 14.45 67.902 14.504 67.938 ;
               RECT 14.45 68.502 14.504 68.538 ;
               RECT 14.45 69.102 14.504 69.138 ;
               RECT 14.45 69.702 14.504 69.738 ;
               RECT 14.45 70.302 14.504 70.338 ;
               RECT 14.45 70.902 14.504 70.938 ;
               RECT 14.45 71.502 14.504 71.538 ;
               RECT 14.45 72.102 14.504 72.138 ;
               RECT 14.45 72.702 14.504 72.738 ;
               RECT 14.45 73.302 14.504 73.338 ;
               RECT 14.45 73.902 14.504 73.938 ;
               RECT 14.45 74.502 14.504 74.538 ;
               RECT 14.45 75.102 14.504 75.138 ;
               RECT 14.45 75.702 14.504 75.738 ;
               RECT 14.45 76.302 14.504 76.338 ;
               RECT 14.45 76.902 14.504 76.938 ;
               RECT 14.45 77.502 14.504 77.538 ;
               RECT 14.45 78.102 14.504 78.138 ;
               RECT 14.45 78.702 14.504 78.738 ;
               RECT 14.45 79.302 14.504 79.338 ;
               RECT 14.45 79.902 14.504 79.938 ;
               RECT 14.45 80.502 14.504 80.538 ;
               RECT 14.45 81.102 14.504 81.138 ;
               RECT 14.45 81.702 14.504 81.738 ;
               RECT 14.45 82.302 14.504 82.338 ;
               RECT 14.45 82.902 14.504 82.938 ;
               RECT 14.45 83.502 14.504 83.538 ;
               RECT 14.45 84.102 14.504 84.138 ;
               RECT 14.45 84.702 14.504 84.738 ;
               RECT 14.45 85.302 14.504 85.338 ;
               RECT 14.45 85.902 14.504 85.938 ;
               RECT 14.45 86.502 14.504 86.538 ;
               RECT 14.45 87.102 14.504 87.138 ;
               RECT 14.45 87.702 14.504 87.738 ;
               RECT 14.45 88.302 14.504 88.338 ;
               RECT 14.45 88.902 14.504 88.938 ;
               RECT 14.45 89.502 14.504 89.538 ;
               RECT 14.45 90.102 14.504 90.138 ;
               RECT 14.45 90.702 14.504 90.738 ;
               RECT 14.45 91.302 14.504 91.338 ;
               RECT 14.45 91.902 14.504 91.938 ;
               RECT 14.45 92.502 14.504 92.538 ;
               RECT 14.45 93.102 14.504 93.138 ;
               RECT 14.45 93.702 14.504 93.738 ;
               RECT 14.45 94.302 14.504 94.338 ;
               RECT 14.45 94.902 14.504 94.938 ;
               RECT 14.45 95.502 14.504 95.538 ;
               RECT 14.45 96.102 14.504 96.138 ;
               RECT 14.45 96.702 14.504 96.738 ;
               RECT 14.45 97.302 14.504 97.338 ;
               RECT 14.45 97.902 14.504 97.938 ;
               RECT 14.45 98.502 14.504 98.538 ;
               RECT 14.45 99.102 14.504 99.138 ;
               RECT 14.45 99.702 14.504 99.738 ;
               RECT 14.45 100.302 14.504 100.338 ;
               RECT 14.45 100.902 14.504 100.938 ;
               RECT 14.45 101.502 14.504 101.538 ;
               RECT 14.45 102.102 14.504 102.138 ;
               RECT 14.45 102.702 14.504 102.738 ;
               RECT 14.45 103.302 14.504 103.338 ;
               RECT 14.45 103.902 14.504 103.938 ;
               RECT 14.45 104.502 14.504 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.658 0.5695 15.71 104.5505 ;
               LAYER v4 ;
               RECT 15.658 0.582 15.71 0.618 ;
               RECT 15.658 1.182 15.71 1.218 ;
               RECT 15.658 1.782 15.71 1.818 ;
               RECT 15.658 2.382 15.71 2.418 ;
               RECT 15.658 2.982 15.71 3.018 ;
               RECT 15.658 3.582 15.71 3.618 ;
               RECT 15.658 4.182 15.71 4.218 ;
               RECT 15.658 4.782 15.71 4.818 ;
               RECT 15.658 5.382 15.71 5.418 ;
               RECT 15.658 5.982 15.71 6.018 ;
               RECT 15.658 6.582 15.71 6.618 ;
               RECT 15.658 7.182 15.71 7.218 ;
               RECT 15.658 7.782 15.71 7.818 ;
               RECT 15.658 8.382 15.71 8.418 ;
               RECT 15.658 8.982 15.71 9.018 ;
               RECT 15.658 9.582 15.71 9.618 ;
               RECT 15.658 10.182 15.71 10.218 ;
               RECT 15.658 10.782 15.71 10.818 ;
               RECT 15.658 11.382 15.71 11.418 ;
               RECT 15.658 11.982 15.71 12.018 ;
               RECT 15.658 12.582 15.71 12.618 ;
               RECT 15.658 13.182 15.71 13.218 ;
               RECT 15.658 13.782 15.71 13.818 ;
               RECT 15.658 14.382 15.71 14.418 ;
               RECT 15.658 14.982 15.71 15.018 ;
               RECT 15.658 15.582 15.71 15.618 ;
               RECT 15.658 16.182 15.71 16.218 ;
               RECT 15.658 16.782 15.71 16.818 ;
               RECT 15.658 17.382 15.71 17.418 ;
               RECT 15.658 17.982 15.71 18.018 ;
               RECT 15.658 18.582 15.71 18.618 ;
               RECT 15.658 19.182 15.71 19.218 ;
               RECT 15.658 19.782 15.71 19.818 ;
               RECT 15.658 20.382 15.71 20.418 ;
               RECT 15.658 20.982 15.71 21.018 ;
               RECT 15.658 21.582 15.71 21.618 ;
               RECT 15.658 22.182 15.71 22.218 ;
               RECT 15.658 22.782 15.71 22.818 ;
               RECT 15.658 23.382 15.71 23.418 ;
               RECT 15.658 23.982 15.71 24.018 ;
               RECT 15.658 24.582 15.71 24.618 ;
               RECT 15.658 25.182 15.71 25.218 ;
               RECT 15.658 25.782 15.71 25.818 ;
               RECT 15.658 26.382 15.71 26.418 ;
               RECT 15.658 26.982 15.71 27.018 ;
               RECT 15.658 27.582 15.71 27.618 ;
               RECT 15.658 28.182 15.71 28.218 ;
               RECT 15.658 28.782 15.71 28.818 ;
               RECT 15.658 29.382 15.71 29.418 ;
               RECT 15.658 29.982 15.71 30.018 ;
               RECT 15.658 30.582 15.71 30.618 ;
               RECT 15.658 31.182 15.71 31.218 ;
               RECT 15.658 31.782 15.71 31.818 ;
               RECT 15.658 32.382 15.71 32.418 ;
               RECT 15.658 32.982 15.71 33.018 ;
               RECT 15.658 33.582 15.71 33.618 ;
               RECT 15.658 34.182 15.71 34.218 ;
               RECT 15.658 34.782 15.71 34.818 ;
               RECT 15.658 35.382 15.71 35.418 ;
               RECT 15.658 35.982 15.71 36.018 ;
               RECT 15.658 36.582 15.71 36.618 ;
               RECT 15.658 37.182 15.71 37.218 ;
               RECT 15.658 37.782 15.71 37.818 ;
               RECT 15.658 38.382 15.71 38.418 ;
               RECT 15.658 38.982 15.71 39.018 ;
               RECT 15.658 39.582 15.71 39.618 ;
               RECT 15.658 40.182 15.71 40.218 ;
               RECT 15.658 40.782 15.71 40.818 ;
               RECT 15.658 41.382 15.71 41.418 ;
               RECT 15.658 41.982 15.71 42.018 ;
               RECT 15.658 42.582 15.71 42.618 ;
               RECT 15.658 43.182 15.71 43.218 ;
               RECT 15.658 43.782 15.71 43.818 ;
               RECT 15.658 44.382 15.71 44.418 ;
               RECT 15.658 44.982 15.71 45.018 ;
               RECT 15.658 45.582 15.71 45.618 ;
               RECT 15.658 46.182 15.71 46.218 ;
               RECT 15.658 46.782 15.71 46.818 ;
               RECT 15.658 47.382 15.71 47.418 ;
               RECT 15.658 47.982 15.71 48.018 ;
               RECT 15.658 48.582 15.71 48.618 ;
               RECT 15.658 48.942 15.71 48.978 ;
               RECT 15.658 49.422 15.71 49.458 ;
               RECT 15.658 49.902 15.71 49.938 ;
               RECT 15.658 50.382 15.71 50.418 ;
               RECT 15.658 50.862 15.71 50.898 ;
               RECT 15.658 51.342 15.71 51.378 ;
               RECT 15.658 51.822 15.71 51.858 ;
               RECT 15.658 52.302 15.71 52.338 ;
               RECT 15.658 52.662 15.71 52.698 ;
               RECT 15.658 52.782 15.71 52.818 ;
               RECT 15.658 53.262 15.71 53.298 ;
               RECT 15.658 53.742 15.71 53.778 ;
               RECT 15.658 54.2275 15.71 54.2525 ;
               RECT 15.658 54.702 15.71 54.738 ;
               RECT 15.658 55.182 15.71 55.218 ;
               RECT 15.658 55.6675 15.71 55.6925 ;
               RECT 15.658 56.142 15.71 56.178 ;
               RECT 15.658 56.502 15.71 56.538 ;
               RECT 15.658 57.102 15.71 57.138 ;
               RECT 15.658 57.702 15.71 57.738 ;
               RECT 15.658 58.302 15.71 58.338 ;
               RECT 15.658 58.902 15.71 58.938 ;
               RECT 15.658 59.502 15.71 59.538 ;
               RECT 15.658 60.102 15.71 60.138 ;
               RECT 15.658 60.702 15.71 60.738 ;
               RECT 15.658 61.302 15.71 61.338 ;
               RECT 15.658 61.902 15.71 61.938 ;
               RECT 15.658 62.502 15.71 62.538 ;
               RECT 15.658 63.102 15.71 63.138 ;
               RECT 15.658 63.702 15.71 63.738 ;
               RECT 15.658 64.302 15.71 64.338 ;
               RECT 15.658 64.902 15.71 64.938 ;
               RECT 15.658 65.502 15.71 65.538 ;
               RECT 15.658 66.102 15.71 66.138 ;
               RECT 15.658 66.702 15.71 66.738 ;
               RECT 15.658 67.302 15.71 67.338 ;
               RECT 15.658 67.902 15.71 67.938 ;
               RECT 15.658 68.502 15.71 68.538 ;
               RECT 15.658 69.102 15.71 69.138 ;
               RECT 15.658 69.702 15.71 69.738 ;
               RECT 15.658 70.302 15.71 70.338 ;
               RECT 15.658 70.902 15.71 70.938 ;
               RECT 15.658 71.502 15.71 71.538 ;
               RECT 15.658 72.102 15.71 72.138 ;
               RECT 15.658 72.702 15.71 72.738 ;
               RECT 15.658 73.302 15.71 73.338 ;
               RECT 15.658 73.902 15.71 73.938 ;
               RECT 15.658 74.502 15.71 74.538 ;
               RECT 15.658 75.102 15.71 75.138 ;
               RECT 15.658 75.702 15.71 75.738 ;
               RECT 15.658 76.302 15.71 76.338 ;
               RECT 15.658 76.902 15.71 76.938 ;
               RECT 15.658 77.502 15.71 77.538 ;
               RECT 15.658 78.102 15.71 78.138 ;
               RECT 15.658 78.702 15.71 78.738 ;
               RECT 15.658 79.302 15.71 79.338 ;
               RECT 15.658 79.902 15.71 79.938 ;
               RECT 15.658 80.502 15.71 80.538 ;
               RECT 15.658 81.102 15.71 81.138 ;
               RECT 15.658 81.702 15.71 81.738 ;
               RECT 15.658 82.302 15.71 82.338 ;
               RECT 15.658 82.902 15.71 82.938 ;
               RECT 15.658 83.502 15.71 83.538 ;
               RECT 15.658 84.102 15.71 84.138 ;
               RECT 15.658 84.702 15.71 84.738 ;
               RECT 15.658 85.302 15.71 85.338 ;
               RECT 15.658 85.902 15.71 85.938 ;
               RECT 15.658 86.502 15.71 86.538 ;
               RECT 15.658 87.102 15.71 87.138 ;
               RECT 15.658 87.702 15.71 87.738 ;
               RECT 15.658 88.302 15.71 88.338 ;
               RECT 15.658 88.902 15.71 88.938 ;
               RECT 15.658 89.502 15.71 89.538 ;
               RECT 15.658 90.102 15.71 90.138 ;
               RECT 15.658 90.702 15.71 90.738 ;
               RECT 15.658 91.302 15.71 91.338 ;
               RECT 15.658 91.902 15.71 91.938 ;
               RECT 15.658 92.502 15.71 92.538 ;
               RECT 15.658 93.102 15.71 93.138 ;
               RECT 15.658 93.702 15.71 93.738 ;
               RECT 15.658 94.302 15.71 94.338 ;
               RECT 15.658 94.902 15.71 94.938 ;
               RECT 15.658 95.502 15.71 95.538 ;
               RECT 15.658 96.102 15.71 96.138 ;
               RECT 15.658 96.702 15.71 96.738 ;
               RECT 15.658 97.302 15.71 97.338 ;
               RECT 15.658 97.902 15.71 97.938 ;
               RECT 15.658 98.502 15.71 98.538 ;
               RECT 15.658 99.102 15.71 99.138 ;
               RECT 15.658 99.702 15.71 99.738 ;
               RECT 15.658 100.302 15.71 100.338 ;
               RECT 15.658 100.902 15.71 100.938 ;
               RECT 15.658 101.502 15.71 101.538 ;
               RECT 15.658 102.102 15.71 102.138 ;
               RECT 15.658 102.702 15.71 102.738 ;
               RECT 15.658 103.302 15.71 103.338 ;
               RECT 15.658 103.902 15.71 103.938 ;
               RECT 15.658 104.502 15.71 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 15.954 0.5695 16.006 104.5505 ;
               LAYER v4 ;
               RECT 15.954 0.582 16.006 0.618 ;
               RECT 15.954 1.182 16.006 1.218 ;
               RECT 15.954 1.782 16.006 1.818 ;
               RECT 15.954 2.382 16.006 2.418 ;
               RECT 15.954 2.982 16.006 3.018 ;
               RECT 15.954 3.582 16.006 3.618 ;
               RECT 15.954 4.182 16.006 4.218 ;
               RECT 15.954 4.782 16.006 4.818 ;
               RECT 15.954 5.382 16.006 5.418 ;
               RECT 15.954 5.982 16.006 6.018 ;
               RECT 15.954 6.582 16.006 6.618 ;
               RECT 15.954 7.182 16.006 7.218 ;
               RECT 15.954 7.782 16.006 7.818 ;
               RECT 15.954 8.382 16.006 8.418 ;
               RECT 15.954 8.982 16.006 9.018 ;
               RECT 15.954 9.582 16.006 9.618 ;
               RECT 15.954 10.182 16.006 10.218 ;
               RECT 15.954 10.782 16.006 10.818 ;
               RECT 15.954 11.382 16.006 11.418 ;
               RECT 15.954 11.982 16.006 12.018 ;
               RECT 15.954 12.582 16.006 12.618 ;
               RECT 15.954 13.182 16.006 13.218 ;
               RECT 15.954 13.782 16.006 13.818 ;
               RECT 15.954 14.382 16.006 14.418 ;
               RECT 15.954 14.982 16.006 15.018 ;
               RECT 15.954 15.582 16.006 15.618 ;
               RECT 15.954 16.182 16.006 16.218 ;
               RECT 15.954 16.782 16.006 16.818 ;
               RECT 15.954 17.382 16.006 17.418 ;
               RECT 15.954 17.982 16.006 18.018 ;
               RECT 15.954 18.582 16.006 18.618 ;
               RECT 15.954 19.182 16.006 19.218 ;
               RECT 15.954 19.782 16.006 19.818 ;
               RECT 15.954 20.382 16.006 20.418 ;
               RECT 15.954 20.982 16.006 21.018 ;
               RECT 15.954 21.582 16.006 21.618 ;
               RECT 15.954 22.182 16.006 22.218 ;
               RECT 15.954 22.782 16.006 22.818 ;
               RECT 15.954 23.382 16.006 23.418 ;
               RECT 15.954 23.982 16.006 24.018 ;
               RECT 15.954 24.582 16.006 24.618 ;
               RECT 15.954 25.182 16.006 25.218 ;
               RECT 15.954 25.782 16.006 25.818 ;
               RECT 15.954 26.382 16.006 26.418 ;
               RECT 15.954 26.982 16.006 27.018 ;
               RECT 15.954 27.582 16.006 27.618 ;
               RECT 15.954 28.182 16.006 28.218 ;
               RECT 15.954 28.782 16.006 28.818 ;
               RECT 15.954 29.382 16.006 29.418 ;
               RECT 15.954 29.982 16.006 30.018 ;
               RECT 15.954 30.582 16.006 30.618 ;
               RECT 15.954 31.182 16.006 31.218 ;
               RECT 15.954 31.782 16.006 31.818 ;
               RECT 15.954 32.382 16.006 32.418 ;
               RECT 15.954 32.982 16.006 33.018 ;
               RECT 15.954 33.582 16.006 33.618 ;
               RECT 15.954 34.182 16.006 34.218 ;
               RECT 15.954 34.782 16.006 34.818 ;
               RECT 15.954 35.382 16.006 35.418 ;
               RECT 15.954 35.982 16.006 36.018 ;
               RECT 15.954 36.582 16.006 36.618 ;
               RECT 15.954 37.182 16.006 37.218 ;
               RECT 15.954 37.782 16.006 37.818 ;
               RECT 15.954 38.382 16.006 38.418 ;
               RECT 15.954 38.982 16.006 39.018 ;
               RECT 15.954 39.582 16.006 39.618 ;
               RECT 15.954 40.182 16.006 40.218 ;
               RECT 15.954 40.782 16.006 40.818 ;
               RECT 15.954 41.382 16.006 41.418 ;
               RECT 15.954 41.982 16.006 42.018 ;
               RECT 15.954 42.582 16.006 42.618 ;
               RECT 15.954 43.182 16.006 43.218 ;
               RECT 15.954 43.782 16.006 43.818 ;
               RECT 15.954 44.382 16.006 44.418 ;
               RECT 15.954 44.982 16.006 45.018 ;
               RECT 15.954 45.582 16.006 45.618 ;
               RECT 15.954 46.182 16.006 46.218 ;
               RECT 15.954 46.782 16.006 46.818 ;
               RECT 15.954 47.382 16.006 47.418 ;
               RECT 15.954 47.982 16.006 48.018 ;
               RECT 15.954 48.582 16.006 48.618 ;
               RECT 15.954 48.942 16.006 48.978 ;
               RECT 15.954 49.422 16.006 49.458 ;
               RECT 15.954 49.902 16.006 49.938 ;
               RECT 15.954 50.382 16.006 50.418 ;
               RECT 15.954 50.862 16.006 50.898 ;
               RECT 15.954 51.342 16.006 51.378 ;
               RECT 15.954 51.822 16.006 51.858 ;
               RECT 15.954 52.302 16.006 52.338 ;
               RECT 15.954 52.662 16.006 52.698 ;
               RECT 15.954 52.782 16.006 52.818 ;
               RECT 15.954 53.2675 16.006 53.2925 ;
               RECT 15.954 53.742 16.006 53.778 ;
               RECT 15.954 54.222 16.006 54.258 ;
               RECT 15.954 54.702 16.006 54.738 ;
               RECT 15.954 55.182 16.006 55.218 ;
               RECT 15.954 55.662 16.006 55.698 ;
               RECT 15.954 56.142 16.006 56.178 ;
               RECT 15.954 56.502 16.006 56.538 ;
               RECT 15.954 57.102 16.006 57.138 ;
               RECT 15.954 57.702 16.006 57.738 ;
               RECT 15.954 58.302 16.006 58.338 ;
               RECT 15.954 58.902 16.006 58.938 ;
               RECT 15.954 59.502 16.006 59.538 ;
               RECT 15.954 60.102 16.006 60.138 ;
               RECT 15.954 60.702 16.006 60.738 ;
               RECT 15.954 61.302 16.006 61.338 ;
               RECT 15.954 61.902 16.006 61.938 ;
               RECT 15.954 62.502 16.006 62.538 ;
               RECT 15.954 63.102 16.006 63.138 ;
               RECT 15.954 63.702 16.006 63.738 ;
               RECT 15.954 64.302 16.006 64.338 ;
               RECT 15.954 64.902 16.006 64.938 ;
               RECT 15.954 65.502 16.006 65.538 ;
               RECT 15.954 66.102 16.006 66.138 ;
               RECT 15.954 66.702 16.006 66.738 ;
               RECT 15.954 67.302 16.006 67.338 ;
               RECT 15.954 67.902 16.006 67.938 ;
               RECT 15.954 68.502 16.006 68.538 ;
               RECT 15.954 69.102 16.006 69.138 ;
               RECT 15.954 69.702 16.006 69.738 ;
               RECT 15.954 70.302 16.006 70.338 ;
               RECT 15.954 70.902 16.006 70.938 ;
               RECT 15.954 71.502 16.006 71.538 ;
               RECT 15.954 72.102 16.006 72.138 ;
               RECT 15.954 72.702 16.006 72.738 ;
               RECT 15.954 73.302 16.006 73.338 ;
               RECT 15.954 73.902 16.006 73.938 ;
               RECT 15.954 74.502 16.006 74.538 ;
               RECT 15.954 75.102 16.006 75.138 ;
               RECT 15.954 75.702 16.006 75.738 ;
               RECT 15.954 76.302 16.006 76.338 ;
               RECT 15.954 76.902 16.006 76.938 ;
               RECT 15.954 77.502 16.006 77.538 ;
               RECT 15.954 78.102 16.006 78.138 ;
               RECT 15.954 78.702 16.006 78.738 ;
               RECT 15.954 79.302 16.006 79.338 ;
               RECT 15.954 79.902 16.006 79.938 ;
               RECT 15.954 80.502 16.006 80.538 ;
               RECT 15.954 81.102 16.006 81.138 ;
               RECT 15.954 81.702 16.006 81.738 ;
               RECT 15.954 82.302 16.006 82.338 ;
               RECT 15.954 82.902 16.006 82.938 ;
               RECT 15.954 83.502 16.006 83.538 ;
               RECT 15.954 84.102 16.006 84.138 ;
               RECT 15.954 84.702 16.006 84.738 ;
               RECT 15.954 85.302 16.006 85.338 ;
               RECT 15.954 85.902 16.006 85.938 ;
               RECT 15.954 86.502 16.006 86.538 ;
               RECT 15.954 87.102 16.006 87.138 ;
               RECT 15.954 87.702 16.006 87.738 ;
               RECT 15.954 88.302 16.006 88.338 ;
               RECT 15.954 88.902 16.006 88.938 ;
               RECT 15.954 89.502 16.006 89.538 ;
               RECT 15.954 90.102 16.006 90.138 ;
               RECT 15.954 90.702 16.006 90.738 ;
               RECT 15.954 91.302 16.006 91.338 ;
               RECT 15.954 91.902 16.006 91.938 ;
               RECT 15.954 92.502 16.006 92.538 ;
               RECT 15.954 93.102 16.006 93.138 ;
               RECT 15.954 93.702 16.006 93.738 ;
               RECT 15.954 94.302 16.006 94.338 ;
               RECT 15.954 94.902 16.006 94.938 ;
               RECT 15.954 95.502 16.006 95.538 ;
               RECT 15.954 96.102 16.006 96.138 ;
               RECT 15.954 96.702 16.006 96.738 ;
               RECT 15.954 97.302 16.006 97.338 ;
               RECT 15.954 97.902 16.006 97.938 ;
               RECT 15.954 98.502 16.006 98.538 ;
               RECT 15.954 99.102 16.006 99.138 ;
               RECT 15.954 99.702 16.006 99.738 ;
               RECT 15.954 100.302 16.006 100.338 ;
               RECT 15.954 100.902 16.006 100.938 ;
               RECT 15.954 101.502 16.006 101.538 ;
               RECT 15.954 102.102 16.006 102.138 ;
               RECT 15.954 102.702 16.006 102.738 ;
               RECT 15.954 103.302 16.006 103.338 ;
               RECT 15.954 103.902 16.006 103.938 ;
               RECT 15.954 104.502 16.006 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.266 0.5695 16.318 104.5505 ;
               LAYER v4 ;
               RECT 16.266 0.582 16.318 0.618 ;
               RECT 16.266 1.182 16.318 1.218 ;
               RECT 16.266 1.782 16.318 1.818 ;
               RECT 16.266 2.382 16.318 2.418 ;
               RECT 16.266 2.982 16.318 3.018 ;
               RECT 16.266 3.582 16.318 3.618 ;
               RECT 16.266 4.182 16.318 4.218 ;
               RECT 16.266 4.782 16.318 4.818 ;
               RECT 16.266 5.382 16.318 5.418 ;
               RECT 16.266 5.982 16.318 6.018 ;
               RECT 16.266 6.582 16.318 6.618 ;
               RECT 16.266 7.182 16.318 7.218 ;
               RECT 16.266 7.782 16.318 7.818 ;
               RECT 16.266 8.382 16.318 8.418 ;
               RECT 16.266 8.982 16.318 9.018 ;
               RECT 16.266 9.582 16.318 9.618 ;
               RECT 16.266 10.182 16.318 10.218 ;
               RECT 16.266 10.782 16.318 10.818 ;
               RECT 16.266 11.382 16.318 11.418 ;
               RECT 16.266 11.982 16.318 12.018 ;
               RECT 16.266 12.582 16.318 12.618 ;
               RECT 16.266 13.182 16.318 13.218 ;
               RECT 16.266 13.782 16.318 13.818 ;
               RECT 16.266 14.382 16.318 14.418 ;
               RECT 16.266 14.982 16.318 15.018 ;
               RECT 16.266 15.582 16.318 15.618 ;
               RECT 16.266 16.182 16.318 16.218 ;
               RECT 16.266 16.782 16.318 16.818 ;
               RECT 16.266 17.382 16.318 17.418 ;
               RECT 16.266 17.982 16.318 18.018 ;
               RECT 16.266 18.582 16.318 18.618 ;
               RECT 16.266 19.182 16.318 19.218 ;
               RECT 16.266 19.782 16.318 19.818 ;
               RECT 16.266 20.382 16.318 20.418 ;
               RECT 16.266 20.982 16.318 21.018 ;
               RECT 16.266 21.582 16.318 21.618 ;
               RECT 16.266 22.182 16.318 22.218 ;
               RECT 16.266 22.782 16.318 22.818 ;
               RECT 16.266 23.382 16.318 23.418 ;
               RECT 16.266 23.982 16.318 24.018 ;
               RECT 16.266 24.582 16.318 24.618 ;
               RECT 16.266 25.182 16.318 25.218 ;
               RECT 16.266 25.782 16.318 25.818 ;
               RECT 16.266 26.382 16.318 26.418 ;
               RECT 16.266 26.982 16.318 27.018 ;
               RECT 16.266 27.582 16.318 27.618 ;
               RECT 16.266 28.182 16.318 28.218 ;
               RECT 16.266 28.782 16.318 28.818 ;
               RECT 16.266 29.382 16.318 29.418 ;
               RECT 16.266 29.982 16.318 30.018 ;
               RECT 16.266 30.582 16.318 30.618 ;
               RECT 16.266 31.182 16.318 31.218 ;
               RECT 16.266 31.782 16.318 31.818 ;
               RECT 16.266 32.382 16.318 32.418 ;
               RECT 16.266 32.982 16.318 33.018 ;
               RECT 16.266 33.582 16.318 33.618 ;
               RECT 16.266 34.182 16.318 34.218 ;
               RECT 16.266 34.782 16.318 34.818 ;
               RECT 16.266 35.382 16.318 35.418 ;
               RECT 16.266 35.982 16.318 36.018 ;
               RECT 16.266 36.582 16.318 36.618 ;
               RECT 16.266 37.182 16.318 37.218 ;
               RECT 16.266 37.782 16.318 37.818 ;
               RECT 16.266 38.382 16.318 38.418 ;
               RECT 16.266 38.982 16.318 39.018 ;
               RECT 16.266 39.582 16.318 39.618 ;
               RECT 16.266 40.182 16.318 40.218 ;
               RECT 16.266 40.782 16.318 40.818 ;
               RECT 16.266 41.382 16.318 41.418 ;
               RECT 16.266 41.982 16.318 42.018 ;
               RECT 16.266 42.582 16.318 42.618 ;
               RECT 16.266 43.182 16.318 43.218 ;
               RECT 16.266 43.782 16.318 43.818 ;
               RECT 16.266 44.382 16.318 44.418 ;
               RECT 16.266 44.982 16.318 45.018 ;
               RECT 16.266 45.582 16.318 45.618 ;
               RECT 16.266 46.182 16.318 46.218 ;
               RECT 16.266 46.782 16.318 46.818 ;
               RECT 16.266 47.382 16.318 47.418 ;
               RECT 16.266 47.982 16.318 48.018 ;
               RECT 16.266 48.582 16.318 48.618 ;
               RECT 16.266 48.942 16.318 48.978 ;
               RECT 16.266 49.902 16.318 49.938 ;
               RECT 16.266 50.382 16.318 50.418 ;
               RECT 16.266 50.862 16.318 50.898 ;
               RECT 16.266 51.342 16.318 51.378 ;
               RECT 16.266 51.822 16.318 51.858 ;
               RECT 16.266 52.302 16.318 52.338 ;
               RECT 16.266 52.662 16.318 52.698 ;
               RECT 16.266 52.782 16.318 52.818 ;
               RECT 16.266 53.262 16.318 53.298 ;
               RECT 16.266 53.742 16.318 53.778 ;
               RECT 16.266 54.222 16.318 54.258 ;
               RECT 16.266 54.702 16.318 54.738 ;
               RECT 16.266 55.662 16.318 55.698 ;
               RECT 16.266 56.142 16.318 56.178 ;
               RECT 16.266 56.502 16.318 56.538 ;
               RECT 16.266 57.102 16.318 57.138 ;
               RECT 16.266 57.702 16.318 57.738 ;
               RECT 16.266 58.302 16.318 58.338 ;
               RECT 16.266 58.902 16.318 58.938 ;
               RECT 16.266 59.502 16.318 59.538 ;
               RECT 16.266 60.102 16.318 60.138 ;
               RECT 16.266 60.702 16.318 60.738 ;
               RECT 16.266 61.302 16.318 61.338 ;
               RECT 16.266 61.902 16.318 61.938 ;
               RECT 16.266 62.502 16.318 62.538 ;
               RECT 16.266 63.102 16.318 63.138 ;
               RECT 16.266 63.702 16.318 63.738 ;
               RECT 16.266 64.302 16.318 64.338 ;
               RECT 16.266 64.902 16.318 64.938 ;
               RECT 16.266 65.502 16.318 65.538 ;
               RECT 16.266 66.102 16.318 66.138 ;
               RECT 16.266 66.702 16.318 66.738 ;
               RECT 16.266 67.302 16.318 67.338 ;
               RECT 16.266 67.902 16.318 67.938 ;
               RECT 16.266 68.502 16.318 68.538 ;
               RECT 16.266 69.102 16.318 69.138 ;
               RECT 16.266 69.702 16.318 69.738 ;
               RECT 16.266 70.302 16.318 70.338 ;
               RECT 16.266 70.902 16.318 70.938 ;
               RECT 16.266 71.502 16.318 71.538 ;
               RECT 16.266 72.102 16.318 72.138 ;
               RECT 16.266 72.702 16.318 72.738 ;
               RECT 16.266 73.302 16.318 73.338 ;
               RECT 16.266 73.902 16.318 73.938 ;
               RECT 16.266 74.502 16.318 74.538 ;
               RECT 16.266 75.102 16.318 75.138 ;
               RECT 16.266 75.702 16.318 75.738 ;
               RECT 16.266 76.302 16.318 76.338 ;
               RECT 16.266 76.902 16.318 76.938 ;
               RECT 16.266 77.502 16.318 77.538 ;
               RECT 16.266 78.102 16.318 78.138 ;
               RECT 16.266 78.702 16.318 78.738 ;
               RECT 16.266 79.302 16.318 79.338 ;
               RECT 16.266 79.902 16.318 79.938 ;
               RECT 16.266 80.502 16.318 80.538 ;
               RECT 16.266 81.102 16.318 81.138 ;
               RECT 16.266 81.702 16.318 81.738 ;
               RECT 16.266 82.302 16.318 82.338 ;
               RECT 16.266 82.902 16.318 82.938 ;
               RECT 16.266 83.502 16.318 83.538 ;
               RECT 16.266 84.102 16.318 84.138 ;
               RECT 16.266 84.702 16.318 84.738 ;
               RECT 16.266 85.302 16.318 85.338 ;
               RECT 16.266 85.902 16.318 85.938 ;
               RECT 16.266 86.502 16.318 86.538 ;
               RECT 16.266 87.102 16.318 87.138 ;
               RECT 16.266 87.702 16.318 87.738 ;
               RECT 16.266 88.302 16.318 88.338 ;
               RECT 16.266 88.902 16.318 88.938 ;
               RECT 16.266 89.502 16.318 89.538 ;
               RECT 16.266 90.102 16.318 90.138 ;
               RECT 16.266 90.702 16.318 90.738 ;
               RECT 16.266 91.302 16.318 91.338 ;
               RECT 16.266 91.902 16.318 91.938 ;
               RECT 16.266 92.502 16.318 92.538 ;
               RECT 16.266 93.102 16.318 93.138 ;
               RECT 16.266 93.702 16.318 93.738 ;
               RECT 16.266 94.302 16.318 94.338 ;
               RECT 16.266 94.902 16.318 94.938 ;
               RECT 16.266 95.502 16.318 95.538 ;
               RECT 16.266 96.102 16.318 96.138 ;
               RECT 16.266 96.702 16.318 96.738 ;
               RECT 16.266 97.302 16.318 97.338 ;
               RECT 16.266 97.902 16.318 97.938 ;
               RECT 16.266 98.502 16.318 98.538 ;
               RECT 16.266 99.102 16.318 99.138 ;
               RECT 16.266 99.702 16.318 99.738 ;
               RECT 16.266 100.302 16.318 100.338 ;
               RECT 16.266 100.902 16.318 100.938 ;
               RECT 16.266 101.502 16.318 101.538 ;
               RECT 16.266 102.102 16.318 102.138 ;
               RECT 16.266 102.702 16.318 102.738 ;
               RECT 16.266 103.302 16.318 103.338 ;
               RECT 16.266 103.902 16.318 103.938 ;
               RECT 16.266 104.502 16.318 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.498 0.5695 16.55 104.5505 ;
               LAYER v4 ;
               RECT 16.498 0.582 16.55 0.618 ;
               RECT 16.498 1.182 16.55 1.218 ;
               RECT 16.498 1.782 16.55 1.818 ;
               RECT 16.498 2.382 16.55 2.418 ;
               RECT 16.498 2.982 16.55 3.018 ;
               RECT 16.498 3.582 16.55 3.618 ;
               RECT 16.498 4.182 16.55 4.218 ;
               RECT 16.498 4.782 16.55 4.818 ;
               RECT 16.498 5.382 16.55 5.418 ;
               RECT 16.498 5.982 16.55 6.018 ;
               RECT 16.498 6.582 16.55 6.618 ;
               RECT 16.498 7.182 16.55 7.218 ;
               RECT 16.498 7.782 16.55 7.818 ;
               RECT 16.498 8.382 16.55 8.418 ;
               RECT 16.498 8.982 16.55 9.018 ;
               RECT 16.498 9.582 16.55 9.618 ;
               RECT 16.498 10.182 16.55 10.218 ;
               RECT 16.498 10.782 16.55 10.818 ;
               RECT 16.498 11.382 16.55 11.418 ;
               RECT 16.498 11.982 16.55 12.018 ;
               RECT 16.498 12.582 16.55 12.618 ;
               RECT 16.498 13.182 16.55 13.218 ;
               RECT 16.498 13.782 16.55 13.818 ;
               RECT 16.498 14.382 16.55 14.418 ;
               RECT 16.498 14.982 16.55 15.018 ;
               RECT 16.498 15.582 16.55 15.618 ;
               RECT 16.498 16.182 16.55 16.218 ;
               RECT 16.498 16.782 16.55 16.818 ;
               RECT 16.498 17.382 16.55 17.418 ;
               RECT 16.498 17.982 16.55 18.018 ;
               RECT 16.498 18.582 16.55 18.618 ;
               RECT 16.498 19.182 16.55 19.218 ;
               RECT 16.498 19.782 16.55 19.818 ;
               RECT 16.498 20.382 16.55 20.418 ;
               RECT 16.498 20.982 16.55 21.018 ;
               RECT 16.498 21.582 16.55 21.618 ;
               RECT 16.498 22.182 16.55 22.218 ;
               RECT 16.498 22.782 16.55 22.818 ;
               RECT 16.498 23.382 16.55 23.418 ;
               RECT 16.498 23.982 16.55 24.018 ;
               RECT 16.498 24.582 16.55 24.618 ;
               RECT 16.498 25.182 16.55 25.218 ;
               RECT 16.498 25.782 16.55 25.818 ;
               RECT 16.498 26.382 16.55 26.418 ;
               RECT 16.498 26.982 16.55 27.018 ;
               RECT 16.498 27.582 16.55 27.618 ;
               RECT 16.498 28.182 16.55 28.218 ;
               RECT 16.498 28.782 16.55 28.818 ;
               RECT 16.498 29.382 16.55 29.418 ;
               RECT 16.498 29.982 16.55 30.018 ;
               RECT 16.498 30.582 16.55 30.618 ;
               RECT 16.498 31.182 16.55 31.218 ;
               RECT 16.498 31.782 16.55 31.818 ;
               RECT 16.498 32.382 16.55 32.418 ;
               RECT 16.498 32.982 16.55 33.018 ;
               RECT 16.498 33.582 16.55 33.618 ;
               RECT 16.498 34.182 16.55 34.218 ;
               RECT 16.498 34.782 16.55 34.818 ;
               RECT 16.498 35.382 16.55 35.418 ;
               RECT 16.498 35.982 16.55 36.018 ;
               RECT 16.498 36.582 16.55 36.618 ;
               RECT 16.498 37.182 16.55 37.218 ;
               RECT 16.498 37.782 16.55 37.818 ;
               RECT 16.498 38.382 16.55 38.418 ;
               RECT 16.498 38.982 16.55 39.018 ;
               RECT 16.498 39.582 16.55 39.618 ;
               RECT 16.498 40.182 16.55 40.218 ;
               RECT 16.498 40.782 16.55 40.818 ;
               RECT 16.498 41.382 16.55 41.418 ;
               RECT 16.498 41.982 16.55 42.018 ;
               RECT 16.498 42.582 16.55 42.618 ;
               RECT 16.498 43.182 16.55 43.218 ;
               RECT 16.498 43.782 16.55 43.818 ;
               RECT 16.498 44.382 16.55 44.418 ;
               RECT 16.498 44.982 16.55 45.018 ;
               RECT 16.498 45.582 16.55 45.618 ;
               RECT 16.498 46.182 16.55 46.218 ;
               RECT 16.498 46.782 16.55 46.818 ;
               RECT 16.498 47.382 16.55 47.418 ;
               RECT 16.498 47.982 16.55 48.018 ;
               RECT 16.498 48.582 16.55 48.618 ;
               RECT 16.498 48.942 16.55 48.978 ;
               RECT 16.498 49.422 16.55 49.458 ;
               RECT 16.498 49.902 16.55 49.938 ;
               RECT 16.498 50.382 16.55 50.418 ;
               RECT 16.498 50.862 16.55 50.898 ;
               RECT 16.498 51.342 16.55 51.378 ;
               RECT 16.498 51.822 16.55 51.858 ;
               RECT 16.498 52.302 16.55 52.338 ;
               RECT 16.498 52.662 16.55 52.698 ;
               RECT 16.498 52.782 16.55 52.818 ;
               RECT 16.498 53.262 16.55 53.298 ;
               RECT 16.498 53.742 16.55 53.778 ;
               RECT 16.498 54.222 16.55 54.258 ;
               RECT 16.498 54.702 16.55 54.738 ;
               RECT 16.498 55.182 16.55 55.218 ;
               RECT 16.498 55.662 16.55 55.698 ;
               RECT 16.498 56.142 16.55 56.178 ;
               RECT 16.498 56.502 16.55 56.538 ;
               RECT 16.498 57.102 16.55 57.138 ;
               RECT 16.498 57.702 16.55 57.738 ;
               RECT 16.498 58.302 16.55 58.338 ;
               RECT 16.498 58.902 16.55 58.938 ;
               RECT 16.498 59.502 16.55 59.538 ;
               RECT 16.498 60.102 16.55 60.138 ;
               RECT 16.498 60.702 16.55 60.738 ;
               RECT 16.498 61.302 16.55 61.338 ;
               RECT 16.498 61.902 16.55 61.938 ;
               RECT 16.498 62.502 16.55 62.538 ;
               RECT 16.498 63.102 16.55 63.138 ;
               RECT 16.498 63.702 16.55 63.738 ;
               RECT 16.498 64.302 16.55 64.338 ;
               RECT 16.498 64.902 16.55 64.938 ;
               RECT 16.498 65.502 16.55 65.538 ;
               RECT 16.498 66.102 16.55 66.138 ;
               RECT 16.498 66.702 16.55 66.738 ;
               RECT 16.498 67.302 16.55 67.338 ;
               RECT 16.498 67.902 16.55 67.938 ;
               RECT 16.498 68.502 16.55 68.538 ;
               RECT 16.498 69.102 16.55 69.138 ;
               RECT 16.498 69.702 16.55 69.738 ;
               RECT 16.498 70.302 16.55 70.338 ;
               RECT 16.498 70.902 16.55 70.938 ;
               RECT 16.498 71.502 16.55 71.538 ;
               RECT 16.498 72.102 16.55 72.138 ;
               RECT 16.498 72.702 16.55 72.738 ;
               RECT 16.498 73.302 16.55 73.338 ;
               RECT 16.498 73.902 16.55 73.938 ;
               RECT 16.498 74.502 16.55 74.538 ;
               RECT 16.498 75.102 16.55 75.138 ;
               RECT 16.498 75.702 16.55 75.738 ;
               RECT 16.498 76.302 16.55 76.338 ;
               RECT 16.498 76.902 16.55 76.938 ;
               RECT 16.498 77.502 16.55 77.538 ;
               RECT 16.498 78.102 16.55 78.138 ;
               RECT 16.498 78.702 16.55 78.738 ;
               RECT 16.498 79.302 16.55 79.338 ;
               RECT 16.498 79.902 16.55 79.938 ;
               RECT 16.498 80.502 16.55 80.538 ;
               RECT 16.498 81.102 16.55 81.138 ;
               RECT 16.498 81.702 16.55 81.738 ;
               RECT 16.498 82.302 16.55 82.338 ;
               RECT 16.498 82.902 16.55 82.938 ;
               RECT 16.498 83.502 16.55 83.538 ;
               RECT 16.498 84.102 16.55 84.138 ;
               RECT 16.498 84.702 16.55 84.738 ;
               RECT 16.498 85.302 16.55 85.338 ;
               RECT 16.498 85.902 16.55 85.938 ;
               RECT 16.498 86.502 16.55 86.538 ;
               RECT 16.498 87.102 16.55 87.138 ;
               RECT 16.498 87.702 16.55 87.738 ;
               RECT 16.498 88.302 16.55 88.338 ;
               RECT 16.498 88.902 16.55 88.938 ;
               RECT 16.498 89.502 16.55 89.538 ;
               RECT 16.498 90.102 16.55 90.138 ;
               RECT 16.498 90.702 16.55 90.738 ;
               RECT 16.498 91.302 16.55 91.338 ;
               RECT 16.498 91.902 16.55 91.938 ;
               RECT 16.498 92.502 16.55 92.538 ;
               RECT 16.498 93.102 16.55 93.138 ;
               RECT 16.498 93.702 16.55 93.738 ;
               RECT 16.498 94.302 16.55 94.338 ;
               RECT 16.498 94.902 16.55 94.938 ;
               RECT 16.498 95.502 16.55 95.538 ;
               RECT 16.498 96.102 16.55 96.138 ;
               RECT 16.498 96.702 16.55 96.738 ;
               RECT 16.498 97.302 16.55 97.338 ;
               RECT 16.498 97.902 16.55 97.938 ;
               RECT 16.498 98.502 16.55 98.538 ;
               RECT 16.498 99.102 16.55 99.138 ;
               RECT 16.498 99.702 16.55 99.738 ;
               RECT 16.498 100.302 16.55 100.338 ;
               RECT 16.498 100.902 16.55 100.938 ;
               RECT 16.498 101.502 16.55 101.538 ;
               RECT 16.498 102.102 16.55 102.138 ;
               RECT 16.498 102.702 16.55 102.738 ;
               RECT 16.498 103.302 16.55 103.338 ;
               RECT 16.498 103.902 16.55 103.938 ;
               RECT 16.498 104.502 16.55 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 16.882 49.153 16.936 55.9925 ;
               LAYER v4 ;
               RECT 16.882 49.422 16.936 49.458 ;
               RECT 16.882 50.3875 16.936 50.4125 ;
               RECT 16.882 50.862 16.936 50.898 ;
               RECT 16.882 51.3475 16.936 51.3725 ;
               RECT 16.882 51.822 16.936 51.858 ;
               RECT 16.882 52.3075 16.936 52.3325 ;
               RECT 16.882 52.662 16.936 52.698 ;
               RECT 16.882 52.782 16.936 52.818 ;
               RECT 16.882 53.262 16.936 53.298 ;
               RECT 16.882 53.7475 16.936 53.7725 ;
               RECT 16.882 54.2275 16.936 54.2525 ;
               RECT 16.882 54.7075 16.936 54.7325 ;
               RECT 16.882 55.182 16.936 55.218 ;
               RECT 16.882 55.662 16.936 55.698 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.204 48.62 17.244 56.5 ;
               LAYER v4 ;
               RECT 17.204 48.942 17.244 48.978 ;
               RECT 17.204 49.422 17.244 49.458 ;
               RECT 17.204 49.7205 17.244 49.7565 ;
               RECT 17.204 49.902 17.244 49.938 ;
               RECT 17.204 50.382 17.244 50.418 ;
               RECT 17.204 50.862 17.244 50.898 ;
               RECT 17.204 51.342 17.244 51.378 ;
               RECT 17.204 51.822 17.244 51.858 ;
               RECT 17.204 52.302 17.244 52.338 ;
               RECT 17.204 52.662 17.244 52.698 ;
               RECT 17.204 52.782 17.244 52.818 ;
               RECT 17.204 53.262 17.244 53.298 ;
               RECT 17.204 53.742 17.244 53.778 ;
               RECT 17.204 54.222 17.244 54.258 ;
               RECT 17.204 54.702 17.244 54.738 ;
               RECT 17.204 55.182 17.244 55.218 ;
               RECT 17.204 55.662 17.244 55.698 ;
               RECT 17.204 56.142 17.244 56.178 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.344 0.5695 17.384 48.94 ;
               LAYER v4 ;
               RECT 17.344 0.582 17.384 0.618 ;
               RECT 17.344 1.182 17.384 1.218 ;
               RECT 17.344 1.782 17.384 1.818 ;
               RECT 17.344 2.382 17.384 2.418 ;
               RECT 17.344 2.982 17.384 3.018 ;
               RECT 17.344 3.582 17.384 3.618 ;
               RECT 17.344 4.182 17.384 4.218 ;
               RECT 17.344 4.782 17.384 4.818 ;
               RECT 17.344 5.382 17.384 5.418 ;
               RECT 17.344 5.982 17.384 6.018 ;
               RECT 17.344 6.582 17.384 6.618 ;
               RECT 17.344 7.182 17.384 7.218 ;
               RECT 17.344 7.782 17.384 7.818 ;
               RECT 17.344 8.382 17.384 8.418 ;
               RECT 17.344 8.982 17.384 9.018 ;
               RECT 17.344 9.582 17.384 9.618 ;
               RECT 17.344 10.182 17.384 10.218 ;
               RECT 17.344 10.782 17.384 10.818 ;
               RECT 17.344 11.382 17.384 11.418 ;
               RECT 17.344 11.982 17.384 12.018 ;
               RECT 17.344 12.582 17.384 12.618 ;
               RECT 17.344 13.182 17.384 13.218 ;
               RECT 17.344 13.782 17.384 13.818 ;
               RECT 17.344 14.382 17.384 14.418 ;
               RECT 17.344 14.982 17.384 15.018 ;
               RECT 17.344 15.582 17.384 15.618 ;
               RECT 17.344 16.182 17.384 16.218 ;
               RECT 17.344 16.782 17.384 16.818 ;
               RECT 17.344 17.382 17.384 17.418 ;
               RECT 17.344 17.982 17.384 18.018 ;
               RECT 17.344 18.582 17.384 18.618 ;
               RECT 17.344 19.182 17.384 19.218 ;
               RECT 17.344 19.782 17.384 19.818 ;
               RECT 17.344 20.382 17.384 20.418 ;
               RECT 17.344 20.982 17.384 21.018 ;
               RECT 17.344 21.582 17.384 21.618 ;
               RECT 17.344 22.182 17.384 22.218 ;
               RECT 17.344 22.782 17.384 22.818 ;
               RECT 17.344 23.382 17.384 23.418 ;
               RECT 17.344 23.982 17.384 24.018 ;
               RECT 17.344 24.582 17.384 24.618 ;
               RECT 17.344 25.182 17.384 25.218 ;
               RECT 17.344 25.782 17.384 25.818 ;
               RECT 17.344 26.382 17.384 26.418 ;
               RECT 17.344 26.982 17.384 27.018 ;
               RECT 17.344 27.582 17.384 27.618 ;
               RECT 17.344 28.182 17.384 28.218 ;
               RECT 17.344 28.782 17.384 28.818 ;
               RECT 17.344 29.382 17.384 29.418 ;
               RECT 17.344 29.982 17.384 30.018 ;
               RECT 17.344 30.582 17.384 30.618 ;
               RECT 17.344 31.182 17.384 31.218 ;
               RECT 17.344 31.782 17.384 31.818 ;
               RECT 17.344 32.382 17.384 32.418 ;
               RECT 17.344 32.982 17.384 33.018 ;
               RECT 17.344 33.582 17.384 33.618 ;
               RECT 17.344 34.182 17.384 34.218 ;
               RECT 17.344 34.782 17.384 34.818 ;
               RECT 17.344 35.382 17.384 35.418 ;
               RECT 17.344 35.982 17.384 36.018 ;
               RECT 17.344 36.582 17.384 36.618 ;
               RECT 17.344 37.182 17.384 37.218 ;
               RECT 17.344 37.782 17.384 37.818 ;
               RECT 17.344 38.382 17.384 38.418 ;
               RECT 17.344 38.982 17.384 39.018 ;
               RECT 17.344 39.582 17.384 39.618 ;
               RECT 17.344 40.182 17.384 40.218 ;
               RECT 17.344 40.782 17.384 40.818 ;
               RECT 17.344 41.382 17.384 41.418 ;
               RECT 17.344 41.982 17.384 42.018 ;
               RECT 17.344 42.582 17.384 42.618 ;
               RECT 17.344 43.182 17.384 43.218 ;
               RECT 17.344 43.782 17.384 43.818 ;
               RECT 17.344 44.382 17.384 44.418 ;
               RECT 17.344 44.982 17.384 45.018 ;
               RECT 17.344 45.582 17.384 45.618 ;
               RECT 17.344 46.182 17.384 46.218 ;
               RECT 17.344 46.782 17.384 46.818 ;
               RECT 17.344 47.382 17.384 47.418 ;
               RECT 17.344 47.982 17.384 48.018 ;
               RECT 17.344 48.582 17.384 48.618 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.344 56.18 17.384 104.5505 ;
               LAYER v4 ;
               RECT 17.344 56.502 17.384 56.538 ;
               RECT 17.344 57.102 17.384 57.138 ;
               RECT 17.344 57.702 17.384 57.738 ;
               RECT 17.344 58.302 17.384 58.338 ;
               RECT 17.344 58.902 17.384 58.938 ;
               RECT 17.344 59.502 17.384 59.538 ;
               RECT 17.344 60.102 17.384 60.138 ;
               RECT 17.344 60.702 17.384 60.738 ;
               RECT 17.344 61.302 17.384 61.338 ;
               RECT 17.344 61.902 17.384 61.938 ;
               RECT 17.344 62.502 17.384 62.538 ;
               RECT 17.344 63.102 17.384 63.138 ;
               RECT 17.344 63.702 17.384 63.738 ;
               RECT 17.344 64.302 17.384 64.338 ;
               RECT 17.344 64.902 17.384 64.938 ;
               RECT 17.344 65.502 17.384 65.538 ;
               RECT 17.344 66.102 17.384 66.138 ;
               RECT 17.344 66.702 17.384 66.738 ;
               RECT 17.344 67.302 17.384 67.338 ;
               RECT 17.344 67.902 17.384 67.938 ;
               RECT 17.344 68.502 17.384 68.538 ;
               RECT 17.344 69.102 17.384 69.138 ;
               RECT 17.344 69.702 17.384 69.738 ;
               RECT 17.344 70.302 17.384 70.338 ;
               RECT 17.344 70.902 17.384 70.938 ;
               RECT 17.344 71.502 17.384 71.538 ;
               RECT 17.344 72.102 17.384 72.138 ;
               RECT 17.344 72.702 17.384 72.738 ;
               RECT 17.344 73.302 17.384 73.338 ;
               RECT 17.344 73.902 17.384 73.938 ;
               RECT 17.344 74.502 17.384 74.538 ;
               RECT 17.344 75.102 17.384 75.138 ;
               RECT 17.344 75.702 17.384 75.738 ;
               RECT 17.344 76.302 17.384 76.338 ;
               RECT 17.344 76.902 17.384 76.938 ;
               RECT 17.344 77.502 17.384 77.538 ;
               RECT 17.344 78.102 17.384 78.138 ;
               RECT 17.344 78.702 17.384 78.738 ;
               RECT 17.344 79.302 17.384 79.338 ;
               RECT 17.344 79.902 17.384 79.938 ;
               RECT 17.344 80.502 17.384 80.538 ;
               RECT 17.344 81.102 17.384 81.138 ;
               RECT 17.344 81.702 17.384 81.738 ;
               RECT 17.344 82.302 17.384 82.338 ;
               RECT 17.344 82.902 17.384 82.938 ;
               RECT 17.344 83.502 17.384 83.538 ;
               RECT 17.344 84.102 17.384 84.138 ;
               RECT 17.344 84.702 17.384 84.738 ;
               RECT 17.344 85.302 17.384 85.338 ;
               RECT 17.344 85.902 17.384 85.938 ;
               RECT 17.344 86.502 17.384 86.538 ;
               RECT 17.344 87.102 17.384 87.138 ;
               RECT 17.344 87.702 17.384 87.738 ;
               RECT 17.344 88.302 17.384 88.338 ;
               RECT 17.344 88.902 17.384 88.938 ;
               RECT 17.344 89.502 17.384 89.538 ;
               RECT 17.344 90.102 17.384 90.138 ;
               RECT 17.344 90.702 17.384 90.738 ;
               RECT 17.344 91.302 17.384 91.338 ;
               RECT 17.344 91.902 17.384 91.938 ;
               RECT 17.344 92.502 17.384 92.538 ;
               RECT 17.344 93.102 17.384 93.138 ;
               RECT 17.344 93.702 17.384 93.738 ;
               RECT 17.344 94.302 17.384 94.338 ;
               RECT 17.344 94.902 17.384 94.938 ;
               RECT 17.344 95.502 17.384 95.538 ;
               RECT 17.344 96.102 17.384 96.138 ;
               RECT 17.344 96.702 17.384 96.738 ;
               RECT 17.344 97.302 17.384 97.338 ;
               RECT 17.344 97.902 17.384 97.938 ;
               RECT 17.344 98.502 17.384 98.538 ;
               RECT 17.344 99.102 17.384 99.138 ;
               RECT 17.344 99.702 17.384 99.738 ;
               RECT 17.344 100.302 17.384 100.338 ;
               RECT 17.344 100.902 17.384 100.938 ;
               RECT 17.344 101.502 17.384 101.538 ;
               RECT 17.344 102.102 17.384 102.138 ;
               RECT 17.344 102.702 17.384 102.738 ;
               RECT 17.344 103.302 17.384 103.338 ;
               RECT 17.344 103.902 17.384 103.938 ;
               RECT 17.344 104.502 17.384 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 17.684 0.5695 17.736 104.5505 ;
               LAYER v4 ;
               RECT 17.684 0.582 17.736 0.618 ;
               RECT 17.684 1.182 17.736 1.218 ;
               RECT 17.684 1.782 17.736 1.818 ;
               RECT 17.684 2.382 17.736 2.418 ;
               RECT 17.684 2.982 17.736 3.018 ;
               RECT 17.684 3.582 17.736 3.618 ;
               RECT 17.684 4.182 17.736 4.218 ;
               RECT 17.684 4.782 17.736 4.818 ;
               RECT 17.684 5.382 17.736 5.418 ;
               RECT 17.684 5.982 17.736 6.018 ;
               RECT 17.684 6.582 17.736 6.618 ;
               RECT 17.684 7.182 17.736 7.218 ;
               RECT 17.684 7.782 17.736 7.818 ;
               RECT 17.684 8.382 17.736 8.418 ;
               RECT 17.684 8.982 17.736 9.018 ;
               RECT 17.684 9.582 17.736 9.618 ;
               RECT 17.684 10.182 17.736 10.218 ;
               RECT 17.684 10.782 17.736 10.818 ;
               RECT 17.684 11.382 17.736 11.418 ;
               RECT 17.684 11.982 17.736 12.018 ;
               RECT 17.684 12.582 17.736 12.618 ;
               RECT 17.684 13.182 17.736 13.218 ;
               RECT 17.684 13.782 17.736 13.818 ;
               RECT 17.684 14.382 17.736 14.418 ;
               RECT 17.684 14.982 17.736 15.018 ;
               RECT 17.684 15.582 17.736 15.618 ;
               RECT 17.684 16.182 17.736 16.218 ;
               RECT 17.684 16.782 17.736 16.818 ;
               RECT 17.684 17.382 17.736 17.418 ;
               RECT 17.684 17.982 17.736 18.018 ;
               RECT 17.684 18.582 17.736 18.618 ;
               RECT 17.684 19.182 17.736 19.218 ;
               RECT 17.684 19.782 17.736 19.818 ;
               RECT 17.684 20.382 17.736 20.418 ;
               RECT 17.684 20.982 17.736 21.018 ;
               RECT 17.684 21.582 17.736 21.618 ;
               RECT 17.684 22.182 17.736 22.218 ;
               RECT 17.684 22.782 17.736 22.818 ;
               RECT 17.684 23.382 17.736 23.418 ;
               RECT 17.684 23.982 17.736 24.018 ;
               RECT 17.684 24.582 17.736 24.618 ;
               RECT 17.684 25.182 17.736 25.218 ;
               RECT 17.684 25.782 17.736 25.818 ;
               RECT 17.684 26.382 17.736 26.418 ;
               RECT 17.684 26.982 17.736 27.018 ;
               RECT 17.684 27.582 17.736 27.618 ;
               RECT 17.684 28.182 17.736 28.218 ;
               RECT 17.684 28.782 17.736 28.818 ;
               RECT 17.684 29.382 17.736 29.418 ;
               RECT 17.684 29.982 17.736 30.018 ;
               RECT 17.684 30.582 17.736 30.618 ;
               RECT 17.684 31.182 17.736 31.218 ;
               RECT 17.684 31.782 17.736 31.818 ;
               RECT 17.684 32.382 17.736 32.418 ;
               RECT 17.684 32.982 17.736 33.018 ;
               RECT 17.684 33.582 17.736 33.618 ;
               RECT 17.684 34.182 17.736 34.218 ;
               RECT 17.684 34.782 17.736 34.818 ;
               RECT 17.684 35.382 17.736 35.418 ;
               RECT 17.684 35.982 17.736 36.018 ;
               RECT 17.684 36.582 17.736 36.618 ;
               RECT 17.684 37.182 17.736 37.218 ;
               RECT 17.684 37.782 17.736 37.818 ;
               RECT 17.684 38.382 17.736 38.418 ;
               RECT 17.684 38.982 17.736 39.018 ;
               RECT 17.684 39.582 17.736 39.618 ;
               RECT 17.684 40.182 17.736 40.218 ;
               RECT 17.684 40.782 17.736 40.818 ;
               RECT 17.684 41.382 17.736 41.418 ;
               RECT 17.684 41.982 17.736 42.018 ;
               RECT 17.684 42.582 17.736 42.618 ;
               RECT 17.684 43.182 17.736 43.218 ;
               RECT 17.684 43.782 17.736 43.818 ;
               RECT 17.684 44.382 17.736 44.418 ;
               RECT 17.684 44.982 17.736 45.018 ;
               RECT 17.684 45.582 17.736 45.618 ;
               RECT 17.684 46.182 17.736 46.218 ;
               RECT 17.684 46.782 17.736 46.818 ;
               RECT 17.684 47.382 17.736 47.418 ;
               RECT 17.684 47.982 17.736 48.018 ;
               RECT 17.684 48.582 17.736 48.618 ;
               RECT 17.684 48.942 17.736 48.978 ;
               RECT 17.684 49.422 17.736 49.458 ;
               RECT 17.684 49.7205 17.736 49.7565 ;
               RECT 17.684 49.902 17.736 49.938 ;
               RECT 17.684 50.382 17.736 50.418 ;
               RECT 17.684 50.862 17.736 50.898 ;
               RECT 17.684 51.342 17.736 51.378 ;
               RECT 17.684 51.822 17.736 51.858 ;
               RECT 17.684 52.302 17.736 52.338 ;
               RECT 17.684 52.782 17.736 52.818 ;
               RECT 17.684 53.262 17.736 53.298 ;
               RECT 17.684 53.742 17.736 53.778 ;
               RECT 17.684 54.222 17.736 54.258 ;
               RECT 17.684 54.702 17.736 54.738 ;
               RECT 17.684 55.182 17.736 55.218 ;
               RECT 17.684 55.662 17.736 55.698 ;
               RECT 17.684 56.142 17.736 56.178 ;
               RECT 17.684 56.502 17.736 56.538 ;
               RECT 17.684 57.102 17.736 57.138 ;
               RECT 17.684 57.702 17.736 57.738 ;
               RECT 17.684 58.302 17.736 58.338 ;
               RECT 17.684 58.902 17.736 58.938 ;
               RECT 17.684 59.502 17.736 59.538 ;
               RECT 17.684 60.102 17.736 60.138 ;
               RECT 17.684 60.702 17.736 60.738 ;
               RECT 17.684 61.302 17.736 61.338 ;
               RECT 17.684 61.902 17.736 61.938 ;
               RECT 17.684 62.502 17.736 62.538 ;
               RECT 17.684 63.102 17.736 63.138 ;
               RECT 17.684 63.702 17.736 63.738 ;
               RECT 17.684 64.302 17.736 64.338 ;
               RECT 17.684 64.902 17.736 64.938 ;
               RECT 17.684 65.502 17.736 65.538 ;
               RECT 17.684 66.102 17.736 66.138 ;
               RECT 17.684 66.702 17.736 66.738 ;
               RECT 17.684 67.302 17.736 67.338 ;
               RECT 17.684 67.902 17.736 67.938 ;
               RECT 17.684 68.502 17.736 68.538 ;
               RECT 17.684 69.102 17.736 69.138 ;
               RECT 17.684 69.702 17.736 69.738 ;
               RECT 17.684 70.302 17.736 70.338 ;
               RECT 17.684 70.902 17.736 70.938 ;
               RECT 17.684 71.502 17.736 71.538 ;
               RECT 17.684 72.102 17.736 72.138 ;
               RECT 17.684 72.702 17.736 72.738 ;
               RECT 17.684 73.302 17.736 73.338 ;
               RECT 17.684 73.902 17.736 73.938 ;
               RECT 17.684 74.502 17.736 74.538 ;
               RECT 17.684 75.102 17.736 75.138 ;
               RECT 17.684 75.702 17.736 75.738 ;
               RECT 17.684 76.302 17.736 76.338 ;
               RECT 17.684 76.902 17.736 76.938 ;
               RECT 17.684 77.502 17.736 77.538 ;
               RECT 17.684 78.102 17.736 78.138 ;
               RECT 17.684 78.702 17.736 78.738 ;
               RECT 17.684 79.302 17.736 79.338 ;
               RECT 17.684 79.902 17.736 79.938 ;
               RECT 17.684 80.502 17.736 80.538 ;
               RECT 17.684 81.102 17.736 81.138 ;
               RECT 17.684 81.702 17.736 81.738 ;
               RECT 17.684 82.302 17.736 82.338 ;
               RECT 17.684 82.902 17.736 82.938 ;
               RECT 17.684 83.502 17.736 83.538 ;
               RECT 17.684 84.102 17.736 84.138 ;
               RECT 17.684 84.702 17.736 84.738 ;
               RECT 17.684 85.302 17.736 85.338 ;
               RECT 17.684 85.902 17.736 85.938 ;
               RECT 17.684 86.502 17.736 86.538 ;
               RECT 17.684 87.102 17.736 87.138 ;
               RECT 17.684 87.702 17.736 87.738 ;
               RECT 17.684 88.302 17.736 88.338 ;
               RECT 17.684 88.902 17.736 88.938 ;
               RECT 17.684 89.502 17.736 89.538 ;
               RECT 17.684 90.102 17.736 90.138 ;
               RECT 17.684 90.702 17.736 90.738 ;
               RECT 17.684 91.302 17.736 91.338 ;
               RECT 17.684 91.902 17.736 91.938 ;
               RECT 17.684 92.502 17.736 92.538 ;
               RECT 17.684 93.102 17.736 93.138 ;
               RECT 17.684 93.702 17.736 93.738 ;
               RECT 17.684 94.302 17.736 94.338 ;
               RECT 17.684 94.902 17.736 94.938 ;
               RECT 17.684 95.502 17.736 95.538 ;
               RECT 17.684 96.102 17.736 96.138 ;
               RECT 17.684 96.702 17.736 96.738 ;
               RECT 17.684 97.302 17.736 97.338 ;
               RECT 17.684 97.902 17.736 97.938 ;
               RECT 17.684 98.502 17.736 98.538 ;
               RECT 17.684 99.102 17.736 99.138 ;
               RECT 17.684 99.702 17.736 99.738 ;
               RECT 17.684 100.302 17.736 100.338 ;
               RECT 17.684 100.902 17.736 100.938 ;
               RECT 17.684 101.502 17.736 101.538 ;
               RECT 17.684 102.102 17.736 102.138 ;
               RECT 17.684 102.702 17.736 102.738 ;
               RECT 17.684 103.302 17.736 103.338 ;
               RECT 17.684 103.902 17.736 103.938 ;
               RECT 17.684 104.502 17.736 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.216 48.62 18.256 56.5 ;
               LAYER v4 ;
               RECT 18.216 48.942 18.256 48.978 ;
               RECT 18.216 49.422 18.256 49.458 ;
               RECT 18.216 49.902 18.256 49.938 ;
               RECT 18.216 50.382 18.256 50.418 ;
               RECT 18.216 50.862 18.256 50.898 ;
               RECT 18.216 51.342 18.256 51.378 ;
               RECT 18.216 51.822 18.256 51.858 ;
               RECT 18.216 52.302 18.256 52.338 ;
               RECT 18.216 52.662 18.256 52.698 ;
               RECT 18.216 52.782 18.256 52.818 ;
               RECT 18.216 53.262 18.256 53.298 ;
               RECT 18.216 54.222 18.256 54.258 ;
               RECT 18.216 54.702 18.256 54.738 ;
               RECT 18.216 55.182 18.256 55.218 ;
               RECT 18.216 55.662 18.256 55.698 ;
               RECT 18.216 56.1475 18.256 56.1725 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.564 0.5695 18.636 104.5505 ;
               LAYER v4 ;
               RECT 18.564 0.5875 18.636 0.6125 ;
               RECT 18.564 1.1875 18.636 1.2125 ;
               RECT 18.564 1.7875 18.636 1.8125 ;
               RECT 18.564 2.3875 18.636 2.4125 ;
               RECT 18.564 2.9875 18.636 3.0125 ;
               RECT 18.564 3.5875 18.636 3.6125 ;
               RECT 18.564 4.1875 18.636 4.2125 ;
               RECT 18.564 4.7875 18.636 4.8125 ;
               RECT 18.564 5.3875 18.636 5.4125 ;
               RECT 18.564 5.9875 18.636 6.0125 ;
               RECT 18.564 6.5875 18.636 6.6125 ;
               RECT 18.564 7.1875 18.636 7.2125 ;
               RECT 18.564 7.7875 18.636 7.8125 ;
               RECT 18.564 8.3875 18.636 8.4125 ;
               RECT 18.564 8.9875 18.636 9.0125 ;
               RECT 18.564 9.5875 18.636 9.6125 ;
               RECT 18.564 10.1875 18.636 10.2125 ;
               RECT 18.564 10.7875 18.636 10.8125 ;
               RECT 18.564 11.3875 18.636 11.4125 ;
               RECT 18.564 11.9875 18.636 12.0125 ;
               RECT 18.564 12.5875 18.636 12.6125 ;
               RECT 18.564 13.1875 18.636 13.2125 ;
               RECT 18.564 13.7875 18.636 13.8125 ;
               RECT 18.564 14.3875 18.636 14.4125 ;
               RECT 18.564 14.9875 18.636 15.0125 ;
               RECT 18.564 15.5875 18.636 15.6125 ;
               RECT 18.564 16.1875 18.636 16.2125 ;
               RECT 18.564 16.7875 18.636 16.8125 ;
               RECT 18.564 17.3875 18.636 17.4125 ;
               RECT 18.564 17.9875 18.636 18.0125 ;
               RECT 18.564 18.5875 18.636 18.6125 ;
               RECT 18.564 19.1875 18.636 19.2125 ;
               RECT 18.564 19.7875 18.636 19.8125 ;
               RECT 18.564 20.3875 18.636 20.4125 ;
               RECT 18.564 20.9875 18.636 21.0125 ;
               RECT 18.564 21.5875 18.636 21.6125 ;
               RECT 18.564 22.1875 18.636 22.2125 ;
               RECT 18.564 22.7875 18.636 22.8125 ;
               RECT 18.564 23.3875 18.636 23.4125 ;
               RECT 18.564 23.9875 18.636 24.0125 ;
               RECT 18.564 24.5875 18.636 24.6125 ;
               RECT 18.564 25.1875 18.636 25.2125 ;
               RECT 18.564 25.7875 18.636 25.8125 ;
               RECT 18.564 26.3875 18.636 26.4125 ;
               RECT 18.564 26.9875 18.636 27.0125 ;
               RECT 18.564 27.5875 18.636 27.6125 ;
               RECT 18.564 28.1875 18.636 28.2125 ;
               RECT 18.564 28.7875 18.636 28.8125 ;
               RECT 18.564 29.3875 18.636 29.4125 ;
               RECT 18.564 29.9875 18.636 30.0125 ;
               RECT 18.564 30.5875 18.636 30.6125 ;
               RECT 18.564 31.1875 18.636 31.2125 ;
               RECT 18.564 31.7875 18.636 31.8125 ;
               RECT 18.564 32.3875 18.636 32.4125 ;
               RECT 18.564 32.9875 18.636 33.0125 ;
               RECT 18.564 33.5875 18.636 33.6125 ;
               RECT 18.564 34.1875 18.636 34.2125 ;
               RECT 18.564 34.7875 18.636 34.8125 ;
               RECT 18.564 35.3875 18.636 35.4125 ;
               RECT 18.564 35.9875 18.636 36.0125 ;
               RECT 18.564 36.5875 18.636 36.6125 ;
               RECT 18.564 37.1875 18.636 37.2125 ;
               RECT 18.564 37.7875 18.636 37.8125 ;
               RECT 18.564 38.3875 18.636 38.4125 ;
               RECT 18.564 38.9875 18.636 39.0125 ;
               RECT 18.564 39.5875 18.636 39.6125 ;
               RECT 18.564 40.1875 18.636 40.2125 ;
               RECT 18.564 40.7875 18.636 40.8125 ;
               RECT 18.564 41.3875 18.636 41.4125 ;
               RECT 18.564 41.9875 18.636 42.0125 ;
               RECT 18.564 42.5875 18.636 42.6125 ;
               RECT 18.564 43.1875 18.636 43.2125 ;
               RECT 18.564 43.7875 18.636 43.8125 ;
               RECT 18.564 44.3875 18.636 44.4125 ;
               RECT 18.564 44.9875 18.636 45.0125 ;
               RECT 18.564 45.5875 18.636 45.6125 ;
               RECT 18.564 46.1875 18.636 46.2125 ;
               RECT 18.564 46.7875 18.636 46.8125 ;
               RECT 18.564 47.3875 18.636 47.4125 ;
               RECT 18.564 47.9875 18.636 48.0125 ;
               RECT 18.564 48.5875 18.636 48.6125 ;
               RECT 18.564 48.9475 18.636 48.9725 ;
               RECT 18.564 49.4275 18.636 49.4525 ;
               RECT 18.564 50.3875 18.636 50.4125 ;
               RECT 18.564 50.8675 18.636 50.8925 ;
               RECT 18.564 51.3475 18.636 51.3725 ;
               RECT 18.564 51.8275 18.636 51.8525 ;
               RECT 18.564 52.3075 18.636 52.3325 ;
               RECT 18.564 52.6675 18.636 52.6925 ;
               RECT 18.564 52.7875 18.636 52.8125 ;
               RECT 18.564 53.2675 18.636 53.2925 ;
               RECT 18.564 53.7475 18.636 53.7725 ;
               RECT 18.564 54.2275 18.636 54.2525 ;
               RECT 18.564 54.7075 18.636 54.7325 ;
               RECT 18.564 55.1875 18.636 55.2125 ;
               RECT 18.564 55.6675 18.636 55.6925 ;
               RECT 18.564 56.1475 18.636 56.1725 ;
               RECT 18.564 56.5075 18.636 56.5325 ;
               RECT 18.564 57.1075 18.636 57.1325 ;
               RECT 18.564 57.7075 18.636 57.7325 ;
               RECT 18.564 58.3075 18.636 58.3325 ;
               RECT 18.564 58.9075 18.636 58.9325 ;
               RECT 18.564 59.5075 18.636 59.5325 ;
               RECT 18.564 60.1075 18.636 60.1325 ;
               RECT 18.564 60.7075 18.636 60.7325 ;
               RECT 18.564 61.3075 18.636 61.3325 ;
               RECT 18.564 61.9075 18.636 61.9325 ;
               RECT 18.564 62.5075 18.636 62.5325 ;
               RECT 18.564 63.1075 18.636 63.1325 ;
               RECT 18.564 63.7075 18.636 63.7325 ;
               RECT 18.564 64.3075 18.636 64.3325 ;
               RECT 18.564 64.9075 18.636 64.9325 ;
               RECT 18.564 65.5075 18.636 65.5325 ;
               RECT 18.564 66.1075 18.636 66.1325 ;
               RECT 18.564 66.7075 18.636 66.7325 ;
               RECT 18.564 67.3075 18.636 67.3325 ;
               RECT 18.564 67.9075 18.636 67.9325 ;
               RECT 18.564 68.5075 18.636 68.5325 ;
               RECT 18.564 69.1075 18.636 69.1325 ;
               RECT 18.564 69.7075 18.636 69.7325 ;
               RECT 18.564 70.3075 18.636 70.3325 ;
               RECT 18.564 70.9075 18.636 70.9325 ;
               RECT 18.564 71.5075 18.636 71.5325 ;
               RECT 18.564 72.1075 18.636 72.1325 ;
               RECT 18.564 72.7075 18.636 72.7325 ;
               RECT 18.564 73.3075 18.636 73.3325 ;
               RECT 18.564 73.9075 18.636 73.9325 ;
               RECT 18.564 74.5075 18.636 74.5325 ;
               RECT 18.564 75.1075 18.636 75.1325 ;
               RECT 18.564 75.7075 18.636 75.7325 ;
               RECT 18.564 76.3075 18.636 76.3325 ;
               RECT 18.564 76.9075 18.636 76.9325 ;
               RECT 18.564 77.5075 18.636 77.5325 ;
               RECT 18.564 78.1075 18.636 78.1325 ;
               RECT 18.564 78.7075 18.636 78.7325 ;
               RECT 18.564 79.3075 18.636 79.3325 ;
               RECT 18.564 79.9075 18.636 79.9325 ;
               RECT 18.564 80.5075 18.636 80.5325 ;
               RECT 18.564 81.1075 18.636 81.1325 ;
               RECT 18.564 81.7075 18.636 81.7325 ;
               RECT 18.564 82.3075 18.636 82.3325 ;
               RECT 18.564 82.9075 18.636 82.9325 ;
               RECT 18.564 83.5075 18.636 83.5325 ;
               RECT 18.564 84.1075 18.636 84.1325 ;
               RECT 18.564 84.7075 18.636 84.7325 ;
               RECT 18.564 85.3075 18.636 85.3325 ;
               RECT 18.564 85.9075 18.636 85.9325 ;
               RECT 18.564 86.5075 18.636 86.5325 ;
               RECT 18.564 87.1075 18.636 87.1325 ;
               RECT 18.564 87.7075 18.636 87.7325 ;
               RECT 18.564 88.3075 18.636 88.3325 ;
               RECT 18.564 88.9075 18.636 88.9325 ;
               RECT 18.564 89.5075 18.636 89.5325 ;
               RECT 18.564 90.1075 18.636 90.1325 ;
               RECT 18.564 90.7075 18.636 90.7325 ;
               RECT 18.564 91.3075 18.636 91.3325 ;
               RECT 18.564 91.9075 18.636 91.9325 ;
               RECT 18.564 92.5075 18.636 92.5325 ;
               RECT 18.564 93.1075 18.636 93.1325 ;
               RECT 18.564 93.7075 18.636 93.7325 ;
               RECT 18.564 94.3075 18.636 94.3325 ;
               RECT 18.564 94.9075 18.636 94.9325 ;
               RECT 18.564 95.5075 18.636 95.5325 ;
               RECT 18.564 96.1075 18.636 96.1325 ;
               RECT 18.564 96.7075 18.636 96.7325 ;
               RECT 18.564 97.3075 18.636 97.3325 ;
               RECT 18.564 97.9075 18.636 97.9325 ;
               RECT 18.564 98.5075 18.636 98.5325 ;
               RECT 18.564 99.1075 18.636 99.1325 ;
               RECT 18.564 99.7075 18.636 99.7325 ;
               RECT 18.564 100.3075 18.636 100.3325 ;
               RECT 18.564 100.9075 18.636 100.9325 ;
               RECT 18.564 101.5075 18.636 101.5325 ;
               RECT 18.564 102.1075 18.636 102.1325 ;
               RECT 18.564 102.7075 18.636 102.7325 ;
               RECT 18.564 103.3075 18.636 103.3325 ;
               RECT 18.564 103.9075 18.636 103.9325 ;
               RECT 18.564 104.5075 18.636 104.5325 ;
          END
          PORT
               LAYER m5 ;
               RECT 18.864 0.5695 18.936 104.5505 ;
               LAYER v4 ;
               RECT 18.864 0.5875 18.936 0.6125 ;
               RECT 18.864 1.1875 18.936 1.2125 ;
               RECT 18.864 1.7875 18.936 1.8125 ;
               RECT 18.864 2.3875 18.936 2.4125 ;
               RECT 18.864 2.9875 18.936 3.0125 ;
               RECT 18.864 3.5875 18.936 3.6125 ;
               RECT 18.864 4.1875 18.936 4.2125 ;
               RECT 18.864 4.7875 18.936 4.8125 ;
               RECT 18.864 5.3875 18.936 5.4125 ;
               RECT 18.864 5.9875 18.936 6.0125 ;
               RECT 18.864 6.5875 18.936 6.6125 ;
               RECT 18.864 7.1875 18.936 7.2125 ;
               RECT 18.864 7.7875 18.936 7.8125 ;
               RECT 18.864 8.3875 18.936 8.4125 ;
               RECT 18.864 8.9875 18.936 9.0125 ;
               RECT 18.864 9.5875 18.936 9.6125 ;
               RECT 18.864 10.1875 18.936 10.2125 ;
               RECT 18.864 10.7875 18.936 10.8125 ;
               RECT 18.864 11.3875 18.936 11.4125 ;
               RECT 18.864 11.9875 18.936 12.0125 ;
               RECT 18.864 12.5875 18.936 12.6125 ;
               RECT 18.864 13.1875 18.936 13.2125 ;
               RECT 18.864 13.7875 18.936 13.8125 ;
               RECT 18.864 14.3875 18.936 14.4125 ;
               RECT 18.864 14.9875 18.936 15.0125 ;
               RECT 18.864 15.5875 18.936 15.6125 ;
               RECT 18.864 16.1875 18.936 16.2125 ;
               RECT 18.864 16.7875 18.936 16.8125 ;
               RECT 18.864 17.3875 18.936 17.4125 ;
               RECT 18.864 17.9875 18.936 18.0125 ;
               RECT 18.864 18.5875 18.936 18.6125 ;
               RECT 18.864 19.1875 18.936 19.2125 ;
               RECT 18.864 19.7875 18.936 19.8125 ;
               RECT 18.864 20.3875 18.936 20.4125 ;
               RECT 18.864 20.9875 18.936 21.0125 ;
               RECT 18.864 21.5875 18.936 21.6125 ;
               RECT 18.864 22.1875 18.936 22.2125 ;
               RECT 18.864 22.7875 18.936 22.8125 ;
               RECT 18.864 23.3875 18.936 23.4125 ;
               RECT 18.864 23.9875 18.936 24.0125 ;
               RECT 18.864 24.5875 18.936 24.6125 ;
               RECT 18.864 25.1875 18.936 25.2125 ;
               RECT 18.864 25.7875 18.936 25.8125 ;
               RECT 18.864 26.3875 18.936 26.4125 ;
               RECT 18.864 26.9875 18.936 27.0125 ;
               RECT 18.864 27.5875 18.936 27.6125 ;
               RECT 18.864 28.1875 18.936 28.2125 ;
               RECT 18.864 28.7875 18.936 28.8125 ;
               RECT 18.864 29.3875 18.936 29.4125 ;
               RECT 18.864 29.9875 18.936 30.0125 ;
               RECT 18.864 30.5875 18.936 30.6125 ;
               RECT 18.864 31.1875 18.936 31.2125 ;
               RECT 18.864 31.7875 18.936 31.8125 ;
               RECT 18.864 32.3875 18.936 32.4125 ;
               RECT 18.864 32.9875 18.936 33.0125 ;
               RECT 18.864 33.5875 18.936 33.6125 ;
               RECT 18.864 34.1875 18.936 34.2125 ;
               RECT 18.864 34.7875 18.936 34.8125 ;
               RECT 18.864 35.3875 18.936 35.4125 ;
               RECT 18.864 35.9875 18.936 36.0125 ;
               RECT 18.864 36.5875 18.936 36.6125 ;
               RECT 18.864 37.1875 18.936 37.2125 ;
               RECT 18.864 37.7875 18.936 37.8125 ;
               RECT 18.864 38.3875 18.936 38.4125 ;
               RECT 18.864 38.9875 18.936 39.0125 ;
               RECT 18.864 39.5875 18.936 39.6125 ;
               RECT 18.864 40.1875 18.936 40.2125 ;
               RECT 18.864 40.7875 18.936 40.8125 ;
               RECT 18.864 41.3875 18.936 41.4125 ;
               RECT 18.864 41.9875 18.936 42.0125 ;
               RECT 18.864 42.5875 18.936 42.6125 ;
               RECT 18.864 43.1875 18.936 43.2125 ;
               RECT 18.864 43.7875 18.936 43.8125 ;
               RECT 18.864 44.3875 18.936 44.4125 ;
               RECT 18.864 44.9875 18.936 45.0125 ;
               RECT 18.864 45.5875 18.936 45.6125 ;
               RECT 18.864 46.1875 18.936 46.2125 ;
               RECT 18.864 46.7875 18.936 46.8125 ;
               RECT 18.864 47.3875 18.936 47.4125 ;
               RECT 18.864 47.9875 18.936 48.0125 ;
               RECT 18.864 48.5875 18.936 48.6125 ;
               RECT 18.864 48.9475 18.936 48.9725 ;
               RECT 18.864 49.4275 18.936 49.4525 ;
               RECT 18.864 49.9075 18.936 49.9325 ;
               RECT 18.864 50.3875 18.936 50.4125 ;
               RECT 18.864 50.8675 18.936 50.8925 ;
               RECT 18.864 51.3475 18.936 51.3725 ;
               RECT 18.864 51.8275 18.936 51.8525 ;
               RECT 18.864 52.3075 18.936 52.3325 ;
               RECT 18.864 52.6675 18.936 52.6925 ;
               RECT 18.864 52.7875 18.936 52.8125 ;
               RECT 18.864 53.2675 18.936 53.2925 ;
               RECT 18.864 53.7475 18.936 53.7725 ;
               RECT 18.864 54.2275 18.936 54.2525 ;
               RECT 18.864 54.7075 18.936 54.7325 ;
               RECT 18.864 55.1875 18.936 55.2125 ;
               RECT 18.864 55.6675 18.936 55.6925 ;
               RECT 18.864 56.1475 18.936 56.1725 ;
               RECT 18.864 56.5075 18.936 56.5325 ;
               RECT 18.864 57.1075 18.936 57.1325 ;
               RECT 18.864 57.7075 18.936 57.7325 ;
               RECT 18.864 58.3075 18.936 58.3325 ;
               RECT 18.864 58.9075 18.936 58.9325 ;
               RECT 18.864 59.5075 18.936 59.5325 ;
               RECT 18.864 60.1075 18.936 60.1325 ;
               RECT 18.864 60.7075 18.936 60.7325 ;
               RECT 18.864 61.3075 18.936 61.3325 ;
               RECT 18.864 61.9075 18.936 61.9325 ;
               RECT 18.864 62.5075 18.936 62.5325 ;
               RECT 18.864 63.1075 18.936 63.1325 ;
               RECT 18.864 63.7075 18.936 63.7325 ;
               RECT 18.864 64.3075 18.936 64.3325 ;
               RECT 18.864 64.9075 18.936 64.9325 ;
               RECT 18.864 65.5075 18.936 65.5325 ;
               RECT 18.864 66.1075 18.936 66.1325 ;
               RECT 18.864 66.7075 18.936 66.7325 ;
               RECT 18.864 67.3075 18.936 67.3325 ;
               RECT 18.864 67.9075 18.936 67.9325 ;
               RECT 18.864 68.5075 18.936 68.5325 ;
               RECT 18.864 69.1075 18.936 69.1325 ;
               RECT 18.864 69.7075 18.936 69.7325 ;
               RECT 18.864 70.3075 18.936 70.3325 ;
               RECT 18.864 70.9075 18.936 70.9325 ;
               RECT 18.864 71.5075 18.936 71.5325 ;
               RECT 18.864 72.1075 18.936 72.1325 ;
               RECT 18.864 72.7075 18.936 72.7325 ;
               RECT 18.864 73.3075 18.936 73.3325 ;
               RECT 18.864 73.9075 18.936 73.9325 ;
               RECT 18.864 74.5075 18.936 74.5325 ;
               RECT 18.864 75.1075 18.936 75.1325 ;
               RECT 18.864 75.7075 18.936 75.7325 ;
               RECT 18.864 76.3075 18.936 76.3325 ;
               RECT 18.864 76.9075 18.936 76.9325 ;
               RECT 18.864 77.5075 18.936 77.5325 ;
               RECT 18.864 78.1075 18.936 78.1325 ;
               RECT 18.864 78.7075 18.936 78.7325 ;
               RECT 18.864 79.3075 18.936 79.3325 ;
               RECT 18.864 79.9075 18.936 79.9325 ;
               RECT 18.864 80.5075 18.936 80.5325 ;
               RECT 18.864 81.1075 18.936 81.1325 ;
               RECT 18.864 81.7075 18.936 81.7325 ;
               RECT 18.864 82.3075 18.936 82.3325 ;
               RECT 18.864 82.9075 18.936 82.9325 ;
               RECT 18.864 83.5075 18.936 83.5325 ;
               RECT 18.864 84.1075 18.936 84.1325 ;
               RECT 18.864 84.7075 18.936 84.7325 ;
               RECT 18.864 85.3075 18.936 85.3325 ;
               RECT 18.864 85.9075 18.936 85.9325 ;
               RECT 18.864 86.5075 18.936 86.5325 ;
               RECT 18.864 87.1075 18.936 87.1325 ;
               RECT 18.864 87.7075 18.936 87.7325 ;
               RECT 18.864 88.3075 18.936 88.3325 ;
               RECT 18.864 88.9075 18.936 88.9325 ;
               RECT 18.864 89.5075 18.936 89.5325 ;
               RECT 18.864 90.1075 18.936 90.1325 ;
               RECT 18.864 90.7075 18.936 90.7325 ;
               RECT 18.864 91.3075 18.936 91.3325 ;
               RECT 18.864 91.9075 18.936 91.9325 ;
               RECT 18.864 92.5075 18.936 92.5325 ;
               RECT 18.864 93.1075 18.936 93.1325 ;
               RECT 18.864 93.7075 18.936 93.7325 ;
               RECT 18.864 94.3075 18.936 94.3325 ;
               RECT 18.864 94.9075 18.936 94.9325 ;
               RECT 18.864 95.5075 18.936 95.5325 ;
               RECT 18.864 96.1075 18.936 96.1325 ;
               RECT 18.864 96.7075 18.936 96.7325 ;
               RECT 18.864 97.3075 18.936 97.3325 ;
               RECT 18.864 97.9075 18.936 97.9325 ;
               RECT 18.864 98.5075 18.936 98.5325 ;
               RECT 18.864 99.1075 18.936 99.1325 ;
               RECT 18.864 99.7075 18.936 99.7325 ;
               RECT 18.864 100.3075 18.936 100.3325 ;
               RECT 18.864 100.9075 18.936 100.9325 ;
               RECT 18.864 101.5075 18.936 101.5325 ;
               RECT 18.864 102.1075 18.936 102.1325 ;
               RECT 18.864 102.7075 18.936 102.7325 ;
               RECT 18.864 103.3075 18.936 103.3325 ;
               RECT 18.864 103.9075 18.936 103.9325 ;
               RECT 18.864 104.5075 18.936 104.5325 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.228 48.64 19.282 56.48 ;
               LAYER v4 ;
               RECT 19.228 48.942 19.282 48.978 ;
               RECT 19.228 49.422 19.282 49.458 ;
               RECT 19.228 49.902 19.282 49.938 ;
               RECT 19.228 50.382 19.282 50.418 ;
               RECT 19.228 50.862 19.282 50.898 ;
               RECT 19.228 51.342 19.282 51.378 ;
               RECT 19.228 51.822 19.282 51.858 ;
               RECT 19.228 52.302 19.282 52.338 ;
               RECT 19.228 52.662 19.282 52.698 ;
               RECT 19.228 52.782 19.282 52.818 ;
               RECT 19.228 53.262 19.282 53.298 ;
               RECT 19.228 53.742 19.282 53.778 ;
               RECT 19.228 54.222 19.282 54.258 ;
               RECT 19.228 54.702 19.282 54.738 ;
               RECT 19.228 55.182 19.282 55.218 ;
               RECT 19.228 55.662 19.282 55.698 ;
               RECT 19.228 56.142 19.282 56.178 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.45 0.5695 19.502 104.5505 ;
               LAYER v4 ;
               RECT 19.45 0.582 19.502 0.618 ;
               RECT 19.45 1.182 19.502 1.218 ;
               RECT 19.45 1.782 19.502 1.818 ;
               RECT 19.45 2.382 19.502 2.418 ;
               RECT 19.45 2.982 19.502 3.018 ;
               RECT 19.45 3.582 19.502 3.618 ;
               RECT 19.45 4.182 19.502 4.218 ;
               RECT 19.45 4.782 19.502 4.818 ;
               RECT 19.45 5.382 19.502 5.418 ;
               RECT 19.45 5.982 19.502 6.018 ;
               RECT 19.45 6.582 19.502 6.618 ;
               RECT 19.45 7.182 19.502 7.218 ;
               RECT 19.45 7.782 19.502 7.818 ;
               RECT 19.45 8.382 19.502 8.418 ;
               RECT 19.45 8.982 19.502 9.018 ;
               RECT 19.45 9.582 19.502 9.618 ;
               RECT 19.45 10.182 19.502 10.218 ;
               RECT 19.45 10.782 19.502 10.818 ;
               RECT 19.45 11.382 19.502 11.418 ;
               RECT 19.45 11.982 19.502 12.018 ;
               RECT 19.45 12.582 19.502 12.618 ;
               RECT 19.45 13.182 19.502 13.218 ;
               RECT 19.45 13.782 19.502 13.818 ;
               RECT 19.45 14.382 19.502 14.418 ;
               RECT 19.45 14.982 19.502 15.018 ;
               RECT 19.45 15.582 19.502 15.618 ;
               RECT 19.45 16.182 19.502 16.218 ;
               RECT 19.45 16.782 19.502 16.818 ;
               RECT 19.45 17.382 19.502 17.418 ;
               RECT 19.45 17.982 19.502 18.018 ;
               RECT 19.45 18.582 19.502 18.618 ;
               RECT 19.45 19.182 19.502 19.218 ;
               RECT 19.45 19.782 19.502 19.818 ;
               RECT 19.45 20.382 19.502 20.418 ;
               RECT 19.45 20.982 19.502 21.018 ;
               RECT 19.45 21.582 19.502 21.618 ;
               RECT 19.45 22.182 19.502 22.218 ;
               RECT 19.45 22.782 19.502 22.818 ;
               RECT 19.45 23.382 19.502 23.418 ;
               RECT 19.45 23.982 19.502 24.018 ;
               RECT 19.45 24.582 19.502 24.618 ;
               RECT 19.45 25.182 19.502 25.218 ;
               RECT 19.45 25.782 19.502 25.818 ;
               RECT 19.45 26.382 19.502 26.418 ;
               RECT 19.45 26.982 19.502 27.018 ;
               RECT 19.45 27.582 19.502 27.618 ;
               RECT 19.45 28.182 19.502 28.218 ;
               RECT 19.45 28.782 19.502 28.818 ;
               RECT 19.45 29.382 19.502 29.418 ;
               RECT 19.45 29.982 19.502 30.018 ;
               RECT 19.45 30.582 19.502 30.618 ;
               RECT 19.45 31.182 19.502 31.218 ;
               RECT 19.45 31.782 19.502 31.818 ;
               RECT 19.45 32.382 19.502 32.418 ;
               RECT 19.45 32.982 19.502 33.018 ;
               RECT 19.45 33.582 19.502 33.618 ;
               RECT 19.45 34.182 19.502 34.218 ;
               RECT 19.45 34.782 19.502 34.818 ;
               RECT 19.45 35.382 19.502 35.418 ;
               RECT 19.45 35.982 19.502 36.018 ;
               RECT 19.45 36.582 19.502 36.618 ;
               RECT 19.45 37.182 19.502 37.218 ;
               RECT 19.45 37.782 19.502 37.818 ;
               RECT 19.45 38.382 19.502 38.418 ;
               RECT 19.45 38.982 19.502 39.018 ;
               RECT 19.45 39.582 19.502 39.618 ;
               RECT 19.45 40.182 19.502 40.218 ;
               RECT 19.45 40.782 19.502 40.818 ;
               RECT 19.45 41.382 19.502 41.418 ;
               RECT 19.45 41.982 19.502 42.018 ;
               RECT 19.45 42.582 19.502 42.618 ;
               RECT 19.45 43.182 19.502 43.218 ;
               RECT 19.45 43.782 19.502 43.818 ;
               RECT 19.45 44.382 19.502 44.418 ;
               RECT 19.45 44.982 19.502 45.018 ;
               RECT 19.45 45.582 19.502 45.618 ;
               RECT 19.45 46.182 19.502 46.218 ;
               RECT 19.45 46.782 19.502 46.818 ;
               RECT 19.45 47.382 19.502 47.418 ;
               RECT 19.45 47.982 19.502 48.018 ;
               RECT 19.45 48.582 19.502 48.618 ;
               RECT 19.45 48.942 19.502 48.978 ;
               RECT 19.45 49.422 19.502 49.458 ;
               RECT 19.45 49.7205 19.502 49.7565 ;
               RECT 19.45 49.902 19.502 49.938 ;
               RECT 19.45 50.382 19.502 50.418 ;
               RECT 19.45 50.862 19.502 50.898 ;
               RECT 19.45 51.342 19.502 51.378 ;
               RECT 19.45 51.822 19.502 51.858 ;
               RECT 19.45 52.302 19.502 52.338 ;
               RECT 19.45 52.662 19.502 52.698 ;
               RECT 19.45 52.782 19.502 52.818 ;
               RECT 19.45 53.262 19.502 53.298 ;
               RECT 19.45 53.742 19.502 53.778 ;
               RECT 19.45 54.222 19.502 54.258 ;
               RECT 19.45 54.702 19.502 54.738 ;
               RECT 19.45 55.182 19.502 55.218 ;
               RECT 19.45 55.662 19.502 55.698 ;
               RECT 19.45 56.142 19.502 56.178 ;
               RECT 19.45 56.502 19.502 56.538 ;
               RECT 19.45 57.102 19.502 57.138 ;
               RECT 19.45 57.702 19.502 57.738 ;
               RECT 19.45 58.302 19.502 58.338 ;
               RECT 19.45 58.902 19.502 58.938 ;
               RECT 19.45 59.502 19.502 59.538 ;
               RECT 19.45 60.102 19.502 60.138 ;
               RECT 19.45 60.702 19.502 60.738 ;
               RECT 19.45 61.302 19.502 61.338 ;
               RECT 19.45 61.902 19.502 61.938 ;
               RECT 19.45 62.502 19.502 62.538 ;
               RECT 19.45 63.102 19.502 63.138 ;
               RECT 19.45 63.702 19.502 63.738 ;
               RECT 19.45 64.302 19.502 64.338 ;
               RECT 19.45 64.902 19.502 64.938 ;
               RECT 19.45 65.502 19.502 65.538 ;
               RECT 19.45 66.102 19.502 66.138 ;
               RECT 19.45 66.702 19.502 66.738 ;
               RECT 19.45 67.302 19.502 67.338 ;
               RECT 19.45 67.902 19.502 67.938 ;
               RECT 19.45 68.502 19.502 68.538 ;
               RECT 19.45 69.102 19.502 69.138 ;
               RECT 19.45 69.702 19.502 69.738 ;
               RECT 19.45 70.302 19.502 70.338 ;
               RECT 19.45 70.902 19.502 70.938 ;
               RECT 19.45 71.502 19.502 71.538 ;
               RECT 19.45 72.102 19.502 72.138 ;
               RECT 19.45 72.702 19.502 72.738 ;
               RECT 19.45 73.302 19.502 73.338 ;
               RECT 19.45 73.902 19.502 73.938 ;
               RECT 19.45 74.502 19.502 74.538 ;
               RECT 19.45 75.102 19.502 75.138 ;
               RECT 19.45 75.702 19.502 75.738 ;
               RECT 19.45 76.302 19.502 76.338 ;
               RECT 19.45 76.902 19.502 76.938 ;
               RECT 19.45 77.502 19.502 77.538 ;
               RECT 19.45 78.102 19.502 78.138 ;
               RECT 19.45 78.702 19.502 78.738 ;
               RECT 19.45 79.302 19.502 79.338 ;
               RECT 19.45 79.902 19.502 79.938 ;
               RECT 19.45 80.502 19.502 80.538 ;
               RECT 19.45 81.102 19.502 81.138 ;
               RECT 19.45 81.702 19.502 81.738 ;
               RECT 19.45 82.302 19.502 82.338 ;
               RECT 19.45 82.902 19.502 82.938 ;
               RECT 19.45 83.502 19.502 83.538 ;
               RECT 19.45 84.102 19.502 84.138 ;
               RECT 19.45 84.702 19.502 84.738 ;
               RECT 19.45 85.302 19.502 85.338 ;
               RECT 19.45 85.902 19.502 85.938 ;
               RECT 19.45 86.502 19.502 86.538 ;
               RECT 19.45 87.102 19.502 87.138 ;
               RECT 19.45 87.702 19.502 87.738 ;
               RECT 19.45 88.302 19.502 88.338 ;
               RECT 19.45 88.902 19.502 88.938 ;
               RECT 19.45 89.502 19.502 89.538 ;
               RECT 19.45 90.102 19.502 90.138 ;
               RECT 19.45 90.702 19.502 90.738 ;
               RECT 19.45 91.302 19.502 91.338 ;
               RECT 19.45 91.902 19.502 91.938 ;
               RECT 19.45 92.502 19.502 92.538 ;
               RECT 19.45 93.102 19.502 93.138 ;
               RECT 19.45 93.702 19.502 93.738 ;
               RECT 19.45 94.302 19.502 94.338 ;
               RECT 19.45 94.902 19.502 94.938 ;
               RECT 19.45 95.502 19.502 95.538 ;
               RECT 19.45 96.102 19.502 96.138 ;
               RECT 19.45 96.702 19.502 96.738 ;
               RECT 19.45 97.302 19.502 97.338 ;
               RECT 19.45 97.902 19.502 97.938 ;
               RECT 19.45 98.502 19.502 98.538 ;
               RECT 19.45 99.102 19.502 99.138 ;
               RECT 19.45 99.702 19.502 99.738 ;
               RECT 19.45 100.302 19.502 100.338 ;
               RECT 19.45 100.902 19.502 100.938 ;
               RECT 19.45 101.502 19.502 101.538 ;
               RECT 19.45 102.102 19.502 102.138 ;
               RECT 19.45 102.702 19.502 102.738 ;
               RECT 19.45 103.302 19.502 103.338 ;
               RECT 19.45 103.902 19.502 103.938 ;
               RECT 19.45 104.502 19.502 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.682 0.5695 19.734 104.5505 ;
               LAYER v4 ;
               RECT 19.682 0.582 19.734 0.618 ;
               RECT 19.682 1.182 19.734 1.218 ;
               RECT 19.682 1.782 19.734 1.818 ;
               RECT 19.682 2.382 19.734 2.418 ;
               RECT 19.682 2.982 19.734 3.018 ;
               RECT 19.682 3.582 19.734 3.618 ;
               RECT 19.682 4.182 19.734 4.218 ;
               RECT 19.682 4.782 19.734 4.818 ;
               RECT 19.682 5.382 19.734 5.418 ;
               RECT 19.682 5.982 19.734 6.018 ;
               RECT 19.682 6.582 19.734 6.618 ;
               RECT 19.682 7.182 19.734 7.218 ;
               RECT 19.682 7.782 19.734 7.818 ;
               RECT 19.682 8.382 19.734 8.418 ;
               RECT 19.682 8.982 19.734 9.018 ;
               RECT 19.682 9.582 19.734 9.618 ;
               RECT 19.682 10.182 19.734 10.218 ;
               RECT 19.682 10.782 19.734 10.818 ;
               RECT 19.682 11.382 19.734 11.418 ;
               RECT 19.682 11.982 19.734 12.018 ;
               RECT 19.682 12.582 19.734 12.618 ;
               RECT 19.682 13.182 19.734 13.218 ;
               RECT 19.682 13.782 19.734 13.818 ;
               RECT 19.682 14.382 19.734 14.418 ;
               RECT 19.682 14.982 19.734 15.018 ;
               RECT 19.682 15.582 19.734 15.618 ;
               RECT 19.682 16.182 19.734 16.218 ;
               RECT 19.682 16.782 19.734 16.818 ;
               RECT 19.682 17.382 19.734 17.418 ;
               RECT 19.682 17.982 19.734 18.018 ;
               RECT 19.682 18.582 19.734 18.618 ;
               RECT 19.682 19.182 19.734 19.218 ;
               RECT 19.682 19.782 19.734 19.818 ;
               RECT 19.682 20.382 19.734 20.418 ;
               RECT 19.682 20.982 19.734 21.018 ;
               RECT 19.682 21.582 19.734 21.618 ;
               RECT 19.682 22.182 19.734 22.218 ;
               RECT 19.682 22.782 19.734 22.818 ;
               RECT 19.682 23.382 19.734 23.418 ;
               RECT 19.682 23.982 19.734 24.018 ;
               RECT 19.682 24.582 19.734 24.618 ;
               RECT 19.682 25.182 19.734 25.218 ;
               RECT 19.682 25.782 19.734 25.818 ;
               RECT 19.682 26.382 19.734 26.418 ;
               RECT 19.682 26.982 19.734 27.018 ;
               RECT 19.682 27.582 19.734 27.618 ;
               RECT 19.682 28.182 19.734 28.218 ;
               RECT 19.682 28.782 19.734 28.818 ;
               RECT 19.682 29.382 19.734 29.418 ;
               RECT 19.682 29.982 19.734 30.018 ;
               RECT 19.682 30.582 19.734 30.618 ;
               RECT 19.682 31.182 19.734 31.218 ;
               RECT 19.682 31.782 19.734 31.818 ;
               RECT 19.682 32.382 19.734 32.418 ;
               RECT 19.682 32.982 19.734 33.018 ;
               RECT 19.682 33.582 19.734 33.618 ;
               RECT 19.682 34.182 19.734 34.218 ;
               RECT 19.682 34.782 19.734 34.818 ;
               RECT 19.682 35.382 19.734 35.418 ;
               RECT 19.682 35.982 19.734 36.018 ;
               RECT 19.682 36.582 19.734 36.618 ;
               RECT 19.682 37.182 19.734 37.218 ;
               RECT 19.682 37.782 19.734 37.818 ;
               RECT 19.682 38.382 19.734 38.418 ;
               RECT 19.682 38.982 19.734 39.018 ;
               RECT 19.682 39.582 19.734 39.618 ;
               RECT 19.682 40.182 19.734 40.218 ;
               RECT 19.682 40.782 19.734 40.818 ;
               RECT 19.682 41.382 19.734 41.418 ;
               RECT 19.682 41.982 19.734 42.018 ;
               RECT 19.682 42.582 19.734 42.618 ;
               RECT 19.682 43.182 19.734 43.218 ;
               RECT 19.682 43.782 19.734 43.818 ;
               RECT 19.682 44.382 19.734 44.418 ;
               RECT 19.682 44.982 19.734 45.018 ;
               RECT 19.682 45.582 19.734 45.618 ;
               RECT 19.682 46.182 19.734 46.218 ;
               RECT 19.682 46.782 19.734 46.818 ;
               RECT 19.682 47.382 19.734 47.418 ;
               RECT 19.682 47.982 19.734 48.018 ;
               RECT 19.682 48.582 19.734 48.618 ;
               RECT 19.682 48.942 19.734 48.978 ;
               RECT 19.682 49.422 19.734 49.458 ;
               RECT 19.682 49.7205 19.734 49.7565 ;
               RECT 19.682 49.902 19.734 49.938 ;
               RECT 19.682 50.382 19.734 50.418 ;
               RECT 19.682 50.862 19.734 50.898 ;
               RECT 19.682 51.342 19.734 51.378 ;
               RECT 19.682 51.822 19.734 51.858 ;
               RECT 19.682 52.302 19.734 52.338 ;
               RECT 19.682 52.782 19.734 52.818 ;
               RECT 19.682 53.262 19.734 53.298 ;
               RECT 19.682 53.742 19.734 53.778 ;
               RECT 19.682 54.222 19.734 54.258 ;
               RECT 19.682 54.702 19.734 54.738 ;
               RECT 19.682 55.662 19.734 55.698 ;
               RECT 19.682 56.502 19.734 56.538 ;
               RECT 19.682 57.102 19.734 57.138 ;
               RECT 19.682 57.702 19.734 57.738 ;
               RECT 19.682 58.302 19.734 58.338 ;
               RECT 19.682 58.902 19.734 58.938 ;
               RECT 19.682 59.502 19.734 59.538 ;
               RECT 19.682 60.102 19.734 60.138 ;
               RECT 19.682 60.702 19.734 60.738 ;
               RECT 19.682 61.302 19.734 61.338 ;
               RECT 19.682 61.902 19.734 61.938 ;
               RECT 19.682 62.502 19.734 62.538 ;
               RECT 19.682 63.102 19.734 63.138 ;
               RECT 19.682 63.702 19.734 63.738 ;
               RECT 19.682 64.302 19.734 64.338 ;
               RECT 19.682 64.902 19.734 64.938 ;
               RECT 19.682 65.502 19.734 65.538 ;
               RECT 19.682 66.102 19.734 66.138 ;
               RECT 19.682 66.702 19.734 66.738 ;
               RECT 19.682 67.302 19.734 67.338 ;
               RECT 19.682 67.902 19.734 67.938 ;
               RECT 19.682 68.502 19.734 68.538 ;
               RECT 19.682 69.102 19.734 69.138 ;
               RECT 19.682 69.702 19.734 69.738 ;
               RECT 19.682 70.302 19.734 70.338 ;
               RECT 19.682 70.902 19.734 70.938 ;
               RECT 19.682 71.502 19.734 71.538 ;
               RECT 19.682 72.102 19.734 72.138 ;
               RECT 19.682 72.702 19.734 72.738 ;
               RECT 19.682 73.302 19.734 73.338 ;
               RECT 19.682 73.902 19.734 73.938 ;
               RECT 19.682 74.502 19.734 74.538 ;
               RECT 19.682 75.102 19.734 75.138 ;
               RECT 19.682 75.702 19.734 75.738 ;
               RECT 19.682 76.302 19.734 76.338 ;
               RECT 19.682 76.902 19.734 76.938 ;
               RECT 19.682 77.502 19.734 77.538 ;
               RECT 19.682 78.102 19.734 78.138 ;
               RECT 19.682 78.702 19.734 78.738 ;
               RECT 19.682 79.302 19.734 79.338 ;
               RECT 19.682 79.902 19.734 79.938 ;
               RECT 19.682 80.502 19.734 80.538 ;
               RECT 19.682 81.102 19.734 81.138 ;
               RECT 19.682 81.702 19.734 81.738 ;
               RECT 19.682 82.302 19.734 82.338 ;
               RECT 19.682 82.902 19.734 82.938 ;
               RECT 19.682 83.502 19.734 83.538 ;
               RECT 19.682 84.102 19.734 84.138 ;
               RECT 19.682 84.702 19.734 84.738 ;
               RECT 19.682 85.302 19.734 85.338 ;
               RECT 19.682 85.902 19.734 85.938 ;
               RECT 19.682 86.502 19.734 86.538 ;
               RECT 19.682 87.102 19.734 87.138 ;
               RECT 19.682 87.702 19.734 87.738 ;
               RECT 19.682 88.302 19.734 88.338 ;
               RECT 19.682 88.902 19.734 88.938 ;
               RECT 19.682 89.502 19.734 89.538 ;
               RECT 19.682 90.102 19.734 90.138 ;
               RECT 19.682 90.702 19.734 90.738 ;
               RECT 19.682 91.302 19.734 91.338 ;
               RECT 19.682 91.902 19.734 91.938 ;
               RECT 19.682 92.502 19.734 92.538 ;
               RECT 19.682 93.102 19.734 93.138 ;
               RECT 19.682 93.702 19.734 93.738 ;
               RECT 19.682 94.302 19.734 94.338 ;
               RECT 19.682 94.902 19.734 94.938 ;
               RECT 19.682 95.502 19.734 95.538 ;
               RECT 19.682 96.102 19.734 96.138 ;
               RECT 19.682 96.702 19.734 96.738 ;
               RECT 19.682 97.302 19.734 97.338 ;
               RECT 19.682 97.902 19.734 97.938 ;
               RECT 19.682 98.502 19.734 98.538 ;
               RECT 19.682 99.102 19.734 99.138 ;
               RECT 19.682 99.702 19.734 99.738 ;
               RECT 19.682 100.302 19.734 100.338 ;
               RECT 19.682 100.902 19.734 100.938 ;
               RECT 19.682 101.502 19.734 101.538 ;
               RECT 19.682 102.102 19.734 102.138 ;
               RECT 19.682 102.702 19.734 102.738 ;
               RECT 19.682 103.302 19.734 103.338 ;
               RECT 19.682 103.902 19.734 103.938 ;
               RECT 19.682 104.502 19.734 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 19.994 0.5695 20.046 104.5505 ;
               LAYER v4 ;
               RECT 19.994 0.582 20.046 0.618 ;
               RECT 19.994 1.182 20.046 1.218 ;
               RECT 19.994 1.782 20.046 1.818 ;
               RECT 19.994 2.382 20.046 2.418 ;
               RECT 19.994 2.982 20.046 3.018 ;
               RECT 19.994 3.582 20.046 3.618 ;
               RECT 19.994 4.182 20.046 4.218 ;
               RECT 19.994 4.782 20.046 4.818 ;
               RECT 19.994 5.382 20.046 5.418 ;
               RECT 19.994 5.982 20.046 6.018 ;
               RECT 19.994 6.582 20.046 6.618 ;
               RECT 19.994 7.182 20.046 7.218 ;
               RECT 19.994 7.782 20.046 7.818 ;
               RECT 19.994 8.382 20.046 8.418 ;
               RECT 19.994 8.982 20.046 9.018 ;
               RECT 19.994 9.582 20.046 9.618 ;
               RECT 19.994 10.182 20.046 10.218 ;
               RECT 19.994 10.782 20.046 10.818 ;
               RECT 19.994 11.382 20.046 11.418 ;
               RECT 19.994 11.982 20.046 12.018 ;
               RECT 19.994 12.582 20.046 12.618 ;
               RECT 19.994 13.182 20.046 13.218 ;
               RECT 19.994 13.782 20.046 13.818 ;
               RECT 19.994 14.382 20.046 14.418 ;
               RECT 19.994 14.982 20.046 15.018 ;
               RECT 19.994 15.582 20.046 15.618 ;
               RECT 19.994 16.182 20.046 16.218 ;
               RECT 19.994 16.782 20.046 16.818 ;
               RECT 19.994 17.382 20.046 17.418 ;
               RECT 19.994 17.982 20.046 18.018 ;
               RECT 19.994 18.582 20.046 18.618 ;
               RECT 19.994 19.182 20.046 19.218 ;
               RECT 19.994 19.782 20.046 19.818 ;
               RECT 19.994 20.382 20.046 20.418 ;
               RECT 19.994 20.982 20.046 21.018 ;
               RECT 19.994 21.582 20.046 21.618 ;
               RECT 19.994 22.182 20.046 22.218 ;
               RECT 19.994 22.782 20.046 22.818 ;
               RECT 19.994 23.382 20.046 23.418 ;
               RECT 19.994 23.982 20.046 24.018 ;
               RECT 19.994 24.582 20.046 24.618 ;
               RECT 19.994 25.182 20.046 25.218 ;
               RECT 19.994 25.782 20.046 25.818 ;
               RECT 19.994 26.382 20.046 26.418 ;
               RECT 19.994 26.982 20.046 27.018 ;
               RECT 19.994 27.582 20.046 27.618 ;
               RECT 19.994 28.182 20.046 28.218 ;
               RECT 19.994 28.782 20.046 28.818 ;
               RECT 19.994 29.382 20.046 29.418 ;
               RECT 19.994 29.982 20.046 30.018 ;
               RECT 19.994 30.582 20.046 30.618 ;
               RECT 19.994 31.182 20.046 31.218 ;
               RECT 19.994 31.782 20.046 31.818 ;
               RECT 19.994 32.382 20.046 32.418 ;
               RECT 19.994 32.982 20.046 33.018 ;
               RECT 19.994 33.582 20.046 33.618 ;
               RECT 19.994 34.182 20.046 34.218 ;
               RECT 19.994 34.782 20.046 34.818 ;
               RECT 19.994 35.382 20.046 35.418 ;
               RECT 19.994 35.982 20.046 36.018 ;
               RECT 19.994 36.582 20.046 36.618 ;
               RECT 19.994 37.182 20.046 37.218 ;
               RECT 19.994 37.782 20.046 37.818 ;
               RECT 19.994 38.382 20.046 38.418 ;
               RECT 19.994 38.982 20.046 39.018 ;
               RECT 19.994 39.582 20.046 39.618 ;
               RECT 19.994 40.182 20.046 40.218 ;
               RECT 19.994 40.782 20.046 40.818 ;
               RECT 19.994 41.382 20.046 41.418 ;
               RECT 19.994 41.982 20.046 42.018 ;
               RECT 19.994 42.582 20.046 42.618 ;
               RECT 19.994 43.182 20.046 43.218 ;
               RECT 19.994 43.782 20.046 43.818 ;
               RECT 19.994 44.382 20.046 44.418 ;
               RECT 19.994 44.982 20.046 45.018 ;
               RECT 19.994 45.582 20.046 45.618 ;
               RECT 19.994 46.182 20.046 46.218 ;
               RECT 19.994 46.782 20.046 46.818 ;
               RECT 19.994 47.382 20.046 47.418 ;
               RECT 19.994 47.982 20.046 48.018 ;
               RECT 19.994 48.582 20.046 48.618 ;
               RECT 19.994 48.942 20.046 48.978 ;
               RECT 19.994 49.422 20.046 49.458 ;
               RECT 19.994 49.902 20.046 49.938 ;
               RECT 19.994 50.382 20.046 50.418 ;
               RECT 19.994 50.862 20.046 50.898 ;
               RECT 19.994 51.342 20.046 51.378 ;
               RECT 19.994 51.822 20.046 51.858 ;
               RECT 19.994 52.302 20.046 52.338 ;
               RECT 19.994 52.662 20.046 52.698 ;
               RECT 19.994 52.782 20.046 52.818 ;
               RECT 19.994 53.2675 20.046 53.2925 ;
               RECT 19.994 53.742 20.046 53.778 ;
               RECT 19.994 54.222 20.046 54.258 ;
               RECT 19.994 54.702 20.046 54.738 ;
               RECT 19.994 55.182 20.046 55.218 ;
               RECT 19.994 55.662 20.046 55.698 ;
               RECT 19.994 56.142 20.046 56.178 ;
               RECT 19.994 56.502 20.046 56.538 ;
               RECT 19.994 57.102 20.046 57.138 ;
               RECT 19.994 57.702 20.046 57.738 ;
               RECT 19.994 58.302 20.046 58.338 ;
               RECT 19.994 58.902 20.046 58.938 ;
               RECT 19.994 59.502 20.046 59.538 ;
               RECT 19.994 60.102 20.046 60.138 ;
               RECT 19.994 60.702 20.046 60.738 ;
               RECT 19.994 61.302 20.046 61.338 ;
               RECT 19.994 61.902 20.046 61.938 ;
               RECT 19.994 62.502 20.046 62.538 ;
               RECT 19.994 63.102 20.046 63.138 ;
               RECT 19.994 63.702 20.046 63.738 ;
               RECT 19.994 64.302 20.046 64.338 ;
               RECT 19.994 64.902 20.046 64.938 ;
               RECT 19.994 65.502 20.046 65.538 ;
               RECT 19.994 66.102 20.046 66.138 ;
               RECT 19.994 66.702 20.046 66.738 ;
               RECT 19.994 67.302 20.046 67.338 ;
               RECT 19.994 67.902 20.046 67.938 ;
               RECT 19.994 68.502 20.046 68.538 ;
               RECT 19.994 69.102 20.046 69.138 ;
               RECT 19.994 69.702 20.046 69.738 ;
               RECT 19.994 70.302 20.046 70.338 ;
               RECT 19.994 70.902 20.046 70.938 ;
               RECT 19.994 71.502 20.046 71.538 ;
               RECT 19.994 72.102 20.046 72.138 ;
               RECT 19.994 72.702 20.046 72.738 ;
               RECT 19.994 73.302 20.046 73.338 ;
               RECT 19.994 73.902 20.046 73.938 ;
               RECT 19.994 74.502 20.046 74.538 ;
               RECT 19.994 75.102 20.046 75.138 ;
               RECT 19.994 75.702 20.046 75.738 ;
               RECT 19.994 76.302 20.046 76.338 ;
               RECT 19.994 76.902 20.046 76.938 ;
               RECT 19.994 77.502 20.046 77.538 ;
               RECT 19.994 78.102 20.046 78.138 ;
               RECT 19.994 78.702 20.046 78.738 ;
               RECT 19.994 79.302 20.046 79.338 ;
               RECT 19.994 79.902 20.046 79.938 ;
               RECT 19.994 80.502 20.046 80.538 ;
               RECT 19.994 81.102 20.046 81.138 ;
               RECT 19.994 81.702 20.046 81.738 ;
               RECT 19.994 82.302 20.046 82.338 ;
               RECT 19.994 82.902 20.046 82.938 ;
               RECT 19.994 83.502 20.046 83.538 ;
               RECT 19.994 84.102 20.046 84.138 ;
               RECT 19.994 84.702 20.046 84.738 ;
               RECT 19.994 85.302 20.046 85.338 ;
               RECT 19.994 85.902 20.046 85.938 ;
               RECT 19.994 86.502 20.046 86.538 ;
               RECT 19.994 87.102 20.046 87.138 ;
               RECT 19.994 87.702 20.046 87.738 ;
               RECT 19.994 88.302 20.046 88.338 ;
               RECT 19.994 88.902 20.046 88.938 ;
               RECT 19.994 89.502 20.046 89.538 ;
               RECT 19.994 90.102 20.046 90.138 ;
               RECT 19.994 90.702 20.046 90.738 ;
               RECT 19.994 91.302 20.046 91.338 ;
               RECT 19.994 91.902 20.046 91.938 ;
               RECT 19.994 92.502 20.046 92.538 ;
               RECT 19.994 93.102 20.046 93.138 ;
               RECT 19.994 93.702 20.046 93.738 ;
               RECT 19.994 94.302 20.046 94.338 ;
               RECT 19.994 94.902 20.046 94.938 ;
               RECT 19.994 95.502 20.046 95.538 ;
               RECT 19.994 96.102 20.046 96.138 ;
               RECT 19.994 96.702 20.046 96.738 ;
               RECT 19.994 97.302 20.046 97.338 ;
               RECT 19.994 97.902 20.046 97.938 ;
               RECT 19.994 98.502 20.046 98.538 ;
               RECT 19.994 99.102 20.046 99.138 ;
               RECT 19.994 99.702 20.046 99.738 ;
               RECT 19.994 100.302 20.046 100.338 ;
               RECT 19.994 100.902 20.046 100.938 ;
               RECT 19.994 101.502 20.046 101.538 ;
               RECT 19.994 102.102 20.046 102.138 ;
               RECT 19.994 102.702 20.046 102.738 ;
               RECT 19.994 103.302 20.046 103.338 ;
               RECT 19.994 103.902 20.046 103.938 ;
               RECT 19.994 104.502 20.046 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 2.174 0.5695 2.226 104.5505 ;
               LAYER v4 ;
               RECT 2.174 0.582 2.226 0.618 ;
               RECT 2.174 1.182 2.226 1.218 ;
               RECT 2.174 1.782 2.226 1.818 ;
               RECT 2.174 2.382 2.226 2.418 ;
               RECT 2.174 2.982 2.226 3.018 ;
               RECT 2.174 3.582 2.226 3.618 ;
               RECT 2.174 4.182 2.226 4.218 ;
               RECT 2.174 4.782 2.226 4.818 ;
               RECT 2.174 5.382 2.226 5.418 ;
               RECT 2.174 5.982 2.226 6.018 ;
               RECT 2.174 6.582 2.226 6.618 ;
               RECT 2.174 7.182 2.226 7.218 ;
               RECT 2.174 7.782 2.226 7.818 ;
               RECT 2.174 8.382 2.226 8.418 ;
               RECT 2.174 8.982 2.226 9.018 ;
               RECT 2.174 9.582 2.226 9.618 ;
               RECT 2.174 10.182 2.226 10.218 ;
               RECT 2.174 10.782 2.226 10.818 ;
               RECT 2.174 11.382 2.226 11.418 ;
               RECT 2.174 11.982 2.226 12.018 ;
               RECT 2.174 12.582 2.226 12.618 ;
               RECT 2.174 13.182 2.226 13.218 ;
               RECT 2.174 13.782 2.226 13.818 ;
               RECT 2.174 14.382 2.226 14.418 ;
               RECT 2.174 14.982 2.226 15.018 ;
               RECT 2.174 15.582 2.226 15.618 ;
               RECT 2.174 16.182 2.226 16.218 ;
               RECT 2.174 16.782 2.226 16.818 ;
               RECT 2.174 17.382 2.226 17.418 ;
               RECT 2.174 17.982 2.226 18.018 ;
               RECT 2.174 18.582 2.226 18.618 ;
               RECT 2.174 19.182 2.226 19.218 ;
               RECT 2.174 19.782 2.226 19.818 ;
               RECT 2.174 20.382 2.226 20.418 ;
               RECT 2.174 20.982 2.226 21.018 ;
               RECT 2.174 21.582 2.226 21.618 ;
               RECT 2.174 22.182 2.226 22.218 ;
               RECT 2.174 22.782 2.226 22.818 ;
               RECT 2.174 23.382 2.226 23.418 ;
               RECT 2.174 23.982 2.226 24.018 ;
               RECT 2.174 24.582 2.226 24.618 ;
               RECT 2.174 25.182 2.226 25.218 ;
               RECT 2.174 25.782 2.226 25.818 ;
               RECT 2.174 26.382 2.226 26.418 ;
               RECT 2.174 26.982 2.226 27.018 ;
               RECT 2.174 27.582 2.226 27.618 ;
               RECT 2.174 28.182 2.226 28.218 ;
               RECT 2.174 28.782 2.226 28.818 ;
               RECT 2.174 29.382 2.226 29.418 ;
               RECT 2.174 29.982 2.226 30.018 ;
               RECT 2.174 30.582 2.226 30.618 ;
               RECT 2.174 31.182 2.226 31.218 ;
               RECT 2.174 31.782 2.226 31.818 ;
               RECT 2.174 32.382 2.226 32.418 ;
               RECT 2.174 32.982 2.226 33.018 ;
               RECT 2.174 33.582 2.226 33.618 ;
               RECT 2.174 34.182 2.226 34.218 ;
               RECT 2.174 34.782 2.226 34.818 ;
               RECT 2.174 35.382 2.226 35.418 ;
               RECT 2.174 35.982 2.226 36.018 ;
               RECT 2.174 36.582 2.226 36.618 ;
               RECT 2.174 37.182 2.226 37.218 ;
               RECT 2.174 37.782 2.226 37.818 ;
               RECT 2.174 38.382 2.226 38.418 ;
               RECT 2.174 38.982 2.226 39.018 ;
               RECT 2.174 39.582 2.226 39.618 ;
               RECT 2.174 40.182 2.226 40.218 ;
               RECT 2.174 40.782 2.226 40.818 ;
               RECT 2.174 41.382 2.226 41.418 ;
               RECT 2.174 41.982 2.226 42.018 ;
               RECT 2.174 42.582 2.226 42.618 ;
               RECT 2.174 43.182 2.226 43.218 ;
               RECT 2.174 43.782 2.226 43.818 ;
               RECT 2.174 44.382 2.226 44.418 ;
               RECT 2.174 44.982 2.226 45.018 ;
               RECT 2.174 45.582 2.226 45.618 ;
               RECT 2.174 46.182 2.226 46.218 ;
               RECT 2.174 46.782 2.226 46.818 ;
               RECT 2.174 47.382 2.226 47.418 ;
               RECT 2.174 47.982 2.226 48.018 ;
               RECT 2.174 48.582 2.226 48.618 ;
               RECT 2.174 48.942 2.226 48.978 ;
               RECT 2.174 48.9475 2.226 48.9725 ;
               RECT 2.174 49.182 2.226 49.218 ;
               RECT 2.174 49.902 2.226 49.938 ;
               RECT 2.174 50.622 2.226 50.658 ;
               RECT 2.174 50.862 2.226 50.898 ;
               RECT 2.174 51.342 2.226 51.378 ;
               RECT 2.174 51.822 2.226 51.858 ;
               RECT 2.174 52.302 2.226 52.338 ;
               RECT 2.174 52.782 2.226 52.818 ;
               RECT 2.174 53.262 2.226 53.298 ;
               RECT 2.174 53.742 2.226 53.778 ;
               RECT 2.174 54.222 2.226 54.258 ;
               RECT 2.174 54.462 2.226 54.498 ;
               RECT 2.174 55.182 2.226 55.218 ;
               RECT 2.174 55.902 2.226 55.938 ;
               RECT 2.174 56.142 2.226 56.178 ;
               RECT 2.174 56.1475 2.226 56.1725 ;
               RECT 2.174 56.502 2.226 56.538 ;
               RECT 2.174 57.102 2.226 57.138 ;
               RECT 2.174 57.702 2.226 57.738 ;
               RECT 2.174 58.302 2.226 58.338 ;
               RECT 2.174 58.902 2.226 58.938 ;
               RECT 2.174 59.502 2.226 59.538 ;
               RECT 2.174 60.102 2.226 60.138 ;
               RECT 2.174 60.702 2.226 60.738 ;
               RECT 2.174 61.302 2.226 61.338 ;
               RECT 2.174 61.902 2.226 61.938 ;
               RECT 2.174 62.502 2.226 62.538 ;
               RECT 2.174 63.102 2.226 63.138 ;
               RECT 2.174 63.702 2.226 63.738 ;
               RECT 2.174 64.302 2.226 64.338 ;
               RECT 2.174 64.902 2.226 64.938 ;
               RECT 2.174 65.502 2.226 65.538 ;
               RECT 2.174 66.102 2.226 66.138 ;
               RECT 2.174 66.702 2.226 66.738 ;
               RECT 2.174 67.302 2.226 67.338 ;
               RECT 2.174 67.902 2.226 67.938 ;
               RECT 2.174 68.502 2.226 68.538 ;
               RECT 2.174 69.102 2.226 69.138 ;
               RECT 2.174 69.702 2.226 69.738 ;
               RECT 2.174 70.302 2.226 70.338 ;
               RECT 2.174 70.902 2.226 70.938 ;
               RECT 2.174 71.502 2.226 71.538 ;
               RECT 2.174 72.102 2.226 72.138 ;
               RECT 2.174 72.702 2.226 72.738 ;
               RECT 2.174 73.302 2.226 73.338 ;
               RECT 2.174 73.902 2.226 73.938 ;
               RECT 2.174 74.502 2.226 74.538 ;
               RECT 2.174 75.102 2.226 75.138 ;
               RECT 2.174 75.702 2.226 75.738 ;
               RECT 2.174 76.302 2.226 76.338 ;
               RECT 2.174 76.902 2.226 76.938 ;
               RECT 2.174 77.502 2.226 77.538 ;
               RECT 2.174 78.102 2.226 78.138 ;
               RECT 2.174 78.702 2.226 78.738 ;
               RECT 2.174 79.302 2.226 79.338 ;
               RECT 2.174 79.902 2.226 79.938 ;
               RECT 2.174 80.502 2.226 80.538 ;
               RECT 2.174 81.102 2.226 81.138 ;
               RECT 2.174 81.702 2.226 81.738 ;
               RECT 2.174 82.302 2.226 82.338 ;
               RECT 2.174 82.902 2.226 82.938 ;
               RECT 2.174 83.502 2.226 83.538 ;
               RECT 2.174 84.102 2.226 84.138 ;
               RECT 2.174 84.702 2.226 84.738 ;
               RECT 2.174 85.302 2.226 85.338 ;
               RECT 2.174 85.902 2.226 85.938 ;
               RECT 2.174 86.502 2.226 86.538 ;
               RECT 2.174 87.102 2.226 87.138 ;
               RECT 2.174 87.702 2.226 87.738 ;
               RECT 2.174 88.302 2.226 88.338 ;
               RECT 2.174 88.902 2.226 88.938 ;
               RECT 2.174 89.502 2.226 89.538 ;
               RECT 2.174 90.102 2.226 90.138 ;
               RECT 2.174 90.702 2.226 90.738 ;
               RECT 2.174 91.302 2.226 91.338 ;
               RECT 2.174 91.902 2.226 91.938 ;
               RECT 2.174 92.502 2.226 92.538 ;
               RECT 2.174 93.102 2.226 93.138 ;
               RECT 2.174 93.702 2.226 93.738 ;
               RECT 2.174 94.302 2.226 94.338 ;
               RECT 2.174 94.902 2.226 94.938 ;
               RECT 2.174 95.502 2.226 95.538 ;
               RECT 2.174 96.102 2.226 96.138 ;
               RECT 2.174 96.702 2.226 96.738 ;
               RECT 2.174 97.302 2.226 97.338 ;
               RECT 2.174 97.902 2.226 97.938 ;
               RECT 2.174 98.502 2.226 98.538 ;
               RECT 2.174 99.102 2.226 99.138 ;
               RECT 2.174 99.702 2.226 99.738 ;
               RECT 2.174 100.302 2.226 100.338 ;
               RECT 2.174 100.902 2.226 100.938 ;
               RECT 2.174 101.502 2.226 101.538 ;
               RECT 2.174 102.102 2.226 102.138 ;
               RECT 2.174 102.702 2.226 102.738 ;
               RECT 2.174 103.302 2.226 103.338 ;
               RECT 2.174 103.902 2.226 103.938 ;
               RECT 2.174 104.502 2.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 2.974 0.5695 3.026 104.5505 ;
               LAYER v4 ;
               RECT 2.974 0.582 3.026 0.618 ;
               RECT 2.974 1.182 3.026 1.218 ;
               RECT 2.974 1.782 3.026 1.818 ;
               RECT 2.974 2.382 3.026 2.418 ;
               RECT 2.974 2.982 3.026 3.018 ;
               RECT 2.974 3.582 3.026 3.618 ;
               RECT 2.974 4.182 3.026 4.218 ;
               RECT 2.974 4.782 3.026 4.818 ;
               RECT 2.974 5.382 3.026 5.418 ;
               RECT 2.974 5.982 3.026 6.018 ;
               RECT 2.974 6.582 3.026 6.618 ;
               RECT 2.974 7.182 3.026 7.218 ;
               RECT 2.974 7.782 3.026 7.818 ;
               RECT 2.974 8.382 3.026 8.418 ;
               RECT 2.974 8.982 3.026 9.018 ;
               RECT 2.974 9.582 3.026 9.618 ;
               RECT 2.974 10.182 3.026 10.218 ;
               RECT 2.974 10.782 3.026 10.818 ;
               RECT 2.974 11.382 3.026 11.418 ;
               RECT 2.974 11.982 3.026 12.018 ;
               RECT 2.974 12.582 3.026 12.618 ;
               RECT 2.974 13.182 3.026 13.218 ;
               RECT 2.974 13.782 3.026 13.818 ;
               RECT 2.974 14.382 3.026 14.418 ;
               RECT 2.974 14.982 3.026 15.018 ;
               RECT 2.974 15.582 3.026 15.618 ;
               RECT 2.974 16.182 3.026 16.218 ;
               RECT 2.974 16.782 3.026 16.818 ;
               RECT 2.974 17.382 3.026 17.418 ;
               RECT 2.974 17.982 3.026 18.018 ;
               RECT 2.974 18.582 3.026 18.618 ;
               RECT 2.974 19.182 3.026 19.218 ;
               RECT 2.974 19.782 3.026 19.818 ;
               RECT 2.974 20.382 3.026 20.418 ;
               RECT 2.974 20.982 3.026 21.018 ;
               RECT 2.974 21.582 3.026 21.618 ;
               RECT 2.974 22.182 3.026 22.218 ;
               RECT 2.974 22.782 3.026 22.818 ;
               RECT 2.974 23.382 3.026 23.418 ;
               RECT 2.974 23.982 3.026 24.018 ;
               RECT 2.974 24.582 3.026 24.618 ;
               RECT 2.974 25.182 3.026 25.218 ;
               RECT 2.974 25.782 3.026 25.818 ;
               RECT 2.974 26.382 3.026 26.418 ;
               RECT 2.974 26.982 3.026 27.018 ;
               RECT 2.974 27.582 3.026 27.618 ;
               RECT 2.974 28.182 3.026 28.218 ;
               RECT 2.974 28.782 3.026 28.818 ;
               RECT 2.974 29.382 3.026 29.418 ;
               RECT 2.974 29.982 3.026 30.018 ;
               RECT 2.974 30.582 3.026 30.618 ;
               RECT 2.974 31.182 3.026 31.218 ;
               RECT 2.974 31.782 3.026 31.818 ;
               RECT 2.974 32.382 3.026 32.418 ;
               RECT 2.974 32.982 3.026 33.018 ;
               RECT 2.974 33.582 3.026 33.618 ;
               RECT 2.974 34.182 3.026 34.218 ;
               RECT 2.974 34.782 3.026 34.818 ;
               RECT 2.974 35.382 3.026 35.418 ;
               RECT 2.974 35.982 3.026 36.018 ;
               RECT 2.974 36.582 3.026 36.618 ;
               RECT 2.974 37.182 3.026 37.218 ;
               RECT 2.974 37.782 3.026 37.818 ;
               RECT 2.974 38.382 3.026 38.418 ;
               RECT 2.974 38.982 3.026 39.018 ;
               RECT 2.974 39.582 3.026 39.618 ;
               RECT 2.974 40.182 3.026 40.218 ;
               RECT 2.974 40.782 3.026 40.818 ;
               RECT 2.974 41.382 3.026 41.418 ;
               RECT 2.974 41.982 3.026 42.018 ;
               RECT 2.974 42.582 3.026 42.618 ;
               RECT 2.974 43.182 3.026 43.218 ;
               RECT 2.974 43.782 3.026 43.818 ;
               RECT 2.974 44.382 3.026 44.418 ;
               RECT 2.974 44.982 3.026 45.018 ;
               RECT 2.974 45.582 3.026 45.618 ;
               RECT 2.974 46.182 3.026 46.218 ;
               RECT 2.974 46.782 3.026 46.818 ;
               RECT 2.974 47.382 3.026 47.418 ;
               RECT 2.974 47.982 3.026 48.018 ;
               RECT 2.974 48.582 3.026 48.618 ;
               RECT 2.974 48.942 3.026 48.978 ;
               RECT 2.974 49.182 3.026 49.218 ;
               RECT 2.974 49.902 3.026 49.938 ;
               RECT 2.974 50.622 3.026 50.658 ;
               RECT 2.974 50.862 3.026 50.898 ;
               RECT 2.974 51.342 3.026 51.378 ;
               RECT 2.974 51.822 3.026 51.858 ;
               RECT 2.974 52.302 3.026 52.338 ;
               RECT 2.974 52.782 3.026 52.818 ;
               RECT 2.974 53.262 3.026 53.298 ;
               RECT 2.974 53.742 3.026 53.778 ;
               RECT 2.974 54.222 3.026 54.258 ;
               RECT 2.974 54.462 3.026 54.498 ;
               RECT 2.974 55.182 3.026 55.218 ;
               RECT 2.974 55.902 3.026 55.938 ;
               RECT 2.974 56.142 3.026 56.178 ;
               RECT 2.974 56.502 3.026 56.538 ;
               RECT 2.974 57.102 3.026 57.138 ;
               RECT 2.974 57.702 3.026 57.738 ;
               RECT 2.974 58.302 3.026 58.338 ;
               RECT 2.974 58.902 3.026 58.938 ;
               RECT 2.974 59.502 3.026 59.538 ;
               RECT 2.974 60.102 3.026 60.138 ;
               RECT 2.974 60.702 3.026 60.738 ;
               RECT 2.974 61.302 3.026 61.338 ;
               RECT 2.974 61.902 3.026 61.938 ;
               RECT 2.974 62.502 3.026 62.538 ;
               RECT 2.974 63.102 3.026 63.138 ;
               RECT 2.974 63.702 3.026 63.738 ;
               RECT 2.974 64.302 3.026 64.338 ;
               RECT 2.974 64.902 3.026 64.938 ;
               RECT 2.974 65.502 3.026 65.538 ;
               RECT 2.974 66.102 3.026 66.138 ;
               RECT 2.974 66.702 3.026 66.738 ;
               RECT 2.974 67.302 3.026 67.338 ;
               RECT 2.974 67.902 3.026 67.938 ;
               RECT 2.974 68.502 3.026 68.538 ;
               RECT 2.974 69.102 3.026 69.138 ;
               RECT 2.974 69.702 3.026 69.738 ;
               RECT 2.974 70.302 3.026 70.338 ;
               RECT 2.974 70.902 3.026 70.938 ;
               RECT 2.974 71.502 3.026 71.538 ;
               RECT 2.974 72.102 3.026 72.138 ;
               RECT 2.974 72.702 3.026 72.738 ;
               RECT 2.974 73.302 3.026 73.338 ;
               RECT 2.974 73.902 3.026 73.938 ;
               RECT 2.974 74.502 3.026 74.538 ;
               RECT 2.974 75.102 3.026 75.138 ;
               RECT 2.974 75.702 3.026 75.738 ;
               RECT 2.974 76.302 3.026 76.338 ;
               RECT 2.974 76.902 3.026 76.938 ;
               RECT 2.974 77.502 3.026 77.538 ;
               RECT 2.974 78.102 3.026 78.138 ;
               RECT 2.974 78.702 3.026 78.738 ;
               RECT 2.974 79.302 3.026 79.338 ;
               RECT 2.974 79.902 3.026 79.938 ;
               RECT 2.974 80.502 3.026 80.538 ;
               RECT 2.974 81.102 3.026 81.138 ;
               RECT 2.974 81.702 3.026 81.738 ;
               RECT 2.974 82.302 3.026 82.338 ;
               RECT 2.974 82.902 3.026 82.938 ;
               RECT 2.974 83.502 3.026 83.538 ;
               RECT 2.974 84.102 3.026 84.138 ;
               RECT 2.974 84.702 3.026 84.738 ;
               RECT 2.974 85.302 3.026 85.338 ;
               RECT 2.974 85.902 3.026 85.938 ;
               RECT 2.974 86.502 3.026 86.538 ;
               RECT 2.974 87.102 3.026 87.138 ;
               RECT 2.974 87.702 3.026 87.738 ;
               RECT 2.974 88.302 3.026 88.338 ;
               RECT 2.974 88.902 3.026 88.938 ;
               RECT 2.974 89.502 3.026 89.538 ;
               RECT 2.974 90.102 3.026 90.138 ;
               RECT 2.974 90.702 3.026 90.738 ;
               RECT 2.974 91.302 3.026 91.338 ;
               RECT 2.974 91.902 3.026 91.938 ;
               RECT 2.974 92.502 3.026 92.538 ;
               RECT 2.974 93.102 3.026 93.138 ;
               RECT 2.974 93.702 3.026 93.738 ;
               RECT 2.974 94.302 3.026 94.338 ;
               RECT 2.974 94.902 3.026 94.938 ;
               RECT 2.974 95.502 3.026 95.538 ;
               RECT 2.974 96.102 3.026 96.138 ;
               RECT 2.974 96.702 3.026 96.738 ;
               RECT 2.974 97.302 3.026 97.338 ;
               RECT 2.974 97.902 3.026 97.938 ;
               RECT 2.974 98.502 3.026 98.538 ;
               RECT 2.974 99.102 3.026 99.138 ;
               RECT 2.974 99.702 3.026 99.738 ;
               RECT 2.974 100.302 3.026 100.338 ;
               RECT 2.974 100.902 3.026 100.938 ;
               RECT 2.974 101.502 3.026 101.538 ;
               RECT 2.974 102.102 3.026 102.138 ;
               RECT 2.974 102.702 3.026 102.738 ;
               RECT 2.974 103.302 3.026 103.338 ;
               RECT 2.974 103.902 3.026 103.938 ;
               RECT 2.974 104.502 3.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 20.29 0.5695 20.342 104.5505 ;
               LAYER v4 ;
               RECT 20.29 0.582 20.342 0.618 ;
               RECT 20.29 1.182 20.342 1.218 ;
               RECT 20.29 1.782 20.342 1.818 ;
               RECT 20.29 2.382 20.342 2.418 ;
               RECT 20.29 2.982 20.342 3.018 ;
               RECT 20.29 3.582 20.342 3.618 ;
               RECT 20.29 4.182 20.342 4.218 ;
               RECT 20.29 4.782 20.342 4.818 ;
               RECT 20.29 5.382 20.342 5.418 ;
               RECT 20.29 5.982 20.342 6.018 ;
               RECT 20.29 6.582 20.342 6.618 ;
               RECT 20.29 7.182 20.342 7.218 ;
               RECT 20.29 7.782 20.342 7.818 ;
               RECT 20.29 8.382 20.342 8.418 ;
               RECT 20.29 8.982 20.342 9.018 ;
               RECT 20.29 9.582 20.342 9.618 ;
               RECT 20.29 10.182 20.342 10.218 ;
               RECT 20.29 10.782 20.342 10.818 ;
               RECT 20.29 11.382 20.342 11.418 ;
               RECT 20.29 11.982 20.342 12.018 ;
               RECT 20.29 12.582 20.342 12.618 ;
               RECT 20.29 13.182 20.342 13.218 ;
               RECT 20.29 13.782 20.342 13.818 ;
               RECT 20.29 14.382 20.342 14.418 ;
               RECT 20.29 14.982 20.342 15.018 ;
               RECT 20.29 15.582 20.342 15.618 ;
               RECT 20.29 16.182 20.342 16.218 ;
               RECT 20.29 16.782 20.342 16.818 ;
               RECT 20.29 17.382 20.342 17.418 ;
               RECT 20.29 17.982 20.342 18.018 ;
               RECT 20.29 18.582 20.342 18.618 ;
               RECT 20.29 19.182 20.342 19.218 ;
               RECT 20.29 19.782 20.342 19.818 ;
               RECT 20.29 20.382 20.342 20.418 ;
               RECT 20.29 20.982 20.342 21.018 ;
               RECT 20.29 21.582 20.342 21.618 ;
               RECT 20.29 22.182 20.342 22.218 ;
               RECT 20.29 22.782 20.342 22.818 ;
               RECT 20.29 23.382 20.342 23.418 ;
               RECT 20.29 23.982 20.342 24.018 ;
               RECT 20.29 24.582 20.342 24.618 ;
               RECT 20.29 25.182 20.342 25.218 ;
               RECT 20.29 25.782 20.342 25.818 ;
               RECT 20.29 26.382 20.342 26.418 ;
               RECT 20.29 26.982 20.342 27.018 ;
               RECT 20.29 27.582 20.342 27.618 ;
               RECT 20.29 28.182 20.342 28.218 ;
               RECT 20.29 28.782 20.342 28.818 ;
               RECT 20.29 29.382 20.342 29.418 ;
               RECT 20.29 29.982 20.342 30.018 ;
               RECT 20.29 30.582 20.342 30.618 ;
               RECT 20.29 31.182 20.342 31.218 ;
               RECT 20.29 31.782 20.342 31.818 ;
               RECT 20.29 32.382 20.342 32.418 ;
               RECT 20.29 32.982 20.342 33.018 ;
               RECT 20.29 33.582 20.342 33.618 ;
               RECT 20.29 34.182 20.342 34.218 ;
               RECT 20.29 34.782 20.342 34.818 ;
               RECT 20.29 35.382 20.342 35.418 ;
               RECT 20.29 35.982 20.342 36.018 ;
               RECT 20.29 36.582 20.342 36.618 ;
               RECT 20.29 37.182 20.342 37.218 ;
               RECT 20.29 37.782 20.342 37.818 ;
               RECT 20.29 38.382 20.342 38.418 ;
               RECT 20.29 38.982 20.342 39.018 ;
               RECT 20.29 39.582 20.342 39.618 ;
               RECT 20.29 40.182 20.342 40.218 ;
               RECT 20.29 40.782 20.342 40.818 ;
               RECT 20.29 41.382 20.342 41.418 ;
               RECT 20.29 41.982 20.342 42.018 ;
               RECT 20.29 42.582 20.342 42.618 ;
               RECT 20.29 43.182 20.342 43.218 ;
               RECT 20.29 43.782 20.342 43.818 ;
               RECT 20.29 44.382 20.342 44.418 ;
               RECT 20.29 44.982 20.342 45.018 ;
               RECT 20.29 45.582 20.342 45.618 ;
               RECT 20.29 46.182 20.342 46.218 ;
               RECT 20.29 46.782 20.342 46.818 ;
               RECT 20.29 47.382 20.342 47.418 ;
               RECT 20.29 47.982 20.342 48.018 ;
               RECT 20.29 48.582 20.342 48.618 ;
               RECT 20.29 48.942 20.342 48.978 ;
               RECT 20.29 49.422 20.342 49.458 ;
               RECT 20.29 49.7205 20.342 49.7565 ;
               RECT 20.29 49.902 20.342 49.938 ;
               RECT 20.29 50.382 20.342 50.418 ;
               RECT 20.29 50.862 20.342 50.898 ;
               RECT 20.29 51.342 20.342 51.378 ;
               RECT 20.29 51.822 20.342 51.858 ;
               RECT 20.29 52.302 20.342 52.338 ;
               RECT 20.29 52.662 20.342 52.698 ;
               RECT 20.29 52.782 20.342 52.818 ;
               RECT 20.29 53.262 20.342 53.298 ;
               RECT 20.29 53.742 20.342 53.778 ;
               RECT 20.29 54.2275 20.342 54.2525 ;
               RECT 20.29 54.702 20.342 54.738 ;
               RECT 20.29 55.182 20.342 55.218 ;
               RECT 20.29 55.6675 20.342 55.6925 ;
               RECT 20.29 56.142 20.342 56.178 ;
               RECT 20.29 56.502 20.342 56.538 ;
               RECT 20.29 57.102 20.342 57.138 ;
               RECT 20.29 57.702 20.342 57.738 ;
               RECT 20.29 58.302 20.342 58.338 ;
               RECT 20.29 58.902 20.342 58.938 ;
               RECT 20.29 59.502 20.342 59.538 ;
               RECT 20.29 60.102 20.342 60.138 ;
               RECT 20.29 60.702 20.342 60.738 ;
               RECT 20.29 61.302 20.342 61.338 ;
               RECT 20.29 61.902 20.342 61.938 ;
               RECT 20.29 62.502 20.342 62.538 ;
               RECT 20.29 63.102 20.342 63.138 ;
               RECT 20.29 63.702 20.342 63.738 ;
               RECT 20.29 64.302 20.342 64.338 ;
               RECT 20.29 64.902 20.342 64.938 ;
               RECT 20.29 65.502 20.342 65.538 ;
               RECT 20.29 66.102 20.342 66.138 ;
               RECT 20.29 66.702 20.342 66.738 ;
               RECT 20.29 67.302 20.342 67.338 ;
               RECT 20.29 67.902 20.342 67.938 ;
               RECT 20.29 68.502 20.342 68.538 ;
               RECT 20.29 69.102 20.342 69.138 ;
               RECT 20.29 69.702 20.342 69.738 ;
               RECT 20.29 70.302 20.342 70.338 ;
               RECT 20.29 70.902 20.342 70.938 ;
               RECT 20.29 71.502 20.342 71.538 ;
               RECT 20.29 72.102 20.342 72.138 ;
               RECT 20.29 72.702 20.342 72.738 ;
               RECT 20.29 73.302 20.342 73.338 ;
               RECT 20.29 73.902 20.342 73.938 ;
               RECT 20.29 74.502 20.342 74.538 ;
               RECT 20.29 75.102 20.342 75.138 ;
               RECT 20.29 75.702 20.342 75.738 ;
               RECT 20.29 76.302 20.342 76.338 ;
               RECT 20.29 76.902 20.342 76.938 ;
               RECT 20.29 77.502 20.342 77.538 ;
               RECT 20.29 78.102 20.342 78.138 ;
               RECT 20.29 78.702 20.342 78.738 ;
               RECT 20.29 79.302 20.342 79.338 ;
               RECT 20.29 79.902 20.342 79.938 ;
               RECT 20.29 80.502 20.342 80.538 ;
               RECT 20.29 81.102 20.342 81.138 ;
               RECT 20.29 81.702 20.342 81.738 ;
               RECT 20.29 82.302 20.342 82.338 ;
               RECT 20.29 82.902 20.342 82.938 ;
               RECT 20.29 83.502 20.342 83.538 ;
               RECT 20.29 84.102 20.342 84.138 ;
               RECT 20.29 84.702 20.342 84.738 ;
               RECT 20.29 85.302 20.342 85.338 ;
               RECT 20.29 85.902 20.342 85.938 ;
               RECT 20.29 86.502 20.342 86.538 ;
               RECT 20.29 87.102 20.342 87.138 ;
               RECT 20.29 87.702 20.342 87.738 ;
               RECT 20.29 88.302 20.342 88.338 ;
               RECT 20.29 88.902 20.342 88.938 ;
               RECT 20.29 89.502 20.342 89.538 ;
               RECT 20.29 90.102 20.342 90.138 ;
               RECT 20.29 90.702 20.342 90.738 ;
               RECT 20.29 91.302 20.342 91.338 ;
               RECT 20.29 91.902 20.342 91.938 ;
               RECT 20.29 92.502 20.342 92.538 ;
               RECT 20.29 93.102 20.342 93.138 ;
               RECT 20.29 93.702 20.342 93.738 ;
               RECT 20.29 94.302 20.342 94.338 ;
               RECT 20.29 94.902 20.342 94.938 ;
               RECT 20.29 95.502 20.342 95.538 ;
               RECT 20.29 96.102 20.342 96.138 ;
               RECT 20.29 96.702 20.342 96.738 ;
               RECT 20.29 97.302 20.342 97.338 ;
               RECT 20.29 97.902 20.342 97.938 ;
               RECT 20.29 98.502 20.342 98.538 ;
               RECT 20.29 99.102 20.342 99.138 ;
               RECT 20.29 99.702 20.342 99.738 ;
               RECT 20.29 100.302 20.342 100.338 ;
               RECT 20.29 100.902 20.342 100.938 ;
               RECT 20.29 101.502 20.342 101.538 ;
               RECT 20.29 102.102 20.342 102.138 ;
               RECT 20.29 102.702 20.342 102.738 ;
               RECT 20.29 103.302 20.342 103.338 ;
               RECT 20.29 103.902 20.342 103.938 ;
               RECT 20.29 104.502 20.342 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 21.496 0.5695 21.55 104.5505 ;
               LAYER v4 ;
               RECT 21.496 0.582 21.55 0.618 ;
               RECT 21.496 1.182 21.55 1.218 ;
               RECT 21.496 1.782 21.55 1.818 ;
               RECT 21.496 2.382 21.55 2.418 ;
               RECT 21.496 2.982 21.55 3.018 ;
               RECT 21.496 3.582 21.55 3.618 ;
               RECT 21.496 4.182 21.55 4.218 ;
               RECT 21.496 4.782 21.55 4.818 ;
               RECT 21.496 5.382 21.55 5.418 ;
               RECT 21.496 5.982 21.55 6.018 ;
               RECT 21.496 6.582 21.55 6.618 ;
               RECT 21.496 7.182 21.55 7.218 ;
               RECT 21.496 7.782 21.55 7.818 ;
               RECT 21.496 8.382 21.55 8.418 ;
               RECT 21.496 8.982 21.55 9.018 ;
               RECT 21.496 9.582 21.55 9.618 ;
               RECT 21.496 10.182 21.55 10.218 ;
               RECT 21.496 10.782 21.55 10.818 ;
               RECT 21.496 11.382 21.55 11.418 ;
               RECT 21.496 11.982 21.55 12.018 ;
               RECT 21.496 12.582 21.55 12.618 ;
               RECT 21.496 13.182 21.55 13.218 ;
               RECT 21.496 13.782 21.55 13.818 ;
               RECT 21.496 14.382 21.55 14.418 ;
               RECT 21.496 14.982 21.55 15.018 ;
               RECT 21.496 15.582 21.55 15.618 ;
               RECT 21.496 16.182 21.55 16.218 ;
               RECT 21.496 16.782 21.55 16.818 ;
               RECT 21.496 17.382 21.55 17.418 ;
               RECT 21.496 17.982 21.55 18.018 ;
               RECT 21.496 18.582 21.55 18.618 ;
               RECT 21.496 19.182 21.55 19.218 ;
               RECT 21.496 19.782 21.55 19.818 ;
               RECT 21.496 20.382 21.55 20.418 ;
               RECT 21.496 20.982 21.55 21.018 ;
               RECT 21.496 21.582 21.55 21.618 ;
               RECT 21.496 22.182 21.55 22.218 ;
               RECT 21.496 22.782 21.55 22.818 ;
               RECT 21.496 23.382 21.55 23.418 ;
               RECT 21.496 23.982 21.55 24.018 ;
               RECT 21.496 24.582 21.55 24.618 ;
               RECT 21.496 25.182 21.55 25.218 ;
               RECT 21.496 25.782 21.55 25.818 ;
               RECT 21.496 26.382 21.55 26.418 ;
               RECT 21.496 26.982 21.55 27.018 ;
               RECT 21.496 27.582 21.55 27.618 ;
               RECT 21.496 28.182 21.55 28.218 ;
               RECT 21.496 28.782 21.55 28.818 ;
               RECT 21.496 29.382 21.55 29.418 ;
               RECT 21.496 29.982 21.55 30.018 ;
               RECT 21.496 30.582 21.55 30.618 ;
               RECT 21.496 31.182 21.55 31.218 ;
               RECT 21.496 31.782 21.55 31.818 ;
               RECT 21.496 32.382 21.55 32.418 ;
               RECT 21.496 32.982 21.55 33.018 ;
               RECT 21.496 33.582 21.55 33.618 ;
               RECT 21.496 34.182 21.55 34.218 ;
               RECT 21.496 34.782 21.55 34.818 ;
               RECT 21.496 35.382 21.55 35.418 ;
               RECT 21.496 35.982 21.55 36.018 ;
               RECT 21.496 36.582 21.55 36.618 ;
               RECT 21.496 37.182 21.55 37.218 ;
               RECT 21.496 37.782 21.55 37.818 ;
               RECT 21.496 38.382 21.55 38.418 ;
               RECT 21.496 38.982 21.55 39.018 ;
               RECT 21.496 39.582 21.55 39.618 ;
               RECT 21.496 40.182 21.55 40.218 ;
               RECT 21.496 40.782 21.55 40.818 ;
               RECT 21.496 41.382 21.55 41.418 ;
               RECT 21.496 41.982 21.55 42.018 ;
               RECT 21.496 42.582 21.55 42.618 ;
               RECT 21.496 43.182 21.55 43.218 ;
               RECT 21.496 43.782 21.55 43.818 ;
               RECT 21.496 44.382 21.55 44.418 ;
               RECT 21.496 44.982 21.55 45.018 ;
               RECT 21.496 45.582 21.55 45.618 ;
               RECT 21.496 46.182 21.55 46.218 ;
               RECT 21.496 46.782 21.55 46.818 ;
               RECT 21.496 47.382 21.55 47.418 ;
               RECT 21.496 47.982 21.55 48.018 ;
               RECT 21.496 48.582 21.55 48.618 ;
               RECT 21.496 48.942 21.55 48.978 ;
               RECT 21.496 49.422 21.55 49.458 ;
               RECT 21.496 49.902 21.55 49.938 ;
               RECT 21.496 50.0835 21.55 50.1195 ;
               RECT 21.496 50.382 21.55 50.418 ;
               RECT 21.496 50.862 21.55 50.898 ;
               RECT 21.496 51.342 21.55 51.378 ;
               RECT 21.496 51.822 21.55 51.858 ;
               RECT 21.496 52.302 21.55 52.338 ;
               RECT 21.496 52.662 21.55 52.698 ;
               RECT 21.496 52.782 21.55 52.818 ;
               RECT 21.496 53.262 21.55 53.298 ;
               RECT 21.496 53.742 21.55 53.778 ;
               RECT 21.496 54.222 21.55 54.258 ;
               RECT 21.496 54.702 21.55 54.738 ;
               RECT 21.496 55.182 21.55 55.218 ;
               RECT 21.496 55.662 21.55 55.698 ;
               RECT 21.496 56.142 21.55 56.178 ;
               RECT 21.496 56.502 21.55 56.538 ;
               RECT 21.496 57.102 21.55 57.138 ;
               RECT 21.496 57.702 21.55 57.738 ;
               RECT 21.496 58.302 21.55 58.338 ;
               RECT 21.496 58.902 21.55 58.938 ;
               RECT 21.496 59.502 21.55 59.538 ;
               RECT 21.496 60.102 21.55 60.138 ;
               RECT 21.496 60.702 21.55 60.738 ;
               RECT 21.496 61.302 21.55 61.338 ;
               RECT 21.496 61.902 21.55 61.938 ;
               RECT 21.496 62.502 21.55 62.538 ;
               RECT 21.496 63.102 21.55 63.138 ;
               RECT 21.496 63.702 21.55 63.738 ;
               RECT 21.496 64.302 21.55 64.338 ;
               RECT 21.496 64.902 21.55 64.938 ;
               RECT 21.496 65.502 21.55 65.538 ;
               RECT 21.496 66.102 21.55 66.138 ;
               RECT 21.496 66.702 21.55 66.738 ;
               RECT 21.496 67.302 21.55 67.338 ;
               RECT 21.496 67.902 21.55 67.938 ;
               RECT 21.496 68.502 21.55 68.538 ;
               RECT 21.496 69.102 21.55 69.138 ;
               RECT 21.496 69.702 21.55 69.738 ;
               RECT 21.496 70.302 21.55 70.338 ;
               RECT 21.496 70.902 21.55 70.938 ;
               RECT 21.496 71.502 21.55 71.538 ;
               RECT 21.496 72.102 21.55 72.138 ;
               RECT 21.496 72.702 21.55 72.738 ;
               RECT 21.496 73.302 21.55 73.338 ;
               RECT 21.496 73.902 21.55 73.938 ;
               RECT 21.496 74.502 21.55 74.538 ;
               RECT 21.496 75.102 21.55 75.138 ;
               RECT 21.496 75.702 21.55 75.738 ;
               RECT 21.496 76.302 21.55 76.338 ;
               RECT 21.496 76.902 21.55 76.938 ;
               RECT 21.496 77.502 21.55 77.538 ;
               RECT 21.496 78.102 21.55 78.138 ;
               RECT 21.496 78.702 21.55 78.738 ;
               RECT 21.496 79.302 21.55 79.338 ;
               RECT 21.496 79.902 21.55 79.938 ;
               RECT 21.496 80.502 21.55 80.538 ;
               RECT 21.496 81.102 21.55 81.138 ;
               RECT 21.496 81.702 21.55 81.738 ;
               RECT 21.496 82.302 21.55 82.338 ;
               RECT 21.496 82.902 21.55 82.938 ;
               RECT 21.496 83.502 21.55 83.538 ;
               RECT 21.496 84.102 21.55 84.138 ;
               RECT 21.496 84.702 21.55 84.738 ;
               RECT 21.496 85.302 21.55 85.338 ;
               RECT 21.496 85.902 21.55 85.938 ;
               RECT 21.496 86.502 21.55 86.538 ;
               RECT 21.496 87.102 21.55 87.138 ;
               RECT 21.496 87.702 21.55 87.738 ;
               RECT 21.496 88.302 21.55 88.338 ;
               RECT 21.496 88.902 21.55 88.938 ;
               RECT 21.496 89.502 21.55 89.538 ;
               RECT 21.496 90.102 21.55 90.138 ;
               RECT 21.496 90.702 21.55 90.738 ;
               RECT 21.496 91.302 21.55 91.338 ;
               RECT 21.496 91.902 21.55 91.938 ;
               RECT 21.496 92.502 21.55 92.538 ;
               RECT 21.496 93.102 21.55 93.138 ;
               RECT 21.496 93.702 21.55 93.738 ;
               RECT 21.496 94.302 21.55 94.338 ;
               RECT 21.496 94.902 21.55 94.938 ;
               RECT 21.496 95.502 21.55 95.538 ;
               RECT 21.496 96.102 21.55 96.138 ;
               RECT 21.496 96.702 21.55 96.738 ;
               RECT 21.496 97.302 21.55 97.338 ;
               RECT 21.496 97.902 21.55 97.938 ;
               RECT 21.496 98.502 21.55 98.538 ;
               RECT 21.496 99.102 21.55 99.138 ;
               RECT 21.496 99.702 21.55 99.738 ;
               RECT 21.496 100.302 21.55 100.338 ;
               RECT 21.496 100.902 21.55 100.938 ;
               RECT 21.496 101.502 21.55 101.538 ;
               RECT 21.496 102.102 21.55 102.138 ;
               RECT 21.496 102.702 21.55 102.738 ;
               RECT 21.496 103.302 21.55 103.338 ;
               RECT 21.496 103.902 21.55 103.938 ;
               RECT 21.496 104.502 21.55 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 22.774 0.5695 22.826 104.5505 ;
               LAYER v4 ;
               RECT 22.774 0.582 22.826 0.618 ;
               RECT 22.774 1.182 22.826 1.218 ;
               RECT 22.774 1.782 22.826 1.818 ;
               RECT 22.774 2.382 22.826 2.418 ;
               RECT 22.774 2.982 22.826 3.018 ;
               RECT 22.774 3.582 22.826 3.618 ;
               RECT 22.774 4.182 22.826 4.218 ;
               RECT 22.774 4.782 22.826 4.818 ;
               RECT 22.774 5.382 22.826 5.418 ;
               RECT 22.774 5.982 22.826 6.018 ;
               RECT 22.774 6.582 22.826 6.618 ;
               RECT 22.774 7.182 22.826 7.218 ;
               RECT 22.774 7.782 22.826 7.818 ;
               RECT 22.774 8.382 22.826 8.418 ;
               RECT 22.774 8.982 22.826 9.018 ;
               RECT 22.774 9.582 22.826 9.618 ;
               RECT 22.774 10.182 22.826 10.218 ;
               RECT 22.774 10.782 22.826 10.818 ;
               RECT 22.774 11.382 22.826 11.418 ;
               RECT 22.774 11.982 22.826 12.018 ;
               RECT 22.774 12.582 22.826 12.618 ;
               RECT 22.774 13.182 22.826 13.218 ;
               RECT 22.774 13.782 22.826 13.818 ;
               RECT 22.774 14.382 22.826 14.418 ;
               RECT 22.774 14.982 22.826 15.018 ;
               RECT 22.774 15.582 22.826 15.618 ;
               RECT 22.774 16.182 22.826 16.218 ;
               RECT 22.774 16.782 22.826 16.818 ;
               RECT 22.774 17.382 22.826 17.418 ;
               RECT 22.774 17.982 22.826 18.018 ;
               RECT 22.774 18.582 22.826 18.618 ;
               RECT 22.774 19.182 22.826 19.218 ;
               RECT 22.774 19.782 22.826 19.818 ;
               RECT 22.774 20.382 22.826 20.418 ;
               RECT 22.774 20.982 22.826 21.018 ;
               RECT 22.774 21.582 22.826 21.618 ;
               RECT 22.774 22.182 22.826 22.218 ;
               RECT 22.774 22.782 22.826 22.818 ;
               RECT 22.774 23.382 22.826 23.418 ;
               RECT 22.774 23.982 22.826 24.018 ;
               RECT 22.774 24.582 22.826 24.618 ;
               RECT 22.774 25.182 22.826 25.218 ;
               RECT 22.774 25.782 22.826 25.818 ;
               RECT 22.774 26.382 22.826 26.418 ;
               RECT 22.774 26.982 22.826 27.018 ;
               RECT 22.774 27.582 22.826 27.618 ;
               RECT 22.774 28.182 22.826 28.218 ;
               RECT 22.774 28.782 22.826 28.818 ;
               RECT 22.774 29.382 22.826 29.418 ;
               RECT 22.774 29.982 22.826 30.018 ;
               RECT 22.774 30.582 22.826 30.618 ;
               RECT 22.774 31.182 22.826 31.218 ;
               RECT 22.774 31.782 22.826 31.818 ;
               RECT 22.774 32.382 22.826 32.418 ;
               RECT 22.774 32.982 22.826 33.018 ;
               RECT 22.774 33.582 22.826 33.618 ;
               RECT 22.774 34.182 22.826 34.218 ;
               RECT 22.774 34.782 22.826 34.818 ;
               RECT 22.774 35.382 22.826 35.418 ;
               RECT 22.774 35.982 22.826 36.018 ;
               RECT 22.774 36.582 22.826 36.618 ;
               RECT 22.774 37.182 22.826 37.218 ;
               RECT 22.774 37.782 22.826 37.818 ;
               RECT 22.774 38.382 22.826 38.418 ;
               RECT 22.774 38.982 22.826 39.018 ;
               RECT 22.774 39.582 22.826 39.618 ;
               RECT 22.774 40.182 22.826 40.218 ;
               RECT 22.774 40.782 22.826 40.818 ;
               RECT 22.774 41.382 22.826 41.418 ;
               RECT 22.774 41.982 22.826 42.018 ;
               RECT 22.774 42.582 22.826 42.618 ;
               RECT 22.774 43.182 22.826 43.218 ;
               RECT 22.774 43.782 22.826 43.818 ;
               RECT 22.774 44.382 22.826 44.418 ;
               RECT 22.774 44.982 22.826 45.018 ;
               RECT 22.774 45.582 22.826 45.618 ;
               RECT 22.774 46.182 22.826 46.218 ;
               RECT 22.774 46.782 22.826 46.818 ;
               RECT 22.774 47.382 22.826 47.418 ;
               RECT 22.774 47.982 22.826 48.018 ;
               RECT 22.774 48.582 22.826 48.618 ;
               RECT 22.774 48.942 22.826 48.978 ;
               RECT 22.774 49.182 22.826 49.218 ;
               RECT 22.774 49.902 22.826 49.938 ;
               RECT 22.774 50.622 22.826 50.658 ;
               RECT 22.774 50.862 22.826 50.898 ;
               RECT 22.774 51.342 22.826 51.378 ;
               RECT 22.774 51.822 22.826 51.858 ;
               RECT 22.774 52.302 22.826 52.338 ;
               RECT 22.774 52.782 22.826 52.818 ;
               RECT 22.774 53.262 22.826 53.298 ;
               RECT 22.774 53.742 22.826 53.778 ;
               RECT 22.774 54.222 22.826 54.258 ;
               RECT 22.774 54.462 22.826 54.498 ;
               RECT 22.774 55.182 22.826 55.218 ;
               RECT 22.774 55.902 22.826 55.938 ;
               RECT 22.774 56.142 22.826 56.178 ;
               RECT 22.774 56.502 22.826 56.538 ;
               RECT 22.774 57.102 22.826 57.138 ;
               RECT 22.774 57.702 22.826 57.738 ;
               RECT 22.774 58.302 22.826 58.338 ;
               RECT 22.774 58.902 22.826 58.938 ;
               RECT 22.774 59.502 22.826 59.538 ;
               RECT 22.774 60.102 22.826 60.138 ;
               RECT 22.774 60.702 22.826 60.738 ;
               RECT 22.774 61.302 22.826 61.338 ;
               RECT 22.774 61.902 22.826 61.938 ;
               RECT 22.774 62.502 22.826 62.538 ;
               RECT 22.774 63.102 22.826 63.138 ;
               RECT 22.774 63.702 22.826 63.738 ;
               RECT 22.774 64.302 22.826 64.338 ;
               RECT 22.774 64.902 22.826 64.938 ;
               RECT 22.774 65.502 22.826 65.538 ;
               RECT 22.774 66.102 22.826 66.138 ;
               RECT 22.774 66.702 22.826 66.738 ;
               RECT 22.774 67.302 22.826 67.338 ;
               RECT 22.774 67.902 22.826 67.938 ;
               RECT 22.774 68.502 22.826 68.538 ;
               RECT 22.774 69.102 22.826 69.138 ;
               RECT 22.774 69.702 22.826 69.738 ;
               RECT 22.774 70.302 22.826 70.338 ;
               RECT 22.774 70.902 22.826 70.938 ;
               RECT 22.774 71.502 22.826 71.538 ;
               RECT 22.774 72.102 22.826 72.138 ;
               RECT 22.774 72.702 22.826 72.738 ;
               RECT 22.774 73.302 22.826 73.338 ;
               RECT 22.774 73.902 22.826 73.938 ;
               RECT 22.774 74.502 22.826 74.538 ;
               RECT 22.774 75.102 22.826 75.138 ;
               RECT 22.774 75.702 22.826 75.738 ;
               RECT 22.774 76.302 22.826 76.338 ;
               RECT 22.774 76.902 22.826 76.938 ;
               RECT 22.774 77.502 22.826 77.538 ;
               RECT 22.774 78.102 22.826 78.138 ;
               RECT 22.774 78.702 22.826 78.738 ;
               RECT 22.774 79.302 22.826 79.338 ;
               RECT 22.774 79.902 22.826 79.938 ;
               RECT 22.774 80.502 22.826 80.538 ;
               RECT 22.774 81.102 22.826 81.138 ;
               RECT 22.774 81.702 22.826 81.738 ;
               RECT 22.774 82.302 22.826 82.338 ;
               RECT 22.774 82.902 22.826 82.938 ;
               RECT 22.774 83.502 22.826 83.538 ;
               RECT 22.774 84.102 22.826 84.138 ;
               RECT 22.774 84.702 22.826 84.738 ;
               RECT 22.774 85.302 22.826 85.338 ;
               RECT 22.774 85.902 22.826 85.938 ;
               RECT 22.774 86.502 22.826 86.538 ;
               RECT 22.774 87.102 22.826 87.138 ;
               RECT 22.774 87.702 22.826 87.738 ;
               RECT 22.774 88.302 22.826 88.338 ;
               RECT 22.774 88.902 22.826 88.938 ;
               RECT 22.774 89.502 22.826 89.538 ;
               RECT 22.774 90.102 22.826 90.138 ;
               RECT 22.774 90.702 22.826 90.738 ;
               RECT 22.774 91.302 22.826 91.338 ;
               RECT 22.774 91.902 22.826 91.938 ;
               RECT 22.774 92.502 22.826 92.538 ;
               RECT 22.774 93.102 22.826 93.138 ;
               RECT 22.774 93.702 22.826 93.738 ;
               RECT 22.774 94.302 22.826 94.338 ;
               RECT 22.774 94.902 22.826 94.938 ;
               RECT 22.774 95.502 22.826 95.538 ;
               RECT 22.774 96.102 22.826 96.138 ;
               RECT 22.774 96.702 22.826 96.738 ;
               RECT 22.774 97.302 22.826 97.338 ;
               RECT 22.774 97.902 22.826 97.938 ;
               RECT 22.774 98.502 22.826 98.538 ;
               RECT 22.774 99.102 22.826 99.138 ;
               RECT 22.774 99.702 22.826 99.738 ;
               RECT 22.774 100.302 22.826 100.338 ;
               RECT 22.774 100.902 22.826 100.938 ;
               RECT 22.774 101.502 22.826 101.538 ;
               RECT 22.774 102.102 22.826 102.138 ;
               RECT 22.774 102.702 22.826 102.738 ;
               RECT 22.774 103.302 22.826 103.338 ;
               RECT 22.774 103.902 22.826 103.938 ;
               RECT 22.774 104.502 22.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 23.574 0.5695 23.626 104.5505 ;
               LAYER v4 ;
               RECT 23.574 0.582 23.626 0.618 ;
               RECT 23.574 1.182 23.626 1.218 ;
               RECT 23.574 1.782 23.626 1.818 ;
               RECT 23.574 2.382 23.626 2.418 ;
               RECT 23.574 2.982 23.626 3.018 ;
               RECT 23.574 3.582 23.626 3.618 ;
               RECT 23.574 4.182 23.626 4.218 ;
               RECT 23.574 4.782 23.626 4.818 ;
               RECT 23.574 5.382 23.626 5.418 ;
               RECT 23.574 5.982 23.626 6.018 ;
               RECT 23.574 6.582 23.626 6.618 ;
               RECT 23.574 7.182 23.626 7.218 ;
               RECT 23.574 7.782 23.626 7.818 ;
               RECT 23.574 8.382 23.626 8.418 ;
               RECT 23.574 8.982 23.626 9.018 ;
               RECT 23.574 9.582 23.626 9.618 ;
               RECT 23.574 10.182 23.626 10.218 ;
               RECT 23.574 10.782 23.626 10.818 ;
               RECT 23.574 11.382 23.626 11.418 ;
               RECT 23.574 11.982 23.626 12.018 ;
               RECT 23.574 12.582 23.626 12.618 ;
               RECT 23.574 13.182 23.626 13.218 ;
               RECT 23.574 13.782 23.626 13.818 ;
               RECT 23.574 14.382 23.626 14.418 ;
               RECT 23.574 14.982 23.626 15.018 ;
               RECT 23.574 15.582 23.626 15.618 ;
               RECT 23.574 16.182 23.626 16.218 ;
               RECT 23.574 16.782 23.626 16.818 ;
               RECT 23.574 17.382 23.626 17.418 ;
               RECT 23.574 17.982 23.626 18.018 ;
               RECT 23.574 18.582 23.626 18.618 ;
               RECT 23.574 19.182 23.626 19.218 ;
               RECT 23.574 19.782 23.626 19.818 ;
               RECT 23.574 20.382 23.626 20.418 ;
               RECT 23.574 20.982 23.626 21.018 ;
               RECT 23.574 21.582 23.626 21.618 ;
               RECT 23.574 22.182 23.626 22.218 ;
               RECT 23.574 22.782 23.626 22.818 ;
               RECT 23.574 23.382 23.626 23.418 ;
               RECT 23.574 23.982 23.626 24.018 ;
               RECT 23.574 24.582 23.626 24.618 ;
               RECT 23.574 25.182 23.626 25.218 ;
               RECT 23.574 25.782 23.626 25.818 ;
               RECT 23.574 26.382 23.626 26.418 ;
               RECT 23.574 26.982 23.626 27.018 ;
               RECT 23.574 27.582 23.626 27.618 ;
               RECT 23.574 28.182 23.626 28.218 ;
               RECT 23.574 28.782 23.626 28.818 ;
               RECT 23.574 29.382 23.626 29.418 ;
               RECT 23.574 29.982 23.626 30.018 ;
               RECT 23.574 30.582 23.626 30.618 ;
               RECT 23.574 31.182 23.626 31.218 ;
               RECT 23.574 31.782 23.626 31.818 ;
               RECT 23.574 32.382 23.626 32.418 ;
               RECT 23.574 32.982 23.626 33.018 ;
               RECT 23.574 33.582 23.626 33.618 ;
               RECT 23.574 34.182 23.626 34.218 ;
               RECT 23.574 34.782 23.626 34.818 ;
               RECT 23.574 35.382 23.626 35.418 ;
               RECT 23.574 35.982 23.626 36.018 ;
               RECT 23.574 36.582 23.626 36.618 ;
               RECT 23.574 37.182 23.626 37.218 ;
               RECT 23.574 37.782 23.626 37.818 ;
               RECT 23.574 38.382 23.626 38.418 ;
               RECT 23.574 38.982 23.626 39.018 ;
               RECT 23.574 39.582 23.626 39.618 ;
               RECT 23.574 40.182 23.626 40.218 ;
               RECT 23.574 40.782 23.626 40.818 ;
               RECT 23.574 41.382 23.626 41.418 ;
               RECT 23.574 41.982 23.626 42.018 ;
               RECT 23.574 42.582 23.626 42.618 ;
               RECT 23.574 43.182 23.626 43.218 ;
               RECT 23.574 43.782 23.626 43.818 ;
               RECT 23.574 44.382 23.626 44.418 ;
               RECT 23.574 44.982 23.626 45.018 ;
               RECT 23.574 45.582 23.626 45.618 ;
               RECT 23.574 46.182 23.626 46.218 ;
               RECT 23.574 46.782 23.626 46.818 ;
               RECT 23.574 47.382 23.626 47.418 ;
               RECT 23.574 47.982 23.626 48.018 ;
               RECT 23.574 48.582 23.626 48.618 ;
               RECT 23.574 48.942 23.626 48.978 ;
               RECT 23.574 49.182 23.626 49.218 ;
               RECT 23.574 49.902 23.626 49.938 ;
               RECT 23.574 50.622 23.626 50.658 ;
               RECT 23.574 50.862 23.626 50.898 ;
               RECT 23.574 51.342 23.626 51.378 ;
               RECT 23.574 51.822 23.626 51.858 ;
               RECT 23.574 52.302 23.626 52.338 ;
               RECT 23.574 52.782 23.626 52.818 ;
               RECT 23.574 53.262 23.626 53.298 ;
               RECT 23.574 53.742 23.626 53.778 ;
               RECT 23.574 54.222 23.626 54.258 ;
               RECT 23.574 54.462 23.626 54.498 ;
               RECT 23.574 55.182 23.626 55.218 ;
               RECT 23.574 55.902 23.626 55.938 ;
               RECT 23.574 56.142 23.626 56.178 ;
               RECT 23.574 56.502 23.626 56.538 ;
               RECT 23.574 57.102 23.626 57.138 ;
               RECT 23.574 57.702 23.626 57.738 ;
               RECT 23.574 58.302 23.626 58.338 ;
               RECT 23.574 58.902 23.626 58.938 ;
               RECT 23.574 59.502 23.626 59.538 ;
               RECT 23.574 60.102 23.626 60.138 ;
               RECT 23.574 60.702 23.626 60.738 ;
               RECT 23.574 61.302 23.626 61.338 ;
               RECT 23.574 61.902 23.626 61.938 ;
               RECT 23.574 62.502 23.626 62.538 ;
               RECT 23.574 63.102 23.626 63.138 ;
               RECT 23.574 63.702 23.626 63.738 ;
               RECT 23.574 64.302 23.626 64.338 ;
               RECT 23.574 64.902 23.626 64.938 ;
               RECT 23.574 65.502 23.626 65.538 ;
               RECT 23.574 66.102 23.626 66.138 ;
               RECT 23.574 66.702 23.626 66.738 ;
               RECT 23.574 67.302 23.626 67.338 ;
               RECT 23.574 67.902 23.626 67.938 ;
               RECT 23.574 68.502 23.626 68.538 ;
               RECT 23.574 69.102 23.626 69.138 ;
               RECT 23.574 69.702 23.626 69.738 ;
               RECT 23.574 70.302 23.626 70.338 ;
               RECT 23.574 70.902 23.626 70.938 ;
               RECT 23.574 71.502 23.626 71.538 ;
               RECT 23.574 72.102 23.626 72.138 ;
               RECT 23.574 72.702 23.626 72.738 ;
               RECT 23.574 73.302 23.626 73.338 ;
               RECT 23.574 73.902 23.626 73.938 ;
               RECT 23.574 74.502 23.626 74.538 ;
               RECT 23.574 75.102 23.626 75.138 ;
               RECT 23.574 75.702 23.626 75.738 ;
               RECT 23.574 76.302 23.626 76.338 ;
               RECT 23.574 76.902 23.626 76.938 ;
               RECT 23.574 77.502 23.626 77.538 ;
               RECT 23.574 78.102 23.626 78.138 ;
               RECT 23.574 78.702 23.626 78.738 ;
               RECT 23.574 79.302 23.626 79.338 ;
               RECT 23.574 79.902 23.626 79.938 ;
               RECT 23.574 80.502 23.626 80.538 ;
               RECT 23.574 81.102 23.626 81.138 ;
               RECT 23.574 81.702 23.626 81.738 ;
               RECT 23.574 82.302 23.626 82.338 ;
               RECT 23.574 82.902 23.626 82.938 ;
               RECT 23.574 83.502 23.626 83.538 ;
               RECT 23.574 84.102 23.626 84.138 ;
               RECT 23.574 84.702 23.626 84.738 ;
               RECT 23.574 85.302 23.626 85.338 ;
               RECT 23.574 85.902 23.626 85.938 ;
               RECT 23.574 86.502 23.626 86.538 ;
               RECT 23.574 87.102 23.626 87.138 ;
               RECT 23.574 87.702 23.626 87.738 ;
               RECT 23.574 88.302 23.626 88.338 ;
               RECT 23.574 88.902 23.626 88.938 ;
               RECT 23.574 89.502 23.626 89.538 ;
               RECT 23.574 90.102 23.626 90.138 ;
               RECT 23.574 90.702 23.626 90.738 ;
               RECT 23.574 91.302 23.626 91.338 ;
               RECT 23.574 91.902 23.626 91.938 ;
               RECT 23.574 92.502 23.626 92.538 ;
               RECT 23.574 93.102 23.626 93.138 ;
               RECT 23.574 93.702 23.626 93.738 ;
               RECT 23.574 94.302 23.626 94.338 ;
               RECT 23.574 94.902 23.626 94.938 ;
               RECT 23.574 95.502 23.626 95.538 ;
               RECT 23.574 96.102 23.626 96.138 ;
               RECT 23.574 96.702 23.626 96.738 ;
               RECT 23.574 97.302 23.626 97.338 ;
               RECT 23.574 97.902 23.626 97.938 ;
               RECT 23.574 98.502 23.626 98.538 ;
               RECT 23.574 99.102 23.626 99.138 ;
               RECT 23.574 99.702 23.626 99.738 ;
               RECT 23.574 100.302 23.626 100.338 ;
               RECT 23.574 100.902 23.626 100.938 ;
               RECT 23.574 101.502 23.626 101.538 ;
               RECT 23.574 102.102 23.626 102.138 ;
               RECT 23.574 102.702 23.626 102.738 ;
               RECT 23.574 103.302 23.626 103.338 ;
               RECT 23.574 103.902 23.626 103.938 ;
               RECT 23.574 104.502 23.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 24.374 0.5695 24.426 104.5505 ;
               LAYER v4 ;
               RECT 24.374 0.582 24.426 0.618 ;
               RECT 24.374 1.182 24.426 1.218 ;
               RECT 24.374 1.782 24.426 1.818 ;
               RECT 24.374 2.382 24.426 2.418 ;
               RECT 24.374 2.982 24.426 3.018 ;
               RECT 24.374 3.582 24.426 3.618 ;
               RECT 24.374 4.182 24.426 4.218 ;
               RECT 24.374 4.782 24.426 4.818 ;
               RECT 24.374 5.382 24.426 5.418 ;
               RECT 24.374 5.982 24.426 6.018 ;
               RECT 24.374 6.582 24.426 6.618 ;
               RECT 24.374 7.182 24.426 7.218 ;
               RECT 24.374 7.782 24.426 7.818 ;
               RECT 24.374 8.382 24.426 8.418 ;
               RECT 24.374 8.982 24.426 9.018 ;
               RECT 24.374 9.582 24.426 9.618 ;
               RECT 24.374 10.182 24.426 10.218 ;
               RECT 24.374 10.782 24.426 10.818 ;
               RECT 24.374 11.382 24.426 11.418 ;
               RECT 24.374 11.982 24.426 12.018 ;
               RECT 24.374 12.582 24.426 12.618 ;
               RECT 24.374 13.182 24.426 13.218 ;
               RECT 24.374 13.782 24.426 13.818 ;
               RECT 24.374 14.382 24.426 14.418 ;
               RECT 24.374 14.982 24.426 15.018 ;
               RECT 24.374 15.582 24.426 15.618 ;
               RECT 24.374 16.182 24.426 16.218 ;
               RECT 24.374 16.782 24.426 16.818 ;
               RECT 24.374 17.382 24.426 17.418 ;
               RECT 24.374 17.982 24.426 18.018 ;
               RECT 24.374 18.582 24.426 18.618 ;
               RECT 24.374 19.182 24.426 19.218 ;
               RECT 24.374 19.782 24.426 19.818 ;
               RECT 24.374 20.382 24.426 20.418 ;
               RECT 24.374 20.982 24.426 21.018 ;
               RECT 24.374 21.582 24.426 21.618 ;
               RECT 24.374 22.182 24.426 22.218 ;
               RECT 24.374 22.782 24.426 22.818 ;
               RECT 24.374 23.382 24.426 23.418 ;
               RECT 24.374 23.982 24.426 24.018 ;
               RECT 24.374 24.582 24.426 24.618 ;
               RECT 24.374 25.182 24.426 25.218 ;
               RECT 24.374 25.782 24.426 25.818 ;
               RECT 24.374 26.382 24.426 26.418 ;
               RECT 24.374 26.982 24.426 27.018 ;
               RECT 24.374 27.582 24.426 27.618 ;
               RECT 24.374 28.182 24.426 28.218 ;
               RECT 24.374 28.782 24.426 28.818 ;
               RECT 24.374 29.382 24.426 29.418 ;
               RECT 24.374 29.982 24.426 30.018 ;
               RECT 24.374 30.582 24.426 30.618 ;
               RECT 24.374 31.182 24.426 31.218 ;
               RECT 24.374 31.782 24.426 31.818 ;
               RECT 24.374 32.382 24.426 32.418 ;
               RECT 24.374 32.982 24.426 33.018 ;
               RECT 24.374 33.582 24.426 33.618 ;
               RECT 24.374 34.182 24.426 34.218 ;
               RECT 24.374 34.782 24.426 34.818 ;
               RECT 24.374 35.382 24.426 35.418 ;
               RECT 24.374 35.982 24.426 36.018 ;
               RECT 24.374 36.582 24.426 36.618 ;
               RECT 24.374 37.182 24.426 37.218 ;
               RECT 24.374 37.782 24.426 37.818 ;
               RECT 24.374 38.382 24.426 38.418 ;
               RECT 24.374 38.982 24.426 39.018 ;
               RECT 24.374 39.582 24.426 39.618 ;
               RECT 24.374 40.182 24.426 40.218 ;
               RECT 24.374 40.782 24.426 40.818 ;
               RECT 24.374 41.382 24.426 41.418 ;
               RECT 24.374 41.982 24.426 42.018 ;
               RECT 24.374 42.582 24.426 42.618 ;
               RECT 24.374 43.182 24.426 43.218 ;
               RECT 24.374 43.782 24.426 43.818 ;
               RECT 24.374 44.382 24.426 44.418 ;
               RECT 24.374 44.982 24.426 45.018 ;
               RECT 24.374 45.582 24.426 45.618 ;
               RECT 24.374 46.182 24.426 46.218 ;
               RECT 24.374 46.782 24.426 46.818 ;
               RECT 24.374 47.382 24.426 47.418 ;
               RECT 24.374 47.982 24.426 48.018 ;
               RECT 24.374 48.582 24.426 48.618 ;
               RECT 24.374 48.942 24.426 48.978 ;
               RECT 24.374 48.9475 24.426 48.9725 ;
               RECT 24.374 49.182 24.426 49.218 ;
               RECT 24.374 49.902 24.426 49.938 ;
               RECT 24.374 50.622 24.426 50.658 ;
               RECT 24.374 50.862 24.426 50.898 ;
               RECT 24.374 51.342 24.426 51.378 ;
               RECT 24.374 51.822 24.426 51.858 ;
               RECT 24.374 52.302 24.426 52.338 ;
               RECT 24.374 52.782 24.426 52.818 ;
               RECT 24.374 53.262 24.426 53.298 ;
               RECT 24.374 53.742 24.426 53.778 ;
               RECT 24.374 54.222 24.426 54.258 ;
               RECT 24.374 54.462 24.426 54.498 ;
               RECT 24.374 55.182 24.426 55.218 ;
               RECT 24.374 55.902 24.426 55.938 ;
               RECT 24.374 56.142 24.426 56.178 ;
               RECT 24.374 56.1475 24.426 56.1725 ;
               RECT 24.374 56.502 24.426 56.538 ;
               RECT 24.374 57.102 24.426 57.138 ;
               RECT 24.374 57.702 24.426 57.738 ;
               RECT 24.374 58.302 24.426 58.338 ;
               RECT 24.374 58.902 24.426 58.938 ;
               RECT 24.374 59.502 24.426 59.538 ;
               RECT 24.374 60.102 24.426 60.138 ;
               RECT 24.374 60.702 24.426 60.738 ;
               RECT 24.374 61.302 24.426 61.338 ;
               RECT 24.374 61.902 24.426 61.938 ;
               RECT 24.374 62.502 24.426 62.538 ;
               RECT 24.374 63.102 24.426 63.138 ;
               RECT 24.374 63.702 24.426 63.738 ;
               RECT 24.374 64.302 24.426 64.338 ;
               RECT 24.374 64.902 24.426 64.938 ;
               RECT 24.374 65.502 24.426 65.538 ;
               RECT 24.374 66.102 24.426 66.138 ;
               RECT 24.374 66.702 24.426 66.738 ;
               RECT 24.374 67.302 24.426 67.338 ;
               RECT 24.374 67.902 24.426 67.938 ;
               RECT 24.374 68.502 24.426 68.538 ;
               RECT 24.374 69.102 24.426 69.138 ;
               RECT 24.374 69.702 24.426 69.738 ;
               RECT 24.374 70.302 24.426 70.338 ;
               RECT 24.374 70.902 24.426 70.938 ;
               RECT 24.374 71.502 24.426 71.538 ;
               RECT 24.374 72.102 24.426 72.138 ;
               RECT 24.374 72.702 24.426 72.738 ;
               RECT 24.374 73.302 24.426 73.338 ;
               RECT 24.374 73.902 24.426 73.938 ;
               RECT 24.374 74.502 24.426 74.538 ;
               RECT 24.374 75.102 24.426 75.138 ;
               RECT 24.374 75.702 24.426 75.738 ;
               RECT 24.374 76.302 24.426 76.338 ;
               RECT 24.374 76.902 24.426 76.938 ;
               RECT 24.374 77.502 24.426 77.538 ;
               RECT 24.374 78.102 24.426 78.138 ;
               RECT 24.374 78.702 24.426 78.738 ;
               RECT 24.374 79.302 24.426 79.338 ;
               RECT 24.374 79.902 24.426 79.938 ;
               RECT 24.374 80.502 24.426 80.538 ;
               RECT 24.374 81.102 24.426 81.138 ;
               RECT 24.374 81.702 24.426 81.738 ;
               RECT 24.374 82.302 24.426 82.338 ;
               RECT 24.374 82.902 24.426 82.938 ;
               RECT 24.374 83.502 24.426 83.538 ;
               RECT 24.374 84.102 24.426 84.138 ;
               RECT 24.374 84.702 24.426 84.738 ;
               RECT 24.374 85.302 24.426 85.338 ;
               RECT 24.374 85.902 24.426 85.938 ;
               RECT 24.374 86.502 24.426 86.538 ;
               RECT 24.374 87.102 24.426 87.138 ;
               RECT 24.374 87.702 24.426 87.738 ;
               RECT 24.374 88.302 24.426 88.338 ;
               RECT 24.374 88.902 24.426 88.938 ;
               RECT 24.374 89.502 24.426 89.538 ;
               RECT 24.374 90.102 24.426 90.138 ;
               RECT 24.374 90.702 24.426 90.738 ;
               RECT 24.374 91.302 24.426 91.338 ;
               RECT 24.374 91.902 24.426 91.938 ;
               RECT 24.374 92.502 24.426 92.538 ;
               RECT 24.374 93.102 24.426 93.138 ;
               RECT 24.374 93.702 24.426 93.738 ;
               RECT 24.374 94.302 24.426 94.338 ;
               RECT 24.374 94.902 24.426 94.938 ;
               RECT 24.374 95.502 24.426 95.538 ;
               RECT 24.374 96.102 24.426 96.138 ;
               RECT 24.374 96.702 24.426 96.738 ;
               RECT 24.374 97.302 24.426 97.338 ;
               RECT 24.374 97.902 24.426 97.938 ;
               RECT 24.374 98.502 24.426 98.538 ;
               RECT 24.374 99.102 24.426 99.138 ;
               RECT 24.374 99.702 24.426 99.738 ;
               RECT 24.374 100.302 24.426 100.338 ;
               RECT 24.374 100.902 24.426 100.938 ;
               RECT 24.374 101.502 24.426 101.538 ;
               RECT 24.374 102.102 24.426 102.138 ;
               RECT 24.374 102.702 24.426 102.738 ;
               RECT 24.374 103.302 24.426 103.338 ;
               RECT 24.374 103.902 24.426 103.938 ;
               RECT 24.374 104.502 24.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 25.174 0.5695 25.226 104.5505 ;
               LAYER v4 ;
               RECT 25.174 0.582 25.226 0.618 ;
               RECT 25.174 1.182 25.226 1.218 ;
               RECT 25.174 1.782 25.226 1.818 ;
               RECT 25.174 2.382 25.226 2.418 ;
               RECT 25.174 2.982 25.226 3.018 ;
               RECT 25.174 3.582 25.226 3.618 ;
               RECT 25.174 4.182 25.226 4.218 ;
               RECT 25.174 4.782 25.226 4.818 ;
               RECT 25.174 5.382 25.226 5.418 ;
               RECT 25.174 5.982 25.226 6.018 ;
               RECT 25.174 6.582 25.226 6.618 ;
               RECT 25.174 7.182 25.226 7.218 ;
               RECT 25.174 7.782 25.226 7.818 ;
               RECT 25.174 8.382 25.226 8.418 ;
               RECT 25.174 8.982 25.226 9.018 ;
               RECT 25.174 9.582 25.226 9.618 ;
               RECT 25.174 10.182 25.226 10.218 ;
               RECT 25.174 10.782 25.226 10.818 ;
               RECT 25.174 11.382 25.226 11.418 ;
               RECT 25.174 11.982 25.226 12.018 ;
               RECT 25.174 12.582 25.226 12.618 ;
               RECT 25.174 13.182 25.226 13.218 ;
               RECT 25.174 13.782 25.226 13.818 ;
               RECT 25.174 14.382 25.226 14.418 ;
               RECT 25.174 14.982 25.226 15.018 ;
               RECT 25.174 15.582 25.226 15.618 ;
               RECT 25.174 16.182 25.226 16.218 ;
               RECT 25.174 16.782 25.226 16.818 ;
               RECT 25.174 17.382 25.226 17.418 ;
               RECT 25.174 17.982 25.226 18.018 ;
               RECT 25.174 18.582 25.226 18.618 ;
               RECT 25.174 19.182 25.226 19.218 ;
               RECT 25.174 19.782 25.226 19.818 ;
               RECT 25.174 20.382 25.226 20.418 ;
               RECT 25.174 20.982 25.226 21.018 ;
               RECT 25.174 21.582 25.226 21.618 ;
               RECT 25.174 22.182 25.226 22.218 ;
               RECT 25.174 22.782 25.226 22.818 ;
               RECT 25.174 23.382 25.226 23.418 ;
               RECT 25.174 23.982 25.226 24.018 ;
               RECT 25.174 24.582 25.226 24.618 ;
               RECT 25.174 25.182 25.226 25.218 ;
               RECT 25.174 25.782 25.226 25.818 ;
               RECT 25.174 26.382 25.226 26.418 ;
               RECT 25.174 26.982 25.226 27.018 ;
               RECT 25.174 27.582 25.226 27.618 ;
               RECT 25.174 28.182 25.226 28.218 ;
               RECT 25.174 28.782 25.226 28.818 ;
               RECT 25.174 29.382 25.226 29.418 ;
               RECT 25.174 29.982 25.226 30.018 ;
               RECT 25.174 30.582 25.226 30.618 ;
               RECT 25.174 31.182 25.226 31.218 ;
               RECT 25.174 31.782 25.226 31.818 ;
               RECT 25.174 32.382 25.226 32.418 ;
               RECT 25.174 32.982 25.226 33.018 ;
               RECT 25.174 33.582 25.226 33.618 ;
               RECT 25.174 34.182 25.226 34.218 ;
               RECT 25.174 34.782 25.226 34.818 ;
               RECT 25.174 35.382 25.226 35.418 ;
               RECT 25.174 35.982 25.226 36.018 ;
               RECT 25.174 36.582 25.226 36.618 ;
               RECT 25.174 37.182 25.226 37.218 ;
               RECT 25.174 37.782 25.226 37.818 ;
               RECT 25.174 38.382 25.226 38.418 ;
               RECT 25.174 38.982 25.226 39.018 ;
               RECT 25.174 39.582 25.226 39.618 ;
               RECT 25.174 40.182 25.226 40.218 ;
               RECT 25.174 40.782 25.226 40.818 ;
               RECT 25.174 41.382 25.226 41.418 ;
               RECT 25.174 41.982 25.226 42.018 ;
               RECT 25.174 42.582 25.226 42.618 ;
               RECT 25.174 43.182 25.226 43.218 ;
               RECT 25.174 43.782 25.226 43.818 ;
               RECT 25.174 44.382 25.226 44.418 ;
               RECT 25.174 44.982 25.226 45.018 ;
               RECT 25.174 45.582 25.226 45.618 ;
               RECT 25.174 46.182 25.226 46.218 ;
               RECT 25.174 46.782 25.226 46.818 ;
               RECT 25.174 47.382 25.226 47.418 ;
               RECT 25.174 47.982 25.226 48.018 ;
               RECT 25.174 48.582 25.226 48.618 ;
               RECT 25.174 48.942 25.226 48.978 ;
               RECT 25.174 49.182 25.226 49.218 ;
               RECT 25.174 49.902 25.226 49.938 ;
               RECT 25.174 50.622 25.226 50.658 ;
               RECT 25.174 50.862 25.226 50.898 ;
               RECT 25.174 51.342 25.226 51.378 ;
               RECT 25.174 51.822 25.226 51.858 ;
               RECT 25.174 52.302 25.226 52.338 ;
               RECT 25.174 52.782 25.226 52.818 ;
               RECT 25.174 53.262 25.226 53.298 ;
               RECT 25.174 53.742 25.226 53.778 ;
               RECT 25.174 54.222 25.226 54.258 ;
               RECT 25.174 54.462 25.226 54.498 ;
               RECT 25.174 55.182 25.226 55.218 ;
               RECT 25.174 55.902 25.226 55.938 ;
               RECT 25.174 56.142 25.226 56.178 ;
               RECT 25.174 56.502 25.226 56.538 ;
               RECT 25.174 57.102 25.226 57.138 ;
               RECT 25.174 57.702 25.226 57.738 ;
               RECT 25.174 58.302 25.226 58.338 ;
               RECT 25.174 58.902 25.226 58.938 ;
               RECT 25.174 59.502 25.226 59.538 ;
               RECT 25.174 60.102 25.226 60.138 ;
               RECT 25.174 60.702 25.226 60.738 ;
               RECT 25.174 61.302 25.226 61.338 ;
               RECT 25.174 61.902 25.226 61.938 ;
               RECT 25.174 62.502 25.226 62.538 ;
               RECT 25.174 63.102 25.226 63.138 ;
               RECT 25.174 63.702 25.226 63.738 ;
               RECT 25.174 64.302 25.226 64.338 ;
               RECT 25.174 64.902 25.226 64.938 ;
               RECT 25.174 65.502 25.226 65.538 ;
               RECT 25.174 66.102 25.226 66.138 ;
               RECT 25.174 66.702 25.226 66.738 ;
               RECT 25.174 67.302 25.226 67.338 ;
               RECT 25.174 67.902 25.226 67.938 ;
               RECT 25.174 68.502 25.226 68.538 ;
               RECT 25.174 69.102 25.226 69.138 ;
               RECT 25.174 69.702 25.226 69.738 ;
               RECT 25.174 70.302 25.226 70.338 ;
               RECT 25.174 70.902 25.226 70.938 ;
               RECT 25.174 71.502 25.226 71.538 ;
               RECT 25.174 72.102 25.226 72.138 ;
               RECT 25.174 72.702 25.226 72.738 ;
               RECT 25.174 73.302 25.226 73.338 ;
               RECT 25.174 73.902 25.226 73.938 ;
               RECT 25.174 74.502 25.226 74.538 ;
               RECT 25.174 75.102 25.226 75.138 ;
               RECT 25.174 75.702 25.226 75.738 ;
               RECT 25.174 76.302 25.226 76.338 ;
               RECT 25.174 76.902 25.226 76.938 ;
               RECT 25.174 77.502 25.226 77.538 ;
               RECT 25.174 78.102 25.226 78.138 ;
               RECT 25.174 78.702 25.226 78.738 ;
               RECT 25.174 79.302 25.226 79.338 ;
               RECT 25.174 79.902 25.226 79.938 ;
               RECT 25.174 80.502 25.226 80.538 ;
               RECT 25.174 81.102 25.226 81.138 ;
               RECT 25.174 81.702 25.226 81.738 ;
               RECT 25.174 82.302 25.226 82.338 ;
               RECT 25.174 82.902 25.226 82.938 ;
               RECT 25.174 83.502 25.226 83.538 ;
               RECT 25.174 84.102 25.226 84.138 ;
               RECT 25.174 84.702 25.226 84.738 ;
               RECT 25.174 85.302 25.226 85.338 ;
               RECT 25.174 85.902 25.226 85.938 ;
               RECT 25.174 86.502 25.226 86.538 ;
               RECT 25.174 87.102 25.226 87.138 ;
               RECT 25.174 87.702 25.226 87.738 ;
               RECT 25.174 88.302 25.226 88.338 ;
               RECT 25.174 88.902 25.226 88.938 ;
               RECT 25.174 89.502 25.226 89.538 ;
               RECT 25.174 90.102 25.226 90.138 ;
               RECT 25.174 90.702 25.226 90.738 ;
               RECT 25.174 91.302 25.226 91.338 ;
               RECT 25.174 91.902 25.226 91.938 ;
               RECT 25.174 92.502 25.226 92.538 ;
               RECT 25.174 93.102 25.226 93.138 ;
               RECT 25.174 93.702 25.226 93.738 ;
               RECT 25.174 94.302 25.226 94.338 ;
               RECT 25.174 94.902 25.226 94.938 ;
               RECT 25.174 95.502 25.226 95.538 ;
               RECT 25.174 96.102 25.226 96.138 ;
               RECT 25.174 96.702 25.226 96.738 ;
               RECT 25.174 97.302 25.226 97.338 ;
               RECT 25.174 97.902 25.226 97.938 ;
               RECT 25.174 98.502 25.226 98.538 ;
               RECT 25.174 99.102 25.226 99.138 ;
               RECT 25.174 99.702 25.226 99.738 ;
               RECT 25.174 100.302 25.226 100.338 ;
               RECT 25.174 100.902 25.226 100.938 ;
               RECT 25.174 101.502 25.226 101.538 ;
               RECT 25.174 102.102 25.226 102.138 ;
               RECT 25.174 102.702 25.226 102.738 ;
               RECT 25.174 103.302 25.226 103.338 ;
               RECT 25.174 103.902 25.226 103.938 ;
               RECT 25.174 104.502 25.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 25.974 0.5695 26.026 104.5505 ;
               LAYER v4 ;
               RECT 25.974 0.582 26.026 0.618 ;
               RECT 25.974 1.182 26.026 1.218 ;
               RECT 25.974 1.782 26.026 1.818 ;
               RECT 25.974 2.382 26.026 2.418 ;
               RECT 25.974 2.982 26.026 3.018 ;
               RECT 25.974 3.582 26.026 3.618 ;
               RECT 25.974 4.182 26.026 4.218 ;
               RECT 25.974 4.782 26.026 4.818 ;
               RECT 25.974 5.382 26.026 5.418 ;
               RECT 25.974 5.982 26.026 6.018 ;
               RECT 25.974 6.582 26.026 6.618 ;
               RECT 25.974 7.182 26.026 7.218 ;
               RECT 25.974 7.782 26.026 7.818 ;
               RECT 25.974 8.382 26.026 8.418 ;
               RECT 25.974 8.982 26.026 9.018 ;
               RECT 25.974 9.582 26.026 9.618 ;
               RECT 25.974 10.182 26.026 10.218 ;
               RECT 25.974 10.782 26.026 10.818 ;
               RECT 25.974 11.382 26.026 11.418 ;
               RECT 25.974 11.982 26.026 12.018 ;
               RECT 25.974 12.582 26.026 12.618 ;
               RECT 25.974 13.182 26.026 13.218 ;
               RECT 25.974 13.782 26.026 13.818 ;
               RECT 25.974 14.382 26.026 14.418 ;
               RECT 25.974 14.982 26.026 15.018 ;
               RECT 25.974 15.582 26.026 15.618 ;
               RECT 25.974 16.182 26.026 16.218 ;
               RECT 25.974 16.782 26.026 16.818 ;
               RECT 25.974 17.382 26.026 17.418 ;
               RECT 25.974 17.982 26.026 18.018 ;
               RECT 25.974 18.582 26.026 18.618 ;
               RECT 25.974 19.182 26.026 19.218 ;
               RECT 25.974 19.782 26.026 19.818 ;
               RECT 25.974 20.382 26.026 20.418 ;
               RECT 25.974 20.982 26.026 21.018 ;
               RECT 25.974 21.582 26.026 21.618 ;
               RECT 25.974 22.182 26.026 22.218 ;
               RECT 25.974 22.782 26.026 22.818 ;
               RECT 25.974 23.382 26.026 23.418 ;
               RECT 25.974 23.982 26.026 24.018 ;
               RECT 25.974 24.582 26.026 24.618 ;
               RECT 25.974 25.182 26.026 25.218 ;
               RECT 25.974 25.782 26.026 25.818 ;
               RECT 25.974 26.382 26.026 26.418 ;
               RECT 25.974 26.982 26.026 27.018 ;
               RECT 25.974 27.582 26.026 27.618 ;
               RECT 25.974 28.182 26.026 28.218 ;
               RECT 25.974 28.782 26.026 28.818 ;
               RECT 25.974 29.382 26.026 29.418 ;
               RECT 25.974 29.982 26.026 30.018 ;
               RECT 25.974 30.582 26.026 30.618 ;
               RECT 25.974 31.182 26.026 31.218 ;
               RECT 25.974 31.782 26.026 31.818 ;
               RECT 25.974 32.382 26.026 32.418 ;
               RECT 25.974 32.982 26.026 33.018 ;
               RECT 25.974 33.582 26.026 33.618 ;
               RECT 25.974 34.182 26.026 34.218 ;
               RECT 25.974 34.782 26.026 34.818 ;
               RECT 25.974 35.382 26.026 35.418 ;
               RECT 25.974 35.982 26.026 36.018 ;
               RECT 25.974 36.582 26.026 36.618 ;
               RECT 25.974 37.182 26.026 37.218 ;
               RECT 25.974 37.782 26.026 37.818 ;
               RECT 25.974 38.382 26.026 38.418 ;
               RECT 25.974 38.982 26.026 39.018 ;
               RECT 25.974 39.582 26.026 39.618 ;
               RECT 25.974 40.182 26.026 40.218 ;
               RECT 25.974 40.782 26.026 40.818 ;
               RECT 25.974 41.382 26.026 41.418 ;
               RECT 25.974 41.982 26.026 42.018 ;
               RECT 25.974 42.582 26.026 42.618 ;
               RECT 25.974 43.182 26.026 43.218 ;
               RECT 25.974 43.782 26.026 43.818 ;
               RECT 25.974 44.382 26.026 44.418 ;
               RECT 25.974 44.982 26.026 45.018 ;
               RECT 25.974 45.582 26.026 45.618 ;
               RECT 25.974 46.182 26.026 46.218 ;
               RECT 25.974 46.782 26.026 46.818 ;
               RECT 25.974 47.382 26.026 47.418 ;
               RECT 25.974 47.982 26.026 48.018 ;
               RECT 25.974 48.582 26.026 48.618 ;
               RECT 25.974 48.942 26.026 48.978 ;
               RECT 25.974 48.9475 26.026 48.9725 ;
               RECT 25.974 49.182 26.026 49.218 ;
               RECT 25.974 49.902 26.026 49.938 ;
               RECT 25.974 50.622 26.026 50.658 ;
               RECT 25.974 50.862 26.026 50.898 ;
               RECT 25.974 51.342 26.026 51.378 ;
               RECT 25.974 51.822 26.026 51.858 ;
               RECT 25.974 52.302 26.026 52.338 ;
               RECT 25.974 52.782 26.026 52.818 ;
               RECT 25.974 53.262 26.026 53.298 ;
               RECT 25.974 53.742 26.026 53.778 ;
               RECT 25.974 54.222 26.026 54.258 ;
               RECT 25.974 54.462 26.026 54.498 ;
               RECT 25.974 55.182 26.026 55.218 ;
               RECT 25.974 55.902 26.026 55.938 ;
               RECT 25.974 56.142 26.026 56.178 ;
               RECT 25.974 56.1475 26.026 56.1725 ;
               RECT 25.974 56.502 26.026 56.538 ;
               RECT 25.974 57.102 26.026 57.138 ;
               RECT 25.974 57.702 26.026 57.738 ;
               RECT 25.974 58.302 26.026 58.338 ;
               RECT 25.974 58.902 26.026 58.938 ;
               RECT 25.974 59.502 26.026 59.538 ;
               RECT 25.974 60.102 26.026 60.138 ;
               RECT 25.974 60.702 26.026 60.738 ;
               RECT 25.974 61.302 26.026 61.338 ;
               RECT 25.974 61.902 26.026 61.938 ;
               RECT 25.974 62.502 26.026 62.538 ;
               RECT 25.974 63.102 26.026 63.138 ;
               RECT 25.974 63.702 26.026 63.738 ;
               RECT 25.974 64.302 26.026 64.338 ;
               RECT 25.974 64.902 26.026 64.938 ;
               RECT 25.974 65.502 26.026 65.538 ;
               RECT 25.974 66.102 26.026 66.138 ;
               RECT 25.974 66.702 26.026 66.738 ;
               RECT 25.974 67.302 26.026 67.338 ;
               RECT 25.974 67.902 26.026 67.938 ;
               RECT 25.974 68.502 26.026 68.538 ;
               RECT 25.974 69.102 26.026 69.138 ;
               RECT 25.974 69.702 26.026 69.738 ;
               RECT 25.974 70.302 26.026 70.338 ;
               RECT 25.974 70.902 26.026 70.938 ;
               RECT 25.974 71.502 26.026 71.538 ;
               RECT 25.974 72.102 26.026 72.138 ;
               RECT 25.974 72.702 26.026 72.738 ;
               RECT 25.974 73.302 26.026 73.338 ;
               RECT 25.974 73.902 26.026 73.938 ;
               RECT 25.974 74.502 26.026 74.538 ;
               RECT 25.974 75.102 26.026 75.138 ;
               RECT 25.974 75.702 26.026 75.738 ;
               RECT 25.974 76.302 26.026 76.338 ;
               RECT 25.974 76.902 26.026 76.938 ;
               RECT 25.974 77.502 26.026 77.538 ;
               RECT 25.974 78.102 26.026 78.138 ;
               RECT 25.974 78.702 26.026 78.738 ;
               RECT 25.974 79.302 26.026 79.338 ;
               RECT 25.974 79.902 26.026 79.938 ;
               RECT 25.974 80.502 26.026 80.538 ;
               RECT 25.974 81.102 26.026 81.138 ;
               RECT 25.974 81.702 26.026 81.738 ;
               RECT 25.974 82.302 26.026 82.338 ;
               RECT 25.974 82.902 26.026 82.938 ;
               RECT 25.974 83.502 26.026 83.538 ;
               RECT 25.974 84.102 26.026 84.138 ;
               RECT 25.974 84.702 26.026 84.738 ;
               RECT 25.974 85.302 26.026 85.338 ;
               RECT 25.974 85.902 26.026 85.938 ;
               RECT 25.974 86.502 26.026 86.538 ;
               RECT 25.974 87.102 26.026 87.138 ;
               RECT 25.974 87.702 26.026 87.738 ;
               RECT 25.974 88.302 26.026 88.338 ;
               RECT 25.974 88.902 26.026 88.938 ;
               RECT 25.974 89.502 26.026 89.538 ;
               RECT 25.974 90.102 26.026 90.138 ;
               RECT 25.974 90.702 26.026 90.738 ;
               RECT 25.974 91.302 26.026 91.338 ;
               RECT 25.974 91.902 26.026 91.938 ;
               RECT 25.974 92.502 26.026 92.538 ;
               RECT 25.974 93.102 26.026 93.138 ;
               RECT 25.974 93.702 26.026 93.738 ;
               RECT 25.974 94.302 26.026 94.338 ;
               RECT 25.974 94.902 26.026 94.938 ;
               RECT 25.974 95.502 26.026 95.538 ;
               RECT 25.974 96.102 26.026 96.138 ;
               RECT 25.974 96.702 26.026 96.738 ;
               RECT 25.974 97.302 26.026 97.338 ;
               RECT 25.974 97.902 26.026 97.938 ;
               RECT 25.974 98.502 26.026 98.538 ;
               RECT 25.974 99.102 26.026 99.138 ;
               RECT 25.974 99.702 26.026 99.738 ;
               RECT 25.974 100.302 26.026 100.338 ;
               RECT 25.974 100.902 26.026 100.938 ;
               RECT 25.974 101.502 26.026 101.538 ;
               RECT 25.974 102.102 26.026 102.138 ;
               RECT 25.974 102.702 26.026 102.738 ;
               RECT 25.974 103.302 26.026 103.338 ;
               RECT 25.974 103.902 26.026 103.938 ;
               RECT 25.974 104.502 26.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 26.774 0.5695 26.826 104.5505 ;
               LAYER v4 ;
               RECT 26.774 0.582 26.826 0.618 ;
               RECT 26.774 1.182 26.826 1.218 ;
               RECT 26.774 1.782 26.826 1.818 ;
               RECT 26.774 2.382 26.826 2.418 ;
               RECT 26.774 2.982 26.826 3.018 ;
               RECT 26.774 3.582 26.826 3.618 ;
               RECT 26.774 4.182 26.826 4.218 ;
               RECT 26.774 4.782 26.826 4.818 ;
               RECT 26.774 5.382 26.826 5.418 ;
               RECT 26.774 5.982 26.826 6.018 ;
               RECT 26.774 6.582 26.826 6.618 ;
               RECT 26.774 7.182 26.826 7.218 ;
               RECT 26.774 7.782 26.826 7.818 ;
               RECT 26.774 8.382 26.826 8.418 ;
               RECT 26.774 8.982 26.826 9.018 ;
               RECT 26.774 9.582 26.826 9.618 ;
               RECT 26.774 10.182 26.826 10.218 ;
               RECT 26.774 10.782 26.826 10.818 ;
               RECT 26.774 11.382 26.826 11.418 ;
               RECT 26.774 11.982 26.826 12.018 ;
               RECT 26.774 12.582 26.826 12.618 ;
               RECT 26.774 13.182 26.826 13.218 ;
               RECT 26.774 13.782 26.826 13.818 ;
               RECT 26.774 14.382 26.826 14.418 ;
               RECT 26.774 14.982 26.826 15.018 ;
               RECT 26.774 15.582 26.826 15.618 ;
               RECT 26.774 16.182 26.826 16.218 ;
               RECT 26.774 16.782 26.826 16.818 ;
               RECT 26.774 17.382 26.826 17.418 ;
               RECT 26.774 17.982 26.826 18.018 ;
               RECT 26.774 18.582 26.826 18.618 ;
               RECT 26.774 19.182 26.826 19.218 ;
               RECT 26.774 19.782 26.826 19.818 ;
               RECT 26.774 20.382 26.826 20.418 ;
               RECT 26.774 20.982 26.826 21.018 ;
               RECT 26.774 21.582 26.826 21.618 ;
               RECT 26.774 22.182 26.826 22.218 ;
               RECT 26.774 22.782 26.826 22.818 ;
               RECT 26.774 23.382 26.826 23.418 ;
               RECT 26.774 23.982 26.826 24.018 ;
               RECT 26.774 24.582 26.826 24.618 ;
               RECT 26.774 25.182 26.826 25.218 ;
               RECT 26.774 25.782 26.826 25.818 ;
               RECT 26.774 26.382 26.826 26.418 ;
               RECT 26.774 26.982 26.826 27.018 ;
               RECT 26.774 27.582 26.826 27.618 ;
               RECT 26.774 28.182 26.826 28.218 ;
               RECT 26.774 28.782 26.826 28.818 ;
               RECT 26.774 29.382 26.826 29.418 ;
               RECT 26.774 29.982 26.826 30.018 ;
               RECT 26.774 30.582 26.826 30.618 ;
               RECT 26.774 31.182 26.826 31.218 ;
               RECT 26.774 31.782 26.826 31.818 ;
               RECT 26.774 32.382 26.826 32.418 ;
               RECT 26.774 32.982 26.826 33.018 ;
               RECT 26.774 33.582 26.826 33.618 ;
               RECT 26.774 34.182 26.826 34.218 ;
               RECT 26.774 34.782 26.826 34.818 ;
               RECT 26.774 35.382 26.826 35.418 ;
               RECT 26.774 35.982 26.826 36.018 ;
               RECT 26.774 36.582 26.826 36.618 ;
               RECT 26.774 37.182 26.826 37.218 ;
               RECT 26.774 37.782 26.826 37.818 ;
               RECT 26.774 38.382 26.826 38.418 ;
               RECT 26.774 38.982 26.826 39.018 ;
               RECT 26.774 39.582 26.826 39.618 ;
               RECT 26.774 40.182 26.826 40.218 ;
               RECT 26.774 40.782 26.826 40.818 ;
               RECT 26.774 41.382 26.826 41.418 ;
               RECT 26.774 41.982 26.826 42.018 ;
               RECT 26.774 42.582 26.826 42.618 ;
               RECT 26.774 43.182 26.826 43.218 ;
               RECT 26.774 43.782 26.826 43.818 ;
               RECT 26.774 44.382 26.826 44.418 ;
               RECT 26.774 44.982 26.826 45.018 ;
               RECT 26.774 45.582 26.826 45.618 ;
               RECT 26.774 46.182 26.826 46.218 ;
               RECT 26.774 46.782 26.826 46.818 ;
               RECT 26.774 47.382 26.826 47.418 ;
               RECT 26.774 47.982 26.826 48.018 ;
               RECT 26.774 48.582 26.826 48.618 ;
               RECT 26.774 48.942 26.826 48.978 ;
               RECT 26.774 49.182 26.826 49.218 ;
               RECT 26.774 49.902 26.826 49.938 ;
               RECT 26.774 50.622 26.826 50.658 ;
               RECT 26.774 50.862 26.826 50.898 ;
               RECT 26.774 51.342 26.826 51.378 ;
               RECT 26.774 51.822 26.826 51.858 ;
               RECT 26.774 52.302 26.826 52.338 ;
               RECT 26.774 52.782 26.826 52.818 ;
               RECT 26.774 53.262 26.826 53.298 ;
               RECT 26.774 53.742 26.826 53.778 ;
               RECT 26.774 54.222 26.826 54.258 ;
               RECT 26.774 54.462 26.826 54.498 ;
               RECT 26.774 55.182 26.826 55.218 ;
               RECT 26.774 55.902 26.826 55.938 ;
               RECT 26.774 56.142 26.826 56.178 ;
               RECT 26.774 56.502 26.826 56.538 ;
               RECT 26.774 57.102 26.826 57.138 ;
               RECT 26.774 57.702 26.826 57.738 ;
               RECT 26.774 58.302 26.826 58.338 ;
               RECT 26.774 58.902 26.826 58.938 ;
               RECT 26.774 59.502 26.826 59.538 ;
               RECT 26.774 60.102 26.826 60.138 ;
               RECT 26.774 60.702 26.826 60.738 ;
               RECT 26.774 61.302 26.826 61.338 ;
               RECT 26.774 61.902 26.826 61.938 ;
               RECT 26.774 62.502 26.826 62.538 ;
               RECT 26.774 63.102 26.826 63.138 ;
               RECT 26.774 63.702 26.826 63.738 ;
               RECT 26.774 64.302 26.826 64.338 ;
               RECT 26.774 64.902 26.826 64.938 ;
               RECT 26.774 65.502 26.826 65.538 ;
               RECT 26.774 66.102 26.826 66.138 ;
               RECT 26.774 66.702 26.826 66.738 ;
               RECT 26.774 67.302 26.826 67.338 ;
               RECT 26.774 67.902 26.826 67.938 ;
               RECT 26.774 68.502 26.826 68.538 ;
               RECT 26.774 69.102 26.826 69.138 ;
               RECT 26.774 69.702 26.826 69.738 ;
               RECT 26.774 70.302 26.826 70.338 ;
               RECT 26.774 70.902 26.826 70.938 ;
               RECT 26.774 71.502 26.826 71.538 ;
               RECT 26.774 72.102 26.826 72.138 ;
               RECT 26.774 72.702 26.826 72.738 ;
               RECT 26.774 73.302 26.826 73.338 ;
               RECT 26.774 73.902 26.826 73.938 ;
               RECT 26.774 74.502 26.826 74.538 ;
               RECT 26.774 75.102 26.826 75.138 ;
               RECT 26.774 75.702 26.826 75.738 ;
               RECT 26.774 76.302 26.826 76.338 ;
               RECT 26.774 76.902 26.826 76.938 ;
               RECT 26.774 77.502 26.826 77.538 ;
               RECT 26.774 78.102 26.826 78.138 ;
               RECT 26.774 78.702 26.826 78.738 ;
               RECT 26.774 79.302 26.826 79.338 ;
               RECT 26.774 79.902 26.826 79.938 ;
               RECT 26.774 80.502 26.826 80.538 ;
               RECT 26.774 81.102 26.826 81.138 ;
               RECT 26.774 81.702 26.826 81.738 ;
               RECT 26.774 82.302 26.826 82.338 ;
               RECT 26.774 82.902 26.826 82.938 ;
               RECT 26.774 83.502 26.826 83.538 ;
               RECT 26.774 84.102 26.826 84.138 ;
               RECT 26.774 84.702 26.826 84.738 ;
               RECT 26.774 85.302 26.826 85.338 ;
               RECT 26.774 85.902 26.826 85.938 ;
               RECT 26.774 86.502 26.826 86.538 ;
               RECT 26.774 87.102 26.826 87.138 ;
               RECT 26.774 87.702 26.826 87.738 ;
               RECT 26.774 88.302 26.826 88.338 ;
               RECT 26.774 88.902 26.826 88.938 ;
               RECT 26.774 89.502 26.826 89.538 ;
               RECT 26.774 90.102 26.826 90.138 ;
               RECT 26.774 90.702 26.826 90.738 ;
               RECT 26.774 91.302 26.826 91.338 ;
               RECT 26.774 91.902 26.826 91.938 ;
               RECT 26.774 92.502 26.826 92.538 ;
               RECT 26.774 93.102 26.826 93.138 ;
               RECT 26.774 93.702 26.826 93.738 ;
               RECT 26.774 94.302 26.826 94.338 ;
               RECT 26.774 94.902 26.826 94.938 ;
               RECT 26.774 95.502 26.826 95.538 ;
               RECT 26.774 96.102 26.826 96.138 ;
               RECT 26.774 96.702 26.826 96.738 ;
               RECT 26.774 97.302 26.826 97.338 ;
               RECT 26.774 97.902 26.826 97.938 ;
               RECT 26.774 98.502 26.826 98.538 ;
               RECT 26.774 99.102 26.826 99.138 ;
               RECT 26.774 99.702 26.826 99.738 ;
               RECT 26.774 100.302 26.826 100.338 ;
               RECT 26.774 100.902 26.826 100.938 ;
               RECT 26.774 101.502 26.826 101.538 ;
               RECT 26.774 102.102 26.826 102.138 ;
               RECT 26.774 102.702 26.826 102.738 ;
               RECT 26.774 103.302 26.826 103.338 ;
               RECT 26.774 103.902 26.826 103.938 ;
               RECT 26.774 104.502 26.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 27.574 0.5695 27.626 104.5505 ;
               LAYER v4 ;
               RECT 27.574 0.582 27.626 0.618 ;
               RECT 27.574 1.182 27.626 1.218 ;
               RECT 27.574 1.782 27.626 1.818 ;
               RECT 27.574 2.382 27.626 2.418 ;
               RECT 27.574 2.982 27.626 3.018 ;
               RECT 27.574 3.582 27.626 3.618 ;
               RECT 27.574 4.182 27.626 4.218 ;
               RECT 27.574 4.782 27.626 4.818 ;
               RECT 27.574 5.382 27.626 5.418 ;
               RECT 27.574 5.982 27.626 6.018 ;
               RECT 27.574 6.582 27.626 6.618 ;
               RECT 27.574 7.182 27.626 7.218 ;
               RECT 27.574 7.782 27.626 7.818 ;
               RECT 27.574 8.382 27.626 8.418 ;
               RECT 27.574 8.982 27.626 9.018 ;
               RECT 27.574 9.582 27.626 9.618 ;
               RECT 27.574 10.182 27.626 10.218 ;
               RECT 27.574 10.782 27.626 10.818 ;
               RECT 27.574 11.382 27.626 11.418 ;
               RECT 27.574 11.982 27.626 12.018 ;
               RECT 27.574 12.582 27.626 12.618 ;
               RECT 27.574 13.182 27.626 13.218 ;
               RECT 27.574 13.782 27.626 13.818 ;
               RECT 27.574 14.382 27.626 14.418 ;
               RECT 27.574 14.982 27.626 15.018 ;
               RECT 27.574 15.582 27.626 15.618 ;
               RECT 27.574 16.182 27.626 16.218 ;
               RECT 27.574 16.782 27.626 16.818 ;
               RECT 27.574 17.382 27.626 17.418 ;
               RECT 27.574 17.982 27.626 18.018 ;
               RECT 27.574 18.582 27.626 18.618 ;
               RECT 27.574 19.182 27.626 19.218 ;
               RECT 27.574 19.782 27.626 19.818 ;
               RECT 27.574 20.382 27.626 20.418 ;
               RECT 27.574 20.982 27.626 21.018 ;
               RECT 27.574 21.582 27.626 21.618 ;
               RECT 27.574 22.182 27.626 22.218 ;
               RECT 27.574 22.782 27.626 22.818 ;
               RECT 27.574 23.382 27.626 23.418 ;
               RECT 27.574 23.982 27.626 24.018 ;
               RECT 27.574 24.582 27.626 24.618 ;
               RECT 27.574 25.182 27.626 25.218 ;
               RECT 27.574 25.782 27.626 25.818 ;
               RECT 27.574 26.382 27.626 26.418 ;
               RECT 27.574 26.982 27.626 27.018 ;
               RECT 27.574 27.582 27.626 27.618 ;
               RECT 27.574 28.182 27.626 28.218 ;
               RECT 27.574 28.782 27.626 28.818 ;
               RECT 27.574 29.382 27.626 29.418 ;
               RECT 27.574 29.982 27.626 30.018 ;
               RECT 27.574 30.582 27.626 30.618 ;
               RECT 27.574 31.182 27.626 31.218 ;
               RECT 27.574 31.782 27.626 31.818 ;
               RECT 27.574 32.382 27.626 32.418 ;
               RECT 27.574 32.982 27.626 33.018 ;
               RECT 27.574 33.582 27.626 33.618 ;
               RECT 27.574 34.182 27.626 34.218 ;
               RECT 27.574 34.782 27.626 34.818 ;
               RECT 27.574 35.382 27.626 35.418 ;
               RECT 27.574 35.982 27.626 36.018 ;
               RECT 27.574 36.582 27.626 36.618 ;
               RECT 27.574 37.182 27.626 37.218 ;
               RECT 27.574 37.782 27.626 37.818 ;
               RECT 27.574 38.382 27.626 38.418 ;
               RECT 27.574 38.982 27.626 39.018 ;
               RECT 27.574 39.582 27.626 39.618 ;
               RECT 27.574 40.182 27.626 40.218 ;
               RECT 27.574 40.782 27.626 40.818 ;
               RECT 27.574 41.382 27.626 41.418 ;
               RECT 27.574 41.982 27.626 42.018 ;
               RECT 27.574 42.582 27.626 42.618 ;
               RECT 27.574 43.182 27.626 43.218 ;
               RECT 27.574 43.782 27.626 43.818 ;
               RECT 27.574 44.382 27.626 44.418 ;
               RECT 27.574 44.982 27.626 45.018 ;
               RECT 27.574 45.582 27.626 45.618 ;
               RECT 27.574 46.182 27.626 46.218 ;
               RECT 27.574 46.782 27.626 46.818 ;
               RECT 27.574 47.382 27.626 47.418 ;
               RECT 27.574 47.982 27.626 48.018 ;
               RECT 27.574 48.582 27.626 48.618 ;
               RECT 27.574 48.942 27.626 48.978 ;
               RECT 27.574 48.9475 27.626 48.9725 ;
               RECT 27.574 49.182 27.626 49.218 ;
               RECT 27.574 49.902 27.626 49.938 ;
               RECT 27.574 50.622 27.626 50.658 ;
               RECT 27.574 50.862 27.626 50.898 ;
               RECT 27.574 51.342 27.626 51.378 ;
               RECT 27.574 51.822 27.626 51.858 ;
               RECT 27.574 52.302 27.626 52.338 ;
               RECT 27.574 52.782 27.626 52.818 ;
               RECT 27.574 53.262 27.626 53.298 ;
               RECT 27.574 53.742 27.626 53.778 ;
               RECT 27.574 54.222 27.626 54.258 ;
               RECT 27.574 54.462 27.626 54.498 ;
               RECT 27.574 55.182 27.626 55.218 ;
               RECT 27.574 55.902 27.626 55.938 ;
               RECT 27.574 56.142 27.626 56.178 ;
               RECT 27.574 56.1475 27.626 56.1725 ;
               RECT 27.574 56.502 27.626 56.538 ;
               RECT 27.574 57.102 27.626 57.138 ;
               RECT 27.574 57.702 27.626 57.738 ;
               RECT 27.574 58.302 27.626 58.338 ;
               RECT 27.574 58.902 27.626 58.938 ;
               RECT 27.574 59.502 27.626 59.538 ;
               RECT 27.574 60.102 27.626 60.138 ;
               RECT 27.574 60.702 27.626 60.738 ;
               RECT 27.574 61.302 27.626 61.338 ;
               RECT 27.574 61.902 27.626 61.938 ;
               RECT 27.574 62.502 27.626 62.538 ;
               RECT 27.574 63.102 27.626 63.138 ;
               RECT 27.574 63.702 27.626 63.738 ;
               RECT 27.574 64.302 27.626 64.338 ;
               RECT 27.574 64.902 27.626 64.938 ;
               RECT 27.574 65.502 27.626 65.538 ;
               RECT 27.574 66.102 27.626 66.138 ;
               RECT 27.574 66.702 27.626 66.738 ;
               RECT 27.574 67.302 27.626 67.338 ;
               RECT 27.574 67.902 27.626 67.938 ;
               RECT 27.574 68.502 27.626 68.538 ;
               RECT 27.574 69.102 27.626 69.138 ;
               RECT 27.574 69.702 27.626 69.738 ;
               RECT 27.574 70.302 27.626 70.338 ;
               RECT 27.574 70.902 27.626 70.938 ;
               RECT 27.574 71.502 27.626 71.538 ;
               RECT 27.574 72.102 27.626 72.138 ;
               RECT 27.574 72.702 27.626 72.738 ;
               RECT 27.574 73.302 27.626 73.338 ;
               RECT 27.574 73.902 27.626 73.938 ;
               RECT 27.574 74.502 27.626 74.538 ;
               RECT 27.574 75.102 27.626 75.138 ;
               RECT 27.574 75.702 27.626 75.738 ;
               RECT 27.574 76.302 27.626 76.338 ;
               RECT 27.574 76.902 27.626 76.938 ;
               RECT 27.574 77.502 27.626 77.538 ;
               RECT 27.574 78.102 27.626 78.138 ;
               RECT 27.574 78.702 27.626 78.738 ;
               RECT 27.574 79.302 27.626 79.338 ;
               RECT 27.574 79.902 27.626 79.938 ;
               RECT 27.574 80.502 27.626 80.538 ;
               RECT 27.574 81.102 27.626 81.138 ;
               RECT 27.574 81.702 27.626 81.738 ;
               RECT 27.574 82.302 27.626 82.338 ;
               RECT 27.574 82.902 27.626 82.938 ;
               RECT 27.574 83.502 27.626 83.538 ;
               RECT 27.574 84.102 27.626 84.138 ;
               RECT 27.574 84.702 27.626 84.738 ;
               RECT 27.574 85.302 27.626 85.338 ;
               RECT 27.574 85.902 27.626 85.938 ;
               RECT 27.574 86.502 27.626 86.538 ;
               RECT 27.574 87.102 27.626 87.138 ;
               RECT 27.574 87.702 27.626 87.738 ;
               RECT 27.574 88.302 27.626 88.338 ;
               RECT 27.574 88.902 27.626 88.938 ;
               RECT 27.574 89.502 27.626 89.538 ;
               RECT 27.574 90.102 27.626 90.138 ;
               RECT 27.574 90.702 27.626 90.738 ;
               RECT 27.574 91.302 27.626 91.338 ;
               RECT 27.574 91.902 27.626 91.938 ;
               RECT 27.574 92.502 27.626 92.538 ;
               RECT 27.574 93.102 27.626 93.138 ;
               RECT 27.574 93.702 27.626 93.738 ;
               RECT 27.574 94.302 27.626 94.338 ;
               RECT 27.574 94.902 27.626 94.938 ;
               RECT 27.574 95.502 27.626 95.538 ;
               RECT 27.574 96.102 27.626 96.138 ;
               RECT 27.574 96.702 27.626 96.738 ;
               RECT 27.574 97.302 27.626 97.338 ;
               RECT 27.574 97.902 27.626 97.938 ;
               RECT 27.574 98.502 27.626 98.538 ;
               RECT 27.574 99.102 27.626 99.138 ;
               RECT 27.574 99.702 27.626 99.738 ;
               RECT 27.574 100.302 27.626 100.338 ;
               RECT 27.574 100.902 27.626 100.938 ;
               RECT 27.574 101.502 27.626 101.538 ;
               RECT 27.574 102.102 27.626 102.138 ;
               RECT 27.574 102.702 27.626 102.738 ;
               RECT 27.574 103.302 27.626 103.338 ;
               RECT 27.574 103.902 27.626 103.938 ;
               RECT 27.574 104.502 27.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 28.374 0.5695 28.426 104.5505 ;
               LAYER v4 ;
               RECT 28.374 0.582 28.426 0.618 ;
               RECT 28.374 1.182 28.426 1.218 ;
               RECT 28.374 1.782 28.426 1.818 ;
               RECT 28.374 2.382 28.426 2.418 ;
               RECT 28.374 2.982 28.426 3.018 ;
               RECT 28.374 3.582 28.426 3.618 ;
               RECT 28.374 4.182 28.426 4.218 ;
               RECT 28.374 4.782 28.426 4.818 ;
               RECT 28.374 5.382 28.426 5.418 ;
               RECT 28.374 5.982 28.426 6.018 ;
               RECT 28.374 6.582 28.426 6.618 ;
               RECT 28.374 7.182 28.426 7.218 ;
               RECT 28.374 7.782 28.426 7.818 ;
               RECT 28.374 8.382 28.426 8.418 ;
               RECT 28.374 8.982 28.426 9.018 ;
               RECT 28.374 9.582 28.426 9.618 ;
               RECT 28.374 10.182 28.426 10.218 ;
               RECT 28.374 10.782 28.426 10.818 ;
               RECT 28.374 11.382 28.426 11.418 ;
               RECT 28.374 11.982 28.426 12.018 ;
               RECT 28.374 12.582 28.426 12.618 ;
               RECT 28.374 13.182 28.426 13.218 ;
               RECT 28.374 13.782 28.426 13.818 ;
               RECT 28.374 14.382 28.426 14.418 ;
               RECT 28.374 14.982 28.426 15.018 ;
               RECT 28.374 15.582 28.426 15.618 ;
               RECT 28.374 16.182 28.426 16.218 ;
               RECT 28.374 16.782 28.426 16.818 ;
               RECT 28.374 17.382 28.426 17.418 ;
               RECT 28.374 17.982 28.426 18.018 ;
               RECT 28.374 18.582 28.426 18.618 ;
               RECT 28.374 19.182 28.426 19.218 ;
               RECT 28.374 19.782 28.426 19.818 ;
               RECT 28.374 20.382 28.426 20.418 ;
               RECT 28.374 20.982 28.426 21.018 ;
               RECT 28.374 21.582 28.426 21.618 ;
               RECT 28.374 22.182 28.426 22.218 ;
               RECT 28.374 22.782 28.426 22.818 ;
               RECT 28.374 23.382 28.426 23.418 ;
               RECT 28.374 23.982 28.426 24.018 ;
               RECT 28.374 24.582 28.426 24.618 ;
               RECT 28.374 25.182 28.426 25.218 ;
               RECT 28.374 25.782 28.426 25.818 ;
               RECT 28.374 26.382 28.426 26.418 ;
               RECT 28.374 26.982 28.426 27.018 ;
               RECT 28.374 27.582 28.426 27.618 ;
               RECT 28.374 28.182 28.426 28.218 ;
               RECT 28.374 28.782 28.426 28.818 ;
               RECT 28.374 29.382 28.426 29.418 ;
               RECT 28.374 29.982 28.426 30.018 ;
               RECT 28.374 30.582 28.426 30.618 ;
               RECT 28.374 31.182 28.426 31.218 ;
               RECT 28.374 31.782 28.426 31.818 ;
               RECT 28.374 32.382 28.426 32.418 ;
               RECT 28.374 32.982 28.426 33.018 ;
               RECT 28.374 33.582 28.426 33.618 ;
               RECT 28.374 34.182 28.426 34.218 ;
               RECT 28.374 34.782 28.426 34.818 ;
               RECT 28.374 35.382 28.426 35.418 ;
               RECT 28.374 35.982 28.426 36.018 ;
               RECT 28.374 36.582 28.426 36.618 ;
               RECT 28.374 37.182 28.426 37.218 ;
               RECT 28.374 37.782 28.426 37.818 ;
               RECT 28.374 38.382 28.426 38.418 ;
               RECT 28.374 38.982 28.426 39.018 ;
               RECT 28.374 39.582 28.426 39.618 ;
               RECT 28.374 40.182 28.426 40.218 ;
               RECT 28.374 40.782 28.426 40.818 ;
               RECT 28.374 41.382 28.426 41.418 ;
               RECT 28.374 41.982 28.426 42.018 ;
               RECT 28.374 42.582 28.426 42.618 ;
               RECT 28.374 43.182 28.426 43.218 ;
               RECT 28.374 43.782 28.426 43.818 ;
               RECT 28.374 44.382 28.426 44.418 ;
               RECT 28.374 44.982 28.426 45.018 ;
               RECT 28.374 45.582 28.426 45.618 ;
               RECT 28.374 46.182 28.426 46.218 ;
               RECT 28.374 46.782 28.426 46.818 ;
               RECT 28.374 47.382 28.426 47.418 ;
               RECT 28.374 47.982 28.426 48.018 ;
               RECT 28.374 48.582 28.426 48.618 ;
               RECT 28.374 48.942 28.426 48.978 ;
               RECT 28.374 49.182 28.426 49.218 ;
               RECT 28.374 49.902 28.426 49.938 ;
               RECT 28.374 50.622 28.426 50.658 ;
               RECT 28.374 50.862 28.426 50.898 ;
               RECT 28.374 51.342 28.426 51.378 ;
               RECT 28.374 51.822 28.426 51.858 ;
               RECT 28.374 52.302 28.426 52.338 ;
               RECT 28.374 52.782 28.426 52.818 ;
               RECT 28.374 53.262 28.426 53.298 ;
               RECT 28.374 53.742 28.426 53.778 ;
               RECT 28.374 54.222 28.426 54.258 ;
               RECT 28.374 54.462 28.426 54.498 ;
               RECT 28.374 55.182 28.426 55.218 ;
               RECT 28.374 55.902 28.426 55.938 ;
               RECT 28.374 56.142 28.426 56.178 ;
               RECT 28.374 56.502 28.426 56.538 ;
               RECT 28.374 57.102 28.426 57.138 ;
               RECT 28.374 57.702 28.426 57.738 ;
               RECT 28.374 58.302 28.426 58.338 ;
               RECT 28.374 58.902 28.426 58.938 ;
               RECT 28.374 59.502 28.426 59.538 ;
               RECT 28.374 60.102 28.426 60.138 ;
               RECT 28.374 60.702 28.426 60.738 ;
               RECT 28.374 61.302 28.426 61.338 ;
               RECT 28.374 61.902 28.426 61.938 ;
               RECT 28.374 62.502 28.426 62.538 ;
               RECT 28.374 63.102 28.426 63.138 ;
               RECT 28.374 63.702 28.426 63.738 ;
               RECT 28.374 64.302 28.426 64.338 ;
               RECT 28.374 64.902 28.426 64.938 ;
               RECT 28.374 65.502 28.426 65.538 ;
               RECT 28.374 66.102 28.426 66.138 ;
               RECT 28.374 66.702 28.426 66.738 ;
               RECT 28.374 67.302 28.426 67.338 ;
               RECT 28.374 67.902 28.426 67.938 ;
               RECT 28.374 68.502 28.426 68.538 ;
               RECT 28.374 69.102 28.426 69.138 ;
               RECT 28.374 69.702 28.426 69.738 ;
               RECT 28.374 70.302 28.426 70.338 ;
               RECT 28.374 70.902 28.426 70.938 ;
               RECT 28.374 71.502 28.426 71.538 ;
               RECT 28.374 72.102 28.426 72.138 ;
               RECT 28.374 72.702 28.426 72.738 ;
               RECT 28.374 73.302 28.426 73.338 ;
               RECT 28.374 73.902 28.426 73.938 ;
               RECT 28.374 74.502 28.426 74.538 ;
               RECT 28.374 75.102 28.426 75.138 ;
               RECT 28.374 75.702 28.426 75.738 ;
               RECT 28.374 76.302 28.426 76.338 ;
               RECT 28.374 76.902 28.426 76.938 ;
               RECT 28.374 77.502 28.426 77.538 ;
               RECT 28.374 78.102 28.426 78.138 ;
               RECT 28.374 78.702 28.426 78.738 ;
               RECT 28.374 79.302 28.426 79.338 ;
               RECT 28.374 79.902 28.426 79.938 ;
               RECT 28.374 80.502 28.426 80.538 ;
               RECT 28.374 81.102 28.426 81.138 ;
               RECT 28.374 81.702 28.426 81.738 ;
               RECT 28.374 82.302 28.426 82.338 ;
               RECT 28.374 82.902 28.426 82.938 ;
               RECT 28.374 83.502 28.426 83.538 ;
               RECT 28.374 84.102 28.426 84.138 ;
               RECT 28.374 84.702 28.426 84.738 ;
               RECT 28.374 85.302 28.426 85.338 ;
               RECT 28.374 85.902 28.426 85.938 ;
               RECT 28.374 86.502 28.426 86.538 ;
               RECT 28.374 87.102 28.426 87.138 ;
               RECT 28.374 87.702 28.426 87.738 ;
               RECT 28.374 88.302 28.426 88.338 ;
               RECT 28.374 88.902 28.426 88.938 ;
               RECT 28.374 89.502 28.426 89.538 ;
               RECT 28.374 90.102 28.426 90.138 ;
               RECT 28.374 90.702 28.426 90.738 ;
               RECT 28.374 91.302 28.426 91.338 ;
               RECT 28.374 91.902 28.426 91.938 ;
               RECT 28.374 92.502 28.426 92.538 ;
               RECT 28.374 93.102 28.426 93.138 ;
               RECT 28.374 93.702 28.426 93.738 ;
               RECT 28.374 94.302 28.426 94.338 ;
               RECT 28.374 94.902 28.426 94.938 ;
               RECT 28.374 95.502 28.426 95.538 ;
               RECT 28.374 96.102 28.426 96.138 ;
               RECT 28.374 96.702 28.426 96.738 ;
               RECT 28.374 97.302 28.426 97.338 ;
               RECT 28.374 97.902 28.426 97.938 ;
               RECT 28.374 98.502 28.426 98.538 ;
               RECT 28.374 99.102 28.426 99.138 ;
               RECT 28.374 99.702 28.426 99.738 ;
               RECT 28.374 100.302 28.426 100.338 ;
               RECT 28.374 100.902 28.426 100.938 ;
               RECT 28.374 101.502 28.426 101.538 ;
               RECT 28.374 102.102 28.426 102.138 ;
               RECT 28.374 102.702 28.426 102.738 ;
               RECT 28.374 103.302 28.426 103.338 ;
               RECT 28.374 103.902 28.426 103.938 ;
               RECT 28.374 104.502 28.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 29.174 0.5695 29.226 104.5505 ;
               LAYER v4 ;
               RECT 29.174 0.582 29.226 0.618 ;
               RECT 29.174 1.182 29.226 1.218 ;
               RECT 29.174 1.782 29.226 1.818 ;
               RECT 29.174 2.382 29.226 2.418 ;
               RECT 29.174 2.982 29.226 3.018 ;
               RECT 29.174 3.582 29.226 3.618 ;
               RECT 29.174 4.182 29.226 4.218 ;
               RECT 29.174 4.782 29.226 4.818 ;
               RECT 29.174 5.382 29.226 5.418 ;
               RECT 29.174 5.982 29.226 6.018 ;
               RECT 29.174 6.582 29.226 6.618 ;
               RECT 29.174 7.182 29.226 7.218 ;
               RECT 29.174 7.782 29.226 7.818 ;
               RECT 29.174 8.382 29.226 8.418 ;
               RECT 29.174 8.982 29.226 9.018 ;
               RECT 29.174 9.582 29.226 9.618 ;
               RECT 29.174 10.182 29.226 10.218 ;
               RECT 29.174 10.782 29.226 10.818 ;
               RECT 29.174 11.382 29.226 11.418 ;
               RECT 29.174 11.982 29.226 12.018 ;
               RECT 29.174 12.582 29.226 12.618 ;
               RECT 29.174 13.182 29.226 13.218 ;
               RECT 29.174 13.782 29.226 13.818 ;
               RECT 29.174 14.382 29.226 14.418 ;
               RECT 29.174 14.982 29.226 15.018 ;
               RECT 29.174 15.582 29.226 15.618 ;
               RECT 29.174 16.182 29.226 16.218 ;
               RECT 29.174 16.782 29.226 16.818 ;
               RECT 29.174 17.382 29.226 17.418 ;
               RECT 29.174 17.982 29.226 18.018 ;
               RECT 29.174 18.582 29.226 18.618 ;
               RECT 29.174 19.182 29.226 19.218 ;
               RECT 29.174 19.782 29.226 19.818 ;
               RECT 29.174 20.382 29.226 20.418 ;
               RECT 29.174 20.982 29.226 21.018 ;
               RECT 29.174 21.582 29.226 21.618 ;
               RECT 29.174 22.182 29.226 22.218 ;
               RECT 29.174 22.782 29.226 22.818 ;
               RECT 29.174 23.382 29.226 23.418 ;
               RECT 29.174 23.982 29.226 24.018 ;
               RECT 29.174 24.582 29.226 24.618 ;
               RECT 29.174 25.182 29.226 25.218 ;
               RECT 29.174 25.782 29.226 25.818 ;
               RECT 29.174 26.382 29.226 26.418 ;
               RECT 29.174 26.982 29.226 27.018 ;
               RECT 29.174 27.582 29.226 27.618 ;
               RECT 29.174 28.182 29.226 28.218 ;
               RECT 29.174 28.782 29.226 28.818 ;
               RECT 29.174 29.382 29.226 29.418 ;
               RECT 29.174 29.982 29.226 30.018 ;
               RECT 29.174 30.582 29.226 30.618 ;
               RECT 29.174 31.182 29.226 31.218 ;
               RECT 29.174 31.782 29.226 31.818 ;
               RECT 29.174 32.382 29.226 32.418 ;
               RECT 29.174 32.982 29.226 33.018 ;
               RECT 29.174 33.582 29.226 33.618 ;
               RECT 29.174 34.182 29.226 34.218 ;
               RECT 29.174 34.782 29.226 34.818 ;
               RECT 29.174 35.382 29.226 35.418 ;
               RECT 29.174 35.982 29.226 36.018 ;
               RECT 29.174 36.582 29.226 36.618 ;
               RECT 29.174 37.182 29.226 37.218 ;
               RECT 29.174 37.782 29.226 37.818 ;
               RECT 29.174 38.382 29.226 38.418 ;
               RECT 29.174 38.982 29.226 39.018 ;
               RECT 29.174 39.582 29.226 39.618 ;
               RECT 29.174 40.182 29.226 40.218 ;
               RECT 29.174 40.782 29.226 40.818 ;
               RECT 29.174 41.382 29.226 41.418 ;
               RECT 29.174 41.982 29.226 42.018 ;
               RECT 29.174 42.582 29.226 42.618 ;
               RECT 29.174 43.182 29.226 43.218 ;
               RECT 29.174 43.782 29.226 43.818 ;
               RECT 29.174 44.382 29.226 44.418 ;
               RECT 29.174 44.982 29.226 45.018 ;
               RECT 29.174 45.582 29.226 45.618 ;
               RECT 29.174 46.182 29.226 46.218 ;
               RECT 29.174 46.782 29.226 46.818 ;
               RECT 29.174 47.382 29.226 47.418 ;
               RECT 29.174 47.982 29.226 48.018 ;
               RECT 29.174 48.582 29.226 48.618 ;
               RECT 29.174 48.942 29.226 48.978 ;
               RECT 29.174 48.9475 29.226 48.9725 ;
               RECT 29.174 49.182 29.226 49.218 ;
               RECT 29.174 49.902 29.226 49.938 ;
               RECT 29.174 50.622 29.226 50.658 ;
               RECT 29.174 50.862 29.226 50.898 ;
               RECT 29.174 51.342 29.226 51.378 ;
               RECT 29.174 51.822 29.226 51.858 ;
               RECT 29.174 52.302 29.226 52.338 ;
               RECT 29.174 52.782 29.226 52.818 ;
               RECT 29.174 53.262 29.226 53.298 ;
               RECT 29.174 53.742 29.226 53.778 ;
               RECT 29.174 54.222 29.226 54.258 ;
               RECT 29.174 54.462 29.226 54.498 ;
               RECT 29.174 55.182 29.226 55.218 ;
               RECT 29.174 55.902 29.226 55.938 ;
               RECT 29.174 56.142 29.226 56.178 ;
               RECT 29.174 56.1475 29.226 56.1725 ;
               RECT 29.174 56.502 29.226 56.538 ;
               RECT 29.174 57.102 29.226 57.138 ;
               RECT 29.174 57.702 29.226 57.738 ;
               RECT 29.174 58.302 29.226 58.338 ;
               RECT 29.174 58.902 29.226 58.938 ;
               RECT 29.174 59.502 29.226 59.538 ;
               RECT 29.174 60.102 29.226 60.138 ;
               RECT 29.174 60.702 29.226 60.738 ;
               RECT 29.174 61.302 29.226 61.338 ;
               RECT 29.174 61.902 29.226 61.938 ;
               RECT 29.174 62.502 29.226 62.538 ;
               RECT 29.174 63.102 29.226 63.138 ;
               RECT 29.174 63.702 29.226 63.738 ;
               RECT 29.174 64.302 29.226 64.338 ;
               RECT 29.174 64.902 29.226 64.938 ;
               RECT 29.174 65.502 29.226 65.538 ;
               RECT 29.174 66.102 29.226 66.138 ;
               RECT 29.174 66.702 29.226 66.738 ;
               RECT 29.174 67.302 29.226 67.338 ;
               RECT 29.174 67.902 29.226 67.938 ;
               RECT 29.174 68.502 29.226 68.538 ;
               RECT 29.174 69.102 29.226 69.138 ;
               RECT 29.174 69.702 29.226 69.738 ;
               RECT 29.174 70.302 29.226 70.338 ;
               RECT 29.174 70.902 29.226 70.938 ;
               RECT 29.174 71.502 29.226 71.538 ;
               RECT 29.174 72.102 29.226 72.138 ;
               RECT 29.174 72.702 29.226 72.738 ;
               RECT 29.174 73.302 29.226 73.338 ;
               RECT 29.174 73.902 29.226 73.938 ;
               RECT 29.174 74.502 29.226 74.538 ;
               RECT 29.174 75.102 29.226 75.138 ;
               RECT 29.174 75.702 29.226 75.738 ;
               RECT 29.174 76.302 29.226 76.338 ;
               RECT 29.174 76.902 29.226 76.938 ;
               RECT 29.174 77.502 29.226 77.538 ;
               RECT 29.174 78.102 29.226 78.138 ;
               RECT 29.174 78.702 29.226 78.738 ;
               RECT 29.174 79.302 29.226 79.338 ;
               RECT 29.174 79.902 29.226 79.938 ;
               RECT 29.174 80.502 29.226 80.538 ;
               RECT 29.174 81.102 29.226 81.138 ;
               RECT 29.174 81.702 29.226 81.738 ;
               RECT 29.174 82.302 29.226 82.338 ;
               RECT 29.174 82.902 29.226 82.938 ;
               RECT 29.174 83.502 29.226 83.538 ;
               RECT 29.174 84.102 29.226 84.138 ;
               RECT 29.174 84.702 29.226 84.738 ;
               RECT 29.174 85.302 29.226 85.338 ;
               RECT 29.174 85.902 29.226 85.938 ;
               RECT 29.174 86.502 29.226 86.538 ;
               RECT 29.174 87.102 29.226 87.138 ;
               RECT 29.174 87.702 29.226 87.738 ;
               RECT 29.174 88.302 29.226 88.338 ;
               RECT 29.174 88.902 29.226 88.938 ;
               RECT 29.174 89.502 29.226 89.538 ;
               RECT 29.174 90.102 29.226 90.138 ;
               RECT 29.174 90.702 29.226 90.738 ;
               RECT 29.174 91.302 29.226 91.338 ;
               RECT 29.174 91.902 29.226 91.938 ;
               RECT 29.174 92.502 29.226 92.538 ;
               RECT 29.174 93.102 29.226 93.138 ;
               RECT 29.174 93.702 29.226 93.738 ;
               RECT 29.174 94.302 29.226 94.338 ;
               RECT 29.174 94.902 29.226 94.938 ;
               RECT 29.174 95.502 29.226 95.538 ;
               RECT 29.174 96.102 29.226 96.138 ;
               RECT 29.174 96.702 29.226 96.738 ;
               RECT 29.174 97.302 29.226 97.338 ;
               RECT 29.174 97.902 29.226 97.938 ;
               RECT 29.174 98.502 29.226 98.538 ;
               RECT 29.174 99.102 29.226 99.138 ;
               RECT 29.174 99.702 29.226 99.738 ;
               RECT 29.174 100.302 29.226 100.338 ;
               RECT 29.174 100.902 29.226 100.938 ;
               RECT 29.174 101.502 29.226 101.538 ;
               RECT 29.174 102.102 29.226 102.138 ;
               RECT 29.174 102.702 29.226 102.738 ;
               RECT 29.174 103.302 29.226 103.338 ;
               RECT 29.174 103.902 29.226 103.938 ;
               RECT 29.174 104.502 29.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 29.974 0.5695 30.026 104.5505 ;
               LAYER v4 ;
               RECT 29.974 0.582 30.026 0.618 ;
               RECT 29.974 1.182 30.026 1.218 ;
               RECT 29.974 1.782 30.026 1.818 ;
               RECT 29.974 2.382 30.026 2.418 ;
               RECT 29.974 2.982 30.026 3.018 ;
               RECT 29.974 3.582 30.026 3.618 ;
               RECT 29.974 4.182 30.026 4.218 ;
               RECT 29.974 4.782 30.026 4.818 ;
               RECT 29.974 5.382 30.026 5.418 ;
               RECT 29.974 5.982 30.026 6.018 ;
               RECT 29.974 6.582 30.026 6.618 ;
               RECT 29.974 7.182 30.026 7.218 ;
               RECT 29.974 7.782 30.026 7.818 ;
               RECT 29.974 8.382 30.026 8.418 ;
               RECT 29.974 8.982 30.026 9.018 ;
               RECT 29.974 9.582 30.026 9.618 ;
               RECT 29.974 10.182 30.026 10.218 ;
               RECT 29.974 10.782 30.026 10.818 ;
               RECT 29.974 11.382 30.026 11.418 ;
               RECT 29.974 11.982 30.026 12.018 ;
               RECT 29.974 12.582 30.026 12.618 ;
               RECT 29.974 13.182 30.026 13.218 ;
               RECT 29.974 13.782 30.026 13.818 ;
               RECT 29.974 14.382 30.026 14.418 ;
               RECT 29.974 14.982 30.026 15.018 ;
               RECT 29.974 15.582 30.026 15.618 ;
               RECT 29.974 16.182 30.026 16.218 ;
               RECT 29.974 16.782 30.026 16.818 ;
               RECT 29.974 17.382 30.026 17.418 ;
               RECT 29.974 17.982 30.026 18.018 ;
               RECT 29.974 18.582 30.026 18.618 ;
               RECT 29.974 19.182 30.026 19.218 ;
               RECT 29.974 19.782 30.026 19.818 ;
               RECT 29.974 20.382 30.026 20.418 ;
               RECT 29.974 20.982 30.026 21.018 ;
               RECT 29.974 21.582 30.026 21.618 ;
               RECT 29.974 22.182 30.026 22.218 ;
               RECT 29.974 22.782 30.026 22.818 ;
               RECT 29.974 23.382 30.026 23.418 ;
               RECT 29.974 23.982 30.026 24.018 ;
               RECT 29.974 24.582 30.026 24.618 ;
               RECT 29.974 25.182 30.026 25.218 ;
               RECT 29.974 25.782 30.026 25.818 ;
               RECT 29.974 26.382 30.026 26.418 ;
               RECT 29.974 26.982 30.026 27.018 ;
               RECT 29.974 27.582 30.026 27.618 ;
               RECT 29.974 28.182 30.026 28.218 ;
               RECT 29.974 28.782 30.026 28.818 ;
               RECT 29.974 29.382 30.026 29.418 ;
               RECT 29.974 29.982 30.026 30.018 ;
               RECT 29.974 30.582 30.026 30.618 ;
               RECT 29.974 31.182 30.026 31.218 ;
               RECT 29.974 31.782 30.026 31.818 ;
               RECT 29.974 32.382 30.026 32.418 ;
               RECT 29.974 32.982 30.026 33.018 ;
               RECT 29.974 33.582 30.026 33.618 ;
               RECT 29.974 34.182 30.026 34.218 ;
               RECT 29.974 34.782 30.026 34.818 ;
               RECT 29.974 35.382 30.026 35.418 ;
               RECT 29.974 35.982 30.026 36.018 ;
               RECT 29.974 36.582 30.026 36.618 ;
               RECT 29.974 37.182 30.026 37.218 ;
               RECT 29.974 37.782 30.026 37.818 ;
               RECT 29.974 38.382 30.026 38.418 ;
               RECT 29.974 38.982 30.026 39.018 ;
               RECT 29.974 39.582 30.026 39.618 ;
               RECT 29.974 40.182 30.026 40.218 ;
               RECT 29.974 40.782 30.026 40.818 ;
               RECT 29.974 41.382 30.026 41.418 ;
               RECT 29.974 41.982 30.026 42.018 ;
               RECT 29.974 42.582 30.026 42.618 ;
               RECT 29.974 43.182 30.026 43.218 ;
               RECT 29.974 43.782 30.026 43.818 ;
               RECT 29.974 44.382 30.026 44.418 ;
               RECT 29.974 44.982 30.026 45.018 ;
               RECT 29.974 45.582 30.026 45.618 ;
               RECT 29.974 46.182 30.026 46.218 ;
               RECT 29.974 46.782 30.026 46.818 ;
               RECT 29.974 47.382 30.026 47.418 ;
               RECT 29.974 47.982 30.026 48.018 ;
               RECT 29.974 48.582 30.026 48.618 ;
               RECT 29.974 48.942 30.026 48.978 ;
               RECT 29.974 49.182 30.026 49.218 ;
               RECT 29.974 49.902 30.026 49.938 ;
               RECT 29.974 50.622 30.026 50.658 ;
               RECT 29.974 50.862 30.026 50.898 ;
               RECT 29.974 51.342 30.026 51.378 ;
               RECT 29.974 51.822 30.026 51.858 ;
               RECT 29.974 52.302 30.026 52.338 ;
               RECT 29.974 52.782 30.026 52.818 ;
               RECT 29.974 53.262 30.026 53.298 ;
               RECT 29.974 53.742 30.026 53.778 ;
               RECT 29.974 54.222 30.026 54.258 ;
               RECT 29.974 54.462 30.026 54.498 ;
               RECT 29.974 55.182 30.026 55.218 ;
               RECT 29.974 55.902 30.026 55.938 ;
               RECT 29.974 56.142 30.026 56.178 ;
               RECT 29.974 56.502 30.026 56.538 ;
               RECT 29.974 57.102 30.026 57.138 ;
               RECT 29.974 57.702 30.026 57.738 ;
               RECT 29.974 58.302 30.026 58.338 ;
               RECT 29.974 58.902 30.026 58.938 ;
               RECT 29.974 59.502 30.026 59.538 ;
               RECT 29.974 60.102 30.026 60.138 ;
               RECT 29.974 60.702 30.026 60.738 ;
               RECT 29.974 61.302 30.026 61.338 ;
               RECT 29.974 61.902 30.026 61.938 ;
               RECT 29.974 62.502 30.026 62.538 ;
               RECT 29.974 63.102 30.026 63.138 ;
               RECT 29.974 63.702 30.026 63.738 ;
               RECT 29.974 64.302 30.026 64.338 ;
               RECT 29.974 64.902 30.026 64.938 ;
               RECT 29.974 65.502 30.026 65.538 ;
               RECT 29.974 66.102 30.026 66.138 ;
               RECT 29.974 66.702 30.026 66.738 ;
               RECT 29.974 67.302 30.026 67.338 ;
               RECT 29.974 67.902 30.026 67.938 ;
               RECT 29.974 68.502 30.026 68.538 ;
               RECT 29.974 69.102 30.026 69.138 ;
               RECT 29.974 69.702 30.026 69.738 ;
               RECT 29.974 70.302 30.026 70.338 ;
               RECT 29.974 70.902 30.026 70.938 ;
               RECT 29.974 71.502 30.026 71.538 ;
               RECT 29.974 72.102 30.026 72.138 ;
               RECT 29.974 72.702 30.026 72.738 ;
               RECT 29.974 73.302 30.026 73.338 ;
               RECT 29.974 73.902 30.026 73.938 ;
               RECT 29.974 74.502 30.026 74.538 ;
               RECT 29.974 75.102 30.026 75.138 ;
               RECT 29.974 75.702 30.026 75.738 ;
               RECT 29.974 76.302 30.026 76.338 ;
               RECT 29.974 76.902 30.026 76.938 ;
               RECT 29.974 77.502 30.026 77.538 ;
               RECT 29.974 78.102 30.026 78.138 ;
               RECT 29.974 78.702 30.026 78.738 ;
               RECT 29.974 79.302 30.026 79.338 ;
               RECT 29.974 79.902 30.026 79.938 ;
               RECT 29.974 80.502 30.026 80.538 ;
               RECT 29.974 81.102 30.026 81.138 ;
               RECT 29.974 81.702 30.026 81.738 ;
               RECT 29.974 82.302 30.026 82.338 ;
               RECT 29.974 82.902 30.026 82.938 ;
               RECT 29.974 83.502 30.026 83.538 ;
               RECT 29.974 84.102 30.026 84.138 ;
               RECT 29.974 84.702 30.026 84.738 ;
               RECT 29.974 85.302 30.026 85.338 ;
               RECT 29.974 85.902 30.026 85.938 ;
               RECT 29.974 86.502 30.026 86.538 ;
               RECT 29.974 87.102 30.026 87.138 ;
               RECT 29.974 87.702 30.026 87.738 ;
               RECT 29.974 88.302 30.026 88.338 ;
               RECT 29.974 88.902 30.026 88.938 ;
               RECT 29.974 89.502 30.026 89.538 ;
               RECT 29.974 90.102 30.026 90.138 ;
               RECT 29.974 90.702 30.026 90.738 ;
               RECT 29.974 91.302 30.026 91.338 ;
               RECT 29.974 91.902 30.026 91.938 ;
               RECT 29.974 92.502 30.026 92.538 ;
               RECT 29.974 93.102 30.026 93.138 ;
               RECT 29.974 93.702 30.026 93.738 ;
               RECT 29.974 94.302 30.026 94.338 ;
               RECT 29.974 94.902 30.026 94.938 ;
               RECT 29.974 95.502 30.026 95.538 ;
               RECT 29.974 96.102 30.026 96.138 ;
               RECT 29.974 96.702 30.026 96.738 ;
               RECT 29.974 97.302 30.026 97.338 ;
               RECT 29.974 97.902 30.026 97.938 ;
               RECT 29.974 98.502 30.026 98.538 ;
               RECT 29.974 99.102 30.026 99.138 ;
               RECT 29.974 99.702 30.026 99.738 ;
               RECT 29.974 100.302 30.026 100.338 ;
               RECT 29.974 100.902 30.026 100.938 ;
               RECT 29.974 101.502 30.026 101.538 ;
               RECT 29.974 102.102 30.026 102.138 ;
               RECT 29.974 102.702 30.026 102.738 ;
               RECT 29.974 103.302 30.026 103.338 ;
               RECT 29.974 103.902 30.026 103.938 ;
               RECT 29.974 104.502 30.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 3.774 0.5695 3.826 104.5505 ;
               LAYER v4 ;
               RECT 3.774 0.582 3.826 0.618 ;
               RECT 3.774 1.182 3.826 1.218 ;
               RECT 3.774 1.782 3.826 1.818 ;
               RECT 3.774 2.382 3.826 2.418 ;
               RECT 3.774 2.982 3.826 3.018 ;
               RECT 3.774 3.582 3.826 3.618 ;
               RECT 3.774 4.182 3.826 4.218 ;
               RECT 3.774 4.782 3.826 4.818 ;
               RECT 3.774 5.382 3.826 5.418 ;
               RECT 3.774 5.982 3.826 6.018 ;
               RECT 3.774 6.582 3.826 6.618 ;
               RECT 3.774 7.182 3.826 7.218 ;
               RECT 3.774 7.782 3.826 7.818 ;
               RECT 3.774 8.382 3.826 8.418 ;
               RECT 3.774 8.982 3.826 9.018 ;
               RECT 3.774 9.582 3.826 9.618 ;
               RECT 3.774 10.182 3.826 10.218 ;
               RECT 3.774 10.782 3.826 10.818 ;
               RECT 3.774 11.382 3.826 11.418 ;
               RECT 3.774 11.982 3.826 12.018 ;
               RECT 3.774 12.582 3.826 12.618 ;
               RECT 3.774 13.182 3.826 13.218 ;
               RECT 3.774 13.782 3.826 13.818 ;
               RECT 3.774 14.382 3.826 14.418 ;
               RECT 3.774 14.982 3.826 15.018 ;
               RECT 3.774 15.582 3.826 15.618 ;
               RECT 3.774 16.182 3.826 16.218 ;
               RECT 3.774 16.782 3.826 16.818 ;
               RECT 3.774 17.382 3.826 17.418 ;
               RECT 3.774 17.982 3.826 18.018 ;
               RECT 3.774 18.582 3.826 18.618 ;
               RECT 3.774 19.182 3.826 19.218 ;
               RECT 3.774 19.782 3.826 19.818 ;
               RECT 3.774 20.382 3.826 20.418 ;
               RECT 3.774 20.982 3.826 21.018 ;
               RECT 3.774 21.582 3.826 21.618 ;
               RECT 3.774 22.182 3.826 22.218 ;
               RECT 3.774 22.782 3.826 22.818 ;
               RECT 3.774 23.382 3.826 23.418 ;
               RECT 3.774 23.982 3.826 24.018 ;
               RECT 3.774 24.582 3.826 24.618 ;
               RECT 3.774 25.182 3.826 25.218 ;
               RECT 3.774 25.782 3.826 25.818 ;
               RECT 3.774 26.382 3.826 26.418 ;
               RECT 3.774 26.982 3.826 27.018 ;
               RECT 3.774 27.582 3.826 27.618 ;
               RECT 3.774 28.182 3.826 28.218 ;
               RECT 3.774 28.782 3.826 28.818 ;
               RECT 3.774 29.382 3.826 29.418 ;
               RECT 3.774 29.982 3.826 30.018 ;
               RECT 3.774 30.582 3.826 30.618 ;
               RECT 3.774 31.182 3.826 31.218 ;
               RECT 3.774 31.782 3.826 31.818 ;
               RECT 3.774 32.382 3.826 32.418 ;
               RECT 3.774 32.982 3.826 33.018 ;
               RECT 3.774 33.582 3.826 33.618 ;
               RECT 3.774 34.182 3.826 34.218 ;
               RECT 3.774 34.782 3.826 34.818 ;
               RECT 3.774 35.382 3.826 35.418 ;
               RECT 3.774 35.982 3.826 36.018 ;
               RECT 3.774 36.582 3.826 36.618 ;
               RECT 3.774 37.182 3.826 37.218 ;
               RECT 3.774 37.782 3.826 37.818 ;
               RECT 3.774 38.382 3.826 38.418 ;
               RECT 3.774 38.982 3.826 39.018 ;
               RECT 3.774 39.582 3.826 39.618 ;
               RECT 3.774 40.182 3.826 40.218 ;
               RECT 3.774 40.782 3.826 40.818 ;
               RECT 3.774 41.382 3.826 41.418 ;
               RECT 3.774 41.982 3.826 42.018 ;
               RECT 3.774 42.582 3.826 42.618 ;
               RECT 3.774 43.182 3.826 43.218 ;
               RECT 3.774 43.782 3.826 43.818 ;
               RECT 3.774 44.382 3.826 44.418 ;
               RECT 3.774 44.982 3.826 45.018 ;
               RECT 3.774 45.582 3.826 45.618 ;
               RECT 3.774 46.182 3.826 46.218 ;
               RECT 3.774 46.782 3.826 46.818 ;
               RECT 3.774 47.382 3.826 47.418 ;
               RECT 3.774 47.982 3.826 48.018 ;
               RECT 3.774 48.582 3.826 48.618 ;
               RECT 3.774 48.942 3.826 48.978 ;
               RECT 3.774 48.9475 3.826 48.9725 ;
               RECT 3.774 49.182 3.826 49.218 ;
               RECT 3.774 49.902 3.826 49.938 ;
               RECT 3.774 50.622 3.826 50.658 ;
               RECT 3.774 50.862 3.826 50.898 ;
               RECT 3.774 51.342 3.826 51.378 ;
               RECT 3.774 51.822 3.826 51.858 ;
               RECT 3.774 52.302 3.826 52.338 ;
               RECT 3.774 52.782 3.826 52.818 ;
               RECT 3.774 53.262 3.826 53.298 ;
               RECT 3.774 53.742 3.826 53.778 ;
               RECT 3.774 54.222 3.826 54.258 ;
               RECT 3.774 54.462 3.826 54.498 ;
               RECT 3.774 55.182 3.826 55.218 ;
               RECT 3.774 55.902 3.826 55.938 ;
               RECT 3.774 56.142 3.826 56.178 ;
               RECT 3.774 56.1475 3.826 56.1725 ;
               RECT 3.774 56.502 3.826 56.538 ;
               RECT 3.774 57.102 3.826 57.138 ;
               RECT 3.774 57.702 3.826 57.738 ;
               RECT 3.774 58.302 3.826 58.338 ;
               RECT 3.774 58.902 3.826 58.938 ;
               RECT 3.774 59.502 3.826 59.538 ;
               RECT 3.774 60.102 3.826 60.138 ;
               RECT 3.774 60.702 3.826 60.738 ;
               RECT 3.774 61.302 3.826 61.338 ;
               RECT 3.774 61.902 3.826 61.938 ;
               RECT 3.774 62.502 3.826 62.538 ;
               RECT 3.774 63.102 3.826 63.138 ;
               RECT 3.774 63.702 3.826 63.738 ;
               RECT 3.774 64.302 3.826 64.338 ;
               RECT 3.774 64.902 3.826 64.938 ;
               RECT 3.774 65.502 3.826 65.538 ;
               RECT 3.774 66.102 3.826 66.138 ;
               RECT 3.774 66.702 3.826 66.738 ;
               RECT 3.774 67.302 3.826 67.338 ;
               RECT 3.774 67.902 3.826 67.938 ;
               RECT 3.774 68.502 3.826 68.538 ;
               RECT 3.774 69.102 3.826 69.138 ;
               RECT 3.774 69.702 3.826 69.738 ;
               RECT 3.774 70.302 3.826 70.338 ;
               RECT 3.774 70.902 3.826 70.938 ;
               RECT 3.774 71.502 3.826 71.538 ;
               RECT 3.774 72.102 3.826 72.138 ;
               RECT 3.774 72.702 3.826 72.738 ;
               RECT 3.774 73.302 3.826 73.338 ;
               RECT 3.774 73.902 3.826 73.938 ;
               RECT 3.774 74.502 3.826 74.538 ;
               RECT 3.774 75.102 3.826 75.138 ;
               RECT 3.774 75.702 3.826 75.738 ;
               RECT 3.774 76.302 3.826 76.338 ;
               RECT 3.774 76.902 3.826 76.938 ;
               RECT 3.774 77.502 3.826 77.538 ;
               RECT 3.774 78.102 3.826 78.138 ;
               RECT 3.774 78.702 3.826 78.738 ;
               RECT 3.774 79.302 3.826 79.338 ;
               RECT 3.774 79.902 3.826 79.938 ;
               RECT 3.774 80.502 3.826 80.538 ;
               RECT 3.774 81.102 3.826 81.138 ;
               RECT 3.774 81.702 3.826 81.738 ;
               RECT 3.774 82.302 3.826 82.338 ;
               RECT 3.774 82.902 3.826 82.938 ;
               RECT 3.774 83.502 3.826 83.538 ;
               RECT 3.774 84.102 3.826 84.138 ;
               RECT 3.774 84.702 3.826 84.738 ;
               RECT 3.774 85.302 3.826 85.338 ;
               RECT 3.774 85.902 3.826 85.938 ;
               RECT 3.774 86.502 3.826 86.538 ;
               RECT 3.774 87.102 3.826 87.138 ;
               RECT 3.774 87.702 3.826 87.738 ;
               RECT 3.774 88.302 3.826 88.338 ;
               RECT 3.774 88.902 3.826 88.938 ;
               RECT 3.774 89.502 3.826 89.538 ;
               RECT 3.774 90.102 3.826 90.138 ;
               RECT 3.774 90.702 3.826 90.738 ;
               RECT 3.774 91.302 3.826 91.338 ;
               RECT 3.774 91.902 3.826 91.938 ;
               RECT 3.774 92.502 3.826 92.538 ;
               RECT 3.774 93.102 3.826 93.138 ;
               RECT 3.774 93.702 3.826 93.738 ;
               RECT 3.774 94.302 3.826 94.338 ;
               RECT 3.774 94.902 3.826 94.938 ;
               RECT 3.774 95.502 3.826 95.538 ;
               RECT 3.774 96.102 3.826 96.138 ;
               RECT 3.774 96.702 3.826 96.738 ;
               RECT 3.774 97.302 3.826 97.338 ;
               RECT 3.774 97.902 3.826 97.938 ;
               RECT 3.774 98.502 3.826 98.538 ;
               RECT 3.774 99.102 3.826 99.138 ;
               RECT 3.774 99.702 3.826 99.738 ;
               RECT 3.774 100.302 3.826 100.338 ;
               RECT 3.774 100.902 3.826 100.938 ;
               RECT 3.774 101.502 3.826 101.538 ;
               RECT 3.774 102.102 3.826 102.138 ;
               RECT 3.774 102.702 3.826 102.738 ;
               RECT 3.774 103.302 3.826 103.338 ;
               RECT 3.774 103.902 3.826 103.938 ;
               RECT 3.774 104.502 3.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 30.774 0.5695 30.826 104.5505 ;
               LAYER v4 ;
               RECT 30.774 0.582 30.826 0.618 ;
               RECT 30.774 1.182 30.826 1.218 ;
               RECT 30.774 1.782 30.826 1.818 ;
               RECT 30.774 2.382 30.826 2.418 ;
               RECT 30.774 2.982 30.826 3.018 ;
               RECT 30.774 3.582 30.826 3.618 ;
               RECT 30.774 4.182 30.826 4.218 ;
               RECT 30.774 4.782 30.826 4.818 ;
               RECT 30.774 5.382 30.826 5.418 ;
               RECT 30.774 5.982 30.826 6.018 ;
               RECT 30.774 6.582 30.826 6.618 ;
               RECT 30.774 7.182 30.826 7.218 ;
               RECT 30.774 7.782 30.826 7.818 ;
               RECT 30.774 8.382 30.826 8.418 ;
               RECT 30.774 8.982 30.826 9.018 ;
               RECT 30.774 9.582 30.826 9.618 ;
               RECT 30.774 10.182 30.826 10.218 ;
               RECT 30.774 10.782 30.826 10.818 ;
               RECT 30.774 11.382 30.826 11.418 ;
               RECT 30.774 11.982 30.826 12.018 ;
               RECT 30.774 12.582 30.826 12.618 ;
               RECT 30.774 13.182 30.826 13.218 ;
               RECT 30.774 13.782 30.826 13.818 ;
               RECT 30.774 14.382 30.826 14.418 ;
               RECT 30.774 14.982 30.826 15.018 ;
               RECT 30.774 15.582 30.826 15.618 ;
               RECT 30.774 16.182 30.826 16.218 ;
               RECT 30.774 16.782 30.826 16.818 ;
               RECT 30.774 17.382 30.826 17.418 ;
               RECT 30.774 17.982 30.826 18.018 ;
               RECT 30.774 18.582 30.826 18.618 ;
               RECT 30.774 19.182 30.826 19.218 ;
               RECT 30.774 19.782 30.826 19.818 ;
               RECT 30.774 20.382 30.826 20.418 ;
               RECT 30.774 20.982 30.826 21.018 ;
               RECT 30.774 21.582 30.826 21.618 ;
               RECT 30.774 22.182 30.826 22.218 ;
               RECT 30.774 22.782 30.826 22.818 ;
               RECT 30.774 23.382 30.826 23.418 ;
               RECT 30.774 23.982 30.826 24.018 ;
               RECT 30.774 24.582 30.826 24.618 ;
               RECT 30.774 25.182 30.826 25.218 ;
               RECT 30.774 25.782 30.826 25.818 ;
               RECT 30.774 26.382 30.826 26.418 ;
               RECT 30.774 26.982 30.826 27.018 ;
               RECT 30.774 27.582 30.826 27.618 ;
               RECT 30.774 28.182 30.826 28.218 ;
               RECT 30.774 28.782 30.826 28.818 ;
               RECT 30.774 29.382 30.826 29.418 ;
               RECT 30.774 29.982 30.826 30.018 ;
               RECT 30.774 30.582 30.826 30.618 ;
               RECT 30.774 31.182 30.826 31.218 ;
               RECT 30.774 31.782 30.826 31.818 ;
               RECT 30.774 32.382 30.826 32.418 ;
               RECT 30.774 32.982 30.826 33.018 ;
               RECT 30.774 33.582 30.826 33.618 ;
               RECT 30.774 34.182 30.826 34.218 ;
               RECT 30.774 34.782 30.826 34.818 ;
               RECT 30.774 35.382 30.826 35.418 ;
               RECT 30.774 35.982 30.826 36.018 ;
               RECT 30.774 36.582 30.826 36.618 ;
               RECT 30.774 37.182 30.826 37.218 ;
               RECT 30.774 37.782 30.826 37.818 ;
               RECT 30.774 38.382 30.826 38.418 ;
               RECT 30.774 38.982 30.826 39.018 ;
               RECT 30.774 39.582 30.826 39.618 ;
               RECT 30.774 40.182 30.826 40.218 ;
               RECT 30.774 40.782 30.826 40.818 ;
               RECT 30.774 41.382 30.826 41.418 ;
               RECT 30.774 41.982 30.826 42.018 ;
               RECT 30.774 42.582 30.826 42.618 ;
               RECT 30.774 43.182 30.826 43.218 ;
               RECT 30.774 43.782 30.826 43.818 ;
               RECT 30.774 44.382 30.826 44.418 ;
               RECT 30.774 44.982 30.826 45.018 ;
               RECT 30.774 45.582 30.826 45.618 ;
               RECT 30.774 46.182 30.826 46.218 ;
               RECT 30.774 46.782 30.826 46.818 ;
               RECT 30.774 47.382 30.826 47.418 ;
               RECT 30.774 47.982 30.826 48.018 ;
               RECT 30.774 48.582 30.826 48.618 ;
               RECT 30.774 48.942 30.826 48.978 ;
               RECT 30.774 48.9475 30.826 48.9725 ;
               RECT 30.774 49.182 30.826 49.218 ;
               RECT 30.774 49.902 30.826 49.938 ;
               RECT 30.774 50.622 30.826 50.658 ;
               RECT 30.774 50.862 30.826 50.898 ;
               RECT 30.774 51.342 30.826 51.378 ;
               RECT 30.774 51.822 30.826 51.858 ;
               RECT 30.774 52.302 30.826 52.338 ;
               RECT 30.774 52.782 30.826 52.818 ;
               RECT 30.774 53.262 30.826 53.298 ;
               RECT 30.774 53.742 30.826 53.778 ;
               RECT 30.774 54.222 30.826 54.258 ;
               RECT 30.774 54.462 30.826 54.498 ;
               RECT 30.774 55.182 30.826 55.218 ;
               RECT 30.774 55.902 30.826 55.938 ;
               RECT 30.774 56.142 30.826 56.178 ;
               RECT 30.774 56.1475 30.826 56.1725 ;
               RECT 30.774 56.502 30.826 56.538 ;
               RECT 30.774 57.102 30.826 57.138 ;
               RECT 30.774 57.702 30.826 57.738 ;
               RECT 30.774 58.302 30.826 58.338 ;
               RECT 30.774 58.902 30.826 58.938 ;
               RECT 30.774 59.502 30.826 59.538 ;
               RECT 30.774 60.102 30.826 60.138 ;
               RECT 30.774 60.702 30.826 60.738 ;
               RECT 30.774 61.302 30.826 61.338 ;
               RECT 30.774 61.902 30.826 61.938 ;
               RECT 30.774 62.502 30.826 62.538 ;
               RECT 30.774 63.102 30.826 63.138 ;
               RECT 30.774 63.702 30.826 63.738 ;
               RECT 30.774 64.302 30.826 64.338 ;
               RECT 30.774 64.902 30.826 64.938 ;
               RECT 30.774 65.502 30.826 65.538 ;
               RECT 30.774 66.102 30.826 66.138 ;
               RECT 30.774 66.702 30.826 66.738 ;
               RECT 30.774 67.302 30.826 67.338 ;
               RECT 30.774 67.902 30.826 67.938 ;
               RECT 30.774 68.502 30.826 68.538 ;
               RECT 30.774 69.102 30.826 69.138 ;
               RECT 30.774 69.702 30.826 69.738 ;
               RECT 30.774 70.302 30.826 70.338 ;
               RECT 30.774 70.902 30.826 70.938 ;
               RECT 30.774 71.502 30.826 71.538 ;
               RECT 30.774 72.102 30.826 72.138 ;
               RECT 30.774 72.702 30.826 72.738 ;
               RECT 30.774 73.302 30.826 73.338 ;
               RECT 30.774 73.902 30.826 73.938 ;
               RECT 30.774 74.502 30.826 74.538 ;
               RECT 30.774 75.102 30.826 75.138 ;
               RECT 30.774 75.702 30.826 75.738 ;
               RECT 30.774 76.302 30.826 76.338 ;
               RECT 30.774 76.902 30.826 76.938 ;
               RECT 30.774 77.502 30.826 77.538 ;
               RECT 30.774 78.102 30.826 78.138 ;
               RECT 30.774 78.702 30.826 78.738 ;
               RECT 30.774 79.302 30.826 79.338 ;
               RECT 30.774 79.902 30.826 79.938 ;
               RECT 30.774 80.502 30.826 80.538 ;
               RECT 30.774 81.102 30.826 81.138 ;
               RECT 30.774 81.702 30.826 81.738 ;
               RECT 30.774 82.302 30.826 82.338 ;
               RECT 30.774 82.902 30.826 82.938 ;
               RECT 30.774 83.502 30.826 83.538 ;
               RECT 30.774 84.102 30.826 84.138 ;
               RECT 30.774 84.702 30.826 84.738 ;
               RECT 30.774 85.302 30.826 85.338 ;
               RECT 30.774 85.902 30.826 85.938 ;
               RECT 30.774 86.502 30.826 86.538 ;
               RECT 30.774 87.102 30.826 87.138 ;
               RECT 30.774 87.702 30.826 87.738 ;
               RECT 30.774 88.302 30.826 88.338 ;
               RECT 30.774 88.902 30.826 88.938 ;
               RECT 30.774 89.502 30.826 89.538 ;
               RECT 30.774 90.102 30.826 90.138 ;
               RECT 30.774 90.702 30.826 90.738 ;
               RECT 30.774 91.302 30.826 91.338 ;
               RECT 30.774 91.902 30.826 91.938 ;
               RECT 30.774 92.502 30.826 92.538 ;
               RECT 30.774 93.102 30.826 93.138 ;
               RECT 30.774 93.702 30.826 93.738 ;
               RECT 30.774 94.302 30.826 94.338 ;
               RECT 30.774 94.902 30.826 94.938 ;
               RECT 30.774 95.502 30.826 95.538 ;
               RECT 30.774 96.102 30.826 96.138 ;
               RECT 30.774 96.702 30.826 96.738 ;
               RECT 30.774 97.302 30.826 97.338 ;
               RECT 30.774 97.902 30.826 97.938 ;
               RECT 30.774 98.502 30.826 98.538 ;
               RECT 30.774 99.102 30.826 99.138 ;
               RECT 30.774 99.702 30.826 99.738 ;
               RECT 30.774 100.302 30.826 100.338 ;
               RECT 30.774 100.902 30.826 100.938 ;
               RECT 30.774 101.502 30.826 101.538 ;
               RECT 30.774 102.102 30.826 102.138 ;
               RECT 30.774 102.702 30.826 102.738 ;
               RECT 30.774 103.302 30.826 103.338 ;
               RECT 30.774 103.902 30.826 103.938 ;
               RECT 30.774 104.502 30.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 31.574 0.5695 31.626 104.5505 ;
               LAYER v4 ;
               RECT 31.574 0.582 31.626 0.618 ;
               RECT 31.574 1.182 31.626 1.218 ;
               RECT 31.574 1.782 31.626 1.818 ;
               RECT 31.574 2.382 31.626 2.418 ;
               RECT 31.574 2.982 31.626 3.018 ;
               RECT 31.574 3.582 31.626 3.618 ;
               RECT 31.574 4.182 31.626 4.218 ;
               RECT 31.574 4.782 31.626 4.818 ;
               RECT 31.574 5.382 31.626 5.418 ;
               RECT 31.574 5.982 31.626 6.018 ;
               RECT 31.574 6.582 31.626 6.618 ;
               RECT 31.574 7.182 31.626 7.218 ;
               RECT 31.574 7.782 31.626 7.818 ;
               RECT 31.574 8.382 31.626 8.418 ;
               RECT 31.574 8.982 31.626 9.018 ;
               RECT 31.574 9.582 31.626 9.618 ;
               RECT 31.574 10.182 31.626 10.218 ;
               RECT 31.574 10.782 31.626 10.818 ;
               RECT 31.574 11.382 31.626 11.418 ;
               RECT 31.574 11.982 31.626 12.018 ;
               RECT 31.574 12.582 31.626 12.618 ;
               RECT 31.574 13.182 31.626 13.218 ;
               RECT 31.574 13.782 31.626 13.818 ;
               RECT 31.574 14.382 31.626 14.418 ;
               RECT 31.574 14.982 31.626 15.018 ;
               RECT 31.574 15.582 31.626 15.618 ;
               RECT 31.574 16.182 31.626 16.218 ;
               RECT 31.574 16.782 31.626 16.818 ;
               RECT 31.574 17.382 31.626 17.418 ;
               RECT 31.574 17.982 31.626 18.018 ;
               RECT 31.574 18.582 31.626 18.618 ;
               RECT 31.574 19.182 31.626 19.218 ;
               RECT 31.574 19.782 31.626 19.818 ;
               RECT 31.574 20.382 31.626 20.418 ;
               RECT 31.574 20.982 31.626 21.018 ;
               RECT 31.574 21.582 31.626 21.618 ;
               RECT 31.574 22.182 31.626 22.218 ;
               RECT 31.574 22.782 31.626 22.818 ;
               RECT 31.574 23.382 31.626 23.418 ;
               RECT 31.574 23.982 31.626 24.018 ;
               RECT 31.574 24.582 31.626 24.618 ;
               RECT 31.574 25.182 31.626 25.218 ;
               RECT 31.574 25.782 31.626 25.818 ;
               RECT 31.574 26.382 31.626 26.418 ;
               RECT 31.574 26.982 31.626 27.018 ;
               RECT 31.574 27.582 31.626 27.618 ;
               RECT 31.574 28.182 31.626 28.218 ;
               RECT 31.574 28.782 31.626 28.818 ;
               RECT 31.574 29.382 31.626 29.418 ;
               RECT 31.574 29.982 31.626 30.018 ;
               RECT 31.574 30.582 31.626 30.618 ;
               RECT 31.574 31.182 31.626 31.218 ;
               RECT 31.574 31.782 31.626 31.818 ;
               RECT 31.574 32.382 31.626 32.418 ;
               RECT 31.574 32.982 31.626 33.018 ;
               RECT 31.574 33.582 31.626 33.618 ;
               RECT 31.574 34.182 31.626 34.218 ;
               RECT 31.574 34.782 31.626 34.818 ;
               RECT 31.574 35.382 31.626 35.418 ;
               RECT 31.574 35.982 31.626 36.018 ;
               RECT 31.574 36.582 31.626 36.618 ;
               RECT 31.574 37.182 31.626 37.218 ;
               RECT 31.574 37.782 31.626 37.818 ;
               RECT 31.574 38.382 31.626 38.418 ;
               RECT 31.574 38.982 31.626 39.018 ;
               RECT 31.574 39.582 31.626 39.618 ;
               RECT 31.574 40.182 31.626 40.218 ;
               RECT 31.574 40.782 31.626 40.818 ;
               RECT 31.574 41.382 31.626 41.418 ;
               RECT 31.574 41.982 31.626 42.018 ;
               RECT 31.574 42.582 31.626 42.618 ;
               RECT 31.574 43.182 31.626 43.218 ;
               RECT 31.574 43.782 31.626 43.818 ;
               RECT 31.574 44.382 31.626 44.418 ;
               RECT 31.574 44.982 31.626 45.018 ;
               RECT 31.574 45.582 31.626 45.618 ;
               RECT 31.574 46.182 31.626 46.218 ;
               RECT 31.574 46.782 31.626 46.818 ;
               RECT 31.574 47.382 31.626 47.418 ;
               RECT 31.574 47.982 31.626 48.018 ;
               RECT 31.574 48.582 31.626 48.618 ;
               RECT 31.574 48.942 31.626 48.978 ;
               RECT 31.574 49.182 31.626 49.218 ;
               RECT 31.574 49.902 31.626 49.938 ;
               RECT 31.574 50.622 31.626 50.658 ;
               RECT 31.574 50.862 31.626 50.898 ;
               RECT 31.574 51.342 31.626 51.378 ;
               RECT 31.574 51.822 31.626 51.858 ;
               RECT 31.574 52.302 31.626 52.338 ;
               RECT 31.574 52.782 31.626 52.818 ;
               RECT 31.574 53.262 31.626 53.298 ;
               RECT 31.574 53.742 31.626 53.778 ;
               RECT 31.574 54.222 31.626 54.258 ;
               RECT 31.574 54.462 31.626 54.498 ;
               RECT 31.574 55.182 31.626 55.218 ;
               RECT 31.574 55.902 31.626 55.938 ;
               RECT 31.574 56.142 31.626 56.178 ;
               RECT 31.574 56.502 31.626 56.538 ;
               RECT 31.574 57.102 31.626 57.138 ;
               RECT 31.574 57.702 31.626 57.738 ;
               RECT 31.574 58.302 31.626 58.338 ;
               RECT 31.574 58.902 31.626 58.938 ;
               RECT 31.574 59.502 31.626 59.538 ;
               RECT 31.574 60.102 31.626 60.138 ;
               RECT 31.574 60.702 31.626 60.738 ;
               RECT 31.574 61.302 31.626 61.338 ;
               RECT 31.574 61.902 31.626 61.938 ;
               RECT 31.574 62.502 31.626 62.538 ;
               RECT 31.574 63.102 31.626 63.138 ;
               RECT 31.574 63.702 31.626 63.738 ;
               RECT 31.574 64.302 31.626 64.338 ;
               RECT 31.574 64.902 31.626 64.938 ;
               RECT 31.574 65.502 31.626 65.538 ;
               RECT 31.574 66.102 31.626 66.138 ;
               RECT 31.574 66.702 31.626 66.738 ;
               RECT 31.574 67.302 31.626 67.338 ;
               RECT 31.574 67.902 31.626 67.938 ;
               RECT 31.574 68.502 31.626 68.538 ;
               RECT 31.574 69.102 31.626 69.138 ;
               RECT 31.574 69.702 31.626 69.738 ;
               RECT 31.574 70.302 31.626 70.338 ;
               RECT 31.574 70.902 31.626 70.938 ;
               RECT 31.574 71.502 31.626 71.538 ;
               RECT 31.574 72.102 31.626 72.138 ;
               RECT 31.574 72.702 31.626 72.738 ;
               RECT 31.574 73.302 31.626 73.338 ;
               RECT 31.574 73.902 31.626 73.938 ;
               RECT 31.574 74.502 31.626 74.538 ;
               RECT 31.574 75.102 31.626 75.138 ;
               RECT 31.574 75.702 31.626 75.738 ;
               RECT 31.574 76.302 31.626 76.338 ;
               RECT 31.574 76.902 31.626 76.938 ;
               RECT 31.574 77.502 31.626 77.538 ;
               RECT 31.574 78.102 31.626 78.138 ;
               RECT 31.574 78.702 31.626 78.738 ;
               RECT 31.574 79.302 31.626 79.338 ;
               RECT 31.574 79.902 31.626 79.938 ;
               RECT 31.574 80.502 31.626 80.538 ;
               RECT 31.574 81.102 31.626 81.138 ;
               RECT 31.574 81.702 31.626 81.738 ;
               RECT 31.574 82.302 31.626 82.338 ;
               RECT 31.574 82.902 31.626 82.938 ;
               RECT 31.574 83.502 31.626 83.538 ;
               RECT 31.574 84.102 31.626 84.138 ;
               RECT 31.574 84.702 31.626 84.738 ;
               RECT 31.574 85.302 31.626 85.338 ;
               RECT 31.574 85.902 31.626 85.938 ;
               RECT 31.574 86.502 31.626 86.538 ;
               RECT 31.574 87.102 31.626 87.138 ;
               RECT 31.574 87.702 31.626 87.738 ;
               RECT 31.574 88.302 31.626 88.338 ;
               RECT 31.574 88.902 31.626 88.938 ;
               RECT 31.574 89.502 31.626 89.538 ;
               RECT 31.574 90.102 31.626 90.138 ;
               RECT 31.574 90.702 31.626 90.738 ;
               RECT 31.574 91.302 31.626 91.338 ;
               RECT 31.574 91.902 31.626 91.938 ;
               RECT 31.574 92.502 31.626 92.538 ;
               RECT 31.574 93.102 31.626 93.138 ;
               RECT 31.574 93.702 31.626 93.738 ;
               RECT 31.574 94.302 31.626 94.338 ;
               RECT 31.574 94.902 31.626 94.938 ;
               RECT 31.574 95.502 31.626 95.538 ;
               RECT 31.574 96.102 31.626 96.138 ;
               RECT 31.574 96.702 31.626 96.738 ;
               RECT 31.574 97.302 31.626 97.338 ;
               RECT 31.574 97.902 31.626 97.938 ;
               RECT 31.574 98.502 31.626 98.538 ;
               RECT 31.574 99.102 31.626 99.138 ;
               RECT 31.574 99.702 31.626 99.738 ;
               RECT 31.574 100.302 31.626 100.338 ;
               RECT 31.574 100.902 31.626 100.938 ;
               RECT 31.574 101.502 31.626 101.538 ;
               RECT 31.574 102.102 31.626 102.138 ;
               RECT 31.574 102.702 31.626 102.738 ;
               RECT 31.574 103.302 31.626 103.338 ;
               RECT 31.574 103.902 31.626 103.938 ;
               RECT 31.574 104.502 31.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 32.374 0.5695 32.426 104.5505 ;
               LAYER v4 ;
               RECT 32.374 0.582 32.426 0.618 ;
               RECT 32.374 1.182 32.426 1.218 ;
               RECT 32.374 1.782 32.426 1.818 ;
               RECT 32.374 2.382 32.426 2.418 ;
               RECT 32.374 2.982 32.426 3.018 ;
               RECT 32.374 3.582 32.426 3.618 ;
               RECT 32.374 4.182 32.426 4.218 ;
               RECT 32.374 4.782 32.426 4.818 ;
               RECT 32.374 5.382 32.426 5.418 ;
               RECT 32.374 5.982 32.426 6.018 ;
               RECT 32.374 6.582 32.426 6.618 ;
               RECT 32.374 7.182 32.426 7.218 ;
               RECT 32.374 7.782 32.426 7.818 ;
               RECT 32.374 8.382 32.426 8.418 ;
               RECT 32.374 8.982 32.426 9.018 ;
               RECT 32.374 9.582 32.426 9.618 ;
               RECT 32.374 10.182 32.426 10.218 ;
               RECT 32.374 10.782 32.426 10.818 ;
               RECT 32.374 11.382 32.426 11.418 ;
               RECT 32.374 11.982 32.426 12.018 ;
               RECT 32.374 12.582 32.426 12.618 ;
               RECT 32.374 13.182 32.426 13.218 ;
               RECT 32.374 13.782 32.426 13.818 ;
               RECT 32.374 14.382 32.426 14.418 ;
               RECT 32.374 14.982 32.426 15.018 ;
               RECT 32.374 15.582 32.426 15.618 ;
               RECT 32.374 16.182 32.426 16.218 ;
               RECT 32.374 16.782 32.426 16.818 ;
               RECT 32.374 17.382 32.426 17.418 ;
               RECT 32.374 17.982 32.426 18.018 ;
               RECT 32.374 18.582 32.426 18.618 ;
               RECT 32.374 19.182 32.426 19.218 ;
               RECT 32.374 19.782 32.426 19.818 ;
               RECT 32.374 20.382 32.426 20.418 ;
               RECT 32.374 20.982 32.426 21.018 ;
               RECT 32.374 21.582 32.426 21.618 ;
               RECT 32.374 22.182 32.426 22.218 ;
               RECT 32.374 22.782 32.426 22.818 ;
               RECT 32.374 23.382 32.426 23.418 ;
               RECT 32.374 23.982 32.426 24.018 ;
               RECT 32.374 24.582 32.426 24.618 ;
               RECT 32.374 25.182 32.426 25.218 ;
               RECT 32.374 25.782 32.426 25.818 ;
               RECT 32.374 26.382 32.426 26.418 ;
               RECT 32.374 26.982 32.426 27.018 ;
               RECT 32.374 27.582 32.426 27.618 ;
               RECT 32.374 28.182 32.426 28.218 ;
               RECT 32.374 28.782 32.426 28.818 ;
               RECT 32.374 29.382 32.426 29.418 ;
               RECT 32.374 29.982 32.426 30.018 ;
               RECT 32.374 30.582 32.426 30.618 ;
               RECT 32.374 31.182 32.426 31.218 ;
               RECT 32.374 31.782 32.426 31.818 ;
               RECT 32.374 32.382 32.426 32.418 ;
               RECT 32.374 32.982 32.426 33.018 ;
               RECT 32.374 33.582 32.426 33.618 ;
               RECT 32.374 34.182 32.426 34.218 ;
               RECT 32.374 34.782 32.426 34.818 ;
               RECT 32.374 35.382 32.426 35.418 ;
               RECT 32.374 35.982 32.426 36.018 ;
               RECT 32.374 36.582 32.426 36.618 ;
               RECT 32.374 37.182 32.426 37.218 ;
               RECT 32.374 37.782 32.426 37.818 ;
               RECT 32.374 38.382 32.426 38.418 ;
               RECT 32.374 38.982 32.426 39.018 ;
               RECT 32.374 39.582 32.426 39.618 ;
               RECT 32.374 40.182 32.426 40.218 ;
               RECT 32.374 40.782 32.426 40.818 ;
               RECT 32.374 41.382 32.426 41.418 ;
               RECT 32.374 41.982 32.426 42.018 ;
               RECT 32.374 42.582 32.426 42.618 ;
               RECT 32.374 43.182 32.426 43.218 ;
               RECT 32.374 43.782 32.426 43.818 ;
               RECT 32.374 44.382 32.426 44.418 ;
               RECT 32.374 44.982 32.426 45.018 ;
               RECT 32.374 45.582 32.426 45.618 ;
               RECT 32.374 46.182 32.426 46.218 ;
               RECT 32.374 46.782 32.426 46.818 ;
               RECT 32.374 47.382 32.426 47.418 ;
               RECT 32.374 47.982 32.426 48.018 ;
               RECT 32.374 48.582 32.426 48.618 ;
               RECT 32.374 48.942 32.426 48.978 ;
               RECT 32.374 48.9475 32.426 48.9725 ;
               RECT 32.374 49.182 32.426 49.218 ;
               RECT 32.374 49.902 32.426 49.938 ;
               RECT 32.374 50.622 32.426 50.658 ;
               RECT 32.374 50.862 32.426 50.898 ;
               RECT 32.374 51.342 32.426 51.378 ;
               RECT 32.374 51.822 32.426 51.858 ;
               RECT 32.374 52.302 32.426 52.338 ;
               RECT 32.374 52.782 32.426 52.818 ;
               RECT 32.374 53.262 32.426 53.298 ;
               RECT 32.374 53.742 32.426 53.778 ;
               RECT 32.374 54.222 32.426 54.258 ;
               RECT 32.374 54.462 32.426 54.498 ;
               RECT 32.374 55.182 32.426 55.218 ;
               RECT 32.374 55.902 32.426 55.938 ;
               RECT 32.374 56.142 32.426 56.178 ;
               RECT 32.374 56.1475 32.426 56.1725 ;
               RECT 32.374 56.502 32.426 56.538 ;
               RECT 32.374 57.102 32.426 57.138 ;
               RECT 32.374 57.702 32.426 57.738 ;
               RECT 32.374 58.302 32.426 58.338 ;
               RECT 32.374 58.902 32.426 58.938 ;
               RECT 32.374 59.502 32.426 59.538 ;
               RECT 32.374 60.102 32.426 60.138 ;
               RECT 32.374 60.702 32.426 60.738 ;
               RECT 32.374 61.302 32.426 61.338 ;
               RECT 32.374 61.902 32.426 61.938 ;
               RECT 32.374 62.502 32.426 62.538 ;
               RECT 32.374 63.102 32.426 63.138 ;
               RECT 32.374 63.702 32.426 63.738 ;
               RECT 32.374 64.302 32.426 64.338 ;
               RECT 32.374 64.902 32.426 64.938 ;
               RECT 32.374 65.502 32.426 65.538 ;
               RECT 32.374 66.102 32.426 66.138 ;
               RECT 32.374 66.702 32.426 66.738 ;
               RECT 32.374 67.302 32.426 67.338 ;
               RECT 32.374 67.902 32.426 67.938 ;
               RECT 32.374 68.502 32.426 68.538 ;
               RECT 32.374 69.102 32.426 69.138 ;
               RECT 32.374 69.702 32.426 69.738 ;
               RECT 32.374 70.302 32.426 70.338 ;
               RECT 32.374 70.902 32.426 70.938 ;
               RECT 32.374 71.502 32.426 71.538 ;
               RECT 32.374 72.102 32.426 72.138 ;
               RECT 32.374 72.702 32.426 72.738 ;
               RECT 32.374 73.302 32.426 73.338 ;
               RECT 32.374 73.902 32.426 73.938 ;
               RECT 32.374 74.502 32.426 74.538 ;
               RECT 32.374 75.102 32.426 75.138 ;
               RECT 32.374 75.702 32.426 75.738 ;
               RECT 32.374 76.302 32.426 76.338 ;
               RECT 32.374 76.902 32.426 76.938 ;
               RECT 32.374 77.502 32.426 77.538 ;
               RECT 32.374 78.102 32.426 78.138 ;
               RECT 32.374 78.702 32.426 78.738 ;
               RECT 32.374 79.302 32.426 79.338 ;
               RECT 32.374 79.902 32.426 79.938 ;
               RECT 32.374 80.502 32.426 80.538 ;
               RECT 32.374 81.102 32.426 81.138 ;
               RECT 32.374 81.702 32.426 81.738 ;
               RECT 32.374 82.302 32.426 82.338 ;
               RECT 32.374 82.902 32.426 82.938 ;
               RECT 32.374 83.502 32.426 83.538 ;
               RECT 32.374 84.102 32.426 84.138 ;
               RECT 32.374 84.702 32.426 84.738 ;
               RECT 32.374 85.302 32.426 85.338 ;
               RECT 32.374 85.902 32.426 85.938 ;
               RECT 32.374 86.502 32.426 86.538 ;
               RECT 32.374 87.102 32.426 87.138 ;
               RECT 32.374 87.702 32.426 87.738 ;
               RECT 32.374 88.302 32.426 88.338 ;
               RECT 32.374 88.902 32.426 88.938 ;
               RECT 32.374 89.502 32.426 89.538 ;
               RECT 32.374 90.102 32.426 90.138 ;
               RECT 32.374 90.702 32.426 90.738 ;
               RECT 32.374 91.302 32.426 91.338 ;
               RECT 32.374 91.902 32.426 91.938 ;
               RECT 32.374 92.502 32.426 92.538 ;
               RECT 32.374 93.102 32.426 93.138 ;
               RECT 32.374 93.702 32.426 93.738 ;
               RECT 32.374 94.302 32.426 94.338 ;
               RECT 32.374 94.902 32.426 94.938 ;
               RECT 32.374 95.502 32.426 95.538 ;
               RECT 32.374 96.102 32.426 96.138 ;
               RECT 32.374 96.702 32.426 96.738 ;
               RECT 32.374 97.302 32.426 97.338 ;
               RECT 32.374 97.902 32.426 97.938 ;
               RECT 32.374 98.502 32.426 98.538 ;
               RECT 32.374 99.102 32.426 99.138 ;
               RECT 32.374 99.702 32.426 99.738 ;
               RECT 32.374 100.302 32.426 100.338 ;
               RECT 32.374 100.902 32.426 100.938 ;
               RECT 32.374 101.502 32.426 101.538 ;
               RECT 32.374 102.102 32.426 102.138 ;
               RECT 32.374 102.702 32.426 102.738 ;
               RECT 32.374 103.302 32.426 103.338 ;
               RECT 32.374 103.902 32.426 103.938 ;
               RECT 32.374 104.502 32.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 33.174 0.5695 33.226 104.5505 ;
               LAYER v4 ;
               RECT 33.174 0.582 33.226 0.618 ;
               RECT 33.174 1.182 33.226 1.218 ;
               RECT 33.174 1.782 33.226 1.818 ;
               RECT 33.174 2.382 33.226 2.418 ;
               RECT 33.174 2.982 33.226 3.018 ;
               RECT 33.174 3.582 33.226 3.618 ;
               RECT 33.174 4.182 33.226 4.218 ;
               RECT 33.174 4.782 33.226 4.818 ;
               RECT 33.174 5.382 33.226 5.418 ;
               RECT 33.174 5.982 33.226 6.018 ;
               RECT 33.174 6.582 33.226 6.618 ;
               RECT 33.174 7.182 33.226 7.218 ;
               RECT 33.174 7.782 33.226 7.818 ;
               RECT 33.174 8.382 33.226 8.418 ;
               RECT 33.174 8.982 33.226 9.018 ;
               RECT 33.174 9.582 33.226 9.618 ;
               RECT 33.174 10.182 33.226 10.218 ;
               RECT 33.174 10.782 33.226 10.818 ;
               RECT 33.174 11.382 33.226 11.418 ;
               RECT 33.174 11.982 33.226 12.018 ;
               RECT 33.174 12.582 33.226 12.618 ;
               RECT 33.174 13.182 33.226 13.218 ;
               RECT 33.174 13.782 33.226 13.818 ;
               RECT 33.174 14.382 33.226 14.418 ;
               RECT 33.174 14.982 33.226 15.018 ;
               RECT 33.174 15.582 33.226 15.618 ;
               RECT 33.174 16.182 33.226 16.218 ;
               RECT 33.174 16.782 33.226 16.818 ;
               RECT 33.174 17.382 33.226 17.418 ;
               RECT 33.174 17.982 33.226 18.018 ;
               RECT 33.174 18.582 33.226 18.618 ;
               RECT 33.174 19.182 33.226 19.218 ;
               RECT 33.174 19.782 33.226 19.818 ;
               RECT 33.174 20.382 33.226 20.418 ;
               RECT 33.174 20.982 33.226 21.018 ;
               RECT 33.174 21.582 33.226 21.618 ;
               RECT 33.174 22.182 33.226 22.218 ;
               RECT 33.174 22.782 33.226 22.818 ;
               RECT 33.174 23.382 33.226 23.418 ;
               RECT 33.174 23.982 33.226 24.018 ;
               RECT 33.174 24.582 33.226 24.618 ;
               RECT 33.174 25.182 33.226 25.218 ;
               RECT 33.174 25.782 33.226 25.818 ;
               RECT 33.174 26.382 33.226 26.418 ;
               RECT 33.174 26.982 33.226 27.018 ;
               RECT 33.174 27.582 33.226 27.618 ;
               RECT 33.174 28.182 33.226 28.218 ;
               RECT 33.174 28.782 33.226 28.818 ;
               RECT 33.174 29.382 33.226 29.418 ;
               RECT 33.174 29.982 33.226 30.018 ;
               RECT 33.174 30.582 33.226 30.618 ;
               RECT 33.174 31.182 33.226 31.218 ;
               RECT 33.174 31.782 33.226 31.818 ;
               RECT 33.174 32.382 33.226 32.418 ;
               RECT 33.174 32.982 33.226 33.018 ;
               RECT 33.174 33.582 33.226 33.618 ;
               RECT 33.174 34.182 33.226 34.218 ;
               RECT 33.174 34.782 33.226 34.818 ;
               RECT 33.174 35.382 33.226 35.418 ;
               RECT 33.174 35.982 33.226 36.018 ;
               RECT 33.174 36.582 33.226 36.618 ;
               RECT 33.174 37.182 33.226 37.218 ;
               RECT 33.174 37.782 33.226 37.818 ;
               RECT 33.174 38.382 33.226 38.418 ;
               RECT 33.174 38.982 33.226 39.018 ;
               RECT 33.174 39.582 33.226 39.618 ;
               RECT 33.174 40.182 33.226 40.218 ;
               RECT 33.174 40.782 33.226 40.818 ;
               RECT 33.174 41.382 33.226 41.418 ;
               RECT 33.174 41.982 33.226 42.018 ;
               RECT 33.174 42.582 33.226 42.618 ;
               RECT 33.174 43.182 33.226 43.218 ;
               RECT 33.174 43.782 33.226 43.818 ;
               RECT 33.174 44.382 33.226 44.418 ;
               RECT 33.174 44.982 33.226 45.018 ;
               RECT 33.174 45.582 33.226 45.618 ;
               RECT 33.174 46.182 33.226 46.218 ;
               RECT 33.174 46.782 33.226 46.818 ;
               RECT 33.174 47.382 33.226 47.418 ;
               RECT 33.174 47.982 33.226 48.018 ;
               RECT 33.174 48.582 33.226 48.618 ;
               RECT 33.174 48.942 33.226 48.978 ;
               RECT 33.174 49.182 33.226 49.218 ;
               RECT 33.174 49.902 33.226 49.938 ;
               RECT 33.174 50.622 33.226 50.658 ;
               RECT 33.174 50.862 33.226 50.898 ;
               RECT 33.174 51.342 33.226 51.378 ;
               RECT 33.174 51.822 33.226 51.858 ;
               RECT 33.174 52.302 33.226 52.338 ;
               RECT 33.174 52.782 33.226 52.818 ;
               RECT 33.174 53.262 33.226 53.298 ;
               RECT 33.174 53.742 33.226 53.778 ;
               RECT 33.174 54.222 33.226 54.258 ;
               RECT 33.174 54.462 33.226 54.498 ;
               RECT 33.174 55.182 33.226 55.218 ;
               RECT 33.174 55.902 33.226 55.938 ;
               RECT 33.174 56.142 33.226 56.178 ;
               RECT 33.174 56.502 33.226 56.538 ;
               RECT 33.174 57.102 33.226 57.138 ;
               RECT 33.174 57.702 33.226 57.738 ;
               RECT 33.174 58.302 33.226 58.338 ;
               RECT 33.174 58.902 33.226 58.938 ;
               RECT 33.174 59.502 33.226 59.538 ;
               RECT 33.174 60.102 33.226 60.138 ;
               RECT 33.174 60.702 33.226 60.738 ;
               RECT 33.174 61.302 33.226 61.338 ;
               RECT 33.174 61.902 33.226 61.938 ;
               RECT 33.174 62.502 33.226 62.538 ;
               RECT 33.174 63.102 33.226 63.138 ;
               RECT 33.174 63.702 33.226 63.738 ;
               RECT 33.174 64.302 33.226 64.338 ;
               RECT 33.174 64.902 33.226 64.938 ;
               RECT 33.174 65.502 33.226 65.538 ;
               RECT 33.174 66.102 33.226 66.138 ;
               RECT 33.174 66.702 33.226 66.738 ;
               RECT 33.174 67.302 33.226 67.338 ;
               RECT 33.174 67.902 33.226 67.938 ;
               RECT 33.174 68.502 33.226 68.538 ;
               RECT 33.174 69.102 33.226 69.138 ;
               RECT 33.174 69.702 33.226 69.738 ;
               RECT 33.174 70.302 33.226 70.338 ;
               RECT 33.174 70.902 33.226 70.938 ;
               RECT 33.174 71.502 33.226 71.538 ;
               RECT 33.174 72.102 33.226 72.138 ;
               RECT 33.174 72.702 33.226 72.738 ;
               RECT 33.174 73.302 33.226 73.338 ;
               RECT 33.174 73.902 33.226 73.938 ;
               RECT 33.174 74.502 33.226 74.538 ;
               RECT 33.174 75.102 33.226 75.138 ;
               RECT 33.174 75.702 33.226 75.738 ;
               RECT 33.174 76.302 33.226 76.338 ;
               RECT 33.174 76.902 33.226 76.938 ;
               RECT 33.174 77.502 33.226 77.538 ;
               RECT 33.174 78.102 33.226 78.138 ;
               RECT 33.174 78.702 33.226 78.738 ;
               RECT 33.174 79.302 33.226 79.338 ;
               RECT 33.174 79.902 33.226 79.938 ;
               RECT 33.174 80.502 33.226 80.538 ;
               RECT 33.174 81.102 33.226 81.138 ;
               RECT 33.174 81.702 33.226 81.738 ;
               RECT 33.174 82.302 33.226 82.338 ;
               RECT 33.174 82.902 33.226 82.938 ;
               RECT 33.174 83.502 33.226 83.538 ;
               RECT 33.174 84.102 33.226 84.138 ;
               RECT 33.174 84.702 33.226 84.738 ;
               RECT 33.174 85.302 33.226 85.338 ;
               RECT 33.174 85.902 33.226 85.938 ;
               RECT 33.174 86.502 33.226 86.538 ;
               RECT 33.174 87.102 33.226 87.138 ;
               RECT 33.174 87.702 33.226 87.738 ;
               RECT 33.174 88.302 33.226 88.338 ;
               RECT 33.174 88.902 33.226 88.938 ;
               RECT 33.174 89.502 33.226 89.538 ;
               RECT 33.174 90.102 33.226 90.138 ;
               RECT 33.174 90.702 33.226 90.738 ;
               RECT 33.174 91.302 33.226 91.338 ;
               RECT 33.174 91.902 33.226 91.938 ;
               RECT 33.174 92.502 33.226 92.538 ;
               RECT 33.174 93.102 33.226 93.138 ;
               RECT 33.174 93.702 33.226 93.738 ;
               RECT 33.174 94.302 33.226 94.338 ;
               RECT 33.174 94.902 33.226 94.938 ;
               RECT 33.174 95.502 33.226 95.538 ;
               RECT 33.174 96.102 33.226 96.138 ;
               RECT 33.174 96.702 33.226 96.738 ;
               RECT 33.174 97.302 33.226 97.338 ;
               RECT 33.174 97.902 33.226 97.938 ;
               RECT 33.174 98.502 33.226 98.538 ;
               RECT 33.174 99.102 33.226 99.138 ;
               RECT 33.174 99.702 33.226 99.738 ;
               RECT 33.174 100.302 33.226 100.338 ;
               RECT 33.174 100.902 33.226 100.938 ;
               RECT 33.174 101.502 33.226 101.538 ;
               RECT 33.174 102.102 33.226 102.138 ;
               RECT 33.174 102.702 33.226 102.738 ;
               RECT 33.174 103.302 33.226 103.338 ;
               RECT 33.174 103.902 33.226 103.938 ;
               RECT 33.174 104.502 33.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 33.974 0.5695 34.026 104.5505 ;
               LAYER v4 ;
               RECT 33.974 0.582 34.026 0.618 ;
               RECT 33.974 1.182 34.026 1.218 ;
               RECT 33.974 1.782 34.026 1.818 ;
               RECT 33.974 2.382 34.026 2.418 ;
               RECT 33.974 2.982 34.026 3.018 ;
               RECT 33.974 3.582 34.026 3.618 ;
               RECT 33.974 4.182 34.026 4.218 ;
               RECT 33.974 4.782 34.026 4.818 ;
               RECT 33.974 5.382 34.026 5.418 ;
               RECT 33.974 5.982 34.026 6.018 ;
               RECT 33.974 6.582 34.026 6.618 ;
               RECT 33.974 7.182 34.026 7.218 ;
               RECT 33.974 7.782 34.026 7.818 ;
               RECT 33.974 8.382 34.026 8.418 ;
               RECT 33.974 8.982 34.026 9.018 ;
               RECT 33.974 9.582 34.026 9.618 ;
               RECT 33.974 10.182 34.026 10.218 ;
               RECT 33.974 10.782 34.026 10.818 ;
               RECT 33.974 11.382 34.026 11.418 ;
               RECT 33.974 11.982 34.026 12.018 ;
               RECT 33.974 12.582 34.026 12.618 ;
               RECT 33.974 13.182 34.026 13.218 ;
               RECT 33.974 13.782 34.026 13.818 ;
               RECT 33.974 14.382 34.026 14.418 ;
               RECT 33.974 14.982 34.026 15.018 ;
               RECT 33.974 15.582 34.026 15.618 ;
               RECT 33.974 16.182 34.026 16.218 ;
               RECT 33.974 16.782 34.026 16.818 ;
               RECT 33.974 17.382 34.026 17.418 ;
               RECT 33.974 17.982 34.026 18.018 ;
               RECT 33.974 18.582 34.026 18.618 ;
               RECT 33.974 19.182 34.026 19.218 ;
               RECT 33.974 19.782 34.026 19.818 ;
               RECT 33.974 20.382 34.026 20.418 ;
               RECT 33.974 20.982 34.026 21.018 ;
               RECT 33.974 21.582 34.026 21.618 ;
               RECT 33.974 22.182 34.026 22.218 ;
               RECT 33.974 22.782 34.026 22.818 ;
               RECT 33.974 23.382 34.026 23.418 ;
               RECT 33.974 23.982 34.026 24.018 ;
               RECT 33.974 24.582 34.026 24.618 ;
               RECT 33.974 25.182 34.026 25.218 ;
               RECT 33.974 25.782 34.026 25.818 ;
               RECT 33.974 26.382 34.026 26.418 ;
               RECT 33.974 26.982 34.026 27.018 ;
               RECT 33.974 27.582 34.026 27.618 ;
               RECT 33.974 28.182 34.026 28.218 ;
               RECT 33.974 28.782 34.026 28.818 ;
               RECT 33.974 29.382 34.026 29.418 ;
               RECT 33.974 29.982 34.026 30.018 ;
               RECT 33.974 30.582 34.026 30.618 ;
               RECT 33.974 31.182 34.026 31.218 ;
               RECT 33.974 31.782 34.026 31.818 ;
               RECT 33.974 32.382 34.026 32.418 ;
               RECT 33.974 32.982 34.026 33.018 ;
               RECT 33.974 33.582 34.026 33.618 ;
               RECT 33.974 34.182 34.026 34.218 ;
               RECT 33.974 34.782 34.026 34.818 ;
               RECT 33.974 35.382 34.026 35.418 ;
               RECT 33.974 35.982 34.026 36.018 ;
               RECT 33.974 36.582 34.026 36.618 ;
               RECT 33.974 37.182 34.026 37.218 ;
               RECT 33.974 37.782 34.026 37.818 ;
               RECT 33.974 38.382 34.026 38.418 ;
               RECT 33.974 38.982 34.026 39.018 ;
               RECT 33.974 39.582 34.026 39.618 ;
               RECT 33.974 40.182 34.026 40.218 ;
               RECT 33.974 40.782 34.026 40.818 ;
               RECT 33.974 41.382 34.026 41.418 ;
               RECT 33.974 41.982 34.026 42.018 ;
               RECT 33.974 42.582 34.026 42.618 ;
               RECT 33.974 43.182 34.026 43.218 ;
               RECT 33.974 43.782 34.026 43.818 ;
               RECT 33.974 44.382 34.026 44.418 ;
               RECT 33.974 44.982 34.026 45.018 ;
               RECT 33.974 45.582 34.026 45.618 ;
               RECT 33.974 46.182 34.026 46.218 ;
               RECT 33.974 46.782 34.026 46.818 ;
               RECT 33.974 47.382 34.026 47.418 ;
               RECT 33.974 47.982 34.026 48.018 ;
               RECT 33.974 48.582 34.026 48.618 ;
               RECT 33.974 48.942 34.026 48.978 ;
               RECT 33.974 48.9475 34.026 48.9725 ;
               RECT 33.974 49.182 34.026 49.218 ;
               RECT 33.974 49.902 34.026 49.938 ;
               RECT 33.974 50.622 34.026 50.658 ;
               RECT 33.974 50.862 34.026 50.898 ;
               RECT 33.974 51.342 34.026 51.378 ;
               RECT 33.974 51.822 34.026 51.858 ;
               RECT 33.974 52.302 34.026 52.338 ;
               RECT 33.974 52.782 34.026 52.818 ;
               RECT 33.974 53.262 34.026 53.298 ;
               RECT 33.974 53.742 34.026 53.778 ;
               RECT 33.974 54.222 34.026 54.258 ;
               RECT 33.974 54.462 34.026 54.498 ;
               RECT 33.974 55.182 34.026 55.218 ;
               RECT 33.974 55.902 34.026 55.938 ;
               RECT 33.974 56.142 34.026 56.178 ;
               RECT 33.974 56.1475 34.026 56.1725 ;
               RECT 33.974 56.502 34.026 56.538 ;
               RECT 33.974 57.102 34.026 57.138 ;
               RECT 33.974 57.702 34.026 57.738 ;
               RECT 33.974 58.302 34.026 58.338 ;
               RECT 33.974 58.902 34.026 58.938 ;
               RECT 33.974 59.502 34.026 59.538 ;
               RECT 33.974 60.102 34.026 60.138 ;
               RECT 33.974 60.702 34.026 60.738 ;
               RECT 33.974 61.302 34.026 61.338 ;
               RECT 33.974 61.902 34.026 61.938 ;
               RECT 33.974 62.502 34.026 62.538 ;
               RECT 33.974 63.102 34.026 63.138 ;
               RECT 33.974 63.702 34.026 63.738 ;
               RECT 33.974 64.302 34.026 64.338 ;
               RECT 33.974 64.902 34.026 64.938 ;
               RECT 33.974 65.502 34.026 65.538 ;
               RECT 33.974 66.102 34.026 66.138 ;
               RECT 33.974 66.702 34.026 66.738 ;
               RECT 33.974 67.302 34.026 67.338 ;
               RECT 33.974 67.902 34.026 67.938 ;
               RECT 33.974 68.502 34.026 68.538 ;
               RECT 33.974 69.102 34.026 69.138 ;
               RECT 33.974 69.702 34.026 69.738 ;
               RECT 33.974 70.302 34.026 70.338 ;
               RECT 33.974 70.902 34.026 70.938 ;
               RECT 33.974 71.502 34.026 71.538 ;
               RECT 33.974 72.102 34.026 72.138 ;
               RECT 33.974 72.702 34.026 72.738 ;
               RECT 33.974 73.302 34.026 73.338 ;
               RECT 33.974 73.902 34.026 73.938 ;
               RECT 33.974 74.502 34.026 74.538 ;
               RECT 33.974 75.102 34.026 75.138 ;
               RECT 33.974 75.702 34.026 75.738 ;
               RECT 33.974 76.302 34.026 76.338 ;
               RECT 33.974 76.902 34.026 76.938 ;
               RECT 33.974 77.502 34.026 77.538 ;
               RECT 33.974 78.102 34.026 78.138 ;
               RECT 33.974 78.702 34.026 78.738 ;
               RECT 33.974 79.302 34.026 79.338 ;
               RECT 33.974 79.902 34.026 79.938 ;
               RECT 33.974 80.502 34.026 80.538 ;
               RECT 33.974 81.102 34.026 81.138 ;
               RECT 33.974 81.702 34.026 81.738 ;
               RECT 33.974 82.302 34.026 82.338 ;
               RECT 33.974 82.902 34.026 82.938 ;
               RECT 33.974 83.502 34.026 83.538 ;
               RECT 33.974 84.102 34.026 84.138 ;
               RECT 33.974 84.702 34.026 84.738 ;
               RECT 33.974 85.302 34.026 85.338 ;
               RECT 33.974 85.902 34.026 85.938 ;
               RECT 33.974 86.502 34.026 86.538 ;
               RECT 33.974 87.102 34.026 87.138 ;
               RECT 33.974 87.702 34.026 87.738 ;
               RECT 33.974 88.302 34.026 88.338 ;
               RECT 33.974 88.902 34.026 88.938 ;
               RECT 33.974 89.502 34.026 89.538 ;
               RECT 33.974 90.102 34.026 90.138 ;
               RECT 33.974 90.702 34.026 90.738 ;
               RECT 33.974 91.302 34.026 91.338 ;
               RECT 33.974 91.902 34.026 91.938 ;
               RECT 33.974 92.502 34.026 92.538 ;
               RECT 33.974 93.102 34.026 93.138 ;
               RECT 33.974 93.702 34.026 93.738 ;
               RECT 33.974 94.302 34.026 94.338 ;
               RECT 33.974 94.902 34.026 94.938 ;
               RECT 33.974 95.502 34.026 95.538 ;
               RECT 33.974 96.102 34.026 96.138 ;
               RECT 33.974 96.702 34.026 96.738 ;
               RECT 33.974 97.302 34.026 97.338 ;
               RECT 33.974 97.902 34.026 97.938 ;
               RECT 33.974 98.502 34.026 98.538 ;
               RECT 33.974 99.102 34.026 99.138 ;
               RECT 33.974 99.702 34.026 99.738 ;
               RECT 33.974 100.302 34.026 100.338 ;
               RECT 33.974 100.902 34.026 100.938 ;
               RECT 33.974 101.502 34.026 101.538 ;
               RECT 33.974 102.102 34.026 102.138 ;
               RECT 33.974 102.702 34.026 102.738 ;
               RECT 33.974 103.302 34.026 103.338 ;
               RECT 33.974 103.902 34.026 103.938 ;
               RECT 33.974 104.502 34.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 34.774 0.5695 34.826 104.5505 ;
               LAYER v4 ;
               RECT 34.774 0.582 34.826 0.618 ;
               RECT 34.774 1.182 34.826 1.218 ;
               RECT 34.774 1.782 34.826 1.818 ;
               RECT 34.774 2.382 34.826 2.418 ;
               RECT 34.774 2.982 34.826 3.018 ;
               RECT 34.774 3.582 34.826 3.618 ;
               RECT 34.774 4.182 34.826 4.218 ;
               RECT 34.774 4.782 34.826 4.818 ;
               RECT 34.774 5.382 34.826 5.418 ;
               RECT 34.774 5.982 34.826 6.018 ;
               RECT 34.774 6.582 34.826 6.618 ;
               RECT 34.774 7.182 34.826 7.218 ;
               RECT 34.774 7.782 34.826 7.818 ;
               RECT 34.774 8.382 34.826 8.418 ;
               RECT 34.774 8.982 34.826 9.018 ;
               RECT 34.774 9.582 34.826 9.618 ;
               RECT 34.774 10.182 34.826 10.218 ;
               RECT 34.774 10.782 34.826 10.818 ;
               RECT 34.774 11.382 34.826 11.418 ;
               RECT 34.774 11.982 34.826 12.018 ;
               RECT 34.774 12.582 34.826 12.618 ;
               RECT 34.774 13.182 34.826 13.218 ;
               RECT 34.774 13.782 34.826 13.818 ;
               RECT 34.774 14.382 34.826 14.418 ;
               RECT 34.774 14.982 34.826 15.018 ;
               RECT 34.774 15.582 34.826 15.618 ;
               RECT 34.774 16.182 34.826 16.218 ;
               RECT 34.774 16.782 34.826 16.818 ;
               RECT 34.774 17.382 34.826 17.418 ;
               RECT 34.774 17.982 34.826 18.018 ;
               RECT 34.774 18.582 34.826 18.618 ;
               RECT 34.774 19.182 34.826 19.218 ;
               RECT 34.774 19.782 34.826 19.818 ;
               RECT 34.774 20.382 34.826 20.418 ;
               RECT 34.774 20.982 34.826 21.018 ;
               RECT 34.774 21.582 34.826 21.618 ;
               RECT 34.774 22.182 34.826 22.218 ;
               RECT 34.774 22.782 34.826 22.818 ;
               RECT 34.774 23.382 34.826 23.418 ;
               RECT 34.774 23.982 34.826 24.018 ;
               RECT 34.774 24.582 34.826 24.618 ;
               RECT 34.774 25.182 34.826 25.218 ;
               RECT 34.774 25.782 34.826 25.818 ;
               RECT 34.774 26.382 34.826 26.418 ;
               RECT 34.774 26.982 34.826 27.018 ;
               RECT 34.774 27.582 34.826 27.618 ;
               RECT 34.774 28.182 34.826 28.218 ;
               RECT 34.774 28.782 34.826 28.818 ;
               RECT 34.774 29.382 34.826 29.418 ;
               RECT 34.774 29.982 34.826 30.018 ;
               RECT 34.774 30.582 34.826 30.618 ;
               RECT 34.774 31.182 34.826 31.218 ;
               RECT 34.774 31.782 34.826 31.818 ;
               RECT 34.774 32.382 34.826 32.418 ;
               RECT 34.774 32.982 34.826 33.018 ;
               RECT 34.774 33.582 34.826 33.618 ;
               RECT 34.774 34.182 34.826 34.218 ;
               RECT 34.774 34.782 34.826 34.818 ;
               RECT 34.774 35.382 34.826 35.418 ;
               RECT 34.774 35.982 34.826 36.018 ;
               RECT 34.774 36.582 34.826 36.618 ;
               RECT 34.774 37.182 34.826 37.218 ;
               RECT 34.774 37.782 34.826 37.818 ;
               RECT 34.774 38.382 34.826 38.418 ;
               RECT 34.774 38.982 34.826 39.018 ;
               RECT 34.774 39.582 34.826 39.618 ;
               RECT 34.774 40.182 34.826 40.218 ;
               RECT 34.774 40.782 34.826 40.818 ;
               RECT 34.774 41.382 34.826 41.418 ;
               RECT 34.774 41.982 34.826 42.018 ;
               RECT 34.774 42.582 34.826 42.618 ;
               RECT 34.774 43.182 34.826 43.218 ;
               RECT 34.774 43.782 34.826 43.818 ;
               RECT 34.774 44.382 34.826 44.418 ;
               RECT 34.774 44.982 34.826 45.018 ;
               RECT 34.774 45.582 34.826 45.618 ;
               RECT 34.774 46.182 34.826 46.218 ;
               RECT 34.774 46.782 34.826 46.818 ;
               RECT 34.774 47.382 34.826 47.418 ;
               RECT 34.774 47.982 34.826 48.018 ;
               RECT 34.774 48.582 34.826 48.618 ;
               RECT 34.774 48.942 34.826 48.978 ;
               RECT 34.774 49.182 34.826 49.218 ;
               RECT 34.774 49.902 34.826 49.938 ;
               RECT 34.774 50.622 34.826 50.658 ;
               RECT 34.774 50.862 34.826 50.898 ;
               RECT 34.774 51.342 34.826 51.378 ;
               RECT 34.774 51.822 34.826 51.858 ;
               RECT 34.774 52.302 34.826 52.338 ;
               RECT 34.774 52.782 34.826 52.818 ;
               RECT 34.774 53.262 34.826 53.298 ;
               RECT 34.774 53.742 34.826 53.778 ;
               RECT 34.774 54.222 34.826 54.258 ;
               RECT 34.774 54.462 34.826 54.498 ;
               RECT 34.774 55.182 34.826 55.218 ;
               RECT 34.774 55.902 34.826 55.938 ;
               RECT 34.774 56.142 34.826 56.178 ;
               RECT 34.774 56.502 34.826 56.538 ;
               RECT 34.774 57.102 34.826 57.138 ;
               RECT 34.774 57.702 34.826 57.738 ;
               RECT 34.774 58.302 34.826 58.338 ;
               RECT 34.774 58.902 34.826 58.938 ;
               RECT 34.774 59.502 34.826 59.538 ;
               RECT 34.774 60.102 34.826 60.138 ;
               RECT 34.774 60.702 34.826 60.738 ;
               RECT 34.774 61.302 34.826 61.338 ;
               RECT 34.774 61.902 34.826 61.938 ;
               RECT 34.774 62.502 34.826 62.538 ;
               RECT 34.774 63.102 34.826 63.138 ;
               RECT 34.774 63.702 34.826 63.738 ;
               RECT 34.774 64.302 34.826 64.338 ;
               RECT 34.774 64.902 34.826 64.938 ;
               RECT 34.774 65.502 34.826 65.538 ;
               RECT 34.774 66.102 34.826 66.138 ;
               RECT 34.774 66.702 34.826 66.738 ;
               RECT 34.774 67.302 34.826 67.338 ;
               RECT 34.774 67.902 34.826 67.938 ;
               RECT 34.774 68.502 34.826 68.538 ;
               RECT 34.774 69.102 34.826 69.138 ;
               RECT 34.774 69.702 34.826 69.738 ;
               RECT 34.774 70.302 34.826 70.338 ;
               RECT 34.774 70.902 34.826 70.938 ;
               RECT 34.774 71.502 34.826 71.538 ;
               RECT 34.774 72.102 34.826 72.138 ;
               RECT 34.774 72.702 34.826 72.738 ;
               RECT 34.774 73.302 34.826 73.338 ;
               RECT 34.774 73.902 34.826 73.938 ;
               RECT 34.774 74.502 34.826 74.538 ;
               RECT 34.774 75.102 34.826 75.138 ;
               RECT 34.774 75.702 34.826 75.738 ;
               RECT 34.774 76.302 34.826 76.338 ;
               RECT 34.774 76.902 34.826 76.938 ;
               RECT 34.774 77.502 34.826 77.538 ;
               RECT 34.774 78.102 34.826 78.138 ;
               RECT 34.774 78.702 34.826 78.738 ;
               RECT 34.774 79.302 34.826 79.338 ;
               RECT 34.774 79.902 34.826 79.938 ;
               RECT 34.774 80.502 34.826 80.538 ;
               RECT 34.774 81.102 34.826 81.138 ;
               RECT 34.774 81.702 34.826 81.738 ;
               RECT 34.774 82.302 34.826 82.338 ;
               RECT 34.774 82.902 34.826 82.938 ;
               RECT 34.774 83.502 34.826 83.538 ;
               RECT 34.774 84.102 34.826 84.138 ;
               RECT 34.774 84.702 34.826 84.738 ;
               RECT 34.774 85.302 34.826 85.338 ;
               RECT 34.774 85.902 34.826 85.938 ;
               RECT 34.774 86.502 34.826 86.538 ;
               RECT 34.774 87.102 34.826 87.138 ;
               RECT 34.774 87.702 34.826 87.738 ;
               RECT 34.774 88.302 34.826 88.338 ;
               RECT 34.774 88.902 34.826 88.938 ;
               RECT 34.774 89.502 34.826 89.538 ;
               RECT 34.774 90.102 34.826 90.138 ;
               RECT 34.774 90.702 34.826 90.738 ;
               RECT 34.774 91.302 34.826 91.338 ;
               RECT 34.774 91.902 34.826 91.938 ;
               RECT 34.774 92.502 34.826 92.538 ;
               RECT 34.774 93.102 34.826 93.138 ;
               RECT 34.774 93.702 34.826 93.738 ;
               RECT 34.774 94.302 34.826 94.338 ;
               RECT 34.774 94.902 34.826 94.938 ;
               RECT 34.774 95.502 34.826 95.538 ;
               RECT 34.774 96.102 34.826 96.138 ;
               RECT 34.774 96.702 34.826 96.738 ;
               RECT 34.774 97.302 34.826 97.338 ;
               RECT 34.774 97.902 34.826 97.938 ;
               RECT 34.774 98.502 34.826 98.538 ;
               RECT 34.774 99.102 34.826 99.138 ;
               RECT 34.774 99.702 34.826 99.738 ;
               RECT 34.774 100.302 34.826 100.338 ;
               RECT 34.774 100.902 34.826 100.938 ;
               RECT 34.774 101.502 34.826 101.538 ;
               RECT 34.774 102.102 34.826 102.138 ;
               RECT 34.774 102.702 34.826 102.738 ;
               RECT 34.774 103.302 34.826 103.338 ;
               RECT 34.774 103.902 34.826 103.938 ;
               RECT 34.774 104.502 34.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 35.574 0.5695 35.626 104.5505 ;
               LAYER v4 ;
               RECT 35.574 0.582 35.626 0.618 ;
               RECT 35.574 1.182 35.626 1.218 ;
               RECT 35.574 1.782 35.626 1.818 ;
               RECT 35.574 2.382 35.626 2.418 ;
               RECT 35.574 2.982 35.626 3.018 ;
               RECT 35.574 3.582 35.626 3.618 ;
               RECT 35.574 4.182 35.626 4.218 ;
               RECT 35.574 4.782 35.626 4.818 ;
               RECT 35.574 5.382 35.626 5.418 ;
               RECT 35.574 5.982 35.626 6.018 ;
               RECT 35.574 6.582 35.626 6.618 ;
               RECT 35.574 7.182 35.626 7.218 ;
               RECT 35.574 7.782 35.626 7.818 ;
               RECT 35.574 8.382 35.626 8.418 ;
               RECT 35.574 8.982 35.626 9.018 ;
               RECT 35.574 9.582 35.626 9.618 ;
               RECT 35.574 10.182 35.626 10.218 ;
               RECT 35.574 10.782 35.626 10.818 ;
               RECT 35.574 11.382 35.626 11.418 ;
               RECT 35.574 11.982 35.626 12.018 ;
               RECT 35.574 12.582 35.626 12.618 ;
               RECT 35.574 13.182 35.626 13.218 ;
               RECT 35.574 13.782 35.626 13.818 ;
               RECT 35.574 14.382 35.626 14.418 ;
               RECT 35.574 14.982 35.626 15.018 ;
               RECT 35.574 15.582 35.626 15.618 ;
               RECT 35.574 16.182 35.626 16.218 ;
               RECT 35.574 16.782 35.626 16.818 ;
               RECT 35.574 17.382 35.626 17.418 ;
               RECT 35.574 17.982 35.626 18.018 ;
               RECT 35.574 18.582 35.626 18.618 ;
               RECT 35.574 19.182 35.626 19.218 ;
               RECT 35.574 19.782 35.626 19.818 ;
               RECT 35.574 20.382 35.626 20.418 ;
               RECT 35.574 20.982 35.626 21.018 ;
               RECT 35.574 21.582 35.626 21.618 ;
               RECT 35.574 22.182 35.626 22.218 ;
               RECT 35.574 22.782 35.626 22.818 ;
               RECT 35.574 23.382 35.626 23.418 ;
               RECT 35.574 23.982 35.626 24.018 ;
               RECT 35.574 24.582 35.626 24.618 ;
               RECT 35.574 25.182 35.626 25.218 ;
               RECT 35.574 25.782 35.626 25.818 ;
               RECT 35.574 26.382 35.626 26.418 ;
               RECT 35.574 26.982 35.626 27.018 ;
               RECT 35.574 27.582 35.626 27.618 ;
               RECT 35.574 28.182 35.626 28.218 ;
               RECT 35.574 28.782 35.626 28.818 ;
               RECT 35.574 29.382 35.626 29.418 ;
               RECT 35.574 29.982 35.626 30.018 ;
               RECT 35.574 30.582 35.626 30.618 ;
               RECT 35.574 31.182 35.626 31.218 ;
               RECT 35.574 31.782 35.626 31.818 ;
               RECT 35.574 32.382 35.626 32.418 ;
               RECT 35.574 32.982 35.626 33.018 ;
               RECT 35.574 33.582 35.626 33.618 ;
               RECT 35.574 34.182 35.626 34.218 ;
               RECT 35.574 34.782 35.626 34.818 ;
               RECT 35.574 35.382 35.626 35.418 ;
               RECT 35.574 35.982 35.626 36.018 ;
               RECT 35.574 36.582 35.626 36.618 ;
               RECT 35.574 37.182 35.626 37.218 ;
               RECT 35.574 37.782 35.626 37.818 ;
               RECT 35.574 38.382 35.626 38.418 ;
               RECT 35.574 38.982 35.626 39.018 ;
               RECT 35.574 39.582 35.626 39.618 ;
               RECT 35.574 40.182 35.626 40.218 ;
               RECT 35.574 40.782 35.626 40.818 ;
               RECT 35.574 41.382 35.626 41.418 ;
               RECT 35.574 41.982 35.626 42.018 ;
               RECT 35.574 42.582 35.626 42.618 ;
               RECT 35.574 43.182 35.626 43.218 ;
               RECT 35.574 43.782 35.626 43.818 ;
               RECT 35.574 44.382 35.626 44.418 ;
               RECT 35.574 44.982 35.626 45.018 ;
               RECT 35.574 45.582 35.626 45.618 ;
               RECT 35.574 46.182 35.626 46.218 ;
               RECT 35.574 46.782 35.626 46.818 ;
               RECT 35.574 47.382 35.626 47.418 ;
               RECT 35.574 47.982 35.626 48.018 ;
               RECT 35.574 48.582 35.626 48.618 ;
               RECT 35.574 48.9475 35.626 48.9725 ;
               RECT 35.574 49.182 35.626 49.218 ;
               RECT 35.574 49.902 35.626 49.938 ;
               RECT 35.574 50.622 35.626 50.658 ;
               RECT 35.574 50.862 35.626 50.898 ;
               RECT 35.574 51.342 35.626 51.378 ;
               RECT 35.574 51.822 35.626 51.858 ;
               RECT 35.574 52.302 35.626 52.338 ;
               RECT 35.574 52.782 35.626 52.818 ;
               RECT 35.574 53.262 35.626 53.298 ;
               RECT 35.574 53.742 35.626 53.778 ;
               RECT 35.574 54.222 35.626 54.258 ;
               RECT 35.574 54.462 35.626 54.498 ;
               RECT 35.574 55.182 35.626 55.218 ;
               RECT 35.574 55.902 35.626 55.938 ;
               RECT 35.574 56.1475 35.626 56.1725 ;
               RECT 35.574 56.502 35.626 56.538 ;
               RECT 35.574 57.102 35.626 57.138 ;
               RECT 35.574 57.702 35.626 57.738 ;
               RECT 35.574 58.302 35.626 58.338 ;
               RECT 35.574 58.902 35.626 58.938 ;
               RECT 35.574 59.502 35.626 59.538 ;
               RECT 35.574 60.102 35.626 60.138 ;
               RECT 35.574 60.702 35.626 60.738 ;
               RECT 35.574 61.302 35.626 61.338 ;
               RECT 35.574 61.902 35.626 61.938 ;
               RECT 35.574 62.502 35.626 62.538 ;
               RECT 35.574 63.102 35.626 63.138 ;
               RECT 35.574 63.702 35.626 63.738 ;
               RECT 35.574 64.302 35.626 64.338 ;
               RECT 35.574 64.902 35.626 64.938 ;
               RECT 35.574 65.502 35.626 65.538 ;
               RECT 35.574 66.102 35.626 66.138 ;
               RECT 35.574 66.702 35.626 66.738 ;
               RECT 35.574 67.302 35.626 67.338 ;
               RECT 35.574 67.902 35.626 67.938 ;
               RECT 35.574 68.502 35.626 68.538 ;
               RECT 35.574 69.102 35.626 69.138 ;
               RECT 35.574 69.702 35.626 69.738 ;
               RECT 35.574 70.302 35.626 70.338 ;
               RECT 35.574 70.902 35.626 70.938 ;
               RECT 35.574 71.502 35.626 71.538 ;
               RECT 35.574 72.102 35.626 72.138 ;
               RECT 35.574 72.702 35.626 72.738 ;
               RECT 35.574 73.302 35.626 73.338 ;
               RECT 35.574 73.902 35.626 73.938 ;
               RECT 35.574 74.502 35.626 74.538 ;
               RECT 35.574 75.102 35.626 75.138 ;
               RECT 35.574 75.702 35.626 75.738 ;
               RECT 35.574 76.302 35.626 76.338 ;
               RECT 35.574 76.902 35.626 76.938 ;
               RECT 35.574 77.502 35.626 77.538 ;
               RECT 35.574 78.102 35.626 78.138 ;
               RECT 35.574 78.702 35.626 78.738 ;
               RECT 35.574 79.302 35.626 79.338 ;
               RECT 35.574 79.902 35.626 79.938 ;
               RECT 35.574 80.502 35.626 80.538 ;
               RECT 35.574 81.102 35.626 81.138 ;
               RECT 35.574 81.702 35.626 81.738 ;
               RECT 35.574 82.302 35.626 82.338 ;
               RECT 35.574 82.902 35.626 82.938 ;
               RECT 35.574 83.502 35.626 83.538 ;
               RECT 35.574 84.102 35.626 84.138 ;
               RECT 35.574 84.702 35.626 84.738 ;
               RECT 35.574 85.302 35.626 85.338 ;
               RECT 35.574 85.902 35.626 85.938 ;
               RECT 35.574 86.502 35.626 86.538 ;
               RECT 35.574 87.102 35.626 87.138 ;
               RECT 35.574 87.702 35.626 87.738 ;
               RECT 35.574 88.302 35.626 88.338 ;
               RECT 35.574 88.902 35.626 88.938 ;
               RECT 35.574 89.502 35.626 89.538 ;
               RECT 35.574 90.102 35.626 90.138 ;
               RECT 35.574 90.702 35.626 90.738 ;
               RECT 35.574 91.302 35.626 91.338 ;
               RECT 35.574 91.902 35.626 91.938 ;
               RECT 35.574 92.502 35.626 92.538 ;
               RECT 35.574 93.102 35.626 93.138 ;
               RECT 35.574 93.702 35.626 93.738 ;
               RECT 35.574 94.302 35.626 94.338 ;
               RECT 35.574 94.902 35.626 94.938 ;
               RECT 35.574 95.502 35.626 95.538 ;
               RECT 35.574 96.102 35.626 96.138 ;
               RECT 35.574 96.702 35.626 96.738 ;
               RECT 35.574 97.302 35.626 97.338 ;
               RECT 35.574 97.902 35.626 97.938 ;
               RECT 35.574 98.502 35.626 98.538 ;
               RECT 35.574 99.102 35.626 99.138 ;
               RECT 35.574 99.702 35.626 99.738 ;
               RECT 35.574 100.302 35.626 100.338 ;
               RECT 35.574 100.902 35.626 100.938 ;
               RECT 35.574 101.502 35.626 101.538 ;
               RECT 35.574 102.102 35.626 102.138 ;
               RECT 35.574 102.702 35.626 102.738 ;
               RECT 35.574 103.302 35.626 103.338 ;
               RECT 35.574 103.902 35.626 103.938 ;
               RECT 35.574 104.502 35.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 4.574 0.5695 4.626 104.5505 ;
               LAYER v4 ;
               RECT 4.574 0.582 4.626 0.618 ;
               RECT 4.574 1.182 4.626 1.218 ;
               RECT 4.574 1.782 4.626 1.818 ;
               RECT 4.574 2.382 4.626 2.418 ;
               RECT 4.574 2.982 4.626 3.018 ;
               RECT 4.574 3.582 4.626 3.618 ;
               RECT 4.574 4.182 4.626 4.218 ;
               RECT 4.574 4.782 4.626 4.818 ;
               RECT 4.574 5.382 4.626 5.418 ;
               RECT 4.574 5.982 4.626 6.018 ;
               RECT 4.574 6.582 4.626 6.618 ;
               RECT 4.574 7.182 4.626 7.218 ;
               RECT 4.574 7.782 4.626 7.818 ;
               RECT 4.574 8.382 4.626 8.418 ;
               RECT 4.574 8.982 4.626 9.018 ;
               RECT 4.574 9.582 4.626 9.618 ;
               RECT 4.574 10.182 4.626 10.218 ;
               RECT 4.574 10.782 4.626 10.818 ;
               RECT 4.574 11.382 4.626 11.418 ;
               RECT 4.574 11.982 4.626 12.018 ;
               RECT 4.574 12.582 4.626 12.618 ;
               RECT 4.574 13.182 4.626 13.218 ;
               RECT 4.574 13.782 4.626 13.818 ;
               RECT 4.574 14.382 4.626 14.418 ;
               RECT 4.574 14.982 4.626 15.018 ;
               RECT 4.574 15.582 4.626 15.618 ;
               RECT 4.574 16.182 4.626 16.218 ;
               RECT 4.574 16.782 4.626 16.818 ;
               RECT 4.574 17.382 4.626 17.418 ;
               RECT 4.574 17.982 4.626 18.018 ;
               RECT 4.574 18.582 4.626 18.618 ;
               RECT 4.574 19.182 4.626 19.218 ;
               RECT 4.574 19.782 4.626 19.818 ;
               RECT 4.574 20.382 4.626 20.418 ;
               RECT 4.574 20.982 4.626 21.018 ;
               RECT 4.574 21.582 4.626 21.618 ;
               RECT 4.574 22.182 4.626 22.218 ;
               RECT 4.574 22.782 4.626 22.818 ;
               RECT 4.574 23.382 4.626 23.418 ;
               RECT 4.574 23.982 4.626 24.018 ;
               RECT 4.574 24.582 4.626 24.618 ;
               RECT 4.574 25.182 4.626 25.218 ;
               RECT 4.574 25.782 4.626 25.818 ;
               RECT 4.574 26.382 4.626 26.418 ;
               RECT 4.574 26.982 4.626 27.018 ;
               RECT 4.574 27.582 4.626 27.618 ;
               RECT 4.574 28.182 4.626 28.218 ;
               RECT 4.574 28.782 4.626 28.818 ;
               RECT 4.574 29.382 4.626 29.418 ;
               RECT 4.574 29.982 4.626 30.018 ;
               RECT 4.574 30.582 4.626 30.618 ;
               RECT 4.574 31.182 4.626 31.218 ;
               RECT 4.574 31.782 4.626 31.818 ;
               RECT 4.574 32.382 4.626 32.418 ;
               RECT 4.574 32.982 4.626 33.018 ;
               RECT 4.574 33.582 4.626 33.618 ;
               RECT 4.574 34.182 4.626 34.218 ;
               RECT 4.574 34.782 4.626 34.818 ;
               RECT 4.574 35.382 4.626 35.418 ;
               RECT 4.574 35.982 4.626 36.018 ;
               RECT 4.574 36.582 4.626 36.618 ;
               RECT 4.574 37.182 4.626 37.218 ;
               RECT 4.574 37.782 4.626 37.818 ;
               RECT 4.574 38.382 4.626 38.418 ;
               RECT 4.574 38.982 4.626 39.018 ;
               RECT 4.574 39.582 4.626 39.618 ;
               RECT 4.574 40.182 4.626 40.218 ;
               RECT 4.574 40.782 4.626 40.818 ;
               RECT 4.574 41.382 4.626 41.418 ;
               RECT 4.574 41.982 4.626 42.018 ;
               RECT 4.574 42.582 4.626 42.618 ;
               RECT 4.574 43.182 4.626 43.218 ;
               RECT 4.574 43.782 4.626 43.818 ;
               RECT 4.574 44.382 4.626 44.418 ;
               RECT 4.574 44.982 4.626 45.018 ;
               RECT 4.574 45.582 4.626 45.618 ;
               RECT 4.574 46.182 4.626 46.218 ;
               RECT 4.574 46.782 4.626 46.818 ;
               RECT 4.574 47.382 4.626 47.418 ;
               RECT 4.574 47.982 4.626 48.018 ;
               RECT 4.574 48.582 4.626 48.618 ;
               RECT 4.574 48.942 4.626 48.978 ;
               RECT 4.574 49.182 4.626 49.218 ;
               RECT 4.574 49.902 4.626 49.938 ;
               RECT 4.574 50.622 4.626 50.658 ;
               RECT 4.574 50.862 4.626 50.898 ;
               RECT 4.574 51.342 4.626 51.378 ;
               RECT 4.574 51.822 4.626 51.858 ;
               RECT 4.574 52.302 4.626 52.338 ;
               RECT 4.574 52.782 4.626 52.818 ;
               RECT 4.574 53.262 4.626 53.298 ;
               RECT 4.574 53.742 4.626 53.778 ;
               RECT 4.574 54.222 4.626 54.258 ;
               RECT 4.574 54.462 4.626 54.498 ;
               RECT 4.574 55.182 4.626 55.218 ;
               RECT 4.574 55.902 4.626 55.938 ;
               RECT 4.574 56.142 4.626 56.178 ;
               RECT 4.574 56.502 4.626 56.538 ;
               RECT 4.574 57.102 4.626 57.138 ;
               RECT 4.574 57.702 4.626 57.738 ;
               RECT 4.574 58.302 4.626 58.338 ;
               RECT 4.574 58.902 4.626 58.938 ;
               RECT 4.574 59.502 4.626 59.538 ;
               RECT 4.574 60.102 4.626 60.138 ;
               RECT 4.574 60.702 4.626 60.738 ;
               RECT 4.574 61.302 4.626 61.338 ;
               RECT 4.574 61.902 4.626 61.938 ;
               RECT 4.574 62.502 4.626 62.538 ;
               RECT 4.574 63.102 4.626 63.138 ;
               RECT 4.574 63.702 4.626 63.738 ;
               RECT 4.574 64.302 4.626 64.338 ;
               RECT 4.574 64.902 4.626 64.938 ;
               RECT 4.574 65.502 4.626 65.538 ;
               RECT 4.574 66.102 4.626 66.138 ;
               RECT 4.574 66.702 4.626 66.738 ;
               RECT 4.574 67.302 4.626 67.338 ;
               RECT 4.574 67.902 4.626 67.938 ;
               RECT 4.574 68.502 4.626 68.538 ;
               RECT 4.574 69.102 4.626 69.138 ;
               RECT 4.574 69.702 4.626 69.738 ;
               RECT 4.574 70.302 4.626 70.338 ;
               RECT 4.574 70.902 4.626 70.938 ;
               RECT 4.574 71.502 4.626 71.538 ;
               RECT 4.574 72.102 4.626 72.138 ;
               RECT 4.574 72.702 4.626 72.738 ;
               RECT 4.574 73.302 4.626 73.338 ;
               RECT 4.574 73.902 4.626 73.938 ;
               RECT 4.574 74.502 4.626 74.538 ;
               RECT 4.574 75.102 4.626 75.138 ;
               RECT 4.574 75.702 4.626 75.738 ;
               RECT 4.574 76.302 4.626 76.338 ;
               RECT 4.574 76.902 4.626 76.938 ;
               RECT 4.574 77.502 4.626 77.538 ;
               RECT 4.574 78.102 4.626 78.138 ;
               RECT 4.574 78.702 4.626 78.738 ;
               RECT 4.574 79.302 4.626 79.338 ;
               RECT 4.574 79.902 4.626 79.938 ;
               RECT 4.574 80.502 4.626 80.538 ;
               RECT 4.574 81.102 4.626 81.138 ;
               RECT 4.574 81.702 4.626 81.738 ;
               RECT 4.574 82.302 4.626 82.338 ;
               RECT 4.574 82.902 4.626 82.938 ;
               RECT 4.574 83.502 4.626 83.538 ;
               RECT 4.574 84.102 4.626 84.138 ;
               RECT 4.574 84.702 4.626 84.738 ;
               RECT 4.574 85.302 4.626 85.338 ;
               RECT 4.574 85.902 4.626 85.938 ;
               RECT 4.574 86.502 4.626 86.538 ;
               RECT 4.574 87.102 4.626 87.138 ;
               RECT 4.574 87.702 4.626 87.738 ;
               RECT 4.574 88.302 4.626 88.338 ;
               RECT 4.574 88.902 4.626 88.938 ;
               RECT 4.574 89.502 4.626 89.538 ;
               RECT 4.574 90.102 4.626 90.138 ;
               RECT 4.574 90.702 4.626 90.738 ;
               RECT 4.574 91.302 4.626 91.338 ;
               RECT 4.574 91.902 4.626 91.938 ;
               RECT 4.574 92.502 4.626 92.538 ;
               RECT 4.574 93.102 4.626 93.138 ;
               RECT 4.574 93.702 4.626 93.738 ;
               RECT 4.574 94.302 4.626 94.338 ;
               RECT 4.574 94.902 4.626 94.938 ;
               RECT 4.574 95.502 4.626 95.538 ;
               RECT 4.574 96.102 4.626 96.138 ;
               RECT 4.574 96.702 4.626 96.738 ;
               RECT 4.574 97.302 4.626 97.338 ;
               RECT 4.574 97.902 4.626 97.938 ;
               RECT 4.574 98.502 4.626 98.538 ;
               RECT 4.574 99.102 4.626 99.138 ;
               RECT 4.574 99.702 4.626 99.738 ;
               RECT 4.574 100.302 4.626 100.338 ;
               RECT 4.574 100.902 4.626 100.938 ;
               RECT 4.574 101.502 4.626 101.538 ;
               RECT 4.574 102.102 4.626 102.138 ;
               RECT 4.574 102.702 4.626 102.738 ;
               RECT 4.574 103.302 4.626 103.338 ;
               RECT 4.574 103.902 4.626 103.938 ;
               RECT 4.574 104.502 4.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 5.374 0.5695 5.426 104.5505 ;
               LAYER v4 ;
               RECT 5.374 0.582 5.426 0.618 ;
               RECT 5.374 1.182 5.426 1.218 ;
               RECT 5.374 1.782 5.426 1.818 ;
               RECT 5.374 2.382 5.426 2.418 ;
               RECT 5.374 2.982 5.426 3.018 ;
               RECT 5.374 3.582 5.426 3.618 ;
               RECT 5.374 4.182 5.426 4.218 ;
               RECT 5.374 4.782 5.426 4.818 ;
               RECT 5.374 5.382 5.426 5.418 ;
               RECT 5.374 5.982 5.426 6.018 ;
               RECT 5.374 6.582 5.426 6.618 ;
               RECT 5.374 7.182 5.426 7.218 ;
               RECT 5.374 7.782 5.426 7.818 ;
               RECT 5.374 8.382 5.426 8.418 ;
               RECT 5.374 8.982 5.426 9.018 ;
               RECT 5.374 9.582 5.426 9.618 ;
               RECT 5.374 10.182 5.426 10.218 ;
               RECT 5.374 10.782 5.426 10.818 ;
               RECT 5.374 11.382 5.426 11.418 ;
               RECT 5.374 11.982 5.426 12.018 ;
               RECT 5.374 12.582 5.426 12.618 ;
               RECT 5.374 13.182 5.426 13.218 ;
               RECT 5.374 13.782 5.426 13.818 ;
               RECT 5.374 14.382 5.426 14.418 ;
               RECT 5.374 14.982 5.426 15.018 ;
               RECT 5.374 15.582 5.426 15.618 ;
               RECT 5.374 16.182 5.426 16.218 ;
               RECT 5.374 16.782 5.426 16.818 ;
               RECT 5.374 17.382 5.426 17.418 ;
               RECT 5.374 17.982 5.426 18.018 ;
               RECT 5.374 18.582 5.426 18.618 ;
               RECT 5.374 19.182 5.426 19.218 ;
               RECT 5.374 19.782 5.426 19.818 ;
               RECT 5.374 20.382 5.426 20.418 ;
               RECT 5.374 20.982 5.426 21.018 ;
               RECT 5.374 21.582 5.426 21.618 ;
               RECT 5.374 22.182 5.426 22.218 ;
               RECT 5.374 22.782 5.426 22.818 ;
               RECT 5.374 23.382 5.426 23.418 ;
               RECT 5.374 23.982 5.426 24.018 ;
               RECT 5.374 24.582 5.426 24.618 ;
               RECT 5.374 25.182 5.426 25.218 ;
               RECT 5.374 25.782 5.426 25.818 ;
               RECT 5.374 26.382 5.426 26.418 ;
               RECT 5.374 26.982 5.426 27.018 ;
               RECT 5.374 27.582 5.426 27.618 ;
               RECT 5.374 28.182 5.426 28.218 ;
               RECT 5.374 28.782 5.426 28.818 ;
               RECT 5.374 29.382 5.426 29.418 ;
               RECT 5.374 29.982 5.426 30.018 ;
               RECT 5.374 30.582 5.426 30.618 ;
               RECT 5.374 31.182 5.426 31.218 ;
               RECT 5.374 31.782 5.426 31.818 ;
               RECT 5.374 32.382 5.426 32.418 ;
               RECT 5.374 32.982 5.426 33.018 ;
               RECT 5.374 33.582 5.426 33.618 ;
               RECT 5.374 34.182 5.426 34.218 ;
               RECT 5.374 34.782 5.426 34.818 ;
               RECT 5.374 35.382 5.426 35.418 ;
               RECT 5.374 35.982 5.426 36.018 ;
               RECT 5.374 36.582 5.426 36.618 ;
               RECT 5.374 37.182 5.426 37.218 ;
               RECT 5.374 37.782 5.426 37.818 ;
               RECT 5.374 38.382 5.426 38.418 ;
               RECT 5.374 38.982 5.426 39.018 ;
               RECT 5.374 39.582 5.426 39.618 ;
               RECT 5.374 40.182 5.426 40.218 ;
               RECT 5.374 40.782 5.426 40.818 ;
               RECT 5.374 41.382 5.426 41.418 ;
               RECT 5.374 41.982 5.426 42.018 ;
               RECT 5.374 42.582 5.426 42.618 ;
               RECT 5.374 43.182 5.426 43.218 ;
               RECT 5.374 43.782 5.426 43.818 ;
               RECT 5.374 44.382 5.426 44.418 ;
               RECT 5.374 44.982 5.426 45.018 ;
               RECT 5.374 45.582 5.426 45.618 ;
               RECT 5.374 46.182 5.426 46.218 ;
               RECT 5.374 46.782 5.426 46.818 ;
               RECT 5.374 47.382 5.426 47.418 ;
               RECT 5.374 47.982 5.426 48.018 ;
               RECT 5.374 48.582 5.426 48.618 ;
               RECT 5.374 48.942 5.426 48.978 ;
               RECT 5.374 48.9475 5.426 48.9725 ;
               RECT 5.374 49.182 5.426 49.218 ;
               RECT 5.374 49.902 5.426 49.938 ;
               RECT 5.374 50.622 5.426 50.658 ;
               RECT 5.374 50.862 5.426 50.898 ;
               RECT 5.374 51.342 5.426 51.378 ;
               RECT 5.374 51.822 5.426 51.858 ;
               RECT 5.374 52.302 5.426 52.338 ;
               RECT 5.374 52.782 5.426 52.818 ;
               RECT 5.374 53.262 5.426 53.298 ;
               RECT 5.374 53.742 5.426 53.778 ;
               RECT 5.374 54.222 5.426 54.258 ;
               RECT 5.374 54.462 5.426 54.498 ;
               RECT 5.374 55.182 5.426 55.218 ;
               RECT 5.374 55.902 5.426 55.938 ;
               RECT 5.374 56.142 5.426 56.178 ;
               RECT 5.374 56.1475 5.426 56.1725 ;
               RECT 5.374 56.502 5.426 56.538 ;
               RECT 5.374 57.102 5.426 57.138 ;
               RECT 5.374 57.702 5.426 57.738 ;
               RECT 5.374 58.302 5.426 58.338 ;
               RECT 5.374 58.902 5.426 58.938 ;
               RECT 5.374 59.502 5.426 59.538 ;
               RECT 5.374 60.102 5.426 60.138 ;
               RECT 5.374 60.702 5.426 60.738 ;
               RECT 5.374 61.302 5.426 61.338 ;
               RECT 5.374 61.902 5.426 61.938 ;
               RECT 5.374 62.502 5.426 62.538 ;
               RECT 5.374 63.102 5.426 63.138 ;
               RECT 5.374 63.702 5.426 63.738 ;
               RECT 5.374 64.302 5.426 64.338 ;
               RECT 5.374 64.902 5.426 64.938 ;
               RECT 5.374 65.502 5.426 65.538 ;
               RECT 5.374 66.102 5.426 66.138 ;
               RECT 5.374 66.702 5.426 66.738 ;
               RECT 5.374 67.302 5.426 67.338 ;
               RECT 5.374 67.902 5.426 67.938 ;
               RECT 5.374 68.502 5.426 68.538 ;
               RECT 5.374 69.102 5.426 69.138 ;
               RECT 5.374 69.702 5.426 69.738 ;
               RECT 5.374 70.302 5.426 70.338 ;
               RECT 5.374 70.902 5.426 70.938 ;
               RECT 5.374 71.502 5.426 71.538 ;
               RECT 5.374 72.102 5.426 72.138 ;
               RECT 5.374 72.702 5.426 72.738 ;
               RECT 5.374 73.302 5.426 73.338 ;
               RECT 5.374 73.902 5.426 73.938 ;
               RECT 5.374 74.502 5.426 74.538 ;
               RECT 5.374 75.102 5.426 75.138 ;
               RECT 5.374 75.702 5.426 75.738 ;
               RECT 5.374 76.302 5.426 76.338 ;
               RECT 5.374 76.902 5.426 76.938 ;
               RECT 5.374 77.502 5.426 77.538 ;
               RECT 5.374 78.102 5.426 78.138 ;
               RECT 5.374 78.702 5.426 78.738 ;
               RECT 5.374 79.302 5.426 79.338 ;
               RECT 5.374 79.902 5.426 79.938 ;
               RECT 5.374 80.502 5.426 80.538 ;
               RECT 5.374 81.102 5.426 81.138 ;
               RECT 5.374 81.702 5.426 81.738 ;
               RECT 5.374 82.302 5.426 82.338 ;
               RECT 5.374 82.902 5.426 82.938 ;
               RECT 5.374 83.502 5.426 83.538 ;
               RECT 5.374 84.102 5.426 84.138 ;
               RECT 5.374 84.702 5.426 84.738 ;
               RECT 5.374 85.302 5.426 85.338 ;
               RECT 5.374 85.902 5.426 85.938 ;
               RECT 5.374 86.502 5.426 86.538 ;
               RECT 5.374 87.102 5.426 87.138 ;
               RECT 5.374 87.702 5.426 87.738 ;
               RECT 5.374 88.302 5.426 88.338 ;
               RECT 5.374 88.902 5.426 88.938 ;
               RECT 5.374 89.502 5.426 89.538 ;
               RECT 5.374 90.102 5.426 90.138 ;
               RECT 5.374 90.702 5.426 90.738 ;
               RECT 5.374 91.302 5.426 91.338 ;
               RECT 5.374 91.902 5.426 91.938 ;
               RECT 5.374 92.502 5.426 92.538 ;
               RECT 5.374 93.102 5.426 93.138 ;
               RECT 5.374 93.702 5.426 93.738 ;
               RECT 5.374 94.302 5.426 94.338 ;
               RECT 5.374 94.902 5.426 94.938 ;
               RECT 5.374 95.502 5.426 95.538 ;
               RECT 5.374 96.102 5.426 96.138 ;
               RECT 5.374 96.702 5.426 96.738 ;
               RECT 5.374 97.302 5.426 97.338 ;
               RECT 5.374 97.902 5.426 97.938 ;
               RECT 5.374 98.502 5.426 98.538 ;
               RECT 5.374 99.102 5.426 99.138 ;
               RECT 5.374 99.702 5.426 99.738 ;
               RECT 5.374 100.302 5.426 100.338 ;
               RECT 5.374 100.902 5.426 100.938 ;
               RECT 5.374 101.502 5.426 101.538 ;
               RECT 5.374 102.102 5.426 102.138 ;
               RECT 5.374 102.702 5.426 102.738 ;
               RECT 5.374 103.302 5.426 103.338 ;
               RECT 5.374 103.902 5.426 103.938 ;
               RECT 5.374 104.502 5.426 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 6.174 0.5695 6.226 104.5505 ;
               LAYER v4 ;
               RECT 6.174 0.582 6.226 0.618 ;
               RECT 6.174 1.182 6.226 1.218 ;
               RECT 6.174 1.782 6.226 1.818 ;
               RECT 6.174 2.382 6.226 2.418 ;
               RECT 6.174 2.982 6.226 3.018 ;
               RECT 6.174 3.582 6.226 3.618 ;
               RECT 6.174 4.182 6.226 4.218 ;
               RECT 6.174 4.782 6.226 4.818 ;
               RECT 6.174 5.382 6.226 5.418 ;
               RECT 6.174 5.982 6.226 6.018 ;
               RECT 6.174 6.582 6.226 6.618 ;
               RECT 6.174 7.182 6.226 7.218 ;
               RECT 6.174 7.782 6.226 7.818 ;
               RECT 6.174 8.382 6.226 8.418 ;
               RECT 6.174 8.982 6.226 9.018 ;
               RECT 6.174 9.582 6.226 9.618 ;
               RECT 6.174 10.182 6.226 10.218 ;
               RECT 6.174 10.782 6.226 10.818 ;
               RECT 6.174 11.382 6.226 11.418 ;
               RECT 6.174 11.982 6.226 12.018 ;
               RECT 6.174 12.582 6.226 12.618 ;
               RECT 6.174 13.182 6.226 13.218 ;
               RECT 6.174 13.782 6.226 13.818 ;
               RECT 6.174 14.382 6.226 14.418 ;
               RECT 6.174 14.982 6.226 15.018 ;
               RECT 6.174 15.582 6.226 15.618 ;
               RECT 6.174 16.182 6.226 16.218 ;
               RECT 6.174 16.782 6.226 16.818 ;
               RECT 6.174 17.382 6.226 17.418 ;
               RECT 6.174 17.982 6.226 18.018 ;
               RECT 6.174 18.582 6.226 18.618 ;
               RECT 6.174 19.182 6.226 19.218 ;
               RECT 6.174 19.782 6.226 19.818 ;
               RECT 6.174 20.382 6.226 20.418 ;
               RECT 6.174 20.982 6.226 21.018 ;
               RECT 6.174 21.582 6.226 21.618 ;
               RECT 6.174 22.182 6.226 22.218 ;
               RECT 6.174 22.782 6.226 22.818 ;
               RECT 6.174 23.382 6.226 23.418 ;
               RECT 6.174 23.982 6.226 24.018 ;
               RECT 6.174 24.582 6.226 24.618 ;
               RECT 6.174 25.182 6.226 25.218 ;
               RECT 6.174 25.782 6.226 25.818 ;
               RECT 6.174 26.382 6.226 26.418 ;
               RECT 6.174 26.982 6.226 27.018 ;
               RECT 6.174 27.582 6.226 27.618 ;
               RECT 6.174 28.182 6.226 28.218 ;
               RECT 6.174 28.782 6.226 28.818 ;
               RECT 6.174 29.382 6.226 29.418 ;
               RECT 6.174 29.982 6.226 30.018 ;
               RECT 6.174 30.582 6.226 30.618 ;
               RECT 6.174 31.182 6.226 31.218 ;
               RECT 6.174 31.782 6.226 31.818 ;
               RECT 6.174 32.382 6.226 32.418 ;
               RECT 6.174 32.982 6.226 33.018 ;
               RECT 6.174 33.582 6.226 33.618 ;
               RECT 6.174 34.182 6.226 34.218 ;
               RECT 6.174 34.782 6.226 34.818 ;
               RECT 6.174 35.382 6.226 35.418 ;
               RECT 6.174 35.982 6.226 36.018 ;
               RECT 6.174 36.582 6.226 36.618 ;
               RECT 6.174 37.182 6.226 37.218 ;
               RECT 6.174 37.782 6.226 37.818 ;
               RECT 6.174 38.382 6.226 38.418 ;
               RECT 6.174 38.982 6.226 39.018 ;
               RECT 6.174 39.582 6.226 39.618 ;
               RECT 6.174 40.182 6.226 40.218 ;
               RECT 6.174 40.782 6.226 40.818 ;
               RECT 6.174 41.382 6.226 41.418 ;
               RECT 6.174 41.982 6.226 42.018 ;
               RECT 6.174 42.582 6.226 42.618 ;
               RECT 6.174 43.182 6.226 43.218 ;
               RECT 6.174 43.782 6.226 43.818 ;
               RECT 6.174 44.382 6.226 44.418 ;
               RECT 6.174 44.982 6.226 45.018 ;
               RECT 6.174 45.582 6.226 45.618 ;
               RECT 6.174 46.182 6.226 46.218 ;
               RECT 6.174 46.782 6.226 46.818 ;
               RECT 6.174 47.382 6.226 47.418 ;
               RECT 6.174 47.982 6.226 48.018 ;
               RECT 6.174 48.582 6.226 48.618 ;
               RECT 6.174 48.942 6.226 48.978 ;
               RECT 6.174 49.182 6.226 49.218 ;
               RECT 6.174 49.902 6.226 49.938 ;
               RECT 6.174 50.622 6.226 50.658 ;
               RECT 6.174 50.862 6.226 50.898 ;
               RECT 6.174 51.342 6.226 51.378 ;
               RECT 6.174 51.822 6.226 51.858 ;
               RECT 6.174 52.302 6.226 52.338 ;
               RECT 6.174 52.782 6.226 52.818 ;
               RECT 6.174 53.262 6.226 53.298 ;
               RECT 6.174 53.742 6.226 53.778 ;
               RECT 6.174 54.222 6.226 54.258 ;
               RECT 6.174 54.462 6.226 54.498 ;
               RECT 6.174 55.182 6.226 55.218 ;
               RECT 6.174 55.902 6.226 55.938 ;
               RECT 6.174 56.142 6.226 56.178 ;
               RECT 6.174 56.502 6.226 56.538 ;
               RECT 6.174 57.102 6.226 57.138 ;
               RECT 6.174 57.702 6.226 57.738 ;
               RECT 6.174 58.302 6.226 58.338 ;
               RECT 6.174 58.902 6.226 58.938 ;
               RECT 6.174 59.502 6.226 59.538 ;
               RECT 6.174 60.102 6.226 60.138 ;
               RECT 6.174 60.702 6.226 60.738 ;
               RECT 6.174 61.302 6.226 61.338 ;
               RECT 6.174 61.902 6.226 61.938 ;
               RECT 6.174 62.502 6.226 62.538 ;
               RECT 6.174 63.102 6.226 63.138 ;
               RECT 6.174 63.702 6.226 63.738 ;
               RECT 6.174 64.302 6.226 64.338 ;
               RECT 6.174 64.902 6.226 64.938 ;
               RECT 6.174 65.502 6.226 65.538 ;
               RECT 6.174 66.102 6.226 66.138 ;
               RECT 6.174 66.702 6.226 66.738 ;
               RECT 6.174 67.302 6.226 67.338 ;
               RECT 6.174 67.902 6.226 67.938 ;
               RECT 6.174 68.502 6.226 68.538 ;
               RECT 6.174 69.102 6.226 69.138 ;
               RECT 6.174 69.702 6.226 69.738 ;
               RECT 6.174 70.302 6.226 70.338 ;
               RECT 6.174 70.902 6.226 70.938 ;
               RECT 6.174 71.502 6.226 71.538 ;
               RECT 6.174 72.102 6.226 72.138 ;
               RECT 6.174 72.702 6.226 72.738 ;
               RECT 6.174 73.302 6.226 73.338 ;
               RECT 6.174 73.902 6.226 73.938 ;
               RECT 6.174 74.502 6.226 74.538 ;
               RECT 6.174 75.102 6.226 75.138 ;
               RECT 6.174 75.702 6.226 75.738 ;
               RECT 6.174 76.302 6.226 76.338 ;
               RECT 6.174 76.902 6.226 76.938 ;
               RECT 6.174 77.502 6.226 77.538 ;
               RECT 6.174 78.102 6.226 78.138 ;
               RECT 6.174 78.702 6.226 78.738 ;
               RECT 6.174 79.302 6.226 79.338 ;
               RECT 6.174 79.902 6.226 79.938 ;
               RECT 6.174 80.502 6.226 80.538 ;
               RECT 6.174 81.102 6.226 81.138 ;
               RECT 6.174 81.702 6.226 81.738 ;
               RECT 6.174 82.302 6.226 82.338 ;
               RECT 6.174 82.902 6.226 82.938 ;
               RECT 6.174 83.502 6.226 83.538 ;
               RECT 6.174 84.102 6.226 84.138 ;
               RECT 6.174 84.702 6.226 84.738 ;
               RECT 6.174 85.302 6.226 85.338 ;
               RECT 6.174 85.902 6.226 85.938 ;
               RECT 6.174 86.502 6.226 86.538 ;
               RECT 6.174 87.102 6.226 87.138 ;
               RECT 6.174 87.702 6.226 87.738 ;
               RECT 6.174 88.302 6.226 88.338 ;
               RECT 6.174 88.902 6.226 88.938 ;
               RECT 6.174 89.502 6.226 89.538 ;
               RECT 6.174 90.102 6.226 90.138 ;
               RECT 6.174 90.702 6.226 90.738 ;
               RECT 6.174 91.302 6.226 91.338 ;
               RECT 6.174 91.902 6.226 91.938 ;
               RECT 6.174 92.502 6.226 92.538 ;
               RECT 6.174 93.102 6.226 93.138 ;
               RECT 6.174 93.702 6.226 93.738 ;
               RECT 6.174 94.302 6.226 94.338 ;
               RECT 6.174 94.902 6.226 94.938 ;
               RECT 6.174 95.502 6.226 95.538 ;
               RECT 6.174 96.102 6.226 96.138 ;
               RECT 6.174 96.702 6.226 96.738 ;
               RECT 6.174 97.302 6.226 97.338 ;
               RECT 6.174 97.902 6.226 97.938 ;
               RECT 6.174 98.502 6.226 98.538 ;
               RECT 6.174 99.102 6.226 99.138 ;
               RECT 6.174 99.702 6.226 99.738 ;
               RECT 6.174 100.302 6.226 100.338 ;
               RECT 6.174 100.902 6.226 100.938 ;
               RECT 6.174 101.502 6.226 101.538 ;
               RECT 6.174 102.102 6.226 102.138 ;
               RECT 6.174 102.702 6.226 102.738 ;
               RECT 6.174 103.302 6.226 103.338 ;
               RECT 6.174 103.902 6.226 103.938 ;
               RECT 6.174 104.502 6.226 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 6.974 0.5695 7.026 104.5505 ;
               LAYER v4 ;
               RECT 6.974 0.582 7.026 0.618 ;
               RECT 6.974 1.182 7.026 1.218 ;
               RECT 6.974 1.782 7.026 1.818 ;
               RECT 6.974 2.382 7.026 2.418 ;
               RECT 6.974 2.982 7.026 3.018 ;
               RECT 6.974 3.582 7.026 3.618 ;
               RECT 6.974 4.182 7.026 4.218 ;
               RECT 6.974 4.782 7.026 4.818 ;
               RECT 6.974 5.382 7.026 5.418 ;
               RECT 6.974 5.982 7.026 6.018 ;
               RECT 6.974 6.582 7.026 6.618 ;
               RECT 6.974 7.182 7.026 7.218 ;
               RECT 6.974 7.782 7.026 7.818 ;
               RECT 6.974 8.382 7.026 8.418 ;
               RECT 6.974 8.982 7.026 9.018 ;
               RECT 6.974 9.582 7.026 9.618 ;
               RECT 6.974 10.182 7.026 10.218 ;
               RECT 6.974 10.782 7.026 10.818 ;
               RECT 6.974 11.382 7.026 11.418 ;
               RECT 6.974 11.982 7.026 12.018 ;
               RECT 6.974 12.582 7.026 12.618 ;
               RECT 6.974 13.182 7.026 13.218 ;
               RECT 6.974 13.782 7.026 13.818 ;
               RECT 6.974 14.382 7.026 14.418 ;
               RECT 6.974 14.982 7.026 15.018 ;
               RECT 6.974 15.582 7.026 15.618 ;
               RECT 6.974 16.182 7.026 16.218 ;
               RECT 6.974 16.782 7.026 16.818 ;
               RECT 6.974 17.382 7.026 17.418 ;
               RECT 6.974 17.982 7.026 18.018 ;
               RECT 6.974 18.582 7.026 18.618 ;
               RECT 6.974 19.182 7.026 19.218 ;
               RECT 6.974 19.782 7.026 19.818 ;
               RECT 6.974 20.382 7.026 20.418 ;
               RECT 6.974 20.982 7.026 21.018 ;
               RECT 6.974 21.582 7.026 21.618 ;
               RECT 6.974 22.182 7.026 22.218 ;
               RECT 6.974 22.782 7.026 22.818 ;
               RECT 6.974 23.382 7.026 23.418 ;
               RECT 6.974 23.982 7.026 24.018 ;
               RECT 6.974 24.582 7.026 24.618 ;
               RECT 6.974 25.182 7.026 25.218 ;
               RECT 6.974 25.782 7.026 25.818 ;
               RECT 6.974 26.382 7.026 26.418 ;
               RECT 6.974 26.982 7.026 27.018 ;
               RECT 6.974 27.582 7.026 27.618 ;
               RECT 6.974 28.182 7.026 28.218 ;
               RECT 6.974 28.782 7.026 28.818 ;
               RECT 6.974 29.382 7.026 29.418 ;
               RECT 6.974 29.982 7.026 30.018 ;
               RECT 6.974 30.582 7.026 30.618 ;
               RECT 6.974 31.182 7.026 31.218 ;
               RECT 6.974 31.782 7.026 31.818 ;
               RECT 6.974 32.382 7.026 32.418 ;
               RECT 6.974 32.982 7.026 33.018 ;
               RECT 6.974 33.582 7.026 33.618 ;
               RECT 6.974 34.182 7.026 34.218 ;
               RECT 6.974 34.782 7.026 34.818 ;
               RECT 6.974 35.382 7.026 35.418 ;
               RECT 6.974 35.982 7.026 36.018 ;
               RECT 6.974 36.582 7.026 36.618 ;
               RECT 6.974 37.182 7.026 37.218 ;
               RECT 6.974 37.782 7.026 37.818 ;
               RECT 6.974 38.382 7.026 38.418 ;
               RECT 6.974 38.982 7.026 39.018 ;
               RECT 6.974 39.582 7.026 39.618 ;
               RECT 6.974 40.182 7.026 40.218 ;
               RECT 6.974 40.782 7.026 40.818 ;
               RECT 6.974 41.382 7.026 41.418 ;
               RECT 6.974 41.982 7.026 42.018 ;
               RECT 6.974 42.582 7.026 42.618 ;
               RECT 6.974 43.182 7.026 43.218 ;
               RECT 6.974 43.782 7.026 43.818 ;
               RECT 6.974 44.382 7.026 44.418 ;
               RECT 6.974 44.982 7.026 45.018 ;
               RECT 6.974 45.582 7.026 45.618 ;
               RECT 6.974 46.182 7.026 46.218 ;
               RECT 6.974 46.782 7.026 46.818 ;
               RECT 6.974 47.382 7.026 47.418 ;
               RECT 6.974 47.982 7.026 48.018 ;
               RECT 6.974 48.582 7.026 48.618 ;
               RECT 6.974 48.942 7.026 48.978 ;
               RECT 6.974 48.9475 7.026 48.9725 ;
               RECT 6.974 49.182 7.026 49.218 ;
               RECT 6.974 49.902 7.026 49.938 ;
               RECT 6.974 50.622 7.026 50.658 ;
               RECT 6.974 50.862 7.026 50.898 ;
               RECT 6.974 51.342 7.026 51.378 ;
               RECT 6.974 51.822 7.026 51.858 ;
               RECT 6.974 52.302 7.026 52.338 ;
               RECT 6.974 52.782 7.026 52.818 ;
               RECT 6.974 53.262 7.026 53.298 ;
               RECT 6.974 53.742 7.026 53.778 ;
               RECT 6.974 54.222 7.026 54.258 ;
               RECT 6.974 54.462 7.026 54.498 ;
               RECT 6.974 55.182 7.026 55.218 ;
               RECT 6.974 55.902 7.026 55.938 ;
               RECT 6.974 56.142 7.026 56.178 ;
               RECT 6.974 56.1475 7.026 56.1725 ;
               RECT 6.974 56.502 7.026 56.538 ;
               RECT 6.974 57.102 7.026 57.138 ;
               RECT 6.974 57.702 7.026 57.738 ;
               RECT 6.974 58.302 7.026 58.338 ;
               RECT 6.974 58.902 7.026 58.938 ;
               RECT 6.974 59.502 7.026 59.538 ;
               RECT 6.974 60.102 7.026 60.138 ;
               RECT 6.974 60.702 7.026 60.738 ;
               RECT 6.974 61.302 7.026 61.338 ;
               RECT 6.974 61.902 7.026 61.938 ;
               RECT 6.974 62.502 7.026 62.538 ;
               RECT 6.974 63.102 7.026 63.138 ;
               RECT 6.974 63.702 7.026 63.738 ;
               RECT 6.974 64.302 7.026 64.338 ;
               RECT 6.974 64.902 7.026 64.938 ;
               RECT 6.974 65.502 7.026 65.538 ;
               RECT 6.974 66.102 7.026 66.138 ;
               RECT 6.974 66.702 7.026 66.738 ;
               RECT 6.974 67.302 7.026 67.338 ;
               RECT 6.974 67.902 7.026 67.938 ;
               RECT 6.974 68.502 7.026 68.538 ;
               RECT 6.974 69.102 7.026 69.138 ;
               RECT 6.974 69.702 7.026 69.738 ;
               RECT 6.974 70.302 7.026 70.338 ;
               RECT 6.974 70.902 7.026 70.938 ;
               RECT 6.974 71.502 7.026 71.538 ;
               RECT 6.974 72.102 7.026 72.138 ;
               RECT 6.974 72.702 7.026 72.738 ;
               RECT 6.974 73.302 7.026 73.338 ;
               RECT 6.974 73.902 7.026 73.938 ;
               RECT 6.974 74.502 7.026 74.538 ;
               RECT 6.974 75.102 7.026 75.138 ;
               RECT 6.974 75.702 7.026 75.738 ;
               RECT 6.974 76.302 7.026 76.338 ;
               RECT 6.974 76.902 7.026 76.938 ;
               RECT 6.974 77.502 7.026 77.538 ;
               RECT 6.974 78.102 7.026 78.138 ;
               RECT 6.974 78.702 7.026 78.738 ;
               RECT 6.974 79.302 7.026 79.338 ;
               RECT 6.974 79.902 7.026 79.938 ;
               RECT 6.974 80.502 7.026 80.538 ;
               RECT 6.974 81.102 7.026 81.138 ;
               RECT 6.974 81.702 7.026 81.738 ;
               RECT 6.974 82.302 7.026 82.338 ;
               RECT 6.974 82.902 7.026 82.938 ;
               RECT 6.974 83.502 7.026 83.538 ;
               RECT 6.974 84.102 7.026 84.138 ;
               RECT 6.974 84.702 7.026 84.738 ;
               RECT 6.974 85.302 7.026 85.338 ;
               RECT 6.974 85.902 7.026 85.938 ;
               RECT 6.974 86.502 7.026 86.538 ;
               RECT 6.974 87.102 7.026 87.138 ;
               RECT 6.974 87.702 7.026 87.738 ;
               RECT 6.974 88.302 7.026 88.338 ;
               RECT 6.974 88.902 7.026 88.938 ;
               RECT 6.974 89.502 7.026 89.538 ;
               RECT 6.974 90.102 7.026 90.138 ;
               RECT 6.974 90.702 7.026 90.738 ;
               RECT 6.974 91.302 7.026 91.338 ;
               RECT 6.974 91.902 7.026 91.938 ;
               RECT 6.974 92.502 7.026 92.538 ;
               RECT 6.974 93.102 7.026 93.138 ;
               RECT 6.974 93.702 7.026 93.738 ;
               RECT 6.974 94.302 7.026 94.338 ;
               RECT 6.974 94.902 7.026 94.938 ;
               RECT 6.974 95.502 7.026 95.538 ;
               RECT 6.974 96.102 7.026 96.138 ;
               RECT 6.974 96.702 7.026 96.738 ;
               RECT 6.974 97.302 7.026 97.338 ;
               RECT 6.974 97.902 7.026 97.938 ;
               RECT 6.974 98.502 7.026 98.538 ;
               RECT 6.974 99.102 7.026 99.138 ;
               RECT 6.974 99.702 7.026 99.738 ;
               RECT 6.974 100.302 7.026 100.338 ;
               RECT 6.974 100.902 7.026 100.938 ;
               RECT 6.974 101.502 7.026 101.538 ;
               RECT 6.974 102.102 7.026 102.138 ;
               RECT 6.974 102.702 7.026 102.738 ;
               RECT 6.974 103.302 7.026 103.338 ;
               RECT 6.974 103.902 7.026 103.938 ;
               RECT 6.974 104.502 7.026 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 7.774 0.5695 7.826 104.5505 ;
               LAYER v4 ;
               RECT 7.774 0.582 7.826 0.618 ;
               RECT 7.774 1.182 7.826 1.218 ;
               RECT 7.774 1.782 7.826 1.818 ;
               RECT 7.774 2.382 7.826 2.418 ;
               RECT 7.774 2.982 7.826 3.018 ;
               RECT 7.774 3.582 7.826 3.618 ;
               RECT 7.774 4.182 7.826 4.218 ;
               RECT 7.774 4.782 7.826 4.818 ;
               RECT 7.774 5.382 7.826 5.418 ;
               RECT 7.774 5.982 7.826 6.018 ;
               RECT 7.774 6.582 7.826 6.618 ;
               RECT 7.774 7.182 7.826 7.218 ;
               RECT 7.774 7.782 7.826 7.818 ;
               RECT 7.774 8.382 7.826 8.418 ;
               RECT 7.774 8.982 7.826 9.018 ;
               RECT 7.774 9.582 7.826 9.618 ;
               RECT 7.774 10.182 7.826 10.218 ;
               RECT 7.774 10.782 7.826 10.818 ;
               RECT 7.774 11.382 7.826 11.418 ;
               RECT 7.774 11.982 7.826 12.018 ;
               RECT 7.774 12.582 7.826 12.618 ;
               RECT 7.774 13.182 7.826 13.218 ;
               RECT 7.774 13.782 7.826 13.818 ;
               RECT 7.774 14.382 7.826 14.418 ;
               RECT 7.774 14.982 7.826 15.018 ;
               RECT 7.774 15.582 7.826 15.618 ;
               RECT 7.774 16.182 7.826 16.218 ;
               RECT 7.774 16.782 7.826 16.818 ;
               RECT 7.774 17.382 7.826 17.418 ;
               RECT 7.774 17.982 7.826 18.018 ;
               RECT 7.774 18.582 7.826 18.618 ;
               RECT 7.774 19.182 7.826 19.218 ;
               RECT 7.774 19.782 7.826 19.818 ;
               RECT 7.774 20.382 7.826 20.418 ;
               RECT 7.774 20.982 7.826 21.018 ;
               RECT 7.774 21.582 7.826 21.618 ;
               RECT 7.774 22.182 7.826 22.218 ;
               RECT 7.774 22.782 7.826 22.818 ;
               RECT 7.774 23.382 7.826 23.418 ;
               RECT 7.774 23.982 7.826 24.018 ;
               RECT 7.774 24.582 7.826 24.618 ;
               RECT 7.774 25.182 7.826 25.218 ;
               RECT 7.774 25.782 7.826 25.818 ;
               RECT 7.774 26.382 7.826 26.418 ;
               RECT 7.774 26.982 7.826 27.018 ;
               RECT 7.774 27.582 7.826 27.618 ;
               RECT 7.774 28.182 7.826 28.218 ;
               RECT 7.774 28.782 7.826 28.818 ;
               RECT 7.774 29.382 7.826 29.418 ;
               RECT 7.774 29.982 7.826 30.018 ;
               RECT 7.774 30.582 7.826 30.618 ;
               RECT 7.774 31.182 7.826 31.218 ;
               RECT 7.774 31.782 7.826 31.818 ;
               RECT 7.774 32.382 7.826 32.418 ;
               RECT 7.774 32.982 7.826 33.018 ;
               RECT 7.774 33.582 7.826 33.618 ;
               RECT 7.774 34.182 7.826 34.218 ;
               RECT 7.774 34.782 7.826 34.818 ;
               RECT 7.774 35.382 7.826 35.418 ;
               RECT 7.774 35.982 7.826 36.018 ;
               RECT 7.774 36.582 7.826 36.618 ;
               RECT 7.774 37.182 7.826 37.218 ;
               RECT 7.774 37.782 7.826 37.818 ;
               RECT 7.774 38.382 7.826 38.418 ;
               RECT 7.774 38.982 7.826 39.018 ;
               RECT 7.774 39.582 7.826 39.618 ;
               RECT 7.774 40.182 7.826 40.218 ;
               RECT 7.774 40.782 7.826 40.818 ;
               RECT 7.774 41.382 7.826 41.418 ;
               RECT 7.774 41.982 7.826 42.018 ;
               RECT 7.774 42.582 7.826 42.618 ;
               RECT 7.774 43.182 7.826 43.218 ;
               RECT 7.774 43.782 7.826 43.818 ;
               RECT 7.774 44.382 7.826 44.418 ;
               RECT 7.774 44.982 7.826 45.018 ;
               RECT 7.774 45.582 7.826 45.618 ;
               RECT 7.774 46.182 7.826 46.218 ;
               RECT 7.774 46.782 7.826 46.818 ;
               RECT 7.774 47.382 7.826 47.418 ;
               RECT 7.774 47.982 7.826 48.018 ;
               RECT 7.774 48.582 7.826 48.618 ;
               RECT 7.774 48.942 7.826 48.978 ;
               RECT 7.774 49.182 7.826 49.218 ;
               RECT 7.774 49.902 7.826 49.938 ;
               RECT 7.774 50.622 7.826 50.658 ;
               RECT 7.774 50.862 7.826 50.898 ;
               RECT 7.774 51.342 7.826 51.378 ;
               RECT 7.774 51.822 7.826 51.858 ;
               RECT 7.774 52.302 7.826 52.338 ;
               RECT 7.774 52.782 7.826 52.818 ;
               RECT 7.774 53.262 7.826 53.298 ;
               RECT 7.774 53.742 7.826 53.778 ;
               RECT 7.774 54.222 7.826 54.258 ;
               RECT 7.774 54.462 7.826 54.498 ;
               RECT 7.774 55.182 7.826 55.218 ;
               RECT 7.774 55.902 7.826 55.938 ;
               RECT 7.774 56.142 7.826 56.178 ;
               RECT 7.774 56.502 7.826 56.538 ;
               RECT 7.774 57.102 7.826 57.138 ;
               RECT 7.774 57.702 7.826 57.738 ;
               RECT 7.774 58.302 7.826 58.338 ;
               RECT 7.774 58.902 7.826 58.938 ;
               RECT 7.774 59.502 7.826 59.538 ;
               RECT 7.774 60.102 7.826 60.138 ;
               RECT 7.774 60.702 7.826 60.738 ;
               RECT 7.774 61.302 7.826 61.338 ;
               RECT 7.774 61.902 7.826 61.938 ;
               RECT 7.774 62.502 7.826 62.538 ;
               RECT 7.774 63.102 7.826 63.138 ;
               RECT 7.774 63.702 7.826 63.738 ;
               RECT 7.774 64.302 7.826 64.338 ;
               RECT 7.774 64.902 7.826 64.938 ;
               RECT 7.774 65.502 7.826 65.538 ;
               RECT 7.774 66.102 7.826 66.138 ;
               RECT 7.774 66.702 7.826 66.738 ;
               RECT 7.774 67.302 7.826 67.338 ;
               RECT 7.774 67.902 7.826 67.938 ;
               RECT 7.774 68.502 7.826 68.538 ;
               RECT 7.774 69.102 7.826 69.138 ;
               RECT 7.774 69.702 7.826 69.738 ;
               RECT 7.774 70.302 7.826 70.338 ;
               RECT 7.774 70.902 7.826 70.938 ;
               RECT 7.774 71.502 7.826 71.538 ;
               RECT 7.774 72.102 7.826 72.138 ;
               RECT 7.774 72.702 7.826 72.738 ;
               RECT 7.774 73.302 7.826 73.338 ;
               RECT 7.774 73.902 7.826 73.938 ;
               RECT 7.774 74.502 7.826 74.538 ;
               RECT 7.774 75.102 7.826 75.138 ;
               RECT 7.774 75.702 7.826 75.738 ;
               RECT 7.774 76.302 7.826 76.338 ;
               RECT 7.774 76.902 7.826 76.938 ;
               RECT 7.774 77.502 7.826 77.538 ;
               RECT 7.774 78.102 7.826 78.138 ;
               RECT 7.774 78.702 7.826 78.738 ;
               RECT 7.774 79.302 7.826 79.338 ;
               RECT 7.774 79.902 7.826 79.938 ;
               RECT 7.774 80.502 7.826 80.538 ;
               RECT 7.774 81.102 7.826 81.138 ;
               RECT 7.774 81.702 7.826 81.738 ;
               RECT 7.774 82.302 7.826 82.338 ;
               RECT 7.774 82.902 7.826 82.938 ;
               RECT 7.774 83.502 7.826 83.538 ;
               RECT 7.774 84.102 7.826 84.138 ;
               RECT 7.774 84.702 7.826 84.738 ;
               RECT 7.774 85.302 7.826 85.338 ;
               RECT 7.774 85.902 7.826 85.938 ;
               RECT 7.774 86.502 7.826 86.538 ;
               RECT 7.774 87.102 7.826 87.138 ;
               RECT 7.774 87.702 7.826 87.738 ;
               RECT 7.774 88.302 7.826 88.338 ;
               RECT 7.774 88.902 7.826 88.938 ;
               RECT 7.774 89.502 7.826 89.538 ;
               RECT 7.774 90.102 7.826 90.138 ;
               RECT 7.774 90.702 7.826 90.738 ;
               RECT 7.774 91.302 7.826 91.338 ;
               RECT 7.774 91.902 7.826 91.938 ;
               RECT 7.774 92.502 7.826 92.538 ;
               RECT 7.774 93.102 7.826 93.138 ;
               RECT 7.774 93.702 7.826 93.738 ;
               RECT 7.774 94.302 7.826 94.338 ;
               RECT 7.774 94.902 7.826 94.938 ;
               RECT 7.774 95.502 7.826 95.538 ;
               RECT 7.774 96.102 7.826 96.138 ;
               RECT 7.774 96.702 7.826 96.738 ;
               RECT 7.774 97.302 7.826 97.338 ;
               RECT 7.774 97.902 7.826 97.938 ;
               RECT 7.774 98.502 7.826 98.538 ;
               RECT 7.774 99.102 7.826 99.138 ;
               RECT 7.774 99.702 7.826 99.738 ;
               RECT 7.774 100.302 7.826 100.338 ;
               RECT 7.774 100.902 7.826 100.938 ;
               RECT 7.774 101.502 7.826 101.538 ;
               RECT 7.774 102.102 7.826 102.138 ;
               RECT 7.774 102.702 7.826 102.738 ;
               RECT 7.774 103.302 7.826 103.338 ;
               RECT 7.774 103.902 7.826 103.938 ;
               RECT 7.774 104.502 7.826 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 8.574 0.5695 8.626 104.5505 ;
               LAYER v4 ;
               RECT 8.574 0.582 8.626 0.618 ;
               RECT 8.574 1.182 8.626 1.218 ;
               RECT 8.574 1.782 8.626 1.818 ;
               RECT 8.574 2.382 8.626 2.418 ;
               RECT 8.574 2.982 8.626 3.018 ;
               RECT 8.574 3.582 8.626 3.618 ;
               RECT 8.574 4.182 8.626 4.218 ;
               RECT 8.574 4.782 8.626 4.818 ;
               RECT 8.574 5.382 8.626 5.418 ;
               RECT 8.574 5.982 8.626 6.018 ;
               RECT 8.574 6.582 8.626 6.618 ;
               RECT 8.574 7.182 8.626 7.218 ;
               RECT 8.574 7.782 8.626 7.818 ;
               RECT 8.574 8.382 8.626 8.418 ;
               RECT 8.574 8.982 8.626 9.018 ;
               RECT 8.574 9.582 8.626 9.618 ;
               RECT 8.574 10.182 8.626 10.218 ;
               RECT 8.574 10.782 8.626 10.818 ;
               RECT 8.574 11.382 8.626 11.418 ;
               RECT 8.574 11.982 8.626 12.018 ;
               RECT 8.574 12.582 8.626 12.618 ;
               RECT 8.574 13.182 8.626 13.218 ;
               RECT 8.574 13.782 8.626 13.818 ;
               RECT 8.574 14.382 8.626 14.418 ;
               RECT 8.574 14.982 8.626 15.018 ;
               RECT 8.574 15.582 8.626 15.618 ;
               RECT 8.574 16.182 8.626 16.218 ;
               RECT 8.574 16.782 8.626 16.818 ;
               RECT 8.574 17.382 8.626 17.418 ;
               RECT 8.574 17.982 8.626 18.018 ;
               RECT 8.574 18.582 8.626 18.618 ;
               RECT 8.574 19.182 8.626 19.218 ;
               RECT 8.574 19.782 8.626 19.818 ;
               RECT 8.574 20.382 8.626 20.418 ;
               RECT 8.574 20.982 8.626 21.018 ;
               RECT 8.574 21.582 8.626 21.618 ;
               RECT 8.574 22.182 8.626 22.218 ;
               RECT 8.574 22.782 8.626 22.818 ;
               RECT 8.574 23.382 8.626 23.418 ;
               RECT 8.574 23.982 8.626 24.018 ;
               RECT 8.574 24.582 8.626 24.618 ;
               RECT 8.574 25.182 8.626 25.218 ;
               RECT 8.574 25.782 8.626 25.818 ;
               RECT 8.574 26.382 8.626 26.418 ;
               RECT 8.574 26.982 8.626 27.018 ;
               RECT 8.574 27.582 8.626 27.618 ;
               RECT 8.574 28.182 8.626 28.218 ;
               RECT 8.574 28.782 8.626 28.818 ;
               RECT 8.574 29.382 8.626 29.418 ;
               RECT 8.574 29.982 8.626 30.018 ;
               RECT 8.574 30.582 8.626 30.618 ;
               RECT 8.574 31.182 8.626 31.218 ;
               RECT 8.574 31.782 8.626 31.818 ;
               RECT 8.574 32.382 8.626 32.418 ;
               RECT 8.574 32.982 8.626 33.018 ;
               RECT 8.574 33.582 8.626 33.618 ;
               RECT 8.574 34.182 8.626 34.218 ;
               RECT 8.574 34.782 8.626 34.818 ;
               RECT 8.574 35.382 8.626 35.418 ;
               RECT 8.574 35.982 8.626 36.018 ;
               RECT 8.574 36.582 8.626 36.618 ;
               RECT 8.574 37.182 8.626 37.218 ;
               RECT 8.574 37.782 8.626 37.818 ;
               RECT 8.574 38.382 8.626 38.418 ;
               RECT 8.574 38.982 8.626 39.018 ;
               RECT 8.574 39.582 8.626 39.618 ;
               RECT 8.574 40.182 8.626 40.218 ;
               RECT 8.574 40.782 8.626 40.818 ;
               RECT 8.574 41.382 8.626 41.418 ;
               RECT 8.574 41.982 8.626 42.018 ;
               RECT 8.574 42.582 8.626 42.618 ;
               RECT 8.574 43.182 8.626 43.218 ;
               RECT 8.574 43.782 8.626 43.818 ;
               RECT 8.574 44.382 8.626 44.418 ;
               RECT 8.574 44.982 8.626 45.018 ;
               RECT 8.574 45.582 8.626 45.618 ;
               RECT 8.574 46.182 8.626 46.218 ;
               RECT 8.574 46.782 8.626 46.818 ;
               RECT 8.574 47.382 8.626 47.418 ;
               RECT 8.574 47.982 8.626 48.018 ;
               RECT 8.574 48.582 8.626 48.618 ;
               RECT 8.574 48.942 8.626 48.978 ;
               RECT 8.574 48.9475 8.626 48.9725 ;
               RECT 8.574 49.182 8.626 49.218 ;
               RECT 8.574 49.902 8.626 49.938 ;
               RECT 8.574 50.622 8.626 50.658 ;
               RECT 8.574 50.862 8.626 50.898 ;
               RECT 8.574 51.342 8.626 51.378 ;
               RECT 8.574 51.822 8.626 51.858 ;
               RECT 8.574 52.302 8.626 52.338 ;
               RECT 8.574 52.782 8.626 52.818 ;
               RECT 8.574 53.262 8.626 53.298 ;
               RECT 8.574 53.742 8.626 53.778 ;
               RECT 8.574 54.222 8.626 54.258 ;
               RECT 8.574 54.462 8.626 54.498 ;
               RECT 8.574 55.182 8.626 55.218 ;
               RECT 8.574 55.902 8.626 55.938 ;
               RECT 8.574 56.142 8.626 56.178 ;
               RECT 8.574 56.1475 8.626 56.1725 ;
               RECT 8.574 56.502 8.626 56.538 ;
               RECT 8.574 57.102 8.626 57.138 ;
               RECT 8.574 57.702 8.626 57.738 ;
               RECT 8.574 58.302 8.626 58.338 ;
               RECT 8.574 58.902 8.626 58.938 ;
               RECT 8.574 59.502 8.626 59.538 ;
               RECT 8.574 60.102 8.626 60.138 ;
               RECT 8.574 60.702 8.626 60.738 ;
               RECT 8.574 61.302 8.626 61.338 ;
               RECT 8.574 61.902 8.626 61.938 ;
               RECT 8.574 62.502 8.626 62.538 ;
               RECT 8.574 63.102 8.626 63.138 ;
               RECT 8.574 63.702 8.626 63.738 ;
               RECT 8.574 64.302 8.626 64.338 ;
               RECT 8.574 64.902 8.626 64.938 ;
               RECT 8.574 65.502 8.626 65.538 ;
               RECT 8.574 66.102 8.626 66.138 ;
               RECT 8.574 66.702 8.626 66.738 ;
               RECT 8.574 67.302 8.626 67.338 ;
               RECT 8.574 67.902 8.626 67.938 ;
               RECT 8.574 68.502 8.626 68.538 ;
               RECT 8.574 69.102 8.626 69.138 ;
               RECT 8.574 69.702 8.626 69.738 ;
               RECT 8.574 70.302 8.626 70.338 ;
               RECT 8.574 70.902 8.626 70.938 ;
               RECT 8.574 71.502 8.626 71.538 ;
               RECT 8.574 72.102 8.626 72.138 ;
               RECT 8.574 72.702 8.626 72.738 ;
               RECT 8.574 73.302 8.626 73.338 ;
               RECT 8.574 73.902 8.626 73.938 ;
               RECT 8.574 74.502 8.626 74.538 ;
               RECT 8.574 75.102 8.626 75.138 ;
               RECT 8.574 75.702 8.626 75.738 ;
               RECT 8.574 76.302 8.626 76.338 ;
               RECT 8.574 76.902 8.626 76.938 ;
               RECT 8.574 77.502 8.626 77.538 ;
               RECT 8.574 78.102 8.626 78.138 ;
               RECT 8.574 78.702 8.626 78.738 ;
               RECT 8.574 79.302 8.626 79.338 ;
               RECT 8.574 79.902 8.626 79.938 ;
               RECT 8.574 80.502 8.626 80.538 ;
               RECT 8.574 81.102 8.626 81.138 ;
               RECT 8.574 81.702 8.626 81.738 ;
               RECT 8.574 82.302 8.626 82.338 ;
               RECT 8.574 82.902 8.626 82.938 ;
               RECT 8.574 83.502 8.626 83.538 ;
               RECT 8.574 84.102 8.626 84.138 ;
               RECT 8.574 84.702 8.626 84.738 ;
               RECT 8.574 85.302 8.626 85.338 ;
               RECT 8.574 85.902 8.626 85.938 ;
               RECT 8.574 86.502 8.626 86.538 ;
               RECT 8.574 87.102 8.626 87.138 ;
               RECT 8.574 87.702 8.626 87.738 ;
               RECT 8.574 88.302 8.626 88.338 ;
               RECT 8.574 88.902 8.626 88.938 ;
               RECT 8.574 89.502 8.626 89.538 ;
               RECT 8.574 90.102 8.626 90.138 ;
               RECT 8.574 90.702 8.626 90.738 ;
               RECT 8.574 91.302 8.626 91.338 ;
               RECT 8.574 91.902 8.626 91.938 ;
               RECT 8.574 92.502 8.626 92.538 ;
               RECT 8.574 93.102 8.626 93.138 ;
               RECT 8.574 93.702 8.626 93.738 ;
               RECT 8.574 94.302 8.626 94.338 ;
               RECT 8.574 94.902 8.626 94.938 ;
               RECT 8.574 95.502 8.626 95.538 ;
               RECT 8.574 96.102 8.626 96.138 ;
               RECT 8.574 96.702 8.626 96.738 ;
               RECT 8.574 97.302 8.626 97.338 ;
               RECT 8.574 97.902 8.626 97.938 ;
               RECT 8.574 98.502 8.626 98.538 ;
               RECT 8.574 99.102 8.626 99.138 ;
               RECT 8.574 99.702 8.626 99.738 ;
               RECT 8.574 100.302 8.626 100.338 ;
               RECT 8.574 100.902 8.626 100.938 ;
               RECT 8.574 101.502 8.626 101.538 ;
               RECT 8.574 102.102 8.626 102.138 ;
               RECT 8.574 102.702 8.626 102.738 ;
               RECT 8.574 103.302 8.626 103.338 ;
               RECT 8.574 103.902 8.626 103.938 ;
               RECT 8.574 104.502 8.626 104.538 ;
          END
          PORT
               LAYER m5 ;
               RECT 9.374 0.5695 9.426 104.5505 ;
               LAYER v4 ;
               RECT 9.374 0.582 9.426 0.618 ;
               RECT 9.374 1.182 9.426 1.218 ;
               RECT 9.374 1.782 9.426 1.818 ;
               RECT 9.374 2.382 9.426 2.418 ;
               RECT 9.374 2.982 9.426 3.018 ;
               RECT 9.374 3.582 9.426 3.618 ;
               RECT 9.374 4.182 9.426 4.218 ;
               RECT 9.374 4.782 9.426 4.818 ;
               RECT 9.374 5.382 9.426 5.418 ;
               RECT 9.374 5.982 9.426 6.018 ;
               RECT 9.374 6.582 9.426 6.618 ;
               RECT 9.374 7.182 9.426 7.218 ;
               RECT 9.374 7.782 9.426 7.818 ;
               RECT 9.374 8.382 9.426 8.418 ;
               RECT 9.374 8.982 9.426 9.018 ;
               RECT 9.374 9.582 9.426 9.618 ;
               RECT 9.374 10.182 9.426 10.218 ;
               RECT 9.374 10.782 9.426 10.818 ;
               RECT 9.374 11.382 9.426 11.418 ;
               RECT 9.374 11.982 9.426 12.018 ;
               RECT 9.374 12.582 9.426 12.618 ;
               RECT 9.374 13.182 9.426 13.218 ;
               RECT 9.374 13.782 9.426 13.818 ;
               RECT 9.374 14.382 9.426 14.418 ;
               RECT 9.374 14.982 9.426 15.018 ;
               RECT 9.374 15.582 9.426 15.618 ;
               RECT 9.374 16.182 9.426 16.218 ;
               RECT 9.374 16.782 9.426 16.818 ;
               RECT 9.374 17.382 9.426 17.418 ;
               RECT 9.374 17.982 9.426 18.018 ;
               RECT 9.374 18.582 9.426 18.618 ;
               RECT 9.374 19.182 9.426 19.218 ;
               RECT 9.374 19.782 9.426 19.818 ;
               RECT 9.374 20.382 9.426 20.418 ;
               RECT 9.374 20.982 9.426 21.018 ;
               RECT 9.374 21.582 9.426 21.618 ;
               RECT 9.374 22.182 9.426 22.218 ;
               RECT 9.374 22.782 9.426 22.818 ;
               RECT 9.374 23.382 9.426 23.418 ;
               RECT 9.374 23.982 9.426 24.018 ;
               RECT 9.374 24.582 9.426 24.618 ;
               RECT 9.374 25.182 9.426 25.218 ;
               RECT 9.374 25.782 9.426 25.818 ;
               RECT 9.374 26.382 9.426 26.418 ;
               RECT 9.374 26.982 9.426 27.018 ;
               RECT 9.374 27.582 9.426 27.618 ;
               RECT 9.374 28.182 9.426 28.218 ;
               RECT 9.374 28.782 9.426 28.818 ;
               RECT 9.374 29.382 9.426 29.418 ;
               RECT 9.374 29.982 9.426 30.018 ;
               RECT 9.374 30.582 9.426 30.618 ;
               RECT 9.374 31.182 9.426 31.218 ;
               RECT 9.374 31.782 9.426 31.818 ;
               RECT 9.374 32.382 9.426 32.418 ;
               RECT 9.374 32.982 9.426 33.018 ;
               RECT 9.374 33.582 9.426 33.618 ;
               RECT 9.374 34.182 9.426 34.218 ;
               RECT 9.374 34.782 9.426 34.818 ;
               RECT 9.374 35.382 9.426 35.418 ;
               RECT 9.374 35.982 9.426 36.018 ;
               RECT 9.374 36.582 9.426 36.618 ;
               RECT 9.374 37.182 9.426 37.218 ;
               RECT 9.374 37.782 9.426 37.818 ;
               RECT 9.374 38.382 9.426 38.418 ;
               RECT 9.374 38.982 9.426 39.018 ;
               RECT 9.374 39.582 9.426 39.618 ;
               RECT 9.374 40.182 9.426 40.218 ;
               RECT 9.374 40.782 9.426 40.818 ;
               RECT 9.374 41.382 9.426 41.418 ;
               RECT 9.374 41.982 9.426 42.018 ;
               RECT 9.374 42.582 9.426 42.618 ;
               RECT 9.374 43.182 9.426 43.218 ;
               RECT 9.374 43.782 9.426 43.818 ;
               RECT 9.374 44.382 9.426 44.418 ;
               RECT 9.374 44.982 9.426 45.018 ;
               RECT 9.374 45.582 9.426 45.618 ;
               RECT 9.374 46.182 9.426 46.218 ;
               RECT 9.374 46.782 9.426 46.818 ;
               RECT 9.374 47.382 9.426 47.418 ;
               RECT 9.374 47.982 9.426 48.018 ;
               RECT 9.374 48.582 9.426 48.618 ;
               RECT 9.374 48.942 9.426 48.978 ;
               RECT 9.374 49.182 9.426 49.218 ;
               RECT 9.374 49.902 9.426 49.938 ;
               RECT 9.374 50.622 9.426 50.658 ;
               RECT 9.374 50.862 9.426 50.898 ;
               RECT 9.374 51.342 9.426 51.378 ;
               RECT 9.374 51.822 9.426 51.858 ;
               RECT 9.374 52.302 9.426 52.338 ;
               RECT 9.374 52.782 9.426 52.818 ;
               RECT 9.374 53.262 9.426 53.298 ;
               RECT 9.374 53.742 9.426 53.778 ;
               RECT 9.374 54.222 9.426 54.258 ;
               RECT 9.374 54.462 9.426 54.498 ;
               RECT 9.374 55.182 9.426 55.218 ;
               RECT 9.374 55.902 9.426 55.938 ;
               RECT 9.374 56.142 9.426 56.178 ;
               RECT 9.374 56.502 9.426 56.538 ;
               RECT 9.374 57.102 9.426 57.138 ;
               RECT 9.374 57.702 9.426 57.738 ;
               RECT 9.374 58.302 9.426 58.338 ;
               RECT 9.374 58.902 9.426 58.938 ;
               RECT 9.374 59.502 9.426 59.538 ;
               RECT 9.374 60.102 9.426 60.138 ;
               RECT 9.374 60.702 9.426 60.738 ;
               RECT 9.374 61.302 9.426 61.338 ;
               RECT 9.374 61.902 9.426 61.938 ;
               RECT 9.374 62.502 9.426 62.538 ;
               RECT 9.374 63.102 9.426 63.138 ;
               RECT 9.374 63.702 9.426 63.738 ;
               RECT 9.374 64.302 9.426 64.338 ;
               RECT 9.374 64.902 9.426 64.938 ;
               RECT 9.374 65.502 9.426 65.538 ;
               RECT 9.374 66.102 9.426 66.138 ;
               RECT 9.374 66.702 9.426 66.738 ;
               RECT 9.374 67.302 9.426 67.338 ;
               RECT 9.374 67.902 9.426 67.938 ;
               RECT 9.374 68.502 9.426 68.538 ;
               RECT 9.374 69.102 9.426 69.138 ;
               RECT 9.374 69.702 9.426 69.738 ;
               RECT 9.374 70.302 9.426 70.338 ;
               RECT 9.374 70.902 9.426 70.938 ;
               RECT 9.374 71.502 9.426 71.538 ;
               RECT 9.374 72.102 9.426 72.138 ;
               RECT 9.374 72.702 9.426 72.738 ;
               RECT 9.374 73.302 9.426 73.338 ;
               RECT 9.374 73.902 9.426 73.938 ;
               RECT 9.374 74.502 9.426 74.538 ;
               RECT 9.374 75.102 9.426 75.138 ;
               RECT 9.374 75.702 9.426 75.738 ;
               RECT 9.374 76.302 9.426 76.338 ;
               RECT 9.374 76.902 9.426 76.938 ;
               RECT 9.374 77.502 9.426 77.538 ;
               RECT 9.374 78.102 9.426 78.138 ;
               RECT 9.374 78.702 9.426 78.738 ;
               RECT 9.374 79.302 9.426 79.338 ;
               RECT 9.374 79.902 9.426 79.938 ;
               RECT 9.374 80.502 9.426 80.538 ;
               RECT 9.374 81.102 9.426 81.138 ;
               RECT 9.374 81.702 9.426 81.738 ;
               RECT 9.374 82.302 9.426 82.338 ;
               RECT 9.374 82.902 9.426 82.938 ;
               RECT 9.374 83.502 9.426 83.538 ;
               RECT 9.374 84.102 9.426 84.138 ;
               RECT 9.374 84.702 9.426 84.738 ;
               RECT 9.374 85.302 9.426 85.338 ;
               RECT 9.374 85.902 9.426 85.938 ;
               RECT 9.374 86.502 9.426 86.538 ;
               RECT 9.374 87.102 9.426 87.138 ;
               RECT 9.374 87.702 9.426 87.738 ;
               RECT 9.374 88.302 9.426 88.338 ;
               RECT 9.374 88.902 9.426 88.938 ;
               RECT 9.374 89.502 9.426 89.538 ;
               RECT 9.374 90.102 9.426 90.138 ;
               RECT 9.374 90.702 9.426 90.738 ;
               RECT 9.374 91.302 9.426 91.338 ;
               RECT 9.374 91.902 9.426 91.938 ;
               RECT 9.374 92.502 9.426 92.538 ;
               RECT 9.374 93.102 9.426 93.138 ;
               RECT 9.374 93.702 9.426 93.738 ;
               RECT 9.374 94.302 9.426 94.338 ;
               RECT 9.374 94.902 9.426 94.938 ;
               RECT 9.374 95.502 9.426 95.538 ;
               RECT 9.374 96.102 9.426 96.138 ;
               RECT 9.374 96.702 9.426 96.738 ;
               RECT 9.374 97.302 9.426 97.338 ;
               RECT 9.374 97.902 9.426 97.938 ;
               RECT 9.374 98.502 9.426 98.538 ;
               RECT 9.374 99.102 9.426 99.138 ;
               RECT 9.374 99.702 9.426 99.738 ;
               RECT 9.374 100.302 9.426 100.338 ;
               RECT 9.374 100.902 9.426 100.938 ;
               RECT 9.374 101.502 9.426 101.538 ;
               RECT 9.374 102.102 9.426 102.138 ;
               RECT 9.374 102.702 9.426 102.738 ;
               RECT 9.374 103.302 9.426 103.338 ;
               RECT 9.374 103.902 9.426 103.938 ;
               RECT 9.374 104.502 9.426 104.538 ;
          END
     END vss
     OBS
          LAYER m0 ;
               RECT 0 0 36.3 105.12 ;
          LAYER m1 ;
               RECT 0 0 36.3 105.12 ;
          LAYER m2 SPACING 0 ;
               RECT -0.0705 -0.038 36.3705 105.158 ;
          LAYER m3 SPACING 0 ;
               RECT -0.035 -0.07 36.335 105.19 ;
          LAYER m4 SPACING 0 ;
               RECT -0.07 -0.038 36.37 105.158 ;
          LAYER m5 SPACING 0 ;
               RECT -0.059 -0.09 36.359 105.21 ;
          LAYER v4 ;
               RECT 0.574 0.281 0.626 0.317 ;
               RECT 0.574 104.803 0.626 104.839 ;
               RECT 0.654 0.806 0.706 0.842 ;
               RECT 0.654 2.006 0.706 2.042 ;
               RECT 0.654 3.206 0.706 3.242 ;
               RECT 0.654 4.406 0.706 4.442 ;
               RECT 0.654 5.606 0.706 5.642 ;
               RECT 0.654 6.806 0.706 6.842 ;
               RECT 0.654 8.006 0.706 8.042 ;
               RECT 0.654 9.206 0.706 9.242 ;
               RECT 0.654 10.406 0.706 10.442 ;
               RECT 0.654 11.606 0.706 11.642 ;
               RECT 0.654 12.806 0.706 12.842 ;
               RECT 0.654 14.006 0.706 14.042 ;
               RECT 0.654 15.206 0.706 15.242 ;
               RECT 0.654 16.406 0.706 16.442 ;
               RECT 0.654 17.606 0.706 17.642 ;
               RECT 0.654 18.806 0.706 18.842 ;
               RECT 0.654 20.006 0.706 20.042 ;
               RECT 0.654 21.206 0.706 21.242 ;
               RECT 0.654 22.406 0.706 22.442 ;
               RECT 0.654 23.606 0.706 23.642 ;
               RECT 0.654 24.806 0.706 24.842 ;
               RECT 0.654 26.006 0.706 26.042 ;
               RECT 0.654 27.206 0.706 27.242 ;
               RECT 0.654 28.406 0.706 28.442 ;
               RECT 0.654 29.606 0.706 29.642 ;
               RECT 0.654 30.806 0.706 30.842 ;
               RECT 0.654 32.006 0.706 32.042 ;
               RECT 0.654 33.206 0.706 33.242 ;
               RECT 0.654 34.406 0.706 34.442 ;
               RECT 0.654 35.606 0.706 35.642 ;
               RECT 0.654 36.806 0.706 36.842 ;
               RECT 0.654 38.006 0.706 38.042 ;
               RECT 0.654 39.206 0.706 39.242 ;
               RECT 0.654 40.406 0.706 40.442 ;
               RECT 0.654 41.606 0.706 41.642 ;
               RECT 0.654 42.806 0.706 42.842 ;
               RECT 0.654 44.006 0.706 44.042 ;
               RECT 0.654 45.206 0.706 45.242 ;
               RECT 0.654 46.406 0.706 46.442 ;
               RECT 0.654 47.606 0.706 47.642 ;
               RECT 0.654 49.422 0.706 49.458 ;
               RECT 0.654 49.662 0.706 49.698 ;
               RECT 0.654 55.422 0.706 55.458 ;
               RECT 0.654 55.662 0.706 55.698 ;
               RECT 0.654 56.726 0.706 56.762 ;
               RECT 0.654 57.926 0.706 57.962 ;
               RECT 0.654 59.126 0.706 59.162 ;
               RECT 0.654 60.326 0.706 60.362 ;
               RECT 0.654 61.526 0.706 61.562 ;
               RECT 0.654 62.726 0.706 62.762 ;
               RECT 0.654 63.926 0.706 63.962 ;
               RECT 0.654 65.126 0.706 65.162 ;
               RECT 0.654 66.326 0.706 66.362 ;
               RECT 0.654 67.526 0.706 67.562 ;
               RECT 0.654 68.726 0.706 68.762 ;
               RECT 0.654 69.926 0.706 69.962 ;
               RECT 0.654 71.126 0.706 71.162 ;
               RECT 0.654 72.326 0.706 72.362 ;
               RECT 0.654 73.526 0.706 73.562 ;
               RECT 0.654 74.726 0.706 74.762 ;
               RECT 0.654 75.926 0.706 75.962 ;
               RECT 0.654 77.126 0.706 77.162 ;
               RECT 0.654 78.326 0.706 78.362 ;
               RECT 0.654 79.526 0.706 79.562 ;
               RECT 0.654 80.726 0.706 80.762 ;
               RECT 0.654 81.926 0.706 81.962 ;
               RECT 0.654 83.126 0.706 83.162 ;
               RECT 0.654 84.326 0.706 84.362 ;
               RECT 0.654 85.526 0.706 85.562 ;
               RECT 0.654 86.726 0.706 86.762 ;
               RECT 0.654 87.926 0.706 87.962 ;
               RECT 0.654 89.126 0.706 89.162 ;
               RECT 0.654 90.326 0.706 90.362 ;
               RECT 0.654 91.526 0.706 91.562 ;
               RECT 0.654 92.726 0.706 92.762 ;
               RECT 0.654 93.926 0.706 93.962 ;
               RECT 0.654 95.126 0.706 95.162 ;
               RECT 0.654 96.326 0.706 96.362 ;
               RECT 0.654 97.526 0.706 97.562 ;
               RECT 0.654 98.726 0.706 98.762 ;
               RECT 0.654 99.926 0.706 99.962 ;
               RECT 0.654 101.126 0.706 101.162 ;
               RECT 0.654 102.326 0.706 102.362 ;
               RECT 0.654 103.526 0.706 103.562 ;
               RECT 0.734 1.558 0.786 1.594 ;
               RECT 0.734 2.758 0.786 2.794 ;
               RECT 0.734 3.958 0.786 3.994 ;
               RECT 0.734 5.158 0.786 5.194 ;
               RECT 0.734 6.358 0.786 6.394 ;
               RECT 0.734 7.558 0.786 7.594 ;
               RECT 0.734 8.758 0.786 8.794 ;
               RECT 0.734 9.958 0.786 9.994 ;
               RECT 0.734 11.158 0.786 11.194 ;
               RECT 0.734 12.358 0.786 12.394 ;
               RECT 0.734 13.558 0.786 13.594 ;
               RECT 0.734 14.758 0.786 14.794 ;
               RECT 0.734 15.958 0.786 15.994 ;
               RECT 0.734 17.158 0.786 17.194 ;
               RECT 0.734 18.358 0.786 18.394 ;
               RECT 0.734 19.558 0.786 19.594 ;
               RECT 0.734 20.758 0.786 20.794 ;
               RECT 0.734 21.958 0.786 21.994 ;
               RECT 0.734 23.158 0.786 23.194 ;
               RECT 0.734 24.358 0.786 24.394 ;
               RECT 0.734 25.558 0.786 25.594 ;
               RECT 0.734 26.758 0.786 26.794 ;
               RECT 0.734 27.958 0.786 27.994 ;
               RECT 0.734 29.158 0.786 29.194 ;
               RECT 0.734 30.358 0.786 30.394 ;
               RECT 0.734 31.558 0.786 31.594 ;
               RECT 0.734 32.758 0.786 32.794 ;
               RECT 0.734 33.958 0.786 33.994 ;
               RECT 0.734 35.158 0.786 35.194 ;
               RECT 0.734 36.358 0.786 36.394 ;
               RECT 0.734 37.558 0.786 37.594 ;
               RECT 0.734 38.758 0.786 38.794 ;
               RECT 0.734 39.958 0.786 39.994 ;
               RECT 0.734 41.158 0.786 41.194 ;
               RECT 0.734 42.358 0.786 42.394 ;
               RECT 0.734 43.558 0.786 43.594 ;
               RECT 0.734 44.758 0.786 44.794 ;
               RECT 0.734 45.958 0.786 45.994 ;
               RECT 0.734 47.158 0.786 47.194 ;
               RECT 0.734 48.358 0.786 48.394 ;
               RECT 0.734 50.142 0.786 50.178 ;
               RECT 0.734 50.382 0.786 50.418 ;
               RECT 0.734 54.702 0.786 54.738 ;
               RECT 0.734 54.942 0.786 54.978 ;
               RECT 0.734 57.478 0.786 57.514 ;
               RECT 0.734 58.678 0.786 58.714 ;
               RECT 0.734 59.878 0.786 59.914 ;
               RECT 0.734 61.078 0.786 61.114 ;
               RECT 0.734 62.278 0.786 62.314 ;
               RECT 0.734 63.478 0.786 63.514 ;
               RECT 0.734 64.678 0.786 64.714 ;
               RECT 0.734 65.878 0.786 65.914 ;
               RECT 0.734 67.078 0.786 67.114 ;
               RECT 0.734 68.278 0.786 68.314 ;
               RECT 0.734 69.478 0.786 69.514 ;
               RECT 0.734 70.678 0.786 70.714 ;
               RECT 0.734 71.878 0.786 71.914 ;
               RECT 0.734 73.078 0.786 73.114 ;
               RECT 0.734 74.278 0.786 74.314 ;
               RECT 0.734 75.478 0.786 75.514 ;
               RECT 0.734 76.678 0.786 76.714 ;
               RECT 0.734 77.878 0.786 77.914 ;
               RECT 0.734 79.078 0.786 79.114 ;
               RECT 0.734 80.278 0.786 80.314 ;
               RECT 0.734 81.478 0.786 81.514 ;
               RECT 0.734 82.678 0.786 82.714 ;
               RECT 0.734 83.878 0.786 83.914 ;
               RECT 0.734 85.078 0.786 85.114 ;
               RECT 0.734 86.278 0.786 86.314 ;
               RECT 0.734 87.478 0.786 87.514 ;
               RECT 0.734 88.678 0.786 88.714 ;
               RECT 0.734 89.878 0.786 89.914 ;
               RECT 0.734 91.078 0.786 91.114 ;
               RECT 0.734 92.278 0.786 92.314 ;
               RECT 0.734 93.478 0.786 93.514 ;
               RECT 0.734 94.678 0.786 94.714 ;
               RECT 0.734 95.878 0.786 95.914 ;
               RECT 0.734 97.078 0.786 97.114 ;
               RECT 0.734 98.278 0.786 98.314 ;
               RECT 0.734 99.478 0.786 99.514 ;
               RECT 0.734 100.678 0.786 100.714 ;
               RECT 0.734 101.878 0.786 101.914 ;
               RECT 0.734 103.078 0.786 103.114 ;
               RECT 0.734 104.278 0.786 104.314 ;
               RECT 0.814 0.806 0.866 0.842 ;
               RECT 0.814 2.006 0.866 2.042 ;
               RECT 0.814 3.206 0.866 3.242 ;
               RECT 0.814 4.406 0.866 4.442 ;
               RECT 0.814 5.606 0.866 5.642 ;
               RECT 0.814 6.806 0.866 6.842 ;
               RECT 0.814 8.006 0.866 8.042 ;
               RECT 0.814 9.206 0.866 9.242 ;
               RECT 0.814 10.406 0.866 10.442 ;
               RECT 0.814 11.606 0.866 11.642 ;
               RECT 0.814 12.806 0.866 12.842 ;
               RECT 0.814 14.006 0.866 14.042 ;
               RECT 0.814 15.206 0.866 15.242 ;
               RECT 0.814 16.406 0.866 16.442 ;
               RECT 0.814 17.606 0.866 17.642 ;
               RECT 0.814 18.806 0.866 18.842 ;
               RECT 0.814 20.006 0.866 20.042 ;
               RECT 0.814 21.206 0.866 21.242 ;
               RECT 0.814 22.406 0.866 22.442 ;
               RECT 0.814 23.606 0.866 23.642 ;
               RECT 0.814 24.806 0.866 24.842 ;
               RECT 0.814 26.006 0.866 26.042 ;
               RECT 0.814 27.206 0.866 27.242 ;
               RECT 0.814 28.406 0.866 28.442 ;
               RECT 0.814 29.606 0.866 29.642 ;
               RECT 0.814 30.806 0.866 30.842 ;
               RECT 0.814 32.006 0.866 32.042 ;
               RECT 0.814 33.206 0.866 33.242 ;
               RECT 0.814 34.406 0.866 34.442 ;
               RECT 0.814 35.606 0.866 35.642 ;
               RECT 0.814 36.806 0.866 36.842 ;
               RECT 0.814 38.006 0.866 38.042 ;
               RECT 0.814 39.206 0.866 39.242 ;
               RECT 0.814 40.406 0.866 40.442 ;
               RECT 0.814 41.606 0.866 41.642 ;
               RECT 0.814 42.806 0.866 42.842 ;
               RECT 0.814 44.006 0.866 44.042 ;
               RECT 0.814 45.206 0.866 45.242 ;
               RECT 0.814 46.406 0.866 46.442 ;
               RECT 0.814 47.606 0.866 47.642 ;
               RECT 0.814 49.422 0.866 49.458 ;
               RECT 0.814 49.662 0.866 49.698 ;
               RECT 0.814 55.422 0.866 55.458 ;
               RECT 0.814 55.662 0.866 55.698 ;
               RECT 0.814 56.726 0.866 56.762 ;
               RECT 0.814 57.926 0.866 57.962 ;
               RECT 0.814 59.126 0.866 59.162 ;
               RECT 0.814 60.326 0.866 60.362 ;
               RECT 0.814 61.526 0.866 61.562 ;
               RECT 0.814 62.726 0.866 62.762 ;
               RECT 0.814 63.926 0.866 63.962 ;
               RECT 0.814 65.126 0.866 65.162 ;
               RECT 0.814 66.326 0.866 66.362 ;
               RECT 0.814 67.526 0.866 67.562 ;
               RECT 0.814 68.726 0.866 68.762 ;
               RECT 0.814 69.926 0.866 69.962 ;
               RECT 0.814 71.126 0.866 71.162 ;
               RECT 0.814 72.326 0.866 72.362 ;
               RECT 0.814 73.526 0.866 73.562 ;
               RECT 0.814 74.726 0.866 74.762 ;
               RECT 0.814 75.926 0.866 75.962 ;
               RECT 0.814 77.126 0.866 77.162 ;
               RECT 0.814 78.326 0.866 78.362 ;
               RECT 0.814 79.526 0.866 79.562 ;
               RECT 0.814 80.726 0.866 80.762 ;
               RECT 0.814 81.926 0.866 81.962 ;
               RECT 0.814 83.126 0.866 83.162 ;
               RECT 0.814 84.326 0.866 84.362 ;
               RECT 0.814 85.526 0.866 85.562 ;
               RECT 0.814 86.726 0.866 86.762 ;
               RECT 0.814 87.926 0.866 87.962 ;
               RECT 0.814 89.126 0.866 89.162 ;
               RECT 0.814 90.326 0.866 90.362 ;
               RECT 0.814 91.526 0.866 91.562 ;
               RECT 0.814 92.726 0.866 92.762 ;
               RECT 0.814 93.926 0.866 93.962 ;
               RECT 0.814 95.126 0.866 95.162 ;
               RECT 0.814 96.326 0.866 96.362 ;
               RECT 0.814 97.526 0.866 97.562 ;
               RECT 0.814 98.726 0.866 98.762 ;
               RECT 0.814 99.926 0.866 99.962 ;
               RECT 0.814 101.126 0.866 101.162 ;
               RECT 0.814 102.326 0.866 102.362 ;
               RECT 0.814 103.526 0.866 103.562 ;
               RECT 0.894 1.558 0.946 1.594 ;
               RECT 0.894 2.758 0.946 2.794 ;
               RECT 0.894 3.958 0.946 3.994 ;
               RECT 0.894 5.158 0.946 5.194 ;
               RECT 0.894 6.358 0.946 6.394 ;
               RECT 0.894 7.558 0.946 7.594 ;
               RECT 0.894 8.758 0.946 8.794 ;
               RECT 0.894 9.958 0.946 9.994 ;
               RECT 0.894 11.158 0.946 11.194 ;
               RECT 0.894 12.358 0.946 12.394 ;
               RECT 0.894 13.558 0.946 13.594 ;
               RECT 0.894 14.758 0.946 14.794 ;
               RECT 0.894 15.958 0.946 15.994 ;
               RECT 0.894 17.158 0.946 17.194 ;
               RECT 0.894 18.358 0.946 18.394 ;
               RECT 0.894 19.558 0.946 19.594 ;
               RECT 0.894 20.758 0.946 20.794 ;
               RECT 0.894 21.958 0.946 21.994 ;
               RECT 0.894 23.158 0.946 23.194 ;
               RECT 0.894 24.358 0.946 24.394 ;
               RECT 0.894 25.558 0.946 25.594 ;
               RECT 0.894 26.758 0.946 26.794 ;
               RECT 0.894 27.958 0.946 27.994 ;
               RECT 0.894 29.158 0.946 29.194 ;
               RECT 0.894 30.358 0.946 30.394 ;
               RECT 0.894 31.558 0.946 31.594 ;
               RECT 0.894 32.758 0.946 32.794 ;
               RECT 0.894 33.958 0.946 33.994 ;
               RECT 0.894 35.158 0.946 35.194 ;
               RECT 0.894 36.358 0.946 36.394 ;
               RECT 0.894 37.558 0.946 37.594 ;
               RECT 0.894 38.758 0.946 38.794 ;
               RECT 0.894 39.958 0.946 39.994 ;
               RECT 0.894 41.158 0.946 41.194 ;
               RECT 0.894 42.358 0.946 42.394 ;
               RECT 0.894 43.558 0.946 43.594 ;
               RECT 0.894 44.758 0.946 44.794 ;
               RECT 0.894 45.958 0.946 45.994 ;
               RECT 0.894 47.158 0.946 47.194 ;
               RECT 0.894 48.358 0.946 48.394 ;
               RECT 0.894 50.142 0.946 50.178 ;
               RECT 0.894 50.382 0.946 50.418 ;
               RECT 0.894 54.702 0.946 54.738 ;
               RECT 0.894 54.942 0.946 54.978 ;
               RECT 0.894 57.478 0.946 57.514 ;
               RECT 0.894 58.678 0.946 58.714 ;
               RECT 0.894 59.878 0.946 59.914 ;
               RECT 0.894 61.078 0.946 61.114 ;
               RECT 0.894 62.278 0.946 62.314 ;
               RECT 0.894 63.478 0.946 63.514 ;
               RECT 0.894 64.678 0.946 64.714 ;
               RECT 0.894 65.878 0.946 65.914 ;
               RECT 0.894 67.078 0.946 67.114 ;
               RECT 0.894 68.278 0.946 68.314 ;
               RECT 0.894 69.478 0.946 69.514 ;
               RECT 0.894 70.678 0.946 70.714 ;
               RECT 0.894 71.878 0.946 71.914 ;
               RECT 0.894 73.078 0.946 73.114 ;
               RECT 0.894 74.278 0.946 74.314 ;
               RECT 0.894 75.478 0.946 75.514 ;
               RECT 0.894 76.678 0.946 76.714 ;
               RECT 0.894 77.878 0.946 77.914 ;
               RECT 0.894 79.078 0.946 79.114 ;
               RECT 0.894 80.278 0.946 80.314 ;
               RECT 0.894 81.478 0.946 81.514 ;
               RECT 0.894 82.678 0.946 82.714 ;
               RECT 0.894 83.878 0.946 83.914 ;
               RECT 0.894 85.078 0.946 85.114 ;
               RECT 0.894 86.278 0.946 86.314 ;
               RECT 0.894 87.478 0.946 87.514 ;
               RECT 0.894 88.678 0.946 88.714 ;
               RECT 0.894 89.878 0.946 89.914 ;
               RECT 0.894 91.078 0.946 91.114 ;
               RECT 0.894 92.278 0.946 92.314 ;
               RECT 0.894 93.478 0.946 93.514 ;
               RECT 0.894 94.678 0.946 94.714 ;
               RECT 0.894 95.878 0.946 95.914 ;
               RECT 0.894 97.078 0.946 97.114 ;
               RECT 0.894 98.278 0.946 98.314 ;
               RECT 0.894 99.478 0.946 99.514 ;
               RECT 0.894 100.678 0.946 100.714 ;
               RECT 0.894 101.878 0.946 101.914 ;
               RECT 0.894 103.078 0.946 103.114 ;
               RECT 0.894 104.278 0.946 104.314 ;
               RECT 0.974 0.281 1.026 0.317 ;
               RECT 0.974 104.803 1.026 104.839 ;
               RECT 1.054 0.806 1.106 0.842 ;
               RECT 1.054 2.006 1.106 2.042 ;
               RECT 1.054 3.206 1.106 3.242 ;
               RECT 1.054 4.406 1.106 4.442 ;
               RECT 1.054 5.606 1.106 5.642 ;
               RECT 1.054 6.806 1.106 6.842 ;
               RECT 1.054 8.006 1.106 8.042 ;
               RECT 1.054 9.206 1.106 9.242 ;
               RECT 1.054 10.406 1.106 10.442 ;
               RECT 1.054 11.606 1.106 11.642 ;
               RECT 1.054 12.806 1.106 12.842 ;
               RECT 1.054 14.006 1.106 14.042 ;
               RECT 1.054 15.206 1.106 15.242 ;
               RECT 1.054 16.406 1.106 16.442 ;
               RECT 1.054 17.606 1.106 17.642 ;
               RECT 1.054 18.806 1.106 18.842 ;
               RECT 1.054 20.006 1.106 20.042 ;
               RECT 1.054 21.206 1.106 21.242 ;
               RECT 1.054 22.406 1.106 22.442 ;
               RECT 1.054 23.606 1.106 23.642 ;
               RECT 1.054 24.806 1.106 24.842 ;
               RECT 1.054 26.006 1.106 26.042 ;
               RECT 1.054 27.206 1.106 27.242 ;
               RECT 1.054 28.406 1.106 28.442 ;
               RECT 1.054 29.606 1.106 29.642 ;
               RECT 1.054 30.806 1.106 30.842 ;
               RECT 1.054 32.006 1.106 32.042 ;
               RECT 1.054 33.206 1.106 33.242 ;
               RECT 1.054 34.406 1.106 34.442 ;
               RECT 1.054 35.606 1.106 35.642 ;
               RECT 1.054 36.806 1.106 36.842 ;
               RECT 1.054 38.006 1.106 38.042 ;
               RECT 1.054 39.206 1.106 39.242 ;
               RECT 1.054 40.406 1.106 40.442 ;
               RECT 1.054 41.606 1.106 41.642 ;
               RECT 1.054 42.806 1.106 42.842 ;
               RECT 1.054 44.006 1.106 44.042 ;
               RECT 1.054 45.206 1.106 45.242 ;
               RECT 1.054 46.406 1.106 46.442 ;
               RECT 1.054 47.606 1.106 47.642 ;
               RECT 1.054 49.422 1.106 49.458 ;
               RECT 1.054 49.662 1.106 49.698 ;
               RECT 1.054 51.102 1.106 51.138 ;
               RECT 1.054 51.582 1.106 51.618 ;
               RECT 1.054 53.502 1.106 53.538 ;
               RECT 1.054 53.982 1.106 54.018 ;
               RECT 1.054 55.422 1.106 55.458 ;
               RECT 1.054 55.662 1.106 55.698 ;
               RECT 1.054 56.726 1.106 56.762 ;
               RECT 1.054 57.926 1.106 57.962 ;
               RECT 1.054 59.126 1.106 59.162 ;
               RECT 1.054 60.326 1.106 60.362 ;
               RECT 1.054 61.526 1.106 61.562 ;
               RECT 1.054 62.726 1.106 62.762 ;
               RECT 1.054 63.926 1.106 63.962 ;
               RECT 1.054 65.126 1.106 65.162 ;
               RECT 1.054 66.326 1.106 66.362 ;
               RECT 1.054 67.526 1.106 67.562 ;
               RECT 1.054 68.726 1.106 68.762 ;
               RECT 1.054 69.926 1.106 69.962 ;
               RECT 1.054 71.126 1.106 71.162 ;
               RECT 1.054 72.326 1.106 72.362 ;
               RECT 1.054 73.526 1.106 73.562 ;
               RECT 1.054 74.726 1.106 74.762 ;
               RECT 1.054 75.926 1.106 75.962 ;
               RECT 1.054 77.126 1.106 77.162 ;
               RECT 1.054 78.326 1.106 78.362 ;
               RECT 1.054 79.526 1.106 79.562 ;
               RECT 1.054 80.726 1.106 80.762 ;
               RECT 1.054 81.926 1.106 81.962 ;
               RECT 1.054 83.126 1.106 83.162 ;
               RECT 1.054 84.326 1.106 84.362 ;
               RECT 1.054 85.526 1.106 85.562 ;
               RECT 1.054 86.726 1.106 86.762 ;
               RECT 1.054 87.926 1.106 87.962 ;
               RECT 1.054 89.126 1.106 89.162 ;
               RECT 1.054 90.326 1.106 90.362 ;
               RECT 1.054 91.526 1.106 91.562 ;
               RECT 1.054 92.726 1.106 92.762 ;
               RECT 1.054 93.926 1.106 93.962 ;
               RECT 1.054 95.126 1.106 95.162 ;
               RECT 1.054 96.326 1.106 96.362 ;
               RECT 1.054 97.526 1.106 97.562 ;
               RECT 1.054 98.726 1.106 98.762 ;
               RECT 1.054 99.926 1.106 99.962 ;
               RECT 1.054 101.126 1.106 101.162 ;
               RECT 1.054 102.326 1.106 102.362 ;
               RECT 1.054 103.526 1.106 103.562 ;
               RECT 1.134 1.558 1.186 1.594 ;
               RECT 1.134 2.758 1.186 2.794 ;
               RECT 1.134 3.958 1.186 3.994 ;
               RECT 1.134 5.158 1.186 5.194 ;
               RECT 1.134 6.358 1.186 6.394 ;
               RECT 1.134 7.558 1.186 7.594 ;
               RECT 1.134 8.758 1.186 8.794 ;
               RECT 1.134 9.958 1.186 9.994 ;
               RECT 1.134 11.158 1.186 11.194 ;
               RECT 1.134 12.358 1.186 12.394 ;
               RECT 1.134 13.558 1.186 13.594 ;
               RECT 1.134 14.758 1.186 14.794 ;
               RECT 1.134 15.958 1.186 15.994 ;
               RECT 1.134 17.158 1.186 17.194 ;
               RECT 1.134 18.358 1.186 18.394 ;
               RECT 1.134 19.558 1.186 19.594 ;
               RECT 1.134 20.758 1.186 20.794 ;
               RECT 1.134 21.958 1.186 21.994 ;
               RECT 1.134 23.158 1.186 23.194 ;
               RECT 1.134 24.358 1.186 24.394 ;
               RECT 1.134 25.558 1.186 25.594 ;
               RECT 1.134 26.758 1.186 26.794 ;
               RECT 1.134 27.958 1.186 27.994 ;
               RECT 1.134 29.158 1.186 29.194 ;
               RECT 1.134 30.358 1.186 30.394 ;
               RECT 1.134 31.558 1.186 31.594 ;
               RECT 1.134 32.758 1.186 32.794 ;
               RECT 1.134 33.958 1.186 33.994 ;
               RECT 1.134 35.158 1.186 35.194 ;
               RECT 1.134 36.358 1.186 36.394 ;
               RECT 1.134 37.558 1.186 37.594 ;
               RECT 1.134 38.758 1.186 38.794 ;
               RECT 1.134 39.958 1.186 39.994 ;
               RECT 1.134 41.158 1.186 41.194 ;
               RECT 1.134 42.358 1.186 42.394 ;
               RECT 1.134 43.558 1.186 43.594 ;
               RECT 1.134 44.758 1.186 44.794 ;
               RECT 1.134 45.958 1.186 45.994 ;
               RECT 1.134 47.158 1.186 47.194 ;
               RECT 1.134 48.358 1.186 48.394 ;
               RECT 1.134 50.142 1.186 50.178 ;
               RECT 1.134 50.382 1.186 50.418 ;
               RECT 1.134 54.702 1.186 54.738 ;
               RECT 1.134 54.942 1.186 54.978 ;
               RECT 1.134 57.478 1.186 57.514 ;
               RECT 1.134 58.678 1.186 58.714 ;
               RECT 1.134 59.878 1.186 59.914 ;
               RECT 1.134 61.078 1.186 61.114 ;
               RECT 1.134 62.278 1.186 62.314 ;
               RECT 1.134 63.478 1.186 63.514 ;
               RECT 1.134 64.678 1.186 64.714 ;
               RECT 1.134 65.878 1.186 65.914 ;
               RECT 1.134 67.078 1.186 67.114 ;
               RECT 1.134 68.278 1.186 68.314 ;
               RECT 1.134 69.478 1.186 69.514 ;
               RECT 1.134 70.678 1.186 70.714 ;
               RECT 1.134 71.878 1.186 71.914 ;
               RECT 1.134 73.078 1.186 73.114 ;
               RECT 1.134 74.278 1.186 74.314 ;
               RECT 1.134 75.478 1.186 75.514 ;
               RECT 1.134 76.678 1.186 76.714 ;
               RECT 1.134 77.878 1.186 77.914 ;
               RECT 1.134 79.078 1.186 79.114 ;
               RECT 1.134 80.278 1.186 80.314 ;
               RECT 1.134 81.478 1.186 81.514 ;
               RECT 1.134 82.678 1.186 82.714 ;
               RECT 1.134 83.878 1.186 83.914 ;
               RECT 1.134 85.078 1.186 85.114 ;
               RECT 1.134 86.278 1.186 86.314 ;
               RECT 1.134 87.478 1.186 87.514 ;
               RECT 1.134 88.678 1.186 88.714 ;
               RECT 1.134 89.878 1.186 89.914 ;
               RECT 1.134 91.078 1.186 91.114 ;
               RECT 1.134 92.278 1.186 92.314 ;
               RECT 1.134 93.478 1.186 93.514 ;
               RECT 1.134 94.678 1.186 94.714 ;
               RECT 1.134 95.878 1.186 95.914 ;
               RECT 1.134 97.078 1.186 97.114 ;
               RECT 1.134 98.278 1.186 98.314 ;
               RECT 1.134 99.478 1.186 99.514 ;
               RECT 1.134 100.678 1.186 100.714 ;
               RECT 1.134 101.878 1.186 101.914 ;
               RECT 1.134 103.078 1.186 103.114 ;
               RECT 1.134 104.278 1.186 104.314 ;
               RECT 1.214 0.806 1.266 0.842 ;
               RECT 1.214 2.006 1.266 2.042 ;
               RECT 1.214 3.206 1.266 3.242 ;
               RECT 1.214 4.406 1.266 4.442 ;
               RECT 1.214 5.606 1.266 5.642 ;
               RECT 1.214 6.806 1.266 6.842 ;
               RECT 1.214 8.006 1.266 8.042 ;
               RECT 1.214 9.206 1.266 9.242 ;
               RECT 1.214 10.406 1.266 10.442 ;
               RECT 1.214 11.606 1.266 11.642 ;
               RECT 1.214 12.806 1.266 12.842 ;
               RECT 1.214 14.006 1.266 14.042 ;
               RECT 1.214 15.206 1.266 15.242 ;
               RECT 1.214 16.406 1.266 16.442 ;
               RECT 1.214 17.606 1.266 17.642 ;
               RECT 1.214 18.806 1.266 18.842 ;
               RECT 1.214 20.006 1.266 20.042 ;
               RECT 1.214 21.206 1.266 21.242 ;
               RECT 1.214 22.406 1.266 22.442 ;
               RECT 1.214 23.606 1.266 23.642 ;
               RECT 1.214 24.806 1.266 24.842 ;
               RECT 1.214 26.006 1.266 26.042 ;
               RECT 1.214 27.206 1.266 27.242 ;
               RECT 1.214 28.406 1.266 28.442 ;
               RECT 1.214 29.606 1.266 29.642 ;
               RECT 1.214 30.806 1.266 30.842 ;
               RECT 1.214 32.006 1.266 32.042 ;
               RECT 1.214 33.206 1.266 33.242 ;
               RECT 1.214 34.406 1.266 34.442 ;
               RECT 1.214 35.606 1.266 35.642 ;
               RECT 1.214 36.806 1.266 36.842 ;
               RECT 1.214 38.006 1.266 38.042 ;
               RECT 1.214 39.206 1.266 39.242 ;
               RECT 1.214 40.406 1.266 40.442 ;
               RECT 1.214 41.606 1.266 41.642 ;
               RECT 1.214 42.806 1.266 42.842 ;
               RECT 1.214 44.006 1.266 44.042 ;
               RECT 1.214 45.206 1.266 45.242 ;
               RECT 1.214 46.406 1.266 46.442 ;
               RECT 1.214 47.606 1.266 47.642 ;
               RECT 1.214 49.422 1.266 49.458 ;
               RECT 1.214 49.662 1.266 49.698 ;
               RECT 1.214 55.422 1.266 55.458 ;
               RECT 1.214 55.662 1.266 55.698 ;
               RECT 1.214 56.726 1.266 56.762 ;
               RECT 1.214 57.926 1.266 57.962 ;
               RECT 1.214 59.126 1.266 59.162 ;
               RECT 1.214 60.326 1.266 60.362 ;
               RECT 1.214 61.526 1.266 61.562 ;
               RECT 1.214 62.726 1.266 62.762 ;
               RECT 1.214 63.926 1.266 63.962 ;
               RECT 1.214 65.126 1.266 65.162 ;
               RECT 1.214 66.326 1.266 66.362 ;
               RECT 1.214 67.526 1.266 67.562 ;
               RECT 1.214 68.726 1.266 68.762 ;
               RECT 1.214 69.926 1.266 69.962 ;
               RECT 1.214 71.126 1.266 71.162 ;
               RECT 1.214 72.326 1.266 72.362 ;
               RECT 1.214 73.526 1.266 73.562 ;
               RECT 1.214 74.726 1.266 74.762 ;
               RECT 1.214 75.926 1.266 75.962 ;
               RECT 1.214 77.126 1.266 77.162 ;
               RECT 1.214 78.326 1.266 78.362 ;
               RECT 1.214 79.526 1.266 79.562 ;
               RECT 1.214 80.726 1.266 80.762 ;
               RECT 1.214 81.926 1.266 81.962 ;
               RECT 1.214 83.126 1.266 83.162 ;
               RECT 1.214 84.326 1.266 84.362 ;
               RECT 1.214 85.526 1.266 85.562 ;
               RECT 1.214 86.726 1.266 86.762 ;
               RECT 1.214 87.926 1.266 87.962 ;
               RECT 1.214 89.126 1.266 89.162 ;
               RECT 1.214 90.326 1.266 90.362 ;
               RECT 1.214 91.526 1.266 91.562 ;
               RECT 1.214 92.726 1.266 92.762 ;
               RECT 1.214 93.926 1.266 93.962 ;
               RECT 1.214 95.126 1.266 95.162 ;
               RECT 1.214 96.326 1.266 96.362 ;
               RECT 1.214 97.526 1.266 97.562 ;
               RECT 1.214 98.726 1.266 98.762 ;
               RECT 1.214 99.926 1.266 99.962 ;
               RECT 1.214 101.126 1.266 101.162 ;
               RECT 1.214 102.326 1.266 102.362 ;
               RECT 1.214 103.526 1.266 103.562 ;
               RECT 1.294 1.558 1.346 1.594 ;
               RECT 1.294 2.758 1.346 2.794 ;
               RECT 1.294 3.958 1.346 3.994 ;
               RECT 1.294 5.158 1.346 5.194 ;
               RECT 1.294 6.358 1.346 6.394 ;
               RECT 1.294 7.558 1.346 7.594 ;
               RECT 1.294 8.758 1.346 8.794 ;
               RECT 1.294 9.958 1.346 9.994 ;
               RECT 1.294 11.158 1.346 11.194 ;
               RECT 1.294 12.358 1.346 12.394 ;
               RECT 1.294 13.558 1.346 13.594 ;
               RECT 1.294 14.758 1.346 14.794 ;
               RECT 1.294 15.958 1.346 15.994 ;
               RECT 1.294 17.158 1.346 17.194 ;
               RECT 1.294 18.358 1.346 18.394 ;
               RECT 1.294 19.558 1.346 19.594 ;
               RECT 1.294 20.758 1.346 20.794 ;
               RECT 1.294 21.958 1.346 21.994 ;
               RECT 1.294 23.158 1.346 23.194 ;
               RECT 1.294 24.358 1.346 24.394 ;
               RECT 1.294 25.558 1.346 25.594 ;
               RECT 1.294 26.758 1.346 26.794 ;
               RECT 1.294 27.958 1.346 27.994 ;
               RECT 1.294 29.158 1.346 29.194 ;
               RECT 1.294 30.358 1.346 30.394 ;
               RECT 1.294 31.558 1.346 31.594 ;
               RECT 1.294 32.758 1.346 32.794 ;
               RECT 1.294 33.958 1.346 33.994 ;
               RECT 1.294 35.158 1.346 35.194 ;
               RECT 1.294 36.358 1.346 36.394 ;
               RECT 1.294 37.558 1.346 37.594 ;
               RECT 1.294 38.758 1.346 38.794 ;
               RECT 1.294 39.958 1.346 39.994 ;
               RECT 1.294 41.158 1.346 41.194 ;
               RECT 1.294 42.358 1.346 42.394 ;
               RECT 1.294 43.558 1.346 43.594 ;
               RECT 1.294 44.758 1.346 44.794 ;
               RECT 1.294 45.958 1.346 45.994 ;
               RECT 1.294 47.158 1.346 47.194 ;
               RECT 1.294 48.358 1.346 48.394 ;
               RECT 1.294 50.142 1.346 50.178 ;
               RECT 1.294 50.382 1.346 50.418 ;
               RECT 1.294 54.702 1.346 54.738 ;
               RECT 1.294 54.942 1.346 54.978 ;
               RECT 1.294 57.478 1.346 57.514 ;
               RECT 1.294 58.678 1.346 58.714 ;
               RECT 1.294 59.878 1.346 59.914 ;
               RECT 1.294 61.078 1.346 61.114 ;
               RECT 1.294 62.278 1.346 62.314 ;
               RECT 1.294 63.478 1.346 63.514 ;
               RECT 1.294 64.678 1.346 64.714 ;
               RECT 1.294 65.878 1.346 65.914 ;
               RECT 1.294 67.078 1.346 67.114 ;
               RECT 1.294 68.278 1.346 68.314 ;
               RECT 1.294 69.478 1.346 69.514 ;
               RECT 1.294 70.678 1.346 70.714 ;
               RECT 1.294 71.878 1.346 71.914 ;
               RECT 1.294 73.078 1.346 73.114 ;
               RECT 1.294 74.278 1.346 74.314 ;
               RECT 1.294 75.478 1.346 75.514 ;
               RECT 1.294 76.678 1.346 76.714 ;
               RECT 1.294 77.878 1.346 77.914 ;
               RECT 1.294 79.078 1.346 79.114 ;
               RECT 1.294 80.278 1.346 80.314 ;
               RECT 1.294 81.478 1.346 81.514 ;
               RECT 1.294 82.678 1.346 82.714 ;
               RECT 1.294 83.878 1.346 83.914 ;
               RECT 1.294 85.078 1.346 85.114 ;
               RECT 1.294 86.278 1.346 86.314 ;
               RECT 1.294 87.478 1.346 87.514 ;
               RECT 1.294 88.678 1.346 88.714 ;
               RECT 1.294 89.878 1.346 89.914 ;
               RECT 1.294 91.078 1.346 91.114 ;
               RECT 1.294 92.278 1.346 92.314 ;
               RECT 1.294 93.478 1.346 93.514 ;
               RECT 1.294 94.678 1.346 94.714 ;
               RECT 1.294 95.878 1.346 95.914 ;
               RECT 1.294 97.078 1.346 97.114 ;
               RECT 1.294 98.278 1.346 98.314 ;
               RECT 1.294 99.478 1.346 99.514 ;
               RECT 1.294 100.678 1.346 100.714 ;
               RECT 1.294 101.878 1.346 101.914 ;
               RECT 1.294 103.078 1.346 103.114 ;
               RECT 1.294 104.278 1.346 104.314 ;
               RECT 1.374 0.281 1.426 0.317 ;
               RECT 1.374 104.803 1.426 104.839 ;
               RECT 1.454 0.806 1.506 0.842 ;
               RECT 1.454 2.006 1.506 2.042 ;
               RECT 1.454 3.206 1.506 3.242 ;
               RECT 1.454 4.406 1.506 4.442 ;
               RECT 1.454 5.606 1.506 5.642 ;
               RECT 1.454 6.806 1.506 6.842 ;
               RECT 1.454 8.006 1.506 8.042 ;
               RECT 1.454 9.206 1.506 9.242 ;
               RECT 1.454 10.406 1.506 10.442 ;
               RECT 1.454 11.606 1.506 11.642 ;
               RECT 1.454 12.806 1.506 12.842 ;
               RECT 1.454 14.006 1.506 14.042 ;
               RECT 1.454 15.206 1.506 15.242 ;
               RECT 1.454 16.406 1.506 16.442 ;
               RECT 1.454 17.606 1.506 17.642 ;
               RECT 1.454 18.806 1.506 18.842 ;
               RECT 1.454 20.006 1.506 20.042 ;
               RECT 1.454 21.206 1.506 21.242 ;
               RECT 1.454 22.406 1.506 22.442 ;
               RECT 1.454 23.606 1.506 23.642 ;
               RECT 1.454 24.806 1.506 24.842 ;
               RECT 1.454 26.006 1.506 26.042 ;
               RECT 1.454 27.206 1.506 27.242 ;
               RECT 1.454 28.406 1.506 28.442 ;
               RECT 1.454 29.606 1.506 29.642 ;
               RECT 1.454 30.806 1.506 30.842 ;
               RECT 1.454 32.006 1.506 32.042 ;
               RECT 1.454 33.206 1.506 33.242 ;
               RECT 1.454 34.406 1.506 34.442 ;
               RECT 1.454 35.606 1.506 35.642 ;
               RECT 1.454 36.806 1.506 36.842 ;
               RECT 1.454 38.006 1.506 38.042 ;
               RECT 1.454 39.206 1.506 39.242 ;
               RECT 1.454 40.406 1.506 40.442 ;
               RECT 1.454 41.606 1.506 41.642 ;
               RECT 1.454 42.806 1.506 42.842 ;
               RECT 1.454 44.006 1.506 44.042 ;
               RECT 1.454 45.206 1.506 45.242 ;
               RECT 1.454 46.406 1.506 46.442 ;
               RECT 1.454 47.606 1.506 47.642 ;
               RECT 1.454 49.422 1.506 49.458 ;
               RECT 1.454 49.662 1.506 49.698 ;
               RECT 1.454 55.422 1.506 55.458 ;
               RECT 1.454 55.662 1.506 55.698 ;
               RECT 1.454 56.726 1.506 56.762 ;
               RECT 1.454 57.926 1.506 57.962 ;
               RECT 1.454 59.126 1.506 59.162 ;
               RECT 1.454 60.326 1.506 60.362 ;
               RECT 1.454 61.526 1.506 61.562 ;
               RECT 1.454 62.726 1.506 62.762 ;
               RECT 1.454 63.926 1.506 63.962 ;
               RECT 1.454 65.126 1.506 65.162 ;
               RECT 1.454 66.326 1.506 66.362 ;
               RECT 1.454 67.526 1.506 67.562 ;
               RECT 1.454 68.726 1.506 68.762 ;
               RECT 1.454 69.926 1.506 69.962 ;
               RECT 1.454 71.126 1.506 71.162 ;
               RECT 1.454 72.326 1.506 72.362 ;
               RECT 1.454 73.526 1.506 73.562 ;
               RECT 1.454 74.726 1.506 74.762 ;
               RECT 1.454 75.926 1.506 75.962 ;
               RECT 1.454 77.126 1.506 77.162 ;
               RECT 1.454 78.326 1.506 78.362 ;
               RECT 1.454 79.526 1.506 79.562 ;
               RECT 1.454 80.726 1.506 80.762 ;
               RECT 1.454 81.926 1.506 81.962 ;
               RECT 1.454 83.126 1.506 83.162 ;
               RECT 1.454 84.326 1.506 84.362 ;
               RECT 1.454 85.526 1.506 85.562 ;
               RECT 1.454 86.726 1.506 86.762 ;
               RECT 1.454 87.926 1.506 87.962 ;
               RECT 1.454 89.126 1.506 89.162 ;
               RECT 1.454 90.326 1.506 90.362 ;
               RECT 1.454 91.526 1.506 91.562 ;
               RECT 1.454 92.726 1.506 92.762 ;
               RECT 1.454 93.926 1.506 93.962 ;
               RECT 1.454 95.126 1.506 95.162 ;
               RECT 1.454 96.326 1.506 96.362 ;
               RECT 1.454 97.526 1.506 97.562 ;
               RECT 1.454 98.726 1.506 98.762 ;
               RECT 1.454 99.926 1.506 99.962 ;
               RECT 1.454 101.126 1.506 101.162 ;
               RECT 1.454 102.326 1.506 102.362 ;
               RECT 1.454 103.526 1.506 103.562 ;
               RECT 1.534 1.558 1.586 1.594 ;
               RECT 1.534 2.758 1.586 2.794 ;
               RECT 1.534 3.958 1.586 3.994 ;
               RECT 1.534 5.158 1.586 5.194 ;
               RECT 1.534 6.358 1.586 6.394 ;
               RECT 1.534 7.558 1.586 7.594 ;
               RECT 1.534 8.758 1.586 8.794 ;
               RECT 1.534 9.958 1.586 9.994 ;
               RECT 1.534 11.158 1.586 11.194 ;
               RECT 1.534 12.358 1.586 12.394 ;
               RECT 1.534 13.558 1.586 13.594 ;
               RECT 1.534 14.758 1.586 14.794 ;
               RECT 1.534 15.958 1.586 15.994 ;
               RECT 1.534 17.158 1.586 17.194 ;
               RECT 1.534 18.358 1.586 18.394 ;
               RECT 1.534 19.558 1.586 19.594 ;
               RECT 1.534 20.758 1.586 20.794 ;
               RECT 1.534 21.958 1.586 21.994 ;
               RECT 1.534 23.158 1.586 23.194 ;
               RECT 1.534 24.358 1.586 24.394 ;
               RECT 1.534 25.558 1.586 25.594 ;
               RECT 1.534 26.758 1.586 26.794 ;
               RECT 1.534 27.958 1.586 27.994 ;
               RECT 1.534 29.158 1.586 29.194 ;
               RECT 1.534 30.358 1.586 30.394 ;
               RECT 1.534 31.558 1.586 31.594 ;
               RECT 1.534 32.758 1.586 32.794 ;
               RECT 1.534 33.958 1.586 33.994 ;
               RECT 1.534 35.158 1.586 35.194 ;
               RECT 1.534 36.358 1.586 36.394 ;
               RECT 1.534 37.558 1.586 37.594 ;
               RECT 1.534 38.758 1.586 38.794 ;
               RECT 1.534 39.958 1.586 39.994 ;
               RECT 1.534 41.158 1.586 41.194 ;
               RECT 1.534 42.358 1.586 42.394 ;
               RECT 1.534 43.558 1.586 43.594 ;
               RECT 1.534 44.758 1.586 44.794 ;
               RECT 1.534 45.958 1.586 45.994 ;
               RECT 1.534 47.158 1.586 47.194 ;
               RECT 1.534 48.358 1.586 48.394 ;
               RECT 1.534 50.142 1.586 50.178 ;
               RECT 1.534 50.382 1.586 50.418 ;
               RECT 1.534 54.702 1.586 54.738 ;
               RECT 1.534 54.942 1.586 54.978 ;
               RECT 1.534 57.478 1.586 57.514 ;
               RECT 1.534 58.678 1.586 58.714 ;
               RECT 1.534 59.878 1.586 59.914 ;
               RECT 1.534 61.078 1.586 61.114 ;
               RECT 1.534 62.278 1.586 62.314 ;
               RECT 1.534 63.478 1.586 63.514 ;
               RECT 1.534 64.678 1.586 64.714 ;
               RECT 1.534 65.878 1.586 65.914 ;
               RECT 1.534 67.078 1.586 67.114 ;
               RECT 1.534 68.278 1.586 68.314 ;
               RECT 1.534 69.478 1.586 69.514 ;
               RECT 1.534 70.678 1.586 70.714 ;
               RECT 1.534 71.878 1.586 71.914 ;
               RECT 1.534 73.078 1.586 73.114 ;
               RECT 1.534 74.278 1.586 74.314 ;
               RECT 1.534 75.478 1.586 75.514 ;
               RECT 1.534 76.678 1.586 76.714 ;
               RECT 1.534 77.878 1.586 77.914 ;
               RECT 1.534 79.078 1.586 79.114 ;
               RECT 1.534 80.278 1.586 80.314 ;
               RECT 1.534 81.478 1.586 81.514 ;
               RECT 1.534 82.678 1.586 82.714 ;
               RECT 1.534 83.878 1.586 83.914 ;
               RECT 1.534 85.078 1.586 85.114 ;
               RECT 1.534 86.278 1.586 86.314 ;
               RECT 1.534 87.478 1.586 87.514 ;
               RECT 1.534 88.678 1.586 88.714 ;
               RECT 1.534 89.878 1.586 89.914 ;
               RECT 1.534 91.078 1.586 91.114 ;
               RECT 1.534 92.278 1.586 92.314 ;
               RECT 1.534 93.478 1.586 93.514 ;
               RECT 1.534 94.678 1.586 94.714 ;
               RECT 1.534 95.878 1.586 95.914 ;
               RECT 1.534 97.078 1.586 97.114 ;
               RECT 1.534 98.278 1.586 98.314 ;
               RECT 1.534 99.478 1.586 99.514 ;
               RECT 1.534 100.678 1.586 100.714 ;
               RECT 1.534 101.878 1.586 101.914 ;
               RECT 1.534 103.078 1.586 103.114 ;
               RECT 1.534 104.278 1.586 104.314 ;
               RECT 1.614 0.806 1.666 0.842 ;
               RECT 1.614 2.006 1.666 2.042 ;
               RECT 1.614 3.206 1.666 3.242 ;
               RECT 1.614 4.406 1.666 4.442 ;
               RECT 1.614 5.606 1.666 5.642 ;
               RECT 1.614 6.806 1.666 6.842 ;
               RECT 1.614 8.006 1.666 8.042 ;
               RECT 1.614 9.206 1.666 9.242 ;
               RECT 1.614 10.406 1.666 10.442 ;
               RECT 1.614 11.606 1.666 11.642 ;
               RECT 1.614 12.806 1.666 12.842 ;
               RECT 1.614 14.006 1.666 14.042 ;
               RECT 1.614 15.206 1.666 15.242 ;
               RECT 1.614 16.406 1.666 16.442 ;
               RECT 1.614 17.606 1.666 17.642 ;
               RECT 1.614 18.806 1.666 18.842 ;
               RECT 1.614 20.006 1.666 20.042 ;
               RECT 1.614 21.206 1.666 21.242 ;
               RECT 1.614 22.406 1.666 22.442 ;
               RECT 1.614 23.606 1.666 23.642 ;
               RECT 1.614 24.806 1.666 24.842 ;
               RECT 1.614 26.006 1.666 26.042 ;
               RECT 1.614 27.206 1.666 27.242 ;
               RECT 1.614 28.406 1.666 28.442 ;
               RECT 1.614 29.606 1.666 29.642 ;
               RECT 1.614 30.806 1.666 30.842 ;
               RECT 1.614 32.006 1.666 32.042 ;
               RECT 1.614 33.206 1.666 33.242 ;
               RECT 1.614 34.406 1.666 34.442 ;
               RECT 1.614 35.606 1.666 35.642 ;
               RECT 1.614 36.806 1.666 36.842 ;
               RECT 1.614 38.006 1.666 38.042 ;
               RECT 1.614 39.206 1.666 39.242 ;
               RECT 1.614 40.406 1.666 40.442 ;
               RECT 1.614 41.606 1.666 41.642 ;
               RECT 1.614 42.806 1.666 42.842 ;
               RECT 1.614 44.006 1.666 44.042 ;
               RECT 1.614 45.206 1.666 45.242 ;
               RECT 1.614 46.406 1.666 46.442 ;
               RECT 1.614 47.606 1.666 47.642 ;
               RECT 1.614 49.422 1.666 49.458 ;
               RECT 1.614 49.662 1.666 49.698 ;
               RECT 1.614 55.422 1.666 55.458 ;
               RECT 1.614 55.662 1.666 55.698 ;
               RECT 1.614 56.726 1.666 56.762 ;
               RECT 1.614 57.926 1.666 57.962 ;
               RECT 1.614 59.126 1.666 59.162 ;
               RECT 1.614 60.326 1.666 60.362 ;
               RECT 1.614 61.526 1.666 61.562 ;
               RECT 1.614 62.726 1.666 62.762 ;
               RECT 1.614 63.926 1.666 63.962 ;
               RECT 1.614 65.126 1.666 65.162 ;
               RECT 1.614 66.326 1.666 66.362 ;
               RECT 1.614 67.526 1.666 67.562 ;
               RECT 1.614 68.726 1.666 68.762 ;
               RECT 1.614 69.926 1.666 69.962 ;
               RECT 1.614 71.126 1.666 71.162 ;
               RECT 1.614 72.326 1.666 72.362 ;
               RECT 1.614 73.526 1.666 73.562 ;
               RECT 1.614 74.726 1.666 74.762 ;
               RECT 1.614 75.926 1.666 75.962 ;
               RECT 1.614 77.126 1.666 77.162 ;
               RECT 1.614 78.326 1.666 78.362 ;
               RECT 1.614 79.526 1.666 79.562 ;
               RECT 1.614 80.726 1.666 80.762 ;
               RECT 1.614 81.926 1.666 81.962 ;
               RECT 1.614 83.126 1.666 83.162 ;
               RECT 1.614 84.326 1.666 84.362 ;
               RECT 1.614 85.526 1.666 85.562 ;
               RECT 1.614 86.726 1.666 86.762 ;
               RECT 1.614 87.926 1.666 87.962 ;
               RECT 1.614 89.126 1.666 89.162 ;
               RECT 1.614 90.326 1.666 90.362 ;
               RECT 1.614 91.526 1.666 91.562 ;
               RECT 1.614 92.726 1.666 92.762 ;
               RECT 1.614 93.926 1.666 93.962 ;
               RECT 1.614 95.126 1.666 95.162 ;
               RECT 1.614 96.326 1.666 96.362 ;
               RECT 1.614 97.526 1.666 97.562 ;
               RECT 1.614 98.726 1.666 98.762 ;
               RECT 1.614 99.926 1.666 99.962 ;
               RECT 1.614 101.126 1.666 101.162 ;
               RECT 1.614 102.326 1.666 102.362 ;
               RECT 1.614 103.526 1.666 103.562 ;
               RECT 1.694 1.558 1.746 1.594 ;
               RECT 1.694 2.758 1.746 2.794 ;
               RECT 1.694 3.958 1.746 3.994 ;
               RECT 1.694 5.158 1.746 5.194 ;
               RECT 1.694 6.358 1.746 6.394 ;
               RECT 1.694 7.558 1.746 7.594 ;
               RECT 1.694 8.758 1.746 8.794 ;
               RECT 1.694 9.958 1.746 9.994 ;
               RECT 1.694 11.158 1.746 11.194 ;
               RECT 1.694 12.358 1.746 12.394 ;
               RECT 1.694 13.558 1.746 13.594 ;
               RECT 1.694 14.758 1.746 14.794 ;
               RECT 1.694 15.958 1.746 15.994 ;
               RECT 1.694 17.158 1.746 17.194 ;
               RECT 1.694 18.358 1.746 18.394 ;
               RECT 1.694 19.558 1.746 19.594 ;
               RECT 1.694 20.758 1.746 20.794 ;
               RECT 1.694 21.958 1.746 21.994 ;
               RECT 1.694 23.158 1.746 23.194 ;
               RECT 1.694 24.358 1.746 24.394 ;
               RECT 1.694 25.558 1.746 25.594 ;
               RECT 1.694 26.758 1.746 26.794 ;
               RECT 1.694 27.958 1.746 27.994 ;
               RECT 1.694 29.158 1.746 29.194 ;
               RECT 1.694 30.358 1.746 30.394 ;
               RECT 1.694 31.558 1.746 31.594 ;
               RECT 1.694 32.758 1.746 32.794 ;
               RECT 1.694 33.958 1.746 33.994 ;
               RECT 1.694 35.158 1.746 35.194 ;
               RECT 1.694 36.358 1.746 36.394 ;
               RECT 1.694 37.558 1.746 37.594 ;
               RECT 1.694 38.758 1.746 38.794 ;
               RECT 1.694 39.958 1.746 39.994 ;
               RECT 1.694 41.158 1.746 41.194 ;
               RECT 1.694 42.358 1.746 42.394 ;
               RECT 1.694 43.558 1.746 43.594 ;
               RECT 1.694 44.758 1.746 44.794 ;
               RECT 1.694 45.958 1.746 45.994 ;
               RECT 1.694 47.158 1.746 47.194 ;
               RECT 1.694 48.358 1.746 48.394 ;
               RECT 1.694 50.142 1.746 50.178 ;
               RECT 1.694 50.382 1.746 50.418 ;
               RECT 1.694 54.702 1.746 54.738 ;
               RECT 1.694 54.942 1.746 54.978 ;
               RECT 1.694 57.478 1.746 57.514 ;
               RECT 1.694 58.678 1.746 58.714 ;
               RECT 1.694 59.878 1.746 59.914 ;
               RECT 1.694 61.078 1.746 61.114 ;
               RECT 1.694 62.278 1.746 62.314 ;
               RECT 1.694 63.478 1.746 63.514 ;
               RECT 1.694 64.678 1.746 64.714 ;
               RECT 1.694 65.878 1.746 65.914 ;
               RECT 1.694 67.078 1.746 67.114 ;
               RECT 1.694 68.278 1.746 68.314 ;
               RECT 1.694 69.478 1.746 69.514 ;
               RECT 1.694 70.678 1.746 70.714 ;
               RECT 1.694 71.878 1.746 71.914 ;
               RECT 1.694 73.078 1.746 73.114 ;
               RECT 1.694 74.278 1.746 74.314 ;
               RECT 1.694 75.478 1.746 75.514 ;
               RECT 1.694 76.678 1.746 76.714 ;
               RECT 1.694 77.878 1.746 77.914 ;
               RECT 1.694 79.078 1.746 79.114 ;
               RECT 1.694 80.278 1.746 80.314 ;
               RECT 1.694 81.478 1.746 81.514 ;
               RECT 1.694 82.678 1.746 82.714 ;
               RECT 1.694 83.878 1.746 83.914 ;
               RECT 1.694 85.078 1.746 85.114 ;
               RECT 1.694 86.278 1.746 86.314 ;
               RECT 1.694 87.478 1.746 87.514 ;
               RECT 1.694 88.678 1.746 88.714 ;
               RECT 1.694 89.878 1.746 89.914 ;
               RECT 1.694 91.078 1.746 91.114 ;
               RECT 1.694 92.278 1.746 92.314 ;
               RECT 1.694 93.478 1.746 93.514 ;
               RECT 1.694 94.678 1.746 94.714 ;
               RECT 1.694 95.878 1.746 95.914 ;
               RECT 1.694 97.078 1.746 97.114 ;
               RECT 1.694 98.278 1.746 98.314 ;
               RECT 1.694 99.478 1.746 99.514 ;
               RECT 1.694 100.678 1.746 100.714 ;
               RECT 1.694 101.878 1.746 101.914 ;
               RECT 1.694 103.078 1.746 103.114 ;
               RECT 1.694 104.278 1.746 104.314 ;
               RECT 1.774 0.281 1.826 0.317 ;
               RECT 1.774 104.803 1.826 104.839 ;
               RECT 1.854 0.806 1.906 0.842 ;
               RECT 1.854 2.006 1.906 2.042 ;
               RECT 1.854 3.206 1.906 3.242 ;
               RECT 1.854 4.406 1.906 4.442 ;
               RECT 1.854 5.606 1.906 5.642 ;
               RECT 1.854 6.806 1.906 6.842 ;
               RECT 1.854 8.006 1.906 8.042 ;
               RECT 1.854 9.206 1.906 9.242 ;
               RECT 1.854 10.406 1.906 10.442 ;
               RECT 1.854 11.606 1.906 11.642 ;
               RECT 1.854 12.806 1.906 12.842 ;
               RECT 1.854 14.006 1.906 14.042 ;
               RECT 1.854 15.206 1.906 15.242 ;
               RECT 1.854 16.406 1.906 16.442 ;
               RECT 1.854 17.606 1.906 17.642 ;
               RECT 1.854 18.806 1.906 18.842 ;
               RECT 1.854 20.006 1.906 20.042 ;
               RECT 1.854 21.206 1.906 21.242 ;
               RECT 1.854 22.406 1.906 22.442 ;
               RECT 1.854 23.606 1.906 23.642 ;
               RECT 1.854 24.806 1.906 24.842 ;
               RECT 1.854 26.006 1.906 26.042 ;
               RECT 1.854 27.206 1.906 27.242 ;
               RECT 1.854 28.406 1.906 28.442 ;
               RECT 1.854 29.606 1.906 29.642 ;
               RECT 1.854 30.806 1.906 30.842 ;
               RECT 1.854 32.006 1.906 32.042 ;
               RECT 1.854 33.206 1.906 33.242 ;
               RECT 1.854 34.406 1.906 34.442 ;
               RECT 1.854 35.606 1.906 35.642 ;
               RECT 1.854 36.806 1.906 36.842 ;
               RECT 1.854 38.006 1.906 38.042 ;
               RECT 1.854 39.206 1.906 39.242 ;
               RECT 1.854 40.406 1.906 40.442 ;
               RECT 1.854 41.606 1.906 41.642 ;
               RECT 1.854 42.806 1.906 42.842 ;
               RECT 1.854 44.006 1.906 44.042 ;
               RECT 1.854 45.206 1.906 45.242 ;
               RECT 1.854 46.406 1.906 46.442 ;
               RECT 1.854 47.606 1.906 47.642 ;
               RECT 1.854 49.422 1.906 49.458 ;
               RECT 1.854 49.662 1.906 49.698 ;
               RECT 1.854 51.102 1.906 51.138 ;
               RECT 1.854 51.582 1.906 51.618 ;
               RECT 1.854 53.502 1.906 53.538 ;
               RECT 1.854 53.982 1.906 54.018 ;
               RECT 1.854 55.422 1.906 55.458 ;
               RECT 1.854 55.662 1.906 55.698 ;
               RECT 1.854 56.726 1.906 56.762 ;
               RECT 1.854 57.926 1.906 57.962 ;
               RECT 1.854 59.126 1.906 59.162 ;
               RECT 1.854 60.326 1.906 60.362 ;
               RECT 1.854 61.526 1.906 61.562 ;
               RECT 1.854 62.726 1.906 62.762 ;
               RECT 1.854 63.926 1.906 63.962 ;
               RECT 1.854 65.126 1.906 65.162 ;
               RECT 1.854 66.326 1.906 66.362 ;
               RECT 1.854 67.526 1.906 67.562 ;
               RECT 1.854 68.726 1.906 68.762 ;
               RECT 1.854 69.926 1.906 69.962 ;
               RECT 1.854 71.126 1.906 71.162 ;
               RECT 1.854 72.326 1.906 72.362 ;
               RECT 1.854 73.526 1.906 73.562 ;
               RECT 1.854 74.726 1.906 74.762 ;
               RECT 1.854 75.926 1.906 75.962 ;
               RECT 1.854 77.126 1.906 77.162 ;
               RECT 1.854 78.326 1.906 78.362 ;
               RECT 1.854 79.526 1.906 79.562 ;
               RECT 1.854 80.726 1.906 80.762 ;
               RECT 1.854 81.926 1.906 81.962 ;
               RECT 1.854 83.126 1.906 83.162 ;
               RECT 1.854 84.326 1.906 84.362 ;
               RECT 1.854 85.526 1.906 85.562 ;
               RECT 1.854 86.726 1.906 86.762 ;
               RECT 1.854 87.926 1.906 87.962 ;
               RECT 1.854 89.126 1.906 89.162 ;
               RECT 1.854 90.326 1.906 90.362 ;
               RECT 1.854 91.526 1.906 91.562 ;
               RECT 1.854 92.726 1.906 92.762 ;
               RECT 1.854 93.926 1.906 93.962 ;
               RECT 1.854 95.126 1.906 95.162 ;
               RECT 1.854 96.326 1.906 96.362 ;
               RECT 1.854 97.526 1.906 97.562 ;
               RECT 1.854 98.726 1.906 98.762 ;
               RECT 1.854 99.926 1.906 99.962 ;
               RECT 1.854 101.126 1.906 101.162 ;
               RECT 1.854 102.326 1.906 102.362 ;
               RECT 1.854 103.526 1.906 103.562 ;
               RECT 1.934 1.558 1.986 1.594 ;
               RECT 1.934 2.758 1.986 2.794 ;
               RECT 1.934 3.958 1.986 3.994 ;
               RECT 1.934 5.158 1.986 5.194 ;
               RECT 1.934 6.358 1.986 6.394 ;
               RECT 1.934 7.558 1.986 7.594 ;
               RECT 1.934 8.758 1.986 8.794 ;
               RECT 1.934 9.958 1.986 9.994 ;
               RECT 1.934 11.158 1.986 11.194 ;
               RECT 1.934 12.358 1.986 12.394 ;
               RECT 1.934 13.558 1.986 13.594 ;
               RECT 1.934 14.758 1.986 14.794 ;
               RECT 1.934 15.958 1.986 15.994 ;
               RECT 1.934 17.158 1.986 17.194 ;
               RECT 1.934 18.358 1.986 18.394 ;
               RECT 1.934 19.558 1.986 19.594 ;
               RECT 1.934 20.758 1.986 20.794 ;
               RECT 1.934 21.958 1.986 21.994 ;
               RECT 1.934 23.158 1.986 23.194 ;
               RECT 1.934 24.358 1.986 24.394 ;
               RECT 1.934 25.558 1.986 25.594 ;
               RECT 1.934 26.758 1.986 26.794 ;
               RECT 1.934 27.958 1.986 27.994 ;
               RECT 1.934 29.158 1.986 29.194 ;
               RECT 1.934 30.358 1.986 30.394 ;
               RECT 1.934 31.558 1.986 31.594 ;
               RECT 1.934 32.758 1.986 32.794 ;
               RECT 1.934 33.958 1.986 33.994 ;
               RECT 1.934 35.158 1.986 35.194 ;
               RECT 1.934 36.358 1.986 36.394 ;
               RECT 1.934 37.558 1.986 37.594 ;
               RECT 1.934 38.758 1.986 38.794 ;
               RECT 1.934 39.958 1.986 39.994 ;
               RECT 1.934 41.158 1.986 41.194 ;
               RECT 1.934 42.358 1.986 42.394 ;
               RECT 1.934 43.558 1.986 43.594 ;
               RECT 1.934 44.758 1.986 44.794 ;
               RECT 1.934 45.958 1.986 45.994 ;
               RECT 1.934 47.158 1.986 47.194 ;
               RECT 1.934 48.358 1.986 48.394 ;
               RECT 1.934 50.142 1.986 50.178 ;
               RECT 1.934 50.382 1.986 50.418 ;
               RECT 1.934 54.702 1.986 54.738 ;
               RECT 1.934 54.942 1.986 54.978 ;
               RECT 1.934 57.478 1.986 57.514 ;
               RECT 1.934 58.678 1.986 58.714 ;
               RECT 1.934 59.878 1.986 59.914 ;
               RECT 1.934 61.078 1.986 61.114 ;
               RECT 1.934 62.278 1.986 62.314 ;
               RECT 1.934 63.478 1.986 63.514 ;
               RECT 1.934 64.678 1.986 64.714 ;
               RECT 1.934 65.878 1.986 65.914 ;
               RECT 1.934 67.078 1.986 67.114 ;
               RECT 1.934 68.278 1.986 68.314 ;
               RECT 1.934 69.478 1.986 69.514 ;
               RECT 1.934 70.678 1.986 70.714 ;
               RECT 1.934 71.878 1.986 71.914 ;
               RECT 1.934 73.078 1.986 73.114 ;
               RECT 1.934 74.278 1.986 74.314 ;
               RECT 1.934 75.478 1.986 75.514 ;
               RECT 1.934 76.678 1.986 76.714 ;
               RECT 1.934 77.878 1.986 77.914 ;
               RECT 1.934 79.078 1.986 79.114 ;
               RECT 1.934 80.278 1.986 80.314 ;
               RECT 1.934 81.478 1.986 81.514 ;
               RECT 1.934 82.678 1.986 82.714 ;
               RECT 1.934 83.878 1.986 83.914 ;
               RECT 1.934 85.078 1.986 85.114 ;
               RECT 1.934 86.278 1.986 86.314 ;
               RECT 1.934 87.478 1.986 87.514 ;
               RECT 1.934 88.678 1.986 88.714 ;
               RECT 1.934 89.878 1.986 89.914 ;
               RECT 1.934 91.078 1.986 91.114 ;
               RECT 1.934 92.278 1.986 92.314 ;
               RECT 1.934 93.478 1.986 93.514 ;
               RECT 1.934 94.678 1.986 94.714 ;
               RECT 1.934 95.878 1.986 95.914 ;
               RECT 1.934 97.078 1.986 97.114 ;
               RECT 1.934 98.278 1.986 98.314 ;
               RECT 1.934 99.478 1.986 99.514 ;
               RECT 1.934 100.678 1.986 100.714 ;
               RECT 1.934 101.878 1.986 101.914 ;
               RECT 1.934 103.078 1.986 103.114 ;
               RECT 1.934 104.278 1.986 104.314 ;
               RECT 2.014 0.806 2.066 0.842 ;
               RECT 2.014 2.006 2.066 2.042 ;
               RECT 2.014 3.206 2.066 3.242 ;
               RECT 2.014 4.406 2.066 4.442 ;
               RECT 2.014 5.606 2.066 5.642 ;
               RECT 2.014 6.806 2.066 6.842 ;
               RECT 2.014 8.006 2.066 8.042 ;
               RECT 2.014 9.206 2.066 9.242 ;
               RECT 2.014 10.406 2.066 10.442 ;
               RECT 2.014 11.606 2.066 11.642 ;
               RECT 2.014 12.806 2.066 12.842 ;
               RECT 2.014 14.006 2.066 14.042 ;
               RECT 2.014 15.206 2.066 15.242 ;
               RECT 2.014 16.406 2.066 16.442 ;
               RECT 2.014 17.606 2.066 17.642 ;
               RECT 2.014 18.806 2.066 18.842 ;
               RECT 2.014 20.006 2.066 20.042 ;
               RECT 2.014 21.206 2.066 21.242 ;
               RECT 2.014 22.406 2.066 22.442 ;
               RECT 2.014 23.606 2.066 23.642 ;
               RECT 2.014 24.806 2.066 24.842 ;
               RECT 2.014 26.006 2.066 26.042 ;
               RECT 2.014 27.206 2.066 27.242 ;
               RECT 2.014 28.406 2.066 28.442 ;
               RECT 2.014 29.606 2.066 29.642 ;
               RECT 2.014 30.806 2.066 30.842 ;
               RECT 2.014 32.006 2.066 32.042 ;
               RECT 2.014 33.206 2.066 33.242 ;
               RECT 2.014 34.406 2.066 34.442 ;
               RECT 2.014 35.606 2.066 35.642 ;
               RECT 2.014 36.806 2.066 36.842 ;
               RECT 2.014 38.006 2.066 38.042 ;
               RECT 2.014 39.206 2.066 39.242 ;
               RECT 2.014 40.406 2.066 40.442 ;
               RECT 2.014 41.606 2.066 41.642 ;
               RECT 2.014 42.806 2.066 42.842 ;
               RECT 2.014 44.006 2.066 44.042 ;
               RECT 2.014 45.206 2.066 45.242 ;
               RECT 2.014 46.406 2.066 46.442 ;
               RECT 2.014 47.606 2.066 47.642 ;
               RECT 2.014 49.422 2.066 49.458 ;
               RECT 2.014 49.662 2.066 49.698 ;
               RECT 2.014 55.422 2.066 55.458 ;
               RECT 2.014 55.662 2.066 55.698 ;
               RECT 2.014 56.726 2.066 56.762 ;
               RECT 2.014 57.926 2.066 57.962 ;
               RECT 2.014 59.126 2.066 59.162 ;
               RECT 2.014 60.326 2.066 60.362 ;
               RECT 2.014 61.526 2.066 61.562 ;
               RECT 2.014 62.726 2.066 62.762 ;
               RECT 2.014 63.926 2.066 63.962 ;
               RECT 2.014 65.126 2.066 65.162 ;
               RECT 2.014 66.326 2.066 66.362 ;
               RECT 2.014 67.526 2.066 67.562 ;
               RECT 2.014 68.726 2.066 68.762 ;
               RECT 2.014 69.926 2.066 69.962 ;
               RECT 2.014 71.126 2.066 71.162 ;
               RECT 2.014 72.326 2.066 72.362 ;
               RECT 2.014 73.526 2.066 73.562 ;
               RECT 2.014 74.726 2.066 74.762 ;
               RECT 2.014 75.926 2.066 75.962 ;
               RECT 2.014 77.126 2.066 77.162 ;
               RECT 2.014 78.326 2.066 78.362 ;
               RECT 2.014 79.526 2.066 79.562 ;
               RECT 2.014 80.726 2.066 80.762 ;
               RECT 2.014 81.926 2.066 81.962 ;
               RECT 2.014 83.126 2.066 83.162 ;
               RECT 2.014 84.326 2.066 84.362 ;
               RECT 2.014 85.526 2.066 85.562 ;
               RECT 2.014 86.726 2.066 86.762 ;
               RECT 2.014 87.926 2.066 87.962 ;
               RECT 2.014 89.126 2.066 89.162 ;
               RECT 2.014 90.326 2.066 90.362 ;
               RECT 2.014 91.526 2.066 91.562 ;
               RECT 2.014 92.726 2.066 92.762 ;
               RECT 2.014 93.926 2.066 93.962 ;
               RECT 2.014 95.126 2.066 95.162 ;
               RECT 2.014 96.326 2.066 96.362 ;
               RECT 2.014 97.526 2.066 97.562 ;
               RECT 2.014 98.726 2.066 98.762 ;
               RECT 2.014 99.926 2.066 99.962 ;
               RECT 2.014 101.126 2.066 101.162 ;
               RECT 2.014 102.326 2.066 102.362 ;
               RECT 2.014 103.526 2.066 103.562 ;
               RECT 2.094 1.558 2.146 1.594 ;
               RECT 2.094 2.758 2.146 2.794 ;
               RECT 2.094 3.958 2.146 3.994 ;
               RECT 2.094 5.158 2.146 5.194 ;
               RECT 2.094 6.358 2.146 6.394 ;
               RECT 2.094 7.558 2.146 7.594 ;
               RECT 2.094 8.758 2.146 8.794 ;
               RECT 2.094 9.958 2.146 9.994 ;
               RECT 2.094 11.158 2.146 11.194 ;
               RECT 2.094 12.358 2.146 12.394 ;
               RECT 2.094 13.558 2.146 13.594 ;
               RECT 2.094 14.758 2.146 14.794 ;
               RECT 2.094 15.958 2.146 15.994 ;
               RECT 2.094 17.158 2.146 17.194 ;
               RECT 2.094 18.358 2.146 18.394 ;
               RECT 2.094 19.558 2.146 19.594 ;
               RECT 2.094 20.758 2.146 20.794 ;
               RECT 2.094 21.958 2.146 21.994 ;
               RECT 2.094 23.158 2.146 23.194 ;
               RECT 2.094 24.358 2.146 24.394 ;
               RECT 2.094 25.558 2.146 25.594 ;
               RECT 2.094 26.758 2.146 26.794 ;
               RECT 2.094 27.958 2.146 27.994 ;
               RECT 2.094 29.158 2.146 29.194 ;
               RECT 2.094 30.358 2.146 30.394 ;
               RECT 2.094 31.558 2.146 31.594 ;
               RECT 2.094 32.758 2.146 32.794 ;
               RECT 2.094 33.958 2.146 33.994 ;
               RECT 2.094 35.158 2.146 35.194 ;
               RECT 2.094 36.358 2.146 36.394 ;
               RECT 2.094 37.558 2.146 37.594 ;
               RECT 2.094 38.758 2.146 38.794 ;
               RECT 2.094 39.958 2.146 39.994 ;
               RECT 2.094 41.158 2.146 41.194 ;
               RECT 2.094 42.358 2.146 42.394 ;
               RECT 2.094 43.558 2.146 43.594 ;
               RECT 2.094 44.758 2.146 44.794 ;
               RECT 2.094 45.958 2.146 45.994 ;
               RECT 2.094 47.158 2.146 47.194 ;
               RECT 2.094 48.358 2.146 48.394 ;
               RECT 2.094 50.142 2.146 50.178 ;
               RECT 2.094 50.382 2.146 50.418 ;
               RECT 2.094 54.702 2.146 54.738 ;
               RECT 2.094 54.942 2.146 54.978 ;
               RECT 2.094 57.478 2.146 57.514 ;
               RECT 2.094 58.678 2.146 58.714 ;
               RECT 2.094 59.878 2.146 59.914 ;
               RECT 2.094 61.078 2.146 61.114 ;
               RECT 2.094 62.278 2.146 62.314 ;
               RECT 2.094 63.478 2.146 63.514 ;
               RECT 2.094 64.678 2.146 64.714 ;
               RECT 2.094 65.878 2.146 65.914 ;
               RECT 2.094 67.078 2.146 67.114 ;
               RECT 2.094 68.278 2.146 68.314 ;
               RECT 2.094 69.478 2.146 69.514 ;
               RECT 2.094 70.678 2.146 70.714 ;
               RECT 2.094 71.878 2.146 71.914 ;
               RECT 2.094 73.078 2.146 73.114 ;
               RECT 2.094 74.278 2.146 74.314 ;
               RECT 2.094 75.478 2.146 75.514 ;
               RECT 2.094 76.678 2.146 76.714 ;
               RECT 2.094 77.878 2.146 77.914 ;
               RECT 2.094 79.078 2.146 79.114 ;
               RECT 2.094 80.278 2.146 80.314 ;
               RECT 2.094 81.478 2.146 81.514 ;
               RECT 2.094 82.678 2.146 82.714 ;
               RECT 2.094 83.878 2.146 83.914 ;
               RECT 2.094 85.078 2.146 85.114 ;
               RECT 2.094 86.278 2.146 86.314 ;
               RECT 2.094 87.478 2.146 87.514 ;
               RECT 2.094 88.678 2.146 88.714 ;
               RECT 2.094 89.878 2.146 89.914 ;
               RECT 2.094 91.078 2.146 91.114 ;
               RECT 2.094 92.278 2.146 92.314 ;
               RECT 2.094 93.478 2.146 93.514 ;
               RECT 2.094 94.678 2.146 94.714 ;
               RECT 2.094 95.878 2.146 95.914 ;
               RECT 2.094 97.078 2.146 97.114 ;
               RECT 2.094 98.278 2.146 98.314 ;
               RECT 2.094 99.478 2.146 99.514 ;
               RECT 2.094 100.678 2.146 100.714 ;
               RECT 2.094 101.878 2.146 101.914 ;
               RECT 2.094 103.078 2.146 103.114 ;
               RECT 2.094 104.278 2.146 104.314 ;
               RECT 2.174 0.281 2.226 0.317 ;
               RECT 2.174 104.803 2.226 104.839 ;
               RECT 2.254 0.806 2.306 0.842 ;
               RECT 2.254 2.006 2.306 2.042 ;
               RECT 2.254 3.206 2.306 3.242 ;
               RECT 2.254 4.406 2.306 4.442 ;
               RECT 2.254 5.606 2.306 5.642 ;
               RECT 2.254 6.806 2.306 6.842 ;
               RECT 2.254 8.006 2.306 8.042 ;
               RECT 2.254 9.206 2.306 9.242 ;
               RECT 2.254 10.406 2.306 10.442 ;
               RECT 2.254 11.606 2.306 11.642 ;
               RECT 2.254 12.806 2.306 12.842 ;
               RECT 2.254 14.006 2.306 14.042 ;
               RECT 2.254 15.206 2.306 15.242 ;
               RECT 2.254 16.406 2.306 16.442 ;
               RECT 2.254 17.606 2.306 17.642 ;
               RECT 2.254 18.806 2.306 18.842 ;
               RECT 2.254 20.006 2.306 20.042 ;
               RECT 2.254 21.206 2.306 21.242 ;
               RECT 2.254 22.406 2.306 22.442 ;
               RECT 2.254 23.606 2.306 23.642 ;
               RECT 2.254 24.806 2.306 24.842 ;
               RECT 2.254 26.006 2.306 26.042 ;
               RECT 2.254 27.206 2.306 27.242 ;
               RECT 2.254 28.406 2.306 28.442 ;
               RECT 2.254 29.606 2.306 29.642 ;
               RECT 2.254 30.806 2.306 30.842 ;
               RECT 2.254 32.006 2.306 32.042 ;
               RECT 2.254 33.206 2.306 33.242 ;
               RECT 2.254 34.406 2.306 34.442 ;
               RECT 2.254 35.606 2.306 35.642 ;
               RECT 2.254 36.806 2.306 36.842 ;
               RECT 2.254 38.006 2.306 38.042 ;
               RECT 2.254 39.206 2.306 39.242 ;
               RECT 2.254 40.406 2.306 40.442 ;
               RECT 2.254 41.606 2.306 41.642 ;
               RECT 2.254 42.806 2.306 42.842 ;
               RECT 2.254 44.006 2.306 44.042 ;
               RECT 2.254 45.206 2.306 45.242 ;
               RECT 2.254 46.406 2.306 46.442 ;
               RECT 2.254 47.606 2.306 47.642 ;
               RECT 2.254 49.422 2.306 49.458 ;
               RECT 2.254 49.662 2.306 49.698 ;
               RECT 2.254 55.422 2.306 55.458 ;
               RECT 2.254 55.662 2.306 55.698 ;
               RECT 2.254 56.726 2.306 56.762 ;
               RECT 2.254 57.926 2.306 57.962 ;
               RECT 2.254 59.126 2.306 59.162 ;
               RECT 2.254 60.326 2.306 60.362 ;
               RECT 2.254 61.526 2.306 61.562 ;
               RECT 2.254 62.726 2.306 62.762 ;
               RECT 2.254 63.926 2.306 63.962 ;
               RECT 2.254 65.126 2.306 65.162 ;
               RECT 2.254 66.326 2.306 66.362 ;
               RECT 2.254 67.526 2.306 67.562 ;
               RECT 2.254 68.726 2.306 68.762 ;
               RECT 2.254 69.926 2.306 69.962 ;
               RECT 2.254 71.126 2.306 71.162 ;
               RECT 2.254 72.326 2.306 72.362 ;
               RECT 2.254 73.526 2.306 73.562 ;
               RECT 2.254 74.726 2.306 74.762 ;
               RECT 2.254 75.926 2.306 75.962 ;
               RECT 2.254 77.126 2.306 77.162 ;
               RECT 2.254 78.326 2.306 78.362 ;
               RECT 2.254 79.526 2.306 79.562 ;
               RECT 2.254 80.726 2.306 80.762 ;
               RECT 2.254 81.926 2.306 81.962 ;
               RECT 2.254 83.126 2.306 83.162 ;
               RECT 2.254 84.326 2.306 84.362 ;
               RECT 2.254 85.526 2.306 85.562 ;
               RECT 2.254 86.726 2.306 86.762 ;
               RECT 2.254 87.926 2.306 87.962 ;
               RECT 2.254 89.126 2.306 89.162 ;
               RECT 2.254 90.326 2.306 90.362 ;
               RECT 2.254 91.526 2.306 91.562 ;
               RECT 2.254 92.726 2.306 92.762 ;
               RECT 2.254 93.926 2.306 93.962 ;
               RECT 2.254 95.126 2.306 95.162 ;
               RECT 2.254 96.326 2.306 96.362 ;
               RECT 2.254 97.526 2.306 97.562 ;
               RECT 2.254 98.726 2.306 98.762 ;
               RECT 2.254 99.926 2.306 99.962 ;
               RECT 2.254 101.126 2.306 101.162 ;
               RECT 2.254 102.326 2.306 102.362 ;
               RECT 2.254 103.526 2.306 103.562 ;
               RECT 2.334 1.558 2.386 1.594 ;
               RECT 2.334 2.758 2.386 2.794 ;
               RECT 2.334 3.958 2.386 3.994 ;
               RECT 2.334 5.158 2.386 5.194 ;
               RECT 2.334 6.358 2.386 6.394 ;
               RECT 2.334 7.558 2.386 7.594 ;
               RECT 2.334 8.758 2.386 8.794 ;
               RECT 2.334 9.958 2.386 9.994 ;
               RECT 2.334 11.158 2.386 11.194 ;
               RECT 2.334 12.358 2.386 12.394 ;
               RECT 2.334 13.558 2.386 13.594 ;
               RECT 2.334 14.758 2.386 14.794 ;
               RECT 2.334 15.958 2.386 15.994 ;
               RECT 2.334 17.158 2.386 17.194 ;
               RECT 2.334 18.358 2.386 18.394 ;
               RECT 2.334 19.558 2.386 19.594 ;
               RECT 2.334 20.758 2.386 20.794 ;
               RECT 2.334 21.958 2.386 21.994 ;
               RECT 2.334 23.158 2.386 23.194 ;
               RECT 2.334 24.358 2.386 24.394 ;
               RECT 2.334 25.558 2.386 25.594 ;
               RECT 2.334 26.758 2.386 26.794 ;
               RECT 2.334 27.958 2.386 27.994 ;
               RECT 2.334 29.158 2.386 29.194 ;
               RECT 2.334 30.358 2.386 30.394 ;
               RECT 2.334 31.558 2.386 31.594 ;
               RECT 2.334 32.758 2.386 32.794 ;
               RECT 2.334 33.958 2.386 33.994 ;
               RECT 2.334 35.158 2.386 35.194 ;
               RECT 2.334 36.358 2.386 36.394 ;
               RECT 2.334 37.558 2.386 37.594 ;
               RECT 2.334 38.758 2.386 38.794 ;
               RECT 2.334 39.958 2.386 39.994 ;
               RECT 2.334 41.158 2.386 41.194 ;
               RECT 2.334 42.358 2.386 42.394 ;
               RECT 2.334 43.558 2.386 43.594 ;
               RECT 2.334 44.758 2.386 44.794 ;
               RECT 2.334 45.958 2.386 45.994 ;
               RECT 2.334 47.158 2.386 47.194 ;
               RECT 2.334 48.358 2.386 48.394 ;
               RECT 2.334 50.142 2.386 50.178 ;
               RECT 2.334 50.382 2.386 50.418 ;
               RECT 2.334 54.702 2.386 54.738 ;
               RECT 2.334 54.942 2.386 54.978 ;
               RECT 2.334 57.478 2.386 57.514 ;
               RECT 2.334 58.678 2.386 58.714 ;
               RECT 2.334 59.878 2.386 59.914 ;
               RECT 2.334 61.078 2.386 61.114 ;
               RECT 2.334 62.278 2.386 62.314 ;
               RECT 2.334 63.478 2.386 63.514 ;
               RECT 2.334 64.678 2.386 64.714 ;
               RECT 2.334 65.878 2.386 65.914 ;
               RECT 2.334 67.078 2.386 67.114 ;
               RECT 2.334 68.278 2.386 68.314 ;
               RECT 2.334 69.478 2.386 69.514 ;
               RECT 2.334 70.678 2.386 70.714 ;
               RECT 2.334 71.878 2.386 71.914 ;
               RECT 2.334 73.078 2.386 73.114 ;
               RECT 2.334 74.278 2.386 74.314 ;
               RECT 2.334 75.478 2.386 75.514 ;
               RECT 2.334 76.678 2.386 76.714 ;
               RECT 2.334 77.878 2.386 77.914 ;
               RECT 2.334 79.078 2.386 79.114 ;
               RECT 2.334 80.278 2.386 80.314 ;
               RECT 2.334 81.478 2.386 81.514 ;
               RECT 2.334 82.678 2.386 82.714 ;
               RECT 2.334 83.878 2.386 83.914 ;
               RECT 2.334 85.078 2.386 85.114 ;
               RECT 2.334 86.278 2.386 86.314 ;
               RECT 2.334 87.478 2.386 87.514 ;
               RECT 2.334 88.678 2.386 88.714 ;
               RECT 2.334 89.878 2.386 89.914 ;
               RECT 2.334 91.078 2.386 91.114 ;
               RECT 2.334 92.278 2.386 92.314 ;
               RECT 2.334 93.478 2.386 93.514 ;
               RECT 2.334 94.678 2.386 94.714 ;
               RECT 2.334 95.878 2.386 95.914 ;
               RECT 2.334 97.078 2.386 97.114 ;
               RECT 2.334 98.278 2.386 98.314 ;
               RECT 2.334 99.478 2.386 99.514 ;
               RECT 2.334 100.678 2.386 100.714 ;
               RECT 2.334 101.878 2.386 101.914 ;
               RECT 2.334 103.078 2.386 103.114 ;
               RECT 2.334 104.278 2.386 104.314 ;
               RECT 2.414 0.806 2.466 0.842 ;
               RECT 2.414 2.006 2.466 2.042 ;
               RECT 2.414 3.206 2.466 3.242 ;
               RECT 2.414 4.406 2.466 4.442 ;
               RECT 2.414 5.606 2.466 5.642 ;
               RECT 2.414 6.806 2.466 6.842 ;
               RECT 2.414 8.006 2.466 8.042 ;
               RECT 2.414 9.206 2.466 9.242 ;
               RECT 2.414 10.406 2.466 10.442 ;
               RECT 2.414 11.606 2.466 11.642 ;
               RECT 2.414 12.806 2.466 12.842 ;
               RECT 2.414 14.006 2.466 14.042 ;
               RECT 2.414 15.206 2.466 15.242 ;
               RECT 2.414 16.406 2.466 16.442 ;
               RECT 2.414 17.606 2.466 17.642 ;
               RECT 2.414 18.806 2.466 18.842 ;
               RECT 2.414 20.006 2.466 20.042 ;
               RECT 2.414 21.206 2.466 21.242 ;
               RECT 2.414 22.406 2.466 22.442 ;
               RECT 2.414 23.606 2.466 23.642 ;
               RECT 2.414 24.806 2.466 24.842 ;
               RECT 2.414 26.006 2.466 26.042 ;
               RECT 2.414 27.206 2.466 27.242 ;
               RECT 2.414 28.406 2.466 28.442 ;
               RECT 2.414 29.606 2.466 29.642 ;
               RECT 2.414 30.806 2.466 30.842 ;
               RECT 2.414 32.006 2.466 32.042 ;
               RECT 2.414 33.206 2.466 33.242 ;
               RECT 2.414 34.406 2.466 34.442 ;
               RECT 2.414 35.606 2.466 35.642 ;
               RECT 2.414 36.806 2.466 36.842 ;
               RECT 2.414 38.006 2.466 38.042 ;
               RECT 2.414 39.206 2.466 39.242 ;
               RECT 2.414 40.406 2.466 40.442 ;
               RECT 2.414 41.606 2.466 41.642 ;
               RECT 2.414 42.806 2.466 42.842 ;
               RECT 2.414 44.006 2.466 44.042 ;
               RECT 2.414 45.206 2.466 45.242 ;
               RECT 2.414 46.406 2.466 46.442 ;
               RECT 2.414 47.606 2.466 47.642 ;
               RECT 2.414 49.422 2.466 49.458 ;
               RECT 2.414 49.662 2.466 49.698 ;
               RECT 2.414 55.422 2.466 55.458 ;
               RECT 2.414 55.662 2.466 55.698 ;
               RECT 2.414 56.726 2.466 56.762 ;
               RECT 2.414 57.926 2.466 57.962 ;
               RECT 2.414 59.126 2.466 59.162 ;
               RECT 2.414 60.326 2.466 60.362 ;
               RECT 2.414 61.526 2.466 61.562 ;
               RECT 2.414 62.726 2.466 62.762 ;
               RECT 2.414 63.926 2.466 63.962 ;
               RECT 2.414 65.126 2.466 65.162 ;
               RECT 2.414 66.326 2.466 66.362 ;
               RECT 2.414 67.526 2.466 67.562 ;
               RECT 2.414 68.726 2.466 68.762 ;
               RECT 2.414 69.926 2.466 69.962 ;
               RECT 2.414 71.126 2.466 71.162 ;
               RECT 2.414 72.326 2.466 72.362 ;
               RECT 2.414 73.526 2.466 73.562 ;
               RECT 2.414 74.726 2.466 74.762 ;
               RECT 2.414 75.926 2.466 75.962 ;
               RECT 2.414 77.126 2.466 77.162 ;
               RECT 2.414 78.326 2.466 78.362 ;
               RECT 2.414 79.526 2.466 79.562 ;
               RECT 2.414 80.726 2.466 80.762 ;
               RECT 2.414 81.926 2.466 81.962 ;
               RECT 2.414 83.126 2.466 83.162 ;
               RECT 2.414 84.326 2.466 84.362 ;
               RECT 2.414 85.526 2.466 85.562 ;
               RECT 2.414 86.726 2.466 86.762 ;
               RECT 2.414 87.926 2.466 87.962 ;
               RECT 2.414 89.126 2.466 89.162 ;
               RECT 2.414 90.326 2.466 90.362 ;
               RECT 2.414 91.526 2.466 91.562 ;
               RECT 2.414 92.726 2.466 92.762 ;
               RECT 2.414 93.926 2.466 93.962 ;
               RECT 2.414 95.126 2.466 95.162 ;
               RECT 2.414 96.326 2.466 96.362 ;
               RECT 2.414 97.526 2.466 97.562 ;
               RECT 2.414 98.726 2.466 98.762 ;
               RECT 2.414 99.926 2.466 99.962 ;
               RECT 2.414 101.126 2.466 101.162 ;
               RECT 2.414 102.326 2.466 102.362 ;
               RECT 2.414 103.526 2.466 103.562 ;
               RECT 2.494 1.558 2.546 1.594 ;
               RECT 2.494 2.758 2.546 2.794 ;
               RECT 2.494 3.958 2.546 3.994 ;
               RECT 2.494 5.158 2.546 5.194 ;
               RECT 2.494 6.358 2.546 6.394 ;
               RECT 2.494 7.558 2.546 7.594 ;
               RECT 2.494 8.758 2.546 8.794 ;
               RECT 2.494 9.958 2.546 9.994 ;
               RECT 2.494 11.158 2.546 11.194 ;
               RECT 2.494 12.358 2.546 12.394 ;
               RECT 2.494 13.558 2.546 13.594 ;
               RECT 2.494 14.758 2.546 14.794 ;
               RECT 2.494 15.958 2.546 15.994 ;
               RECT 2.494 17.158 2.546 17.194 ;
               RECT 2.494 18.358 2.546 18.394 ;
               RECT 2.494 19.558 2.546 19.594 ;
               RECT 2.494 20.758 2.546 20.794 ;
               RECT 2.494 21.958 2.546 21.994 ;
               RECT 2.494 23.158 2.546 23.194 ;
               RECT 2.494 24.358 2.546 24.394 ;
               RECT 2.494 25.558 2.546 25.594 ;
               RECT 2.494 26.758 2.546 26.794 ;
               RECT 2.494 27.958 2.546 27.994 ;
               RECT 2.494 29.158 2.546 29.194 ;
               RECT 2.494 30.358 2.546 30.394 ;
               RECT 2.494 31.558 2.546 31.594 ;
               RECT 2.494 32.758 2.546 32.794 ;
               RECT 2.494 33.958 2.546 33.994 ;
               RECT 2.494 35.158 2.546 35.194 ;
               RECT 2.494 36.358 2.546 36.394 ;
               RECT 2.494 37.558 2.546 37.594 ;
               RECT 2.494 38.758 2.546 38.794 ;
               RECT 2.494 39.958 2.546 39.994 ;
               RECT 2.494 41.158 2.546 41.194 ;
               RECT 2.494 42.358 2.546 42.394 ;
               RECT 2.494 43.558 2.546 43.594 ;
               RECT 2.494 44.758 2.546 44.794 ;
               RECT 2.494 45.958 2.546 45.994 ;
               RECT 2.494 47.158 2.546 47.194 ;
               RECT 2.494 48.358 2.546 48.394 ;
               RECT 2.494 50.142 2.546 50.178 ;
               RECT 2.494 50.382 2.546 50.418 ;
               RECT 2.494 54.702 2.546 54.738 ;
               RECT 2.494 54.942 2.546 54.978 ;
               RECT 2.494 57.478 2.546 57.514 ;
               RECT 2.494 58.678 2.546 58.714 ;
               RECT 2.494 59.878 2.546 59.914 ;
               RECT 2.494 61.078 2.546 61.114 ;
               RECT 2.494 62.278 2.546 62.314 ;
               RECT 2.494 63.478 2.546 63.514 ;
               RECT 2.494 64.678 2.546 64.714 ;
               RECT 2.494 65.878 2.546 65.914 ;
               RECT 2.494 67.078 2.546 67.114 ;
               RECT 2.494 68.278 2.546 68.314 ;
               RECT 2.494 69.478 2.546 69.514 ;
               RECT 2.494 70.678 2.546 70.714 ;
               RECT 2.494 71.878 2.546 71.914 ;
               RECT 2.494 73.078 2.546 73.114 ;
               RECT 2.494 74.278 2.546 74.314 ;
               RECT 2.494 75.478 2.546 75.514 ;
               RECT 2.494 76.678 2.546 76.714 ;
               RECT 2.494 77.878 2.546 77.914 ;
               RECT 2.494 79.078 2.546 79.114 ;
               RECT 2.494 80.278 2.546 80.314 ;
               RECT 2.494 81.478 2.546 81.514 ;
               RECT 2.494 82.678 2.546 82.714 ;
               RECT 2.494 83.878 2.546 83.914 ;
               RECT 2.494 85.078 2.546 85.114 ;
               RECT 2.494 86.278 2.546 86.314 ;
               RECT 2.494 87.478 2.546 87.514 ;
               RECT 2.494 88.678 2.546 88.714 ;
               RECT 2.494 89.878 2.546 89.914 ;
               RECT 2.494 91.078 2.546 91.114 ;
               RECT 2.494 92.278 2.546 92.314 ;
               RECT 2.494 93.478 2.546 93.514 ;
               RECT 2.494 94.678 2.546 94.714 ;
               RECT 2.494 95.878 2.546 95.914 ;
               RECT 2.494 97.078 2.546 97.114 ;
               RECT 2.494 98.278 2.546 98.314 ;
               RECT 2.494 99.478 2.546 99.514 ;
               RECT 2.494 100.678 2.546 100.714 ;
               RECT 2.494 101.878 2.546 101.914 ;
               RECT 2.494 103.078 2.546 103.114 ;
               RECT 2.494 104.278 2.546 104.314 ;
               RECT 2.574 0.281 2.626 0.317 ;
               RECT 2.574 104.803 2.626 104.839 ;
               RECT 2.654 0.806 2.706 0.842 ;
               RECT 2.654 2.006 2.706 2.042 ;
               RECT 2.654 3.206 2.706 3.242 ;
               RECT 2.654 4.406 2.706 4.442 ;
               RECT 2.654 5.606 2.706 5.642 ;
               RECT 2.654 6.806 2.706 6.842 ;
               RECT 2.654 8.006 2.706 8.042 ;
               RECT 2.654 9.206 2.706 9.242 ;
               RECT 2.654 10.406 2.706 10.442 ;
               RECT 2.654 11.606 2.706 11.642 ;
               RECT 2.654 12.806 2.706 12.842 ;
               RECT 2.654 14.006 2.706 14.042 ;
               RECT 2.654 15.206 2.706 15.242 ;
               RECT 2.654 16.406 2.706 16.442 ;
               RECT 2.654 17.606 2.706 17.642 ;
               RECT 2.654 18.806 2.706 18.842 ;
               RECT 2.654 20.006 2.706 20.042 ;
               RECT 2.654 21.206 2.706 21.242 ;
               RECT 2.654 22.406 2.706 22.442 ;
               RECT 2.654 23.606 2.706 23.642 ;
               RECT 2.654 24.806 2.706 24.842 ;
               RECT 2.654 26.006 2.706 26.042 ;
               RECT 2.654 27.206 2.706 27.242 ;
               RECT 2.654 28.406 2.706 28.442 ;
               RECT 2.654 29.606 2.706 29.642 ;
               RECT 2.654 30.806 2.706 30.842 ;
               RECT 2.654 32.006 2.706 32.042 ;
               RECT 2.654 33.206 2.706 33.242 ;
               RECT 2.654 34.406 2.706 34.442 ;
               RECT 2.654 35.606 2.706 35.642 ;
               RECT 2.654 36.806 2.706 36.842 ;
               RECT 2.654 38.006 2.706 38.042 ;
               RECT 2.654 39.206 2.706 39.242 ;
               RECT 2.654 40.406 2.706 40.442 ;
               RECT 2.654 41.606 2.706 41.642 ;
               RECT 2.654 42.806 2.706 42.842 ;
               RECT 2.654 44.006 2.706 44.042 ;
               RECT 2.654 45.206 2.706 45.242 ;
               RECT 2.654 46.406 2.706 46.442 ;
               RECT 2.654 47.606 2.706 47.642 ;
               RECT 2.654 49.422 2.706 49.458 ;
               RECT 2.654 49.662 2.706 49.698 ;
               RECT 2.654 51.102 2.706 51.138 ;
               RECT 2.654 51.582 2.706 51.618 ;
               RECT 2.654 53.502 2.706 53.538 ;
               RECT 2.654 53.982 2.706 54.018 ;
               RECT 2.654 55.422 2.706 55.458 ;
               RECT 2.654 55.662 2.706 55.698 ;
               RECT 2.654 56.726 2.706 56.762 ;
               RECT 2.654 57.926 2.706 57.962 ;
               RECT 2.654 59.126 2.706 59.162 ;
               RECT 2.654 60.326 2.706 60.362 ;
               RECT 2.654 61.526 2.706 61.562 ;
               RECT 2.654 62.726 2.706 62.762 ;
               RECT 2.654 63.926 2.706 63.962 ;
               RECT 2.654 65.126 2.706 65.162 ;
               RECT 2.654 66.326 2.706 66.362 ;
               RECT 2.654 67.526 2.706 67.562 ;
               RECT 2.654 68.726 2.706 68.762 ;
               RECT 2.654 69.926 2.706 69.962 ;
               RECT 2.654 71.126 2.706 71.162 ;
               RECT 2.654 72.326 2.706 72.362 ;
               RECT 2.654 73.526 2.706 73.562 ;
               RECT 2.654 74.726 2.706 74.762 ;
               RECT 2.654 75.926 2.706 75.962 ;
               RECT 2.654 77.126 2.706 77.162 ;
               RECT 2.654 78.326 2.706 78.362 ;
               RECT 2.654 79.526 2.706 79.562 ;
               RECT 2.654 80.726 2.706 80.762 ;
               RECT 2.654 81.926 2.706 81.962 ;
               RECT 2.654 83.126 2.706 83.162 ;
               RECT 2.654 84.326 2.706 84.362 ;
               RECT 2.654 85.526 2.706 85.562 ;
               RECT 2.654 86.726 2.706 86.762 ;
               RECT 2.654 87.926 2.706 87.962 ;
               RECT 2.654 89.126 2.706 89.162 ;
               RECT 2.654 90.326 2.706 90.362 ;
               RECT 2.654 91.526 2.706 91.562 ;
               RECT 2.654 92.726 2.706 92.762 ;
               RECT 2.654 93.926 2.706 93.962 ;
               RECT 2.654 95.126 2.706 95.162 ;
               RECT 2.654 96.326 2.706 96.362 ;
               RECT 2.654 97.526 2.706 97.562 ;
               RECT 2.654 98.726 2.706 98.762 ;
               RECT 2.654 99.926 2.706 99.962 ;
               RECT 2.654 101.126 2.706 101.162 ;
               RECT 2.654 102.326 2.706 102.362 ;
               RECT 2.654 103.526 2.706 103.562 ;
               RECT 2.734 1.558 2.786 1.594 ;
               RECT 2.734 2.758 2.786 2.794 ;
               RECT 2.734 3.958 2.786 3.994 ;
               RECT 2.734 5.158 2.786 5.194 ;
               RECT 2.734 6.358 2.786 6.394 ;
               RECT 2.734 7.558 2.786 7.594 ;
               RECT 2.734 8.758 2.786 8.794 ;
               RECT 2.734 9.958 2.786 9.994 ;
               RECT 2.734 11.158 2.786 11.194 ;
               RECT 2.734 12.358 2.786 12.394 ;
               RECT 2.734 13.558 2.786 13.594 ;
               RECT 2.734 14.758 2.786 14.794 ;
               RECT 2.734 15.958 2.786 15.994 ;
               RECT 2.734 17.158 2.786 17.194 ;
               RECT 2.734 18.358 2.786 18.394 ;
               RECT 2.734 19.558 2.786 19.594 ;
               RECT 2.734 20.758 2.786 20.794 ;
               RECT 2.734 21.958 2.786 21.994 ;
               RECT 2.734 23.158 2.786 23.194 ;
               RECT 2.734 24.358 2.786 24.394 ;
               RECT 2.734 25.558 2.786 25.594 ;
               RECT 2.734 26.758 2.786 26.794 ;
               RECT 2.734 27.958 2.786 27.994 ;
               RECT 2.734 29.158 2.786 29.194 ;
               RECT 2.734 30.358 2.786 30.394 ;
               RECT 2.734 31.558 2.786 31.594 ;
               RECT 2.734 32.758 2.786 32.794 ;
               RECT 2.734 33.958 2.786 33.994 ;
               RECT 2.734 35.158 2.786 35.194 ;
               RECT 2.734 36.358 2.786 36.394 ;
               RECT 2.734 37.558 2.786 37.594 ;
               RECT 2.734 38.758 2.786 38.794 ;
               RECT 2.734 39.958 2.786 39.994 ;
               RECT 2.734 41.158 2.786 41.194 ;
               RECT 2.734 42.358 2.786 42.394 ;
               RECT 2.734 43.558 2.786 43.594 ;
               RECT 2.734 44.758 2.786 44.794 ;
               RECT 2.734 45.958 2.786 45.994 ;
               RECT 2.734 47.158 2.786 47.194 ;
               RECT 2.734 48.358 2.786 48.394 ;
               RECT 2.734 50.142 2.786 50.178 ;
               RECT 2.734 50.382 2.786 50.418 ;
               RECT 2.734 54.702 2.786 54.738 ;
               RECT 2.734 54.942 2.786 54.978 ;
               RECT 2.734 57.478 2.786 57.514 ;
               RECT 2.734 58.678 2.786 58.714 ;
               RECT 2.734 59.878 2.786 59.914 ;
               RECT 2.734 61.078 2.786 61.114 ;
               RECT 2.734 62.278 2.786 62.314 ;
               RECT 2.734 63.478 2.786 63.514 ;
               RECT 2.734 64.678 2.786 64.714 ;
               RECT 2.734 65.878 2.786 65.914 ;
               RECT 2.734 67.078 2.786 67.114 ;
               RECT 2.734 68.278 2.786 68.314 ;
               RECT 2.734 69.478 2.786 69.514 ;
               RECT 2.734 70.678 2.786 70.714 ;
               RECT 2.734 71.878 2.786 71.914 ;
               RECT 2.734 73.078 2.786 73.114 ;
               RECT 2.734 74.278 2.786 74.314 ;
               RECT 2.734 75.478 2.786 75.514 ;
               RECT 2.734 76.678 2.786 76.714 ;
               RECT 2.734 77.878 2.786 77.914 ;
               RECT 2.734 79.078 2.786 79.114 ;
               RECT 2.734 80.278 2.786 80.314 ;
               RECT 2.734 81.478 2.786 81.514 ;
               RECT 2.734 82.678 2.786 82.714 ;
               RECT 2.734 83.878 2.786 83.914 ;
               RECT 2.734 85.078 2.786 85.114 ;
               RECT 2.734 86.278 2.786 86.314 ;
               RECT 2.734 87.478 2.786 87.514 ;
               RECT 2.734 88.678 2.786 88.714 ;
               RECT 2.734 89.878 2.786 89.914 ;
               RECT 2.734 91.078 2.786 91.114 ;
               RECT 2.734 92.278 2.786 92.314 ;
               RECT 2.734 93.478 2.786 93.514 ;
               RECT 2.734 94.678 2.786 94.714 ;
               RECT 2.734 95.878 2.786 95.914 ;
               RECT 2.734 97.078 2.786 97.114 ;
               RECT 2.734 98.278 2.786 98.314 ;
               RECT 2.734 99.478 2.786 99.514 ;
               RECT 2.734 100.678 2.786 100.714 ;
               RECT 2.734 101.878 2.786 101.914 ;
               RECT 2.734 103.078 2.786 103.114 ;
               RECT 2.734 104.278 2.786 104.314 ;
               RECT 2.814 0.806 2.866 0.842 ;
               RECT 2.814 2.006 2.866 2.042 ;
               RECT 2.814 3.206 2.866 3.242 ;
               RECT 2.814 4.406 2.866 4.442 ;
               RECT 2.814 5.606 2.866 5.642 ;
               RECT 2.814 6.806 2.866 6.842 ;
               RECT 2.814 8.006 2.866 8.042 ;
               RECT 2.814 9.206 2.866 9.242 ;
               RECT 2.814 10.406 2.866 10.442 ;
               RECT 2.814 11.606 2.866 11.642 ;
               RECT 2.814 12.806 2.866 12.842 ;
               RECT 2.814 14.006 2.866 14.042 ;
               RECT 2.814 15.206 2.866 15.242 ;
               RECT 2.814 16.406 2.866 16.442 ;
               RECT 2.814 17.606 2.866 17.642 ;
               RECT 2.814 18.806 2.866 18.842 ;
               RECT 2.814 20.006 2.866 20.042 ;
               RECT 2.814 21.206 2.866 21.242 ;
               RECT 2.814 22.406 2.866 22.442 ;
               RECT 2.814 23.606 2.866 23.642 ;
               RECT 2.814 24.806 2.866 24.842 ;
               RECT 2.814 26.006 2.866 26.042 ;
               RECT 2.814 27.206 2.866 27.242 ;
               RECT 2.814 28.406 2.866 28.442 ;
               RECT 2.814 29.606 2.866 29.642 ;
               RECT 2.814 30.806 2.866 30.842 ;
               RECT 2.814 32.006 2.866 32.042 ;
               RECT 2.814 33.206 2.866 33.242 ;
               RECT 2.814 34.406 2.866 34.442 ;
               RECT 2.814 35.606 2.866 35.642 ;
               RECT 2.814 36.806 2.866 36.842 ;
               RECT 2.814 38.006 2.866 38.042 ;
               RECT 2.814 39.206 2.866 39.242 ;
               RECT 2.814 40.406 2.866 40.442 ;
               RECT 2.814 41.606 2.866 41.642 ;
               RECT 2.814 42.806 2.866 42.842 ;
               RECT 2.814 44.006 2.866 44.042 ;
               RECT 2.814 45.206 2.866 45.242 ;
               RECT 2.814 46.406 2.866 46.442 ;
               RECT 2.814 47.606 2.866 47.642 ;
               RECT 2.814 49.422 2.866 49.458 ;
               RECT 2.814 49.662 2.866 49.698 ;
               RECT 2.814 55.422 2.866 55.458 ;
               RECT 2.814 55.662 2.866 55.698 ;
               RECT 2.814 56.726 2.866 56.762 ;
               RECT 2.814 57.926 2.866 57.962 ;
               RECT 2.814 59.126 2.866 59.162 ;
               RECT 2.814 60.326 2.866 60.362 ;
               RECT 2.814 61.526 2.866 61.562 ;
               RECT 2.814 62.726 2.866 62.762 ;
               RECT 2.814 63.926 2.866 63.962 ;
               RECT 2.814 65.126 2.866 65.162 ;
               RECT 2.814 66.326 2.866 66.362 ;
               RECT 2.814 67.526 2.866 67.562 ;
               RECT 2.814 68.726 2.866 68.762 ;
               RECT 2.814 69.926 2.866 69.962 ;
               RECT 2.814 71.126 2.866 71.162 ;
               RECT 2.814 72.326 2.866 72.362 ;
               RECT 2.814 73.526 2.866 73.562 ;
               RECT 2.814 74.726 2.866 74.762 ;
               RECT 2.814 75.926 2.866 75.962 ;
               RECT 2.814 77.126 2.866 77.162 ;
               RECT 2.814 78.326 2.866 78.362 ;
               RECT 2.814 79.526 2.866 79.562 ;
               RECT 2.814 80.726 2.866 80.762 ;
               RECT 2.814 81.926 2.866 81.962 ;
               RECT 2.814 83.126 2.866 83.162 ;
               RECT 2.814 84.326 2.866 84.362 ;
               RECT 2.814 85.526 2.866 85.562 ;
               RECT 2.814 86.726 2.866 86.762 ;
               RECT 2.814 87.926 2.866 87.962 ;
               RECT 2.814 89.126 2.866 89.162 ;
               RECT 2.814 90.326 2.866 90.362 ;
               RECT 2.814 91.526 2.866 91.562 ;
               RECT 2.814 92.726 2.866 92.762 ;
               RECT 2.814 93.926 2.866 93.962 ;
               RECT 2.814 95.126 2.866 95.162 ;
               RECT 2.814 96.326 2.866 96.362 ;
               RECT 2.814 97.526 2.866 97.562 ;
               RECT 2.814 98.726 2.866 98.762 ;
               RECT 2.814 99.926 2.866 99.962 ;
               RECT 2.814 101.126 2.866 101.162 ;
               RECT 2.814 102.326 2.866 102.362 ;
               RECT 2.814 103.526 2.866 103.562 ;
               RECT 2.894 1.558 2.946 1.594 ;
               RECT 2.894 2.758 2.946 2.794 ;
               RECT 2.894 3.958 2.946 3.994 ;
               RECT 2.894 5.158 2.946 5.194 ;
               RECT 2.894 6.358 2.946 6.394 ;
               RECT 2.894 7.558 2.946 7.594 ;
               RECT 2.894 8.758 2.946 8.794 ;
               RECT 2.894 9.958 2.946 9.994 ;
               RECT 2.894 11.158 2.946 11.194 ;
               RECT 2.894 12.358 2.946 12.394 ;
               RECT 2.894 13.558 2.946 13.594 ;
               RECT 2.894 14.758 2.946 14.794 ;
               RECT 2.894 15.958 2.946 15.994 ;
               RECT 2.894 17.158 2.946 17.194 ;
               RECT 2.894 18.358 2.946 18.394 ;
               RECT 2.894 19.558 2.946 19.594 ;
               RECT 2.894 20.758 2.946 20.794 ;
               RECT 2.894 21.958 2.946 21.994 ;
               RECT 2.894 23.158 2.946 23.194 ;
               RECT 2.894 24.358 2.946 24.394 ;
               RECT 2.894 25.558 2.946 25.594 ;
               RECT 2.894 26.758 2.946 26.794 ;
               RECT 2.894 27.958 2.946 27.994 ;
               RECT 2.894 29.158 2.946 29.194 ;
               RECT 2.894 30.358 2.946 30.394 ;
               RECT 2.894 31.558 2.946 31.594 ;
               RECT 2.894 32.758 2.946 32.794 ;
               RECT 2.894 33.958 2.946 33.994 ;
               RECT 2.894 35.158 2.946 35.194 ;
               RECT 2.894 36.358 2.946 36.394 ;
               RECT 2.894 37.558 2.946 37.594 ;
               RECT 2.894 38.758 2.946 38.794 ;
               RECT 2.894 39.958 2.946 39.994 ;
               RECT 2.894 41.158 2.946 41.194 ;
               RECT 2.894 42.358 2.946 42.394 ;
               RECT 2.894 43.558 2.946 43.594 ;
               RECT 2.894 44.758 2.946 44.794 ;
               RECT 2.894 45.958 2.946 45.994 ;
               RECT 2.894 47.158 2.946 47.194 ;
               RECT 2.894 48.358 2.946 48.394 ;
               RECT 2.894 50.142 2.946 50.178 ;
               RECT 2.894 50.382 2.946 50.418 ;
               RECT 2.894 54.702 2.946 54.738 ;
               RECT 2.894 54.942 2.946 54.978 ;
               RECT 2.894 57.478 2.946 57.514 ;
               RECT 2.894 58.678 2.946 58.714 ;
               RECT 2.894 59.878 2.946 59.914 ;
               RECT 2.894 61.078 2.946 61.114 ;
               RECT 2.894 62.278 2.946 62.314 ;
               RECT 2.894 63.478 2.946 63.514 ;
               RECT 2.894 64.678 2.946 64.714 ;
               RECT 2.894 65.878 2.946 65.914 ;
               RECT 2.894 67.078 2.946 67.114 ;
               RECT 2.894 68.278 2.946 68.314 ;
               RECT 2.894 69.478 2.946 69.514 ;
               RECT 2.894 70.678 2.946 70.714 ;
               RECT 2.894 71.878 2.946 71.914 ;
               RECT 2.894 73.078 2.946 73.114 ;
               RECT 2.894 74.278 2.946 74.314 ;
               RECT 2.894 75.478 2.946 75.514 ;
               RECT 2.894 76.678 2.946 76.714 ;
               RECT 2.894 77.878 2.946 77.914 ;
               RECT 2.894 79.078 2.946 79.114 ;
               RECT 2.894 80.278 2.946 80.314 ;
               RECT 2.894 81.478 2.946 81.514 ;
               RECT 2.894 82.678 2.946 82.714 ;
               RECT 2.894 83.878 2.946 83.914 ;
               RECT 2.894 85.078 2.946 85.114 ;
               RECT 2.894 86.278 2.946 86.314 ;
               RECT 2.894 87.478 2.946 87.514 ;
               RECT 2.894 88.678 2.946 88.714 ;
               RECT 2.894 89.878 2.946 89.914 ;
               RECT 2.894 91.078 2.946 91.114 ;
               RECT 2.894 92.278 2.946 92.314 ;
               RECT 2.894 93.478 2.946 93.514 ;
               RECT 2.894 94.678 2.946 94.714 ;
               RECT 2.894 95.878 2.946 95.914 ;
               RECT 2.894 97.078 2.946 97.114 ;
               RECT 2.894 98.278 2.946 98.314 ;
               RECT 2.894 99.478 2.946 99.514 ;
               RECT 2.894 100.678 2.946 100.714 ;
               RECT 2.894 101.878 2.946 101.914 ;
               RECT 2.894 103.078 2.946 103.114 ;
               RECT 2.894 104.278 2.946 104.314 ;
               RECT 2.974 0.281 3.026 0.317 ;
               RECT 2.974 104.803 3.026 104.839 ;
               RECT 3.054 0.806 3.106 0.842 ;
               RECT 3.054 2.006 3.106 2.042 ;
               RECT 3.054 3.206 3.106 3.242 ;
               RECT 3.054 4.406 3.106 4.442 ;
               RECT 3.054 5.606 3.106 5.642 ;
               RECT 3.054 6.806 3.106 6.842 ;
               RECT 3.054 8.006 3.106 8.042 ;
               RECT 3.054 9.206 3.106 9.242 ;
               RECT 3.054 10.406 3.106 10.442 ;
               RECT 3.054 11.606 3.106 11.642 ;
               RECT 3.054 12.806 3.106 12.842 ;
               RECT 3.054 14.006 3.106 14.042 ;
               RECT 3.054 15.206 3.106 15.242 ;
               RECT 3.054 16.406 3.106 16.442 ;
               RECT 3.054 17.606 3.106 17.642 ;
               RECT 3.054 18.806 3.106 18.842 ;
               RECT 3.054 20.006 3.106 20.042 ;
               RECT 3.054 21.206 3.106 21.242 ;
               RECT 3.054 22.406 3.106 22.442 ;
               RECT 3.054 23.606 3.106 23.642 ;
               RECT 3.054 24.806 3.106 24.842 ;
               RECT 3.054 26.006 3.106 26.042 ;
               RECT 3.054 27.206 3.106 27.242 ;
               RECT 3.054 28.406 3.106 28.442 ;
               RECT 3.054 29.606 3.106 29.642 ;
               RECT 3.054 30.806 3.106 30.842 ;
               RECT 3.054 32.006 3.106 32.042 ;
               RECT 3.054 33.206 3.106 33.242 ;
               RECT 3.054 34.406 3.106 34.442 ;
               RECT 3.054 35.606 3.106 35.642 ;
               RECT 3.054 36.806 3.106 36.842 ;
               RECT 3.054 38.006 3.106 38.042 ;
               RECT 3.054 39.206 3.106 39.242 ;
               RECT 3.054 40.406 3.106 40.442 ;
               RECT 3.054 41.606 3.106 41.642 ;
               RECT 3.054 42.806 3.106 42.842 ;
               RECT 3.054 44.006 3.106 44.042 ;
               RECT 3.054 45.206 3.106 45.242 ;
               RECT 3.054 46.406 3.106 46.442 ;
               RECT 3.054 47.606 3.106 47.642 ;
               RECT 3.054 49.422 3.106 49.458 ;
               RECT 3.054 49.662 3.106 49.698 ;
               RECT 3.054 55.422 3.106 55.458 ;
               RECT 3.054 55.662 3.106 55.698 ;
               RECT 3.054 56.726 3.106 56.762 ;
               RECT 3.054 57.926 3.106 57.962 ;
               RECT 3.054 59.126 3.106 59.162 ;
               RECT 3.054 60.326 3.106 60.362 ;
               RECT 3.054 61.526 3.106 61.562 ;
               RECT 3.054 62.726 3.106 62.762 ;
               RECT 3.054 63.926 3.106 63.962 ;
               RECT 3.054 65.126 3.106 65.162 ;
               RECT 3.054 66.326 3.106 66.362 ;
               RECT 3.054 67.526 3.106 67.562 ;
               RECT 3.054 68.726 3.106 68.762 ;
               RECT 3.054 69.926 3.106 69.962 ;
               RECT 3.054 71.126 3.106 71.162 ;
               RECT 3.054 72.326 3.106 72.362 ;
               RECT 3.054 73.526 3.106 73.562 ;
               RECT 3.054 74.726 3.106 74.762 ;
               RECT 3.054 75.926 3.106 75.962 ;
               RECT 3.054 77.126 3.106 77.162 ;
               RECT 3.054 78.326 3.106 78.362 ;
               RECT 3.054 79.526 3.106 79.562 ;
               RECT 3.054 80.726 3.106 80.762 ;
               RECT 3.054 81.926 3.106 81.962 ;
               RECT 3.054 83.126 3.106 83.162 ;
               RECT 3.054 84.326 3.106 84.362 ;
               RECT 3.054 85.526 3.106 85.562 ;
               RECT 3.054 86.726 3.106 86.762 ;
               RECT 3.054 87.926 3.106 87.962 ;
               RECT 3.054 89.126 3.106 89.162 ;
               RECT 3.054 90.326 3.106 90.362 ;
               RECT 3.054 91.526 3.106 91.562 ;
               RECT 3.054 92.726 3.106 92.762 ;
               RECT 3.054 93.926 3.106 93.962 ;
               RECT 3.054 95.126 3.106 95.162 ;
               RECT 3.054 96.326 3.106 96.362 ;
               RECT 3.054 97.526 3.106 97.562 ;
               RECT 3.054 98.726 3.106 98.762 ;
               RECT 3.054 99.926 3.106 99.962 ;
               RECT 3.054 101.126 3.106 101.162 ;
               RECT 3.054 102.326 3.106 102.362 ;
               RECT 3.054 103.526 3.106 103.562 ;
               RECT 3.134 1.558 3.186 1.594 ;
               RECT 3.134 2.758 3.186 2.794 ;
               RECT 3.134 3.958 3.186 3.994 ;
               RECT 3.134 5.158 3.186 5.194 ;
               RECT 3.134 6.358 3.186 6.394 ;
               RECT 3.134 7.558 3.186 7.594 ;
               RECT 3.134 8.758 3.186 8.794 ;
               RECT 3.134 9.958 3.186 9.994 ;
               RECT 3.134 11.158 3.186 11.194 ;
               RECT 3.134 12.358 3.186 12.394 ;
               RECT 3.134 13.558 3.186 13.594 ;
               RECT 3.134 14.758 3.186 14.794 ;
               RECT 3.134 15.958 3.186 15.994 ;
               RECT 3.134 17.158 3.186 17.194 ;
               RECT 3.134 18.358 3.186 18.394 ;
               RECT 3.134 19.558 3.186 19.594 ;
               RECT 3.134 20.758 3.186 20.794 ;
               RECT 3.134 21.958 3.186 21.994 ;
               RECT 3.134 23.158 3.186 23.194 ;
               RECT 3.134 24.358 3.186 24.394 ;
               RECT 3.134 25.558 3.186 25.594 ;
               RECT 3.134 26.758 3.186 26.794 ;
               RECT 3.134 27.958 3.186 27.994 ;
               RECT 3.134 29.158 3.186 29.194 ;
               RECT 3.134 30.358 3.186 30.394 ;
               RECT 3.134 31.558 3.186 31.594 ;
               RECT 3.134 32.758 3.186 32.794 ;
               RECT 3.134 33.958 3.186 33.994 ;
               RECT 3.134 35.158 3.186 35.194 ;
               RECT 3.134 36.358 3.186 36.394 ;
               RECT 3.134 37.558 3.186 37.594 ;
               RECT 3.134 38.758 3.186 38.794 ;
               RECT 3.134 39.958 3.186 39.994 ;
               RECT 3.134 41.158 3.186 41.194 ;
               RECT 3.134 42.358 3.186 42.394 ;
               RECT 3.134 43.558 3.186 43.594 ;
               RECT 3.134 44.758 3.186 44.794 ;
               RECT 3.134 45.958 3.186 45.994 ;
               RECT 3.134 47.158 3.186 47.194 ;
               RECT 3.134 48.358 3.186 48.394 ;
               RECT 3.134 50.142 3.186 50.178 ;
               RECT 3.134 50.382 3.186 50.418 ;
               RECT 3.134 54.702 3.186 54.738 ;
               RECT 3.134 54.942 3.186 54.978 ;
               RECT 3.134 57.478 3.186 57.514 ;
               RECT 3.134 58.678 3.186 58.714 ;
               RECT 3.134 59.878 3.186 59.914 ;
               RECT 3.134 61.078 3.186 61.114 ;
               RECT 3.134 62.278 3.186 62.314 ;
               RECT 3.134 63.478 3.186 63.514 ;
               RECT 3.134 64.678 3.186 64.714 ;
               RECT 3.134 65.878 3.186 65.914 ;
               RECT 3.134 67.078 3.186 67.114 ;
               RECT 3.134 68.278 3.186 68.314 ;
               RECT 3.134 69.478 3.186 69.514 ;
               RECT 3.134 70.678 3.186 70.714 ;
               RECT 3.134 71.878 3.186 71.914 ;
               RECT 3.134 73.078 3.186 73.114 ;
               RECT 3.134 74.278 3.186 74.314 ;
               RECT 3.134 75.478 3.186 75.514 ;
               RECT 3.134 76.678 3.186 76.714 ;
               RECT 3.134 77.878 3.186 77.914 ;
               RECT 3.134 79.078 3.186 79.114 ;
               RECT 3.134 80.278 3.186 80.314 ;
               RECT 3.134 81.478 3.186 81.514 ;
               RECT 3.134 82.678 3.186 82.714 ;
               RECT 3.134 83.878 3.186 83.914 ;
               RECT 3.134 85.078 3.186 85.114 ;
               RECT 3.134 86.278 3.186 86.314 ;
               RECT 3.134 87.478 3.186 87.514 ;
               RECT 3.134 88.678 3.186 88.714 ;
               RECT 3.134 89.878 3.186 89.914 ;
               RECT 3.134 91.078 3.186 91.114 ;
               RECT 3.134 92.278 3.186 92.314 ;
               RECT 3.134 93.478 3.186 93.514 ;
               RECT 3.134 94.678 3.186 94.714 ;
               RECT 3.134 95.878 3.186 95.914 ;
               RECT 3.134 97.078 3.186 97.114 ;
               RECT 3.134 98.278 3.186 98.314 ;
               RECT 3.134 99.478 3.186 99.514 ;
               RECT 3.134 100.678 3.186 100.714 ;
               RECT 3.134 101.878 3.186 101.914 ;
               RECT 3.134 103.078 3.186 103.114 ;
               RECT 3.134 104.278 3.186 104.314 ;
               RECT 3.214 0.806 3.266 0.842 ;
               RECT 3.214 2.006 3.266 2.042 ;
               RECT 3.214 3.206 3.266 3.242 ;
               RECT 3.214 4.406 3.266 4.442 ;
               RECT 3.214 5.606 3.266 5.642 ;
               RECT 3.214 6.806 3.266 6.842 ;
               RECT 3.214 8.006 3.266 8.042 ;
               RECT 3.214 9.206 3.266 9.242 ;
               RECT 3.214 10.406 3.266 10.442 ;
               RECT 3.214 11.606 3.266 11.642 ;
               RECT 3.214 12.806 3.266 12.842 ;
               RECT 3.214 14.006 3.266 14.042 ;
               RECT 3.214 15.206 3.266 15.242 ;
               RECT 3.214 16.406 3.266 16.442 ;
               RECT 3.214 17.606 3.266 17.642 ;
               RECT 3.214 18.806 3.266 18.842 ;
               RECT 3.214 20.006 3.266 20.042 ;
               RECT 3.214 21.206 3.266 21.242 ;
               RECT 3.214 22.406 3.266 22.442 ;
               RECT 3.214 23.606 3.266 23.642 ;
               RECT 3.214 24.806 3.266 24.842 ;
               RECT 3.214 26.006 3.266 26.042 ;
               RECT 3.214 27.206 3.266 27.242 ;
               RECT 3.214 28.406 3.266 28.442 ;
               RECT 3.214 29.606 3.266 29.642 ;
               RECT 3.214 30.806 3.266 30.842 ;
               RECT 3.214 32.006 3.266 32.042 ;
               RECT 3.214 33.206 3.266 33.242 ;
               RECT 3.214 34.406 3.266 34.442 ;
               RECT 3.214 35.606 3.266 35.642 ;
               RECT 3.214 36.806 3.266 36.842 ;
               RECT 3.214 38.006 3.266 38.042 ;
               RECT 3.214 39.206 3.266 39.242 ;
               RECT 3.214 40.406 3.266 40.442 ;
               RECT 3.214 41.606 3.266 41.642 ;
               RECT 3.214 42.806 3.266 42.842 ;
               RECT 3.214 44.006 3.266 44.042 ;
               RECT 3.214 45.206 3.266 45.242 ;
               RECT 3.214 46.406 3.266 46.442 ;
               RECT 3.214 47.606 3.266 47.642 ;
               RECT 3.214 49.422 3.266 49.458 ;
               RECT 3.214 49.662 3.266 49.698 ;
               RECT 3.214 55.422 3.266 55.458 ;
               RECT 3.214 55.662 3.266 55.698 ;
               RECT 3.214 56.726 3.266 56.762 ;
               RECT 3.214 57.926 3.266 57.962 ;
               RECT 3.214 59.126 3.266 59.162 ;
               RECT 3.214 60.326 3.266 60.362 ;
               RECT 3.214 61.526 3.266 61.562 ;
               RECT 3.214 62.726 3.266 62.762 ;
               RECT 3.214 63.926 3.266 63.962 ;
               RECT 3.214 65.126 3.266 65.162 ;
               RECT 3.214 66.326 3.266 66.362 ;
               RECT 3.214 67.526 3.266 67.562 ;
               RECT 3.214 68.726 3.266 68.762 ;
               RECT 3.214 69.926 3.266 69.962 ;
               RECT 3.214 71.126 3.266 71.162 ;
               RECT 3.214 72.326 3.266 72.362 ;
               RECT 3.214 73.526 3.266 73.562 ;
               RECT 3.214 74.726 3.266 74.762 ;
               RECT 3.214 75.926 3.266 75.962 ;
               RECT 3.214 77.126 3.266 77.162 ;
               RECT 3.214 78.326 3.266 78.362 ;
               RECT 3.214 79.526 3.266 79.562 ;
               RECT 3.214 80.726 3.266 80.762 ;
               RECT 3.214 81.926 3.266 81.962 ;
               RECT 3.214 83.126 3.266 83.162 ;
               RECT 3.214 84.326 3.266 84.362 ;
               RECT 3.214 85.526 3.266 85.562 ;
               RECT 3.214 86.726 3.266 86.762 ;
               RECT 3.214 87.926 3.266 87.962 ;
               RECT 3.214 89.126 3.266 89.162 ;
               RECT 3.214 90.326 3.266 90.362 ;
               RECT 3.214 91.526 3.266 91.562 ;
               RECT 3.214 92.726 3.266 92.762 ;
               RECT 3.214 93.926 3.266 93.962 ;
               RECT 3.214 95.126 3.266 95.162 ;
               RECT 3.214 96.326 3.266 96.362 ;
               RECT 3.214 97.526 3.266 97.562 ;
               RECT 3.214 98.726 3.266 98.762 ;
               RECT 3.214 99.926 3.266 99.962 ;
               RECT 3.214 101.126 3.266 101.162 ;
               RECT 3.214 102.326 3.266 102.362 ;
               RECT 3.214 103.526 3.266 103.562 ;
               RECT 3.294 1.558 3.346 1.594 ;
               RECT 3.294 2.758 3.346 2.794 ;
               RECT 3.294 3.958 3.346 3.994 ;
               RECT 3.294 5.158 3.346 5.194 ;
               RECT 3.294 6.358 3.346 6.394 ;
               RECT 3.294 7.558 3.346 7.594 ;
               RECT 3.294 8.758 3.346 8.794 ;
               RECT 3.294 9.958 3.346 9.994 ;
               RECT 3.294 11.158 3.346 11.194 ;
               RECT 3.294 12.358 3.346 12.394 ;
               RECT 3.294 13.558 3.346 13.594 ;
               RECT 3.294 14.758 3.346 14.794 ;
               RECT 3.294 15.958 3.346 15.994 ;
               RECT 3.294 17.158 3.346 17.194 ;
               RECT 3.294 18.358 3.346 18.394 ;
               RECT 3.294 19.558 3.346 19.594 ;
               RECT 3.294 20.758 3.346 20.794 ;
               RECT 3.294 21.958 3.346 21.994 ;
               RECT 3.294 23.158 3.346 23.194 ;
               RECT 3.294 24.358 3.346 24.394 ;
               RECT 3.294 25.558 3.346 25.594 ;
               RECT 3.294 26.758 3.346 26.794 ;
               RECT 3.294 27.958 3.346 27.994 ;
               RECT 3.294 29.158 3.346 29.194 ;
               RECT 3.294 30.358 3.346 30.394 ;
               RECT 3.294 31.558 3.346 31.594 ;
               RECT 3.294 32.758 3.346 32.794 ;
               RECT 3.294 33.958 3.346 33.994 ;
               RECT 3.294 35.158 3.346 35.194 ;
               RECT 3.294 36.358 3.346 36.394 ;
               RECT 3.294 37.558 3.346 37.594 ;
               RECT 3.294 38.758 3.346 38.794 ;
               RECT 3.294 39.958 3.346 39.994 ;
               RECT 3.294 41.158 3.346 41.194 ;
               RECT 3.294 42.358 3.346 42.394 ;
               RECT 3.294 43.558 3.346 43.594 ;
               RECT 3.294 44.758 3.346 44.794 ;
               RECT 3.294 45.958 3.346 45.994 ;
               RECT 3.294 47.158 3.346 47.194 ;
               RECT 3.294 48.358 3.346 48.394 ;
               RECT 3.294 50.142 3.346 50.178 ;
               RECT 3.294 50.382 3.346 50.418 ;
               RECT 3.294 54.702 3.346 54.738 ;
               RECT 3.294 54.942 3.346 54.978 ;
               RECT 3.294 57.478 3.346 57.514 ;
               RECT 3.294 58.678 3.346 58.714 ;
               RECT 3.294 59.878 3.346 59.914 ;
               RECT 3.294 61.078 3.346 61.114 ;
               RECT 3.294 62.278 3.346 62.314 ;
               RECT 3.294 63.478 3.346 63.514 ;
               RECT 3.294 64.678 3.346 64.714 ;
               RECT 3.294 65.878 3.346 65.914 ;
               RECT 3.294 67.078 3.346 67.114 ;
               RECT 3.294 68.278 3.346 68.314 ;
               RECT 3.294 69.478 3.346 69.514 ;
               RECT 3.294 70.678 3.346 70.714 ;
               RECT 3.294 71.878 3.346 71.914 ;
               RECT 3.294 73.078 3.346 73.114 ;
               RECT 3.294 74.278 3.346 74.314 ;
               RECT 3.294 75.478 3.346 75.514 ;
               RECT 3.294 76.678 3.346 76.714 ;
               RECT 3.294 77.878 3.346 77.914 ;
               RECT 3.294 79.078 3.346 79.114 ;
               RECT 3.294 80.278 3.346 80.314 ;
               RECT 3.294 81.478 3.346 81.514 ;
               RECT 3.294 82.678 3.346 82.714 ;
               RECT 3.294 83.878 3.346 83.914 ;
               RECT 3.294 85.078 3.346 85.114 ;
               RECT 3.294 86.278 3.346 86.314 ;
               RECT 3.294 87.478 3.346 87.514 ;
               RECT 3.294 88.678 3.346 88.714 ;
               RECT 3.294 89.878 3.346 89.914 ;
               RECT 3.294 91.078 3.346 91.114 ;
               RECT 3.294 92.278 3.346 92.314 ;
               RECT 3.294 93.478 3.346 93.514 ;
               RECT 3.294 94.678 3.346 94.714 ;
               RECT 3.294 95.878 3.346 95.914 ;
               RECT 3.294 97.078 3.346 97.114 ;
               RECT 3.294 98.278 3.346 98.314 ;
               RECT 3.294 99.478 3.346 99.514 ;
               RECT 3.294 100.678 3.346 100.714 ;
               RECT 3.294 101.878 3.346 101.914 ;
               RECT 3.294 103.078 3.346 103.114 ;
               RECT 3.294 104.278 3.346 104.314 ;
               RECT 3.374 0.281 3.426 0.317 ;
               RECT 3.374 104.803 3.426 104.839 ;
               RECT 3.454 0.806 3.506 0.842 ;
               RECT 3.454 2.006 3.506 2.042 ;
               RECT 3.454 3.206 3.506 3.242 ;
               RECT 3.454 4.406 3.506 4.442 ;
               RECT 3.454 5.606 3.506 5.642 ;
               RECT 3.454 6.806 3.506 6.842 ;
               RECT 3.454 8.006 3.506 8.042 ;
               RECT 3.454 9.206 3.506 9.242 ;
               RECT 3.454 10.406 3.506 10.442 ;
               RECT 3.454 11.606 3.506 11.642 ;
               RECT 3.454 12.806 3.506 12.842 ;
               RECT 3.454 14.006 3.506 14.042 ;
               RECT 3.454 15.206 3.506 15.242 ;
               RECT 3.454 16.406 3.506 16.442 ;
               RECT 3.454 17.606 3.506 17.642 ;
               RECT 3.454 18.806 3.506 18.842 ;
               RECT 3.454 20.006 3.506 20.042 ;
               RECT 3.454 21.206 3.506 21.242 ;
               RECT 3.454 22.406 3.506 22.442 ;
               RECT 3.454 23.606 3.506 23.642 ;
               RECT 3.454 24.806 3.506 24.842 ;
               RECT 3.454 26.006 3.506 26.042 ;
               RECT 3.454 27.206 3.506 27.242 ;
               RECT 3.454 28.406 3.506 28.442 ;
               RECT 3.454 29.606 3.506 29.642 ;
               RECT 3.454 30.806 3.506 30.842 ;
               RECT 3.454 32.006 3.506 32.042 ;
               RECT 3.454 33.206 3.506 33.242 ;
               RECT 3.454 34.406 3.506 34.442 ;
               RECT 3.454 35.606 3.506 35.642 ;
               RECT 3.454 36.806 3.506 36.842 ;
               RECT 3.454 38.006 3.506 38.042 ;
               RECT 3.454 39.206 3.506 39.242 ;
               RECT 3.454 40.406 3.506 40.442 ;
               RECT 3.454 41.606 3.506 41.642 ;
               RECT 3.454 42.806 3.506 42.842 ;
               RECT 3.454 44.006 3.506 44.042 ;
               RECT 3.454 45.206 3.506 45.242 ;
               RECT 3.454 46.406 3.506 46.442 ;
               RECT 3.454 47.606 3.506 47.642 ;
               RECT 3.454 49.422 3.506 49.458 ;
               RECT 3.454 49.662 3.506 49.698 ;
               RECT 3.454 51.102 3.506 51.138 ;
               RECT 3.454 51.582 3.506 51.618 ;
               RECT 3.454 53.502 3.506 53.538 ;
               RECT 3.454 53.982 3.506 54.018 ;
               RECT 3.454 55.422 3.506 55.458 ;
               RECT 3.454 55.662 3.506 55.698 ;
               RECT 3.454 56.726 3.506 56.762 ;
               RECT 3.454 57.926 3.506 57.962 ;
               RECT 3.454 59.126 3.506 59.162 ;
               RECT 3.454 60.326 3.506 60.362 ;
               RECT 3.454 61.526 3.506 61.562 ;
               RECT 3.454 62.726 3.506 62.762 ;
               RECT 3.454 63.926 3.506 63.962 ;
               RECT 3.454 65.126 3.506 65.162 ;
               RECT 3.454 66.326 3.506 66.362 ;
               RECT 3.454 67.526 3.506 67.562 ;
               RECT 3.454 68.726 3.506 68.762 ;
               RECT 3.454 69.926 3.506 69.962 ;
               RECT 3.454 71.126 3.506 71.162 ;
               RECT 3.454 72.326 3.506 72.362 ;
               RECT 3.454 73.526 3.506 73.562 ;
               RECT 3.454 74.726 3.506 74.762 ;
               RECT 3.454 75.926 3.506 75.962 ;
               RECT 3.454 77.126 3.506 77.162 ;
               RECT 3.454 78.326 3.506 78.362 ;
               RECT 3.454 79.526 3.506 79.562 ;
               RECT 3.454 80.726 3.506 80.762 ;
               RECT 3.454 81.926 3.506 81.962 ;
               RECT 3.454 83.126 3.506 83.162 ;
               RECT 3.454 84.326 3.506 84.362 ;
               RECT 3.454 85.526 3.506 85.562 ;
               RECT 3.454 86.726 3.506 86.762 ;
               RECT 3.454 87.926 3.506 87.962 ;
               RECT 3.454 89.126 3.506 89.162 ;
               RECT 3.454 90.326 3.506 90.362 ;
               RECT 3.454 91.526 3.506 91.562 ;
               RECT 3.454 92.726 3.506 92.762 ;
               RECT 3.454 93.926 3.506 93.962 ;
               RECT 3.454 95.126 3.506 95.162 ;
               RECT 3.454 96.326 3.506 96.362 ;
               RECT 3.454 97.526 3.506 97.562 ;
               RECT 3.454 98.726 3.506 98.762 ;
               RECT 3.454 99.926 3.506 99.962 ;
               RECT 3.454 101.126 3.506 101.162 ;
               RECT 3.454 102.326 3.506 102.362 ;
               RECT 3.454 103.526 3.506 103.562 ;
               RECT 3.534 1.558 3.586 1.594 ;
               RECT 3.534 2.758 3.586 2.794 ;
               RECT 3.534 3.958 3.586 3.994 ;
               RECT 3.534 5.158 3.586 5.194 ;
               RECT 3.534 6.358 3.586 6.394 ;
               RECT 3.534 7.558 3.586 7.594 ;
               RECT 3.534 8.758 3.586 8.794 ;
               RECT 3.534 9.958 3.586 9.994 ;
               RECT 3.534 11.158 3.586 11.194 ;
               RECT 3.534 12.358 3.586 12.394 ;
               RECT 3.534 13.558 3.586 13.594 ;
               RECT 3.534 14.758 3.586 14.794 ;
               RECT 3.534 15.958 3.586 15.994 ;
               RECT 3.534 17.158 3.586 17.194 ;
               RECT 3.534 18.358 3.586 18.394 ;
               RECT 3.534 19.558 3.586 19.594 ;
               RECT 3.534 20.758 3.586 20.794 ;
               RECT 3.534 21.958 3.586 21.994 ;
               RECT 3.534 23.158 3.586 23.194 ;
               RECT 3.534 24.358 3.586 24.394 ;
               RECT 3.534 25.558 3.586 25.594 ;
               RECT 3.534 26.758 3.586 26.794 ;
               RECT 3.534 27.958 3.586 27.994 ;
               RECT 3.534 29.158 3.586 29.194 ;
               RECT 3.534 30.358 3.586 30.394 ;
               RECT 3.534 31.558 3.586 31.594 ;
               RECT 3.534 32.758 3.586 32.794 ;
               RECT 3.534 33.958 3.586 33.994 ;
               RECT 3.534 35.158 3.586 35.194 ;
               RECT 3.534 36.358 3.586 36.394 ;
               RECT 3.534 37.558 3.586 37.594 ;
               RECT 3.534 38.758 3.586 38.794 ;
               RECT 3.534 39.958 3.586 39.994 ;
               RECT 3.534 41.158 3.586 41.194 ;
               RECT 3.534 42.358 3.586 42.394 ;
               RECT 3.534 43.558 3.586 43.594 ;
               RECT 3.534 44.758 3.586 44.794 ;
               RECT 3.534 45.958 3.586 45.994 ;
               RECT 3.534 47.158 3.586 47.194 ;
               RECT 3.534 48.358 3.586 48.394 ;
               RECT 3.534 50.142 3.586 50.178 ;
               RECT 3.534 50.382 3.586 50.418 ;
               RECT 3.534 54.702 3.586 54.738 ;
               RECT 3.534 54.942 3.586 54.978 ;
               RECT 3.534 57.478 3.586 57.514 ;
               RECT 3.534 58.678 3.586 58.714 ;
               RECT 3.534 59.878 3.586 59.914 ;
               RECT 3.534 61.078 3.586 61.114 ;
               RECT 3.534 62.278 3.586 62.314 ;
               RECT 3.534 63.478 3.586 63.514 ;
               RECT 3.534 64.678 3.586 64.714 ;
               RECT 3.534 65.878 3.586 65.914 ;
               RECT 3.534 67.078 3.586 67.114 ;
               RECT 3.534 68.278 3.586 68.314 ;
               RECT 3.534 69.478 3.586 69.514 ;
               RECT 3.534 70.678 3.586 70.714 ;
               RECT 3.534 71.878 3.586 71.914 ;
               RECT 3.534 73.078 3.586 73.114 ;
               RECT 3.534 74.278 3.586 74.314 ;
               RECT 3.534 75.478 3.586 75.514 ;
               RECT 3.534 76.678 3.586 76.714 ;
               RECT 3.534 77.878 3.586 77.914 ;
               RECT 3.534 79.078 3.586 79.114 ;
               RECT 3.534 80.278 3.586 80.314 ;
               RECT 3.534 81.478 3.586 81.514 ;
               RECT 3.534 82.678 3.586 82.714 ;
               RECT 3.534 83.878 3.586 83.914 ;
               RECT 3.534 85.078 3.586 85.114 ;
               RECT 3.534 86.278 3.586 86.314 ;
               RECT 3.534 87.478 3.586 87.514 ;
               RECT 3.534 88.678 3.586 88.714 ;
               RECT 3.534 89.878 3.586 89.914 ;
               RECT 3.534 91.078 3.586 91.114 ;
               RECT 3.534 92.278 3.586 92.314 ;
               RECT 3.534 93.478 3.586 93.514 ;
               RECT 3.534 94.678 3.586 94.714 ;
               RECT 3.534 95.878 3.586 95.914 ;
               RECT 3.534 97.078 3.586 97.114 ;
               RECT 3.534 98.278 3.586 98.314 ;
               RECT 3.534 99.478 3.586 99.514 ;
               RECT 3.534 100.678 3.586 100.714 ;
               RECT 3.534 101.878 3.586 101.914 ;
               RECT 3.534 103.078 3.586 103.114 ;
               RECT 3.534 104.278 3.586 104.314 ;
               RECT 3.614 0.806 3.666 0.842 ;
               RECT 3.614 2.006 3.666 2.042 ;
               RECT 3.614 3.206 3.666 3.242 ;
               RECT 3.614 4.406 3.666 4.442 ;
               RECT 3.614 5.606 3.666 5.642 ;
               RECT 3.614 6.806 3.666 6.842 ;
               RECT 3.614 8.006 3.666 8.042 ;
               RECT 3.614 9.206 3.666 9.242 ;
               RECT 3.614 10.406 3.666 10.442 ;
               RECT 3.614 11.606 3.666 11.642 ;
               RECT 3.614 12.806 3.666 12.842 ;
               RECT 3.614 14.006 3.666 14.042 ;
               RECT 3.614 15.206 3.666 15.242 ;
               RECT 3.614 16.406 3.666 16.442 ;
               RECT 3.614 17.606 3.666 17.642 ;
               RECT 3.614 18.806 3.666 18.842 ;
               RECT 3.614 20.006 3.666 20.042 ;
               RECT 3.614 21.206 3.666 21.242 ;
               RECT 3.614 22.406 3.666 22.442 ;
               RECT 3.614 23.606 3.666 23.642 ;
               RECT 3.614 24.806 3.666 24.842 ;
               RECT 3.614 26.006 3.666 26.042 ;
               RECT 3.614 27.206 3.666 27.242 ;
               RECT 3.614 28.406 3.666 28.442 ;
               RECT 3.614 29.606 3.666 29.642 ;
               RECT 3.614 30.806 3.666 30.842 ;
               RECT 3.614 32.006 3.666 32.042 ;
               RECT 3.614 33.206 3.666 33.242 ;
               RECT 3.614 34.406 3.666 34.442 ;
               RECT 3.614 35.606 3.666 35.642 ;
               RECT 3.614 36.806 3.666 36.842 ;
               RECT 3.614 38.006 3.666 38.042 ;
               RECT 3.614 39.206 3.666 39.242 ;
               RECT 3.614 40.406 3.666 40.442 ;
               RECT 3.614 41.606 3.666 41.642 ;
               RECT 3.614 42.806 3.666 42.842 ;
               RECT 3.614 44.006 3.666 44.042 ;
               RECT 3.614 45.206 3.666 45.242 ;
               RECT 3.614 46.406 3.666 46.442 ;
               RECT 3.614 47.606 3.666 47.642 ;
               RECT 3.614 49.422 3.666 49.458 ;
               RECT 3.614 49.662 3.666 49.698 ;
               RECT 3.614 55.422 3.666 55.458 ;
               RECT 3.614 55.662 3.666 55.698 ;
               RECT 3.614 56.726 3.666 56.762 ;
               RECT 3.614 57.926 3.666 57.962 ;
               RECT 3.614 59.126 3.666 59.162 ;
               RECT 3.614 60.326 3.666 60.362 ;
               RECT 3.614 61.526 3.666 61.562 ;
               RECT 3.614 62.726 3.666 62.762 ;
               RECT 3.614 63.926 3.666 63.962 ;
               RECT 3.614 65.126 3.666 65.162 ;
               RECT 3.614 66.326 3.666 66.362 ;
               RECT 3.614 67.526 3.666 67.562 ;
               RECT 3.614 68.726 3.666 68.762 ;
               RECT 3.614 69.926 3.666 69.962 ;
               RECT 3.614 71.126 3.666 71.162 ;
               RECT 3.614 72.326 3.666 72.362 ;
               RECT 3.614 73.526 3.666 73.562 ;
               RECT 3.614 74.726 3.666 74.762 ;
               RECT 3.614 75.926 3.666 75.962 ;
               RECT 3.614 77.126 3.666 77.162 ;
               RECT 3.614 78.326 3.666 78.362 ;
               RECT 3.614 79.526 3.666 79.562 ;
               RECT 3.614 80.726 3.666 80.762 ;
               RECT 3.614 81.926 3.666 81.962 ;
               RECT 3.614 83.126 3.666 83.162 ;
               RECT 3.614 84.326 3.666 84.362 ;
               RECT 3.614 85.526 3.666 85.562 ;
               RECT 3.614 86.726 3.666 86.762 ;
               RECT 3.614 87.926 3.666 87.962 ;
               RECT 3.614 89.126 3.666 89.162 ;
               RECT 3.614 90.326 3.666 90.362 ;
               RECT 3.614 91.526 3.666 91.562 ;
               RECT 3.614 92.726 3.666 92.762 ;
               RECT 3.614 93.926 3.666 93.962 ;
               RECT 3.614 95.126 3.666 95.162 ;
               RECT 3.614 96.326 3.666 96.362 ;
               RECT 3.614 97.526 3.666 97.562 ;
               RECT 3.614 98.726 3.666 98.762 ;
               RECT 3.614 99.926 3.666 99.962 ;
               RECT 3.614 101.126 3.666 101.162 ;
               RECT 3.614 102.326 3.666 102.362 ;
               RECT 3.614 103.526 3.666 103.562 ;
               RECT 3.694 1.558 3.746 1.594 ;
               RECT 3.694 2.758 3.746 2.794 ;
               RECT 3.694 3.958 3.746 3.994 ;
               RECT 3.694 5.158 3.746 5.194 ;
               RECT 3.694 6.358 3.746 6.394 ;
               RECT 3.694 7.558 3.746 7.594 ;
               RECT 3.694 8.758 3.746 8.794 ;
               RECT 3.694 9.958 3.746 9.994 ;
               RECT 3.694 11.158 3.746 11.194 ;
               RECT 3.694 12.358 3.746 12.394 ;
               RECT 3.694 13.558 3.746 13.594 ;
               RECT 3.694 14.758 3.746 14.794 ;
               RECT 3.694 15.958 3.746 15.994 ;
               RECT 3.694 17.158 3.746 17.194 ;
               RECT 3.694 18.358 3.746 18.394 ;
               RECT 3.694 19.558 3.746 19.594 ;
               RECT 3.694 20.758 3.746 20.794 ;
               RECT 3.694 21.958 3.746 21.994 ;
               RECT 3.694 23.158 3.746 23.194 ;
               RECT 3.694 24.358 3.746 24.394 ;
               RECT 3.694 25.558 3.746 25.594 ;
               RECT 3.694 26.758 3.746 26.794 ;
               RECT 3.694 27.958 3.746 27.994 ;
               RECT 3.694 29.158 3.746 29.194 ;
               RECT 3.694 30.358 3.746 30.394 ;
               RECT 3.694 31.558 3.746 31.594 ;
               RECT 3.694 32.758 3.746 32.794 ;
               RECT 3.694 33.958 3.746 33.994 ;
               RECT 3.694 35.158 3.746 35.194 ;
               RECT 3.694 36.358 3.746 36.394 ;
               RECT 3.694 37.558 3.746 37.594 ;
               RECT 3.694 38.758 3.746 38.794 ;
               RECT 3.694 39.958 3.746 39.994 ;
               RECT 3.694 41.158 3.746 41.194 ;
               RECT 3.694 42.358 3.746 42.394 ;
               RECT 3.694 43.558 3.746 43.594 ;
               RECT 3.694 44.758 3.746 44.794 ;
               RECT 3.694 45.958 3.746 45.994 ;
               RECT 3.694 47.158 3.746 47.194 ;
               RECT 3.694 48.358 3.746 48.394 ;
               RECT 3.694 50.142 3.746 50.178 ;
               RECT 3.694 50.382 3.746 50.418 ;
               RECT 3.694 54.702 3.746 54.738 ;
               RECT 3.694 54.942 3.746 54.978 ;
               RECT 3.694 57.478 3.746 57.514 ;
               RECT 3.694 58.678 3.746 58.714 ;
               RECT 3.694 59.878 3.746 59.914 ;
               RECT 3.694 61.078 3.746 61.114 ;
               RECT 3.694 62.278 3.746 62.314 ;
               RECT 3.694 63.478 3.746 63.514 ;
               RECT 3.694 64.678 3.746 64.714 ;
               RECT 3.694 65.878 3.746 65.914 ;
               RECT 3.694 67.078 3.746 67.114 ;
               RECT 3.694 68.278 3.746 68.314 ;
               RECT 3.694 69.478 3.746 69.514 ;
               RECT 3.694 70.678 3.746 70.714 ;
               RECT 3.694 71.878 3.746 71.914 ;
               RECT 3.694 73.078 3.746 73.114 ;
               RECT 3.694 74.278 3.746 74.314 ;
               RECT 3.694 75.478 3.746 75.514 ;
               RECT 3.694 76.678 3.746 76.714 ;
               RECT 3.694 77.878 3.746 77.914 ;
               RECT 3.694 79.078 3.746 79.114 ;
               RECT 3.694 80.278 3.746 80.314 ;
               RECT 3.694 81.478 3.746 81.514 ;
               RECT 3.694 82.678 3.746 82.714 ;
               RECT 3.694 83.878 3.746 83.914 ;
               RECT 3.694 85.078 3.746 85.114 ;
               RECT 3.694 86.278 3.746 86.314 ;
               RECT 3.694 87.478 3.746 87.514 ;
               RECT 3.694 88.678 3.746 88.714 ;
               RECT 3.694 89.878 3.746 89.914 ;
               RECT 3.694 91.078 3.746 91.114 ;
               RECT 3.694 92.278 3.746 92.314 ;
               RECT 3.694 93.478 3.746 93.514 ;
               RECT 3.694 94.678 3.746 94.714 ;
               RECT 3.694 95.878 3.746 95.914 ;
               RECT 3.694 97.078 3.746 97.114 ;
               RECT 3.694 98.278 3.746 98.314 ;
               RECT 3.694 99.478 3.746 99.514 ;
               RECT 3.694 100.678 3.746 100.714 ;
               RECT 3.694 101.878 3.746 101.914 ;
               RECT 3.694 103.078 3.746 103.114 ;
               RECT 3.694 104.278 3.746 104.314 ;
               RECT 3.774 0.281 3.826 0.317 ;
               RECT 3.774 104.803 3.826 104.839 ;
               RECT 3.854 0.806 3.906 0.842 ;
               RECT 3.854 2.006 3.906 2.042 ;
               RECT 3.854 3.206 3.906 3.242 ;
               RECT 3.854 4.406 3.906 4.442 ;
               RECT 3.854 5.606 3.906 5.642 ;
               RECT 3.854 6.806 3.906 6.842 ;
               RECT 3.854 8.006 3.906 8.042 ;
               RECT 3.854 9.206 3.906 9.242 ;
               RECT 3.854 10.406 3.906 10.442 ;
               RECT 3.854 11.606 3.906 11.642 ;
               RECT 3.854 12.806 3.906 12.842 ;
               RECT 3.854 14.006 3.906 14.042 ;
               RECT 3.854 15.206 3.906 15.242 ;
               RECT 3.854 16.406 3.906 16.442 ;
               RECT 3.854 17.606 3.906 17.642 ;
               RECT 3.854 18.806 3.906 18.842 ;
               RECT 3.854 20.006 3.906 20.042 ;
               RECT 3.854 21.206 3.906 21.242 ;
               RECT 3.854 22.406 3.906 22.442 ;
               RECT 3.854 23.606 3.906 23.642 ;
               RECT 3.854 24.806 3.906 24.842 ;
               RECT 3.854 26.006 3.906 26.042 ;
               RECT 3.854 27.206 3.906 27.242 ;
               RECT 3.854 28.406 3.906 28.442 ;
               RECT 3.854 29.606 3.906 29.642 ;
               RECT 3.854 30.806 3.906 30.842 ;
               RECT 3.854 32.006 3.906 32.042 ;
               RECT 3.854 33.206 3.906 33.242 ;
               RECT 3.854 34.406 3.906 34.442 ;
               RECT 3.854 35.606 3.906 35.642 ;
               RECT 3.854 36.806 3.906 36.842 ;
               RECT 3.854 38.006 3.906 38.042 ;
               RECT 3.854 39.206 3.906 39.242 ;
               RECT 3.854 40.406 3.906 40.442 ;
               RECT 3.854 41.606 3.906 41.642 ;
               RECT 3.854 42.806 3.906 42.842 ;
               RECT 3.854 44.006 3.906 44.042 ;
               RECT 3.854 45.206 3.906 45.242 ;
               RECT 3.854 46.406 3.906 46.442 ;
               RECT 3.854 47.606 3.906 47.642 ;
               RECT 3.854 49.422 3.906 49.458 ;
               RECT 3.854 49.662 3.906 49.698 ;
               RECT 3.854 55.422 3.906 55.458 ;
               RECT 3.854 55.662 3.906 55.698 ;
               RECT 3.854 56.726 3.906 56.762 ;
               RECT 3.854 57.926 3.906 57.962 ;
               RECT 3.854 59.126 3.906 59.162 ;
               RECT 3.854 60.326 3.906 60.362 ;
               RECT 3.854 61.526 3.906 61.562 ;
               RECT 3.854 62.726 3.906 62.762 ;
               RECT 3.854 63.926 3.906 63.962 ;
               RECT 3.854 65.126 3.906 65.162 ;
               RECT 3.854 66.326 3.906 66.362 ;
               RECT 3.854 67.526 3.906 67.562 ;
               RECT 3.854 68.726 3.906 68.762 ;
               RECT 3.854 69.926 3.906 69.962 ;
               RECT 3.854 71.126 3.906 71.162 ;
               RECT 3.854 72.326 3.906 72.362 ;
               RECT 3.854 73.526 3.906 73.562 ;
               RECT 3.854 74.726 3.906 74.762 ;
               RECT 3.854 75.926 3.906 75.962 ;
               RECT 3.854 77.126 3.906 77.162 ;
               RECT 3.854 78.326 3.906 78.362 ;
               RECT 3.854 79.526 3.906 79.562 ;
               RECT 3.854 80.726 3.906 80.762 ;
               RECT 3.854 81.926 3.906 81.962 ;
               RECT 3.854 83.126 3.906 83.162 ;
               RECT 3.854 84.326 3.906 84.362 ;
               RECT 3.854 85.526 3.906 85.562 ;
               RECT 3.854 86.726 3.906 86.762 ;
               RECT 3.854 87.926 3.906 87.962 ;
               RECT 3.854 89.126 3.906 89.162 ;
               RECT 3.854 90.326 3.906 90.362 ;
               RECT 3.854 91.526 3.906 91.562 ;
               RECT 3.854 92.726 3.906 92.762 ;
               RECT 3.854 93.926 3.906 93.962 ;
               RECT 3.854 95.126 3.906 95.162 ;
               RECT 3.854 96.326 3.906 96.362 ;
               RECT 3.854 97.526 3.906 97.562 ;
               RECT 3.854 98.726 3.906 98.762 ;
               RECT 3.854 99.926 3.906 99.962 ;
               RECT 3.854 101.126 3.906 101.162 ;
               RECT 3.854 102.326 3.906 102.362 ;
               RECT 3.854 103.526 3.906 103.562 ;
               RECT 3.934 1.558 3.986 1.594 ;
               RECT 3.934 2.758 3.986 2.794 ;
               RECT 3.934 3.958 3.986 3.994 ;
               RECT 3.934 5.158 3.986 5.194 ;
               RECT 3.934 6.358 3.986 6.394 ;
               RECT 3.934 7.558 3.986 7.594 ;
               RECT 3.934 8.758 3.986 8.794 ;
               RECT 3.934 9.958 3.986 9.994 ;
               RECT 3.934 11.158 3.986 11.194 ;
               RECT 3.934 12.358 3.986 12.394 ;
               RECT 3.934 13.558 3.986 13.594 ;
               RECT 3.934 14.758 3.986 14.794 ;
               RECT 3.934 15.958 3.986 15.994 ;
               RECT 3.934 17.158 3.986 17.194 ;
               RECT 3.934 18.358 3.986 18.394 ;
               RECT 3.934 19.558 3.986 19.594 ;
               RECT 3.934 20.758 3.986 20.794 ;
               RECT 3.934 21.958 3.986 21.994 ;
               RECT 3.934 23.158 3.986 23.194 ;
               RECT 3.934 24.358 3.986 24.394 ;
               RECT 3.934 25.558 3.986 25.594 ;
               RECT 3.934 26.758 3.986 26.794 ;
               RECT 3.934 27.958 3.986 27.994 ;
               RECT 3.934 29.158 3.986 29.194 ;
               RECT 3.934 30.358 3.986 30.394 ;
               RECT 3.934 31.558 3.986 31.594 ;
               RECT 3.934 32.758 3.986 32.794 ;
               RECT 3.934 33.958 3.986 33.994 ;
               RECT 3.934 35.158 3.986 35.194 ;
               RECT 3.934 36.358 3.986 36.394 ;
               RECT 3.934 37.558 3.986 37.594 ;
               RECT 3.934 38.758 3.986 38.794 ;
               RECT 3.934 39.958 3.986 39.994 ;
               RECT 3.934 41.158 3.986 41.194 ;
               RECT 3.934 42.358 3.986 42.394 ;
               RECT 3.934 43.558 3.986 43.594 ;
               RECT 3.934 44.758 3.986 44.794 ;
               RECT 3.934 45.958 3.986 45.994 ;
               RECT 3.934 47.158 3.986 47.194 ;
               RECT 3.934 48.358 3.986 48.394 ;
               RECT 3.934 50.142 3.986 50.178 ;
               RECT 3.934 50.382 3.986 50.418 ;
               RECT 3.934 54.702 3.986 54.738 ;
               RECT 3.934 54.942 3.986 54.978 ;
               RECT 3.934 57.478 3.986 57.514 ;
               RECT 3.934 58.678 3.986 58.714 ;
               RECT 3.934 59.878 3.986 59.914 ;
               RECT 3.934 61.078 3.986 61.114 ;
               RECT 3.934 62.278 3.986 62.314 ;
               RECT 3.934 63.478 3.986 63.514 ;
               RECT 3.934 64.678 3.986 64.714 ;
               RECT 3.934 65.878 3.986 65.914 ;
               RECT 3.934 67.078 3.986 67.114 ;
               RECT 3.934 68.278 3.986 68.314 ;
               RECT 3.934 69.478 3.986 69.514 ;
               RECT 3.934 70.678 3.986 70.714 ;
               RECT 3.934 71.878 3.986 71.914 ;
               RECT 3.934 73.078 3.986 73.114 ;
               RECT 3.934 74.278 3.986 74.314 ;
               RECT 3.934 75.478 3.986 75.514 ;
               RECT 3.934 76.678 3.986 76.714 ;
               RECT 3.934 77.878 3.986 77.914 ;
               RECT 3.934 79.078 3.986 79.114 ;
               RECT 3.934 80.278 3.986 80.314 ;
               RECT 3.934 81.478 3.986 81.514 ;
               RECT 3.934 82.678 3.986 82.714 ;
               RECT 3.934 83.878 3.986 83.914 ;
               RECT 3.934 85.078 3.986 85.114 ;
               RECT 3.934 86.278 3.986 86.314 ;
               RECT 3.934 87.478 3.986 87.514 ;
               RECT 3.934 88.678 3.986 88.714 ;
               RECT 3.934 89.878 3.986 89.914 ;
               RECT 3.934 91.078 3.986 91.114 ;
               RECT 3.934 92.278 3.986 92.314 ;
               RECT 3.934 93.478 3.986 93.514 ;
               RECT 3.934 94.678 3.986 94.714 ;
               RECT 3.934 95.878 3.986 95.914 ;
               RECT 3.934 97.078 3.986 97.114 ;
               RECT 3.934 98.278 3.986 98.314 ;
               RECT 3.934 99.478 3.986 99.514 ;
               RECT 3.934 100.678 3.986 100.714 ;
               RECT 3.934 101.878 3.986 101.914 ;
               RECT 3.934 103.078 3.986 103.114 ;
               RECT 3.934 104.278 3.986 104.314 ;
               RECT 4.014 0.806 4.066 0.842 ;
               RECT 4.014 2.006 4.066 2.042 ;
               RECT 4.014 3.206 4.066 3.242 ;
               RECT 4.014 4.406 4.066 4.442 ;
               RECT 4.014 5.606 4.066 5.642 ;
               RECT 4.014 6.806 4.066 6.842 ;
               RECT 4.014 8.006 4.066 8.042 ;
               RECT 4.014 9.206 4.066 9.242 ;
               RECT 4.014 10.406 4.066 10.442 ;
               RECT 4.014 11.606 4.066 11.642 ;
               RECT 4.014 12.806 4.066 12.842 ;
               RECT 4.014 14.006 4.066 14.042 ;
               RECT 4.014 15.206 4.066 15.242 ;
               RECT 4.014 16.406 4.066 16.442 ;
               RECT 4.014 17.606 4.066 17.642 ;
               RECT 4.014 18.806 4.066 18.842 ;
               RECT 4.014 20.006 4.066 20.042 ;
               RECT 4.014 21.206 4.066 21.242 ;
               RECT 4.014 22.406 4.066 22.442 ;
               RECT 4.014 23.606 4.066 23.642 ;
               RECT 4.014 24.806 4.066 24.842 ;
               RECT 4.014 26.006 4.066 26.042 ;
               RECT 4.014 27.206 4.066 27.242 ;
               RECT 4.014 28.406 4.066 28.442 ;
               RECT 4.014 29.606 4.066 29.642 ;
               RECT 4.014 30.806 4.066 30.842 ;
               RECT 4.014 32.006 4.066 32.042 ;
               RECT 4.014 33.206 4.066 33.242 ;
               RECT 4.014 34.406 4.066 34.442 ;
               RECT 4.014 35.606 4.066 35.642 ;
               RECT 4.014 36.806 4.066 36.842 ;
               RECT 4.014 38.006 4.066 38.042 ;
               RECT 4.014 39.206 4.066 39.242 ;
               RECT 4.014 40.406 4.066 40.442 ;
               RECT 4.014 41.606 4.066 41.642 ;
               RECT 4.014 42.806 4.066 42.842 ;
               RECT 4.014 44.006 4.066 44.042 ;
               RECT 4.014 45.206 4.066 45.242 ;
               RECT 4.014 46.406 4.066 46.442 ;
               RECT 4.014 47.606 4.066 47.642 ;
               RECT 4.014 49.422 4.066 49.458 ;
               RECT 4.014 49.662 4.066 49.698 ;
               RECT 4.014 55.422 4.066 55.458 ;
               RECT 4.014 55.662 4.066 55.698 ;
               RECT 4.014 56.726 4.066 56.762 ;
               RECT 4.014 57.926 4.066 57.962 ;
               RECT 4.014 59.126 4.066 59.162 ;
               RECT 4.014 60.326 4.066 60.362 ;
               RECT 4.014 61.526 4.066 61.562 ;
               RECT 4.014 62.726 4.066 62.762 ;
               RECT 4.014 63.926 4.066 63.962 ;
               RECT 4.014 65.126 4.066 65.162 ;
               RECT 4.014 66.326 4.066 66.362 ;
               RECT 4.014 67.526 4.066 67.562 ;
               RECT 4.014 68.726 4.066 68.762 ;
               RECT 4.014 69.926 4.066 69.962 ;
               RECT 4.014 71.126 4.066 71.162 ;
               RECT 4.014 72.326 4.066 72.362 ;
               RECT 4.014 73.526 4.066 73.562 ;
               RECT 4.014 74.726 4.066 74.762 ;
               RECT 4.014 75.926 4.066 75.962 ;
               RECT 4.014 77.126 4.066 77.162 ;
               RECT 4.014 78.326 4.066 78.362 ;
               RECT 4.014 79.526 4.066 79.562 ;
               RECT 4.014 80.726 4.066 80.762 ;
               RECT 4.014 81.926 4.066 81.962 ;
               RECT 4.014 83.126 4.066 83.162 ;
               RECT 4.014 84.326 4.066 84.362 ;
               RECT 4.014 85.526 4.066 85.562 ;
               RECT 4.014 86.726 4.066 86.762 ;
               RECT 4.014 87.926 4.066 87.962 ;
               RECT 4.014 89.126 4.066 89.162 ;
               RECT 4.014 90.326 4.066 90.362 ;
               RECT 4.014 91.526 4.066 91.562 ;
               RECT 4.014 92.726 4.066 92.762 ;
               RECT 4.014 93.926 4.066 93.962 ;
               RECT 4.014 95.126 4.066 95.162 ;
               RECT 4.014 96.326 4.066 96.362 ;
               RECT 4.014 97.526 4.066 97.562 ;
               RECT 4.014 98.726 4.066 98.762 ;
               RECT 4.014 99.926 4.066 99.962 ;
               RECT 4.014 101.126 4.066 101.162 ;
               RECT 4.014 102.326 4.066 102.362 ;
               RECT 4.014 103.526 4.066 103.562 ;
               RECT 4.094 1.558 4.146 1.594 ;
               RECT 4.094 2.758 4.146 2.794 ;
               RECT 4.094 3.958 4.146 3.994 ;
               RECT 4.094 5.158 4.146 5.194 ;
               RECT 4.094 6.358 4.146 6.394 ;
               RECT 4.094 7.558 4.146 7.594 ;
               RECT 4.094 8.758 4.146 8.794 ;
               RECT 4.094 9.958 4.146 9.994 ;
               RECT 4.094 11.158 4.146 11.194 ;
               RECT 4.094 12.358 4.146 12.394 ;
               RECT 4.094 13.558 4.146 13.594 ;
               RECT 4.094 14.758 4.146 14.794 ;
               RECT 4.094 15.958 4.146 15.994 ;
               RECT 4.094 17.158 4.146 17.194 ;
               RECT 4.094 18.358 4.146 18.394 ;
               RECT 4.094 19.558 4.146 19.594 ;
               RECT 4.094 20.758 4.146 20.794 ;
               RECT 4.094 21.958 4.146 21.994 ;
               RECT 4.094 23.158 4.146 23.194 ;
               RECT 4.094 24.358 4.146 24.394 ;
               RECT 4.094 25.558 4.146 25.594 ;
               RECT 4.094 26.758 4.146 26.794 ;
               RECT 4.094 27.958 4.146 27.994 ;
               RECT 4.094 29.158 4.146 29.194 ;
               RECT 4.094 30.358 4.146 30.394 ;
               RECT 4.094 31.558 4.146 31.594 ;
               RECT 4.094 32.758 4.146 32.794 ;
               RECT 4.094 33.958 4.146 33.994 ;
               RECT 4.094 35.158 4.146 35.194 ;
               RECT 4.094 36.358 4.146 36.394 ;
               RECT 4.094 37.558 4.146 37.594 ;
               RECT 4.094 38.758 4.146 38.794 ;
               RECT 4.094 39.958 4.146 39.994 ;
               RECT 4.094 41.158 4.146 41.194 ;
               RECT 4.094 42.358 4.146 42.394 ;
               RECT 4.094 43.558 4.146 43.594 ;
               RECT 4.094 44.758 4.146 44.794 ;
               RECT 4.094 45.958 4.146 45.994 ;
               RECT 4.094 47.158 4.146 47.194 ;
               RECT 4.094 48.358 4.146 48.394 ;
               RECT 4.094 50.142 4.146 50.178 ;
               RECT 4.094 50.382 4.146 50.418 ;
               RECT 4.094 54.702 4.146 54.738 ;
               RECT 4.094 54.942 4.146 54.978 ;
               RECT 4.094 57.478 4.146 57.514 ;
               RECT 4.094 58.678 4.146 58.714 ;
               RECT 4.094 59.878 4.146 59.914 ;
               RECT 4.094 61.078 4.146 61.114 ;
               RECT 4.094 62.278 4.146 62.314 ;
               RECT 4.094 63.478 4.146 63.514 ;
               RECT 4.094 64.678 4.146 64.714 ;
               RECT 4.094 65.878 4.146 65.914 ;
               RECT 4.094 67.078 4.146 67.114 ;
               RECT 4.094 68.278 4.146 68.314 ;
               RECT 4.094 69.478 4.146 69.514 ;
               RECT 4.094 70.678 4.146 70.714 ;
               RECT 4.094 71.878 4.146 71.914 ;
               RECT 4.094 73.078 4.146 73.114 ;
               RECT 4.094 74.278 4.146 74.314 ;
               RECT 4.094 75.478 4.146 75.514 ;
               RECT 4.094 76.678 4.146 76.714 ;
               RECT 4.094 77.878 4.146 77.914 ;
               RECT 4.094 79.078 4.146 79.114 ;
               RECT 4.094 80.278 4.146 80.314 ;
               RECT 4.094 81.478 4.146 81.514 ;
               RECT 4.094 82.678 4.146 82.714 ;
               RECT 4.094 83.878 4.146 83.914 ;
               RECT 4.094 85.078 4.146 85.114 ;
               RECT 4.094 86.278 4.146 86.314 ;
               RECT 4.094 87.478 4.146 87.514 ;
               RECT 4.094 88.678 4.146 88.714 ;
               RECT 4.094 89.878 4.146 89.914 ;
               RECT 4.094 91.078 4.146 91.114 ;
               RECT 4.094 92.278 4.146 92.314 ;
               RECT 4.094 93.478 4.146 93.514 ;
               RECT 4.094 94.678 4.146 94.714 ;
               RECT 4.094 95.878 4.146 95.914 ;
               RECT 4.094 97.078 4.146 97.114 ;
               RECT 4.094 98.278 4.146 98.314 ;
               RECT 4.094 99.478 4.146 99.514 ;
               RECT 4.094 100.678 4.146 100.714 ;
               RECT 4.094 101.878 4.146 101.914 ;
               RECT 4.094 103.078 4.146 103.114 ;
               RECT 4.094 104.278 4.146 104.314 ;
               RECT 4.174 0.281 4.226 0.317 ;
               RECT 4.174 104.803 4.226 104.839 ;
               RECT 4.254 0.806 4.306 0.842 ;
               RECT 4.254 2.006 4.306 2.042 ;
               RECT 4.254 3.206 4.306 3.242 ;
               RECT 4.254 4.406 4.306 4.442 ;
               RECT 4.254 5.606 4.306 5.642 ;
               RECT 4.254 6.806 4.306 6.842 ;
               RECT 4.254 8.006 4.306 8.042 ;
               RECT 4.254 9.206 4.306 9.242 ;
               RECT 4.254 10.406 4.306 10.442 ;
               RECT 4.254 11.606 4.306 11.642 ;
               RECT 4.254 12.806 4.306 12.842 ;
               RECT 4.254 14.006 4.306 14.042 ;
               RECT 4.254 15.206 4.306 15.242 ;
               RECT 4.254 16.406 4.306 16.442 ;
               RECT 4.254 17.606 4.306 17.642 ;
               RECT 4.254 18.806 4.306 18.842 ;
               RECT 4.254 20.006 4.306 20.042 ;
               RECT 4.254 21.206 4.306 21.242 ;
               RECT 4.254 22.406 4.306 22.442 ;
               RECT 4.254 23.606 4.306 23.642 ;
               RECT 4.254 24.806 4.306 24.842 ;
               RECT 4.254 26.006 4.306 26.042 ;
               RECT 4.254 27.206 4.306 27.242 ;
               RECT 4.254 28.406 4.306 28.442 ;
               RECT 4.254 29.606 4.306 29.642 ;
               RECT 4.254 30.806 4.306 30.842 ;
               RECT 4.254 32.006 4.306 32.042 ;
               RECT 4.254 33.206 4.306 33.242 ;
               RECT 4.254 34.406 4.306 34.442 ;
               RECT 4.254 35.606 4.306 35.642 ;
               RECT 4.254 36.806 4.306 36.842 ;
               RECT 4.254 38.006 4.306 38.042 ;
               RECT 4.254 39.206 4.306 39.242 ;
               RECT 4.254 40.406 4.306 40.442 ;
               RECT 4.254 41.606 4.306 41.642 ;
               RECT 4.254 42.806 4.306 42.842 ;
               RECT 4.254 44.006 4.306 44.042 ;
               RECT 4.254 45.206 4.306 45.242 ;
               RECT 4.254 46.406 4.306 46.442 ;
               RECT 4.254 47.606 4.306 47.642 ;
               RECT 4.254 49.422 4.306 49.458 ;
               RECT 4.254 49.662 4.306 49.698 ;
               RECT 4.254 51.102 4.306 51.138 ;
               RECT 4.254 51.582 4.306 51.618 ;
               RECT 4.254 53.502 4.306 53.538 ;
               RECT 4.254 53.982 4.306 54.018 ;
               RECT 4.254 55.422 4.306 55.458 ;
               RECT 4.254 55.662 4.306 55.698 ;
               RECT 4.254 56.726 4.306 56.762 ;
               RECT 4.254 57.926 4.306 57.962 ;
               RECT 4.254 59.126 4.306 59.162 ;
               RECT 4.254 60.326 4.306 60.362 ;
               RECT 4.254 61.526 4.306 61.562 ;
               RECT 4.254 62.726 4.306 62.762 ;
               RECT 4.254 63.926 4.306 63.962 ;
               RECT 4.254 65.126 4.306 65.162 ;
               RECT 4.254 66.326 4.306 66.362 ;
               RECT 4.254 67.526 4.306 67.562 ;
               RECT 4.254 68.726 4.306 68.762 ;
               RECT 4.254 69.926 4.306 69.962 ;
               RECT 4.254 71.126 4.306 71.162 ;
               RECT 4.254 72.326 4.306 72.362 ;
               RECT 4.254 73.526 4.306 73.562 ;
               RECT 4.254 74.726 4.306 74.762 ;
               RECT 4.254 75.926 4.306 75.962 ;
               RECT 4.254 77.126 4.306 77.162 ;
               RECT 4.254 78.326 4.306 78.362 ;
               RECT 4.254 79.526 4.306 79.562 ;
               RECT 4.254 80.726 4.306 80.762 ;
               RECT 4.254 81.926 4.306 81.962 ;
               RECT 4.254 83.126 4.306 83.162 ;
               RECT 4.254 84.326 4.306 84.362 ;
               RECT 4.254 85.526 4.306 85.562 ;
               RECT 4.254 86.726 4.306 86.762 ;
               RECT 4.254 87.926 4.306 87.962 ;
               RECT 4.254 89.126 4.306 89.162 ;
               RECT 4.254 90.326 4.306 90.362 ;
               RECT 4.254 91.526 4.306 91.562 ;
               RECT 4.254 92.726 4.306 92.762 ;
               RECT 4.254 93.926 4.306 93.962 ;
               RECT 4.254 95.126 4.306 95.162 ;
               RECT 4.254 96.326 4.306 96.362 ;
               RECT 4.254 97.526 4.306 97.562 ;
               RECT 4.254 98.726 4.306 98.762 ;
               RECT 4.254 99.926 4.306 99.962 ;
               RECT 4.254 101.126 4.306 101.162 ;
               RECT 4.254 102.326 4.306 102.362 ;
               RECT 4.254 103.526 4.306 103.562 ;
               RECT 4.334 1.558 4.386 1.594 ;
               RECT 4.334 2.758 4.386 2.794 ;
               RECT 4.334 3.958 4.386 3.994 ;
               RECT 4.334 5.158 4.386 5.194 ;
               RECT 4.334 6.358 4.386 6.394 ;
               RECT 4.334 7.558 4.386 7.594 ;
               RECT 4.334 8.758 4.386 8.794 ;
               RECT 4.334 9.958 4.386 9.994 ;
               RECT 4.334 11.158 4.386 11.194 ;
               RECT 4.334 12.358 4.386 12.394 ;
               RECT 4.334 13.558 4.386 13.594 ;
               RECT 4.334 14.758 4.386 14.794 ;
               RECT 4.334 15.958 4.386 15.994 ;
               RECT 4.334 17.158 4.386 17.194 ;
               RECT 4.334 18.358 4.386 18.394 ;
               RECT 4.334 19.558 4.386 19.594 ;
               RECT 4.334 20.758 4.386 20.794 ;
               RECT 4.334 21.958 4.386 21.994 ;
               RECT 4.334 23.158 4.386 23.194 ;
               RECT 4.334 24.358 4.386 24.394 ;
               RECT 4.334 25.558 4.386 25.594 ;
               RECT 4.334 26.758 4.386 26.794 ;
               RECT 4.334 27.958 4.386 27.994 ;
               RECT 4.334 29.158 4.386 29.194 ;
               RECT 4.334 30.358 4.386 30.394 ;
               RECT 4.334 31.558 4.386 31.594 ;
               RECT 4.334 32.758 4.386 32.794 ;
               RECT 4.334 33.958 4.386 33.994 ;
               RECT 4.334 35.158 4.386 35.194 ;
               RECT 4.334 36.358 4.386 36.394 ;
               RECT 4.334 37.558 4.386 37.594 ;
               RECT 4.334 38.758 4.386 38.794 ;
               RECT 4.334 39.958 4.386 39.994 ;
               RECT 4.334 41.158 4.386 41.194 ;
               RECT 4.334 42.358 4.386 42.394 ;
               RECT 4.334 43.558 4.386 43.594 ;
               RECT 4.334 44.758 4.386 44.794 ;
               RECT 4.334 45.958 4.386 45.994 ;
               RECT 4.334 47.158 4.386 47.194 ;
               RECT 4.334 48.358 4.386 48.394 ;
               RECT 4.334 50.142 4.386 50.178 ;
               RECT 4.334 50.382 4.386 50.418 ;
               RECT 4.334 54.702 4.386 54.738 ;
               RECT 4.334 54.942 4.386 54.978 ;
               RECT 4.334 57.478 4.386 57.514 ;
               RECT 4.334 58.678 4.386 58.714 ;
               RECT 4.334 59.878 4.386 59.914 ;
               RECT 4.334 61.078 4.386 61.114 ;
               RECT 4.334 62.278 4.386 62.314 ;
               RECT 4.334 63.478 4.386 63.514 ;
               RECT 4.334 64.678 4.386 64.714 ;
               RECT 4.334 65.878 4.386 65.914 ;
               RECT 4.334 67.078 4.386 67.114 ;
               RECT 4.334 68.278 4.386 68.314 ;
               RECT 4.334 69.478 4.386 69.514 ;
               RECT 4.334 70.678 4.386 70.714 ;
               RECT 4.334 71.878 4.386 71.914 ;
               RECT 4.334 73.078 4.386 73.114 ;
               RECT 4.334 74.278 4.386 74.314 ;
               RECT 4.334 75.478 4.386 75.514 ;
               RECT 4.334 76.678 4.386 76.714 ;
               RECT 4.334 77.878 4.386 77.914 ;
               RECT 4.334 79.078 4.386 79.114 ;
               RECT 4.334 80.278 4.386 80.314 ;
               RECT 4.334 81.478 4.386 81.514 ;
               RECT 4.334 82.678 4.386 82.714 ;
               RECT 4.334 83.878 4.386 83.914 ;
               RECT 4.334 85.078 4.386 85.114 ;
               RECT 4.334 86.278 4.386 86.314 ;
               RECT 4.334 87.478 4.386 87.514 ;
               RECT 4.334 88.678 4.386 88.714 ;
               RECT 4.334 89.878 4.386 89.914 ;
               RECT 4.334 91.078 4.386 91.114 ;
               RECT 4.334 92.278 4.386 92.314 ;
               RECT 4.334 93.478 4.386 93.514 ;
               RECT 4.334 94.678 4.386 94.714 ;
               RECT 4.334 95.878 4.386 95.914 ;
               RECT 4.334 97.078 4.386 97.114 ;
               RECT 4.334 98.278 4.386 98.314 ;
               RECT 4.334 99.478 4.386 99.514 ;
               RECT 4.334 100.678 4.386 100.714 ;
               RECT 4.334 101.878 4.386 101.914 ;
               RECT 4.334 103.078 4.386 103.114 ;
               RECT 4.334 104.278 4.386 104.314 ;
               RECT 4.414 0.806 4.466 0.842 ;
               RECT 4.414 2.006 4.466 2.042 ;
               RECT 4.414 3.206 4.466 3.242 ;
               RECT 4.414 4.406 4.466 4.442 ;
               RECT 4.414 5.606 4.466 5.642 ;
               RECT 4.414 6.806 4.466 6.842 ;
               RECT 4.414 8.006 4.466 8.042 ;
               RECT 4.414 9.206 4.466 9.242 ;
               RECT 4.414 10.406 4.466 10.442 ;
               RECT 4.414 11.606 4.466 11.642 ;
               RECT 4.414 12.806 4.466 12.842 ;
               RECT 4.414 14.006 4.466 14.042 ;
               RECT 4.414 15.206 4.466 15.242 ;
               RECT 4.414 16.406 4.466 16.442 ;
               RECT 4.414 17.606 4.466 17.642 ;
               RECT 4.414 18.806 4.466 18.842 ;
               RECT 4.414 20.006 4.466 20.042 ;
               RECT 4.414 21.206 4.466 21.242 ;
               RECT 4.414 22.406 4.466 22.442 ;
               RECT 4.414 23.606 4.466 23.642 ;
               RECT 4.414 24.806 4.466 24.842 ;
               RECT 4.414 26.006 4.466 26.042 ;
               RECT 4.414 27.206 4.466 27.242 ;
               RECT 4.414 28.406 4.466 28.442 ;
               RECT 4.414 29.606 4.466 29.642 ;
               RECT 4.414 30.806 4.466 30.842 ;
               RECT 4.414 32.006 4.466 32.042 ;
               RECT 4.414 33.206 4.466 33.242 ;
               RECT 4.414 34.406 4.466 34.442 ;
               RECT 4.414 35.606 4.466 35.642 ;
               RECT 4.414 36.806 4.466 36.842 ;
               RECT 4.414 38.006 4.466 38.042 ;
               RECT 4.414 39.206 4.466 39.242 ;
               RECT 4.414 40.406 4.466 40.442 ;
               RECT 4.414 41.606 4.466 41.642 ;
               RECT 4.414 42.806 4.466 42.842 ;
               RECT 4.414 44.006 4.466 44.042 ;
               RECT 4.414 45.206 4.466 45.242 ;
               RECT 4.414 46.406 4.466 46.442 ;
               RECT 4.414 47.606 4.466 47.642 ;
               RECT 4.414 49.422 4.466 49.458 ;
               RECT 4.414 49.662 4.466 49.698 ;
               RECT 4.414 55.422 4.466 55.458 ;
               RECT 4.414 55.662 4.466 55.698 ;
               RECT 4.414 56.726 4.466 56.762 ;
               RECT 4.414 57.926 4.466 57.962 ;
               RECT 4.414 59.126 4.466 59.162 ;
               RECT 4.414 60.326 4.466 60.362 ;
               RECT 4.414 61.526 4.466 61.562 ;
               RECT 4.414 62.726 4.466 62.762 ;
               RECT 4.414 63.926 4.466 63.962 ;
               RECT 4.414 65.126 4.466 65.162 ;
               RECT 4.414 66.326 4.466 66.362 ;
               RECT 4.414 67.526 4.466 67.562 ;
               RECT 4.414 68.726 4.466 68.762 ;
               RECT 4.414 69.926 4.466 69.962 ;
               RECT 4.414 71.126 4.466 71.162 ;
               RECT 4.414 72.326 4.466 72.362 ;
               RECT 4.414 73.526 4.466 73.562 ;
               RECT 4.414 74.726 4.466 74.762 ;
               RECT 4.414 75.926 4.466 75.962 ;
               RECT 4.414 77.126 4.466 77.162 ;
               RECT 4.414 78.326 4.466 78.362 ;
               RECT 4.414 79.526 4.466 79.562 ;
               RECT 4.414 80.726 4.466 80.762 ;
               RECT 4.414 81.926 4.466 81.962 ;
               RECT 4.414 83.126 4.466 83.162 ;
               RECT 4.414 84.326 4.466 84.362 ;
               RECT 4.414 85.526 4.466 85.562 ;
               RECT 4.414 86.726 4.466 86.762 ;
               RECT 4.414 87.926 4.466 87.962 ;
               RECT 4.414 89.126 4.466 89.162 ;
               RECT 4.414 90.326 4.466 90.362 ;
               RECT 4.414 91.526 4.466 91.562 ;
               RECT 4.414 92.726 4.466 92.762 ;
               RECT 4.414 93.926 4.466 93.962 ;
               RECT 4.414 95.126 4.466 95.162 ;
               RECT 4.414 96.326 4.466 96.362 ;
               RECT 4.414 97.526 4.466 97.562 ;
               RECT 4.414 98.726 4.466 98.762 ;
               RECT 4.414 99.926 4.466 99.962 ;
               RECT 4.414 101.126 4.466 101.162 ;
               RECT 4.414 102.326 4.466 102.362 ;
               RECT 4.414 103.526 4.466 103.562 ;
               RECT 4.494 1.558 4.546 1.594 ;
               RECT 4.494 2.758 4.546 2.794 ;
               RECT 4.494 3.958 4.546 3.994 ;
               RECT 4.494 5.158 4.546 5.194 ;
               RECT 4.494 6.358 4.546 6.394 ;
               RECT 4.494 7.558 4.546 7.594 ;
               RECT 4.494 8.758 4.546 8.794 ;
               RECT 4.494 9.958 4.546 9.994 ;
               RECT 4.494 11.158 4.546 11.194 ;
               RECT 4.494 12.358 4.546 12.394 ;
               RECT 4.494 13.558 4.546 13.594 ;
               RECT 4.494 14.758 4.546 14.794 ;
               RECT 4.494 15.958 4.546 15.994 ;
               RECT 4.494 17.158 4.546 17.194 ;
               RECT 4.494 18.358 4.546 18.394 ;
               RECT 4.494 19.558 4.546 19.594 ;
               RECT 4.494 20.758 4.546 20.794 ;
               RECT 4.494 21.958 4.546 21.994 ;
               RECT 4.494 23.158 4.546 23.194 ;
               RECT 4.494 24.358 4.546 24.394 ;
               RECT 4.494 25.558 4.546 25.594 ;
               RECT 4.494 26.758 4.546 26.794 ;
               RECT 4.494 27.958 4.546 27.994 ;
               RECT 4.494 29.158 4.546 29.194 ;
               RECT 4.494 30.358 4.546 30.394 ;
               RECT 4.494 31.558 4.546 31.594 ;
               RECT 4.494 32.758 4.546 32.794 ;
               RECT 4.494 33.958 4.546 33.994 ;
               RECT 4.494 35.158 4.546 35.194 ;
               RECT 4.494 36.358 4.546 36.394 ;
               RECT 4.494 37.558 4.546 37.594 ;
               RECT 4.494 38.758 4.546 38.794 ;
               RECT 4.494 39.958 4.546 39.994 ;
               RECT 4.494 41.158 4.546 41.194 ;
               RECT 4.494 42.358 4.546 42.394 ;
               RECT 4.494 43.558 4.546 43.594 ;
               RECT 4.494 44.758 4.546 44.794 ;
               RECT 4.494 45.958 4.546 45.994 ;
               RECT 4.494 47.158 4.546 47.194 ;
               RECT 4.494 48.358 4.546 48.394 ;
               RECT 4.494 50.142 4.546 50.178 ;
               RECT 4.494 50.382 4.546 50.418 ;
               RECT 4.494 54.702 4.546 54.738 ;
               RECT 4.494 54.942 4.546 54.978 ;
               RECT 4.494 57.478 4.546 57.514 ;
               RECT 4.494 58.678 4.546 58.714 ;
               RECT 4.494 59.878 4.546 59.914 ;
               RECT 4.494 61.078 4.546 61.114 ;
               RECT 4.494 62.278 4.546 62.314 ;
               RECT 4.494 63.478 4.546 63.514 ;
               RECT 4.494 64.678 4.546 64.714 ;
               RECT 4.494 65.878 4.546 65.914 ;
               RECT 4.494 67.078 4.546 67.114 ;
               RECT 4.494 68.278 4.546 68.314 ;
               RECT 4.494 69.478 4.546 69.514 ;
               RECT 4.494 70.678 4.546 70.714 ;
               RECT 4.494 71.878 4.546 71.914 ;
               RECT 4.494 73.078 4.546 73.114 ;
               RECT 4.494 74.278 4.546 74.314 ;
               RECT 4.494 75.478 4.546 75.514 ;
               RECT 4.494 76.678 4.546 76.714 ;
               RECT 4.494 77.878 4.546 77.914 ;
               RECT 4.494 79.078 4.546 79.114 ;
               RECT 4.494 80.278 4.546 80.314 ;
               RECT 4.494 81.478 4.546 81.514 ;
               RECT 4.494 82.678 4.546 82.714 ;
               RECT 4.494 83.878 4.546 83.914 ;
               RECT 4.494 85.078 4.546 85.114 ;
               RECT 4.494 86.278 4.546 86.314 ;
               RECT 4.494 87.478 4.546 87.514 ;
               RECT 4.494 88.678 4.546 88.714 ;
               RECT 4.494 89.878 4.546 89.914 ;
               RECT 4.494 91.078 4.546 91.114 ;
               RECT 4.494 92.278 4.546 92.314 ;
               RECT 4.494 93.478 4.546 93.514 ;
               RECT 4.494 94.678 4.546 94.714 ;
               RECT 4.494 95.878 4.546 95.914 ;
               RECT 4.494 97.078 4.546 97.114 ;
               RECT 4.494 98.278 4.546 98.314 ;
               RECT 4.494 99.478 4.546 99.514 ;
               RECT 4.494 100.678 4.546 100.714 ;
               RECT 4.494 101.878 4.546 101.914 ;
               RECT 4.494 103.078 4.546 103.114 ;
               RECT 4.494 104.278 4.546 104.314 ;
               RECT 4.574 0.281 4.626 0.317 ;
               RECT 4.574 104.803 4.626 104.839 ;
               RECT 4.654 0.806 4.706 0.842 ;
               RECT 4.654 2.006 4.706 2.042 ;
               RECT 4.654 3.206 4.706 3.242 ;
               RECT 4.654 4.406 4.706 4.442 ;
               RECT 4.654 5.606 4.706 5.642 ;
               RECT 4.654 6.806 4.706 6.842 ;
               RECT 4.654 8.006 4.706 8.042 ;
               RECT 4.654 9.206 4.706 9.242 ;
               RECT 4.654 10.406 4.706 10.442 ;
               RECT 4.654 11.606 4.706 11.642 ;
               RECT 4.654 12.806 4.706 12.842 ;
               RECT 4.654 14.006 4.706 14.042 ;
               RECT 4.654 15.206 4.706 15.242 ;
               RECT 4.654 16.406 4.706 16.442 ;
               RECT 4.654 17.606 4.706 17.642 ;
               RECT 4.654 18.806 4.706 18.842 ;
               RECT 4.654 20.006 4.706 20.042 ;
               RECT 4.654 21.206 4.706 21.242 ;
               RECT 4.654 22.406 4.706 22.442 ;
               RECT 4.654 23.606 4.706 23.642 ;
               RECT 4.654 24.806 4.706 24.842 ;
               RECT 4.654 26.006 4.706 26.042 ;
               RECT 4.654 27.206 4.706 27.242 ;
               RECT 4.654 28.406 4.706 28.442 ;
               RECT 4.654 29.606 4.706 29.642 ;
               RECT 4.654 30.806 4.706 30.842 ;
               RECT 4.654 32.006 4.706 32.042 ;
               RECT 4.654 33.206 4.706 33.242 ;
               RECT 4.654 34.406 4.706 34.442 ;
               RECT 4.654 35.606 4.706 35.642 ;
               RECT 4.654 36.806 4.706 36.842 ;
               RECT 4.654 38.006 4.706 38.042 ;
               RECT 4.654 39.206 4.706 39.242 ;
               RECT 4.654 40.406 4.706 40.442 ;
               RECT 4.654 41.606 4.706 41.642 ;
               RECT 4.654 42.806 4.706 42.842 ;
               RECT 4.654 44.006 4.706 44.042 ;
               RECT 4.654 45.206 4.706 45.242 ;
               RECT 4.654 46.406 4.706 46.442 ;
               RECT 4.654 47.606 4.706 47.642 ;
               RECT 4.654 49.422 4.706 49.458 ;
               RECT 4.654 49.662 4.706 49.698 ;
               RECT 4.654 55.422 4.706 55.458 ;
               RECT 4.654 55.662 4.706 55.698 ;
               RECT 4.654 56.726 4.706 56.762 ;
               RECT 4.654 57.926 4.706 57.962 ;
               RECT 4.654 59.126 4.706 59.162 ;
               RECT 4.654 60.326 4.706 60.362 ;
               RECT 4.654 61.526 4.706 61.562 ;
               RECT 4.654 62.726 4.706 62.762 ;
               RECT 4.654 63.926 4.706 63.962 ;
               RECT 4.654 65.126 4.706 65.162 ;
               RECT 4.654 66.326 4.706 66.362 ;
               RECT 4.654 67.526 4.706 67.562 ;
               RECT 4.654 68.726 4.706 68.762 ;
               RECT 4.654 69.926 4.706 69.962 ;
               RECT 4.654 71.126 4.706 71.162 ;
               RECT 4.654 72.326 4.706 72.362 ;
               RECT 4.654 73.526 4.706 73.562 ;
               RECT 4.654 74.726 4.706 74.762 ;
               RECT 4.654 75.926 4.706 75.962 ;
               RECT 4.654 77.126 4.706 77.162 ;
               RECT 4.654 78.326 4.706 78.362 ;
               RECT 4.654 79.526 4.706 79.562 ;
               RECT 4.654 80.726 4.706 80.762 ;
               RECT 4.654 81.926 4.706 81.962 ;
               RECT 4.654 83.126 4.706 83.162 ;
               RECT 4.654 84.326 4.706 84.362 ;
               RECT 4.654 85.526 4.706 85.562 ;
               RECT 4.654 86.726 4.706 86.762 ;
               RECT 4.654 87.926 4.706 87.962 ;
               RECT 4.654 89.126 4.706 89.162 ;
               RECT 4.654 90.326 4.706 90.362 ;
               RECT 4.654 91.526 4.706 91.562 ;
               RECT 4.654 92.726 4.706 92.762 ;
               RECT 4.654 93.926 4.706 93.962 ;
               RECT 4.654 95.126 4.706 95.162 ;
               RECT 4.654 96.326 4.706 96.362 ;
               RECT 4.654 97.526 4.706 97.562 ;
               RECT 4.654 98.726 4.706 98.762 ;
               RECT 4.654 99.926 4.706 99.962 ;
               RECT 4.654 101.126 4.706 101.162 ;
               RECT 4.654 102.326 4.706 102.362 ;
               RECT 4.654 103.526 4.706 103.562 ;
               RECT 4.734 1.558 4.786 1.594 ;
               RECT 4.734 2.758 4.786 2.794 ;
               RECT 4.734 3.958 4.786 3.994 ;
               RECT 4.734 5.158 4.786 5.194 ;
               RECT 4.734 6.358 4.786 6.394 ;
               RECT 4.734 7.558 4.786 7.594 ;
               RECT 4.734 8.758 4.786 8.794 ;
               RECT 4.734 9.958 4.786 9.994 ;
               RECT 4.734 11.158 4.786 11.194 ;
               RECT 4.734 12.358 4.786 12.394 ;
               RECT 4.734 13.558 4.786 13.594 ;
               RECT 4.734 14.758 4.786 14.794 ;
               RECT 4.734 15.958 4.786 15.994 ;
               RECT 4.734 17.158 4.786 17.194 ;
               RECT 4.734 18.358 4.786 18.394 ;
               RECT 4.734 19.558 4.786 19.594 ;
               RECT 4.734 20.758 4.786 20.794 ;
               RECT 4.734 21.958 4.786 21.994 ;
               RECT 4.734 23.158 4.786 23.194 ;
               RECT 4.734 24.358 4.786 24.394 ;
               RECT 4.734 25.558 4.786 25.594 ;
               RECT 4.734 26.758 4.786 26.794 ;
               RECT 4.734 27.958 4.786 27.994 ;
               RECT 4.734 29.158 4.786 29.194 ;
               RECT 4.734 30.358 4.786 30.394 ;
               RECT 4.734 31.558 4.786 31.594 ;
               RECT 4.734 32.758 4.786 32.794 ;
               RECT 4.734 33.958 4.786 33.994 ;
               RECT 4.734 35.158 4.786 35.194 ;
               RECT 4.734 36.358 4.786 36.394 ;
               RECT 4.734 37.558 4.786 37.594 ;
               RECT 4.734 38.758 4.786 38.794 ;
               RECT 4.734 39.958 4.786 39.994 ;
               RECT 4.734 41.158 4.786 41.194 ;
               RECT 4.734 42.358 4.786 42.394 ;
               RECT 4.734 43.558 4.786 43.594 ;
               RECT 4.734 44.758 4.786 44.794 ;
               RECT 4.734 45.958 4.786 45.994 ;
               RECT 4.734 47.158 4.786 47.194 ;
               RECT 4.734 48.358 4.786 48.394 ;
               RECT 4.734 50.142 4.786 50.178 ;
               RECT 4.734 50.382 4.786 50.418 ;
               RECT 4.734 54.702 4.786 54.738 ;
               RECT 4.734 54.942 4.786 54.978 ;
               RECT 4.734 57.478 4.786 57.514 ;
               RECT 4.734 58.678 4.786 58.714 ;
               RECT 4.734 59.878 4.786 59.914 ;
               RECT 4.734 61.078 4.786 61.114 ;
               RECT 4.734 62.278 4.786 62.314 ;
               RECT 4.734 63.478 4.786 63.514 ;
               RECT 4.734 64.678 4.786 64.714 ;
               RECT 4.734 65.878 4.786 65.914 ;
               RECT 4.734 67.078 4.786 67.114 ;
               RECT 4.734 68.278 4.786 68.314 ;
               RECT 4.734 69.478 4.786 69.514 ;
               RECT 4.734 70.678 4.786 70.714 ;
               RECT 4.734 71.878 4.786 71.914 ;
               RECT 4.734 73.078 4.786 73.114 ;
               RECT 4.734 74.278 4.786 74.314 ;
               RECT 4.734 75.478 4.786 75.514 ;
               RECT 4.734 76.678 4.786 76.714 ;
               RECT 4.734 77.878 4.786 77.914 ;
               RECT 4.734 79.078 4.786 79.114 ;
               RECT 4.734 80.278 4.786 80.314 ;
               RECT 4.734 81.478 4.786 81.514 ;
               RECT 4.734 82.678 4.786 82.714 ;
               RECT 4.734 83.878 4.786 83.914 ;
               RECT 4.734 85.078 4.786 85.114 ;
               RECT 4.734 86.278 4.786 86.314 ;
               RECT 4.734 87.478 4.786 87.514 ;
               RECT 4.734 88.678 4.786 88.714 ;
               RECT 4.734 89.878 4.786 89.914 ;
               RECT 4.734 91.078 4.786 91.114 ;
               RECT 4.734 92.278 4.786 92.314 ;
               RECT 4.734 93.478 4.786 93.514 ;
               RECT 4.734 94.678 4.786 94.714 ;
               RECT 4.734 95.878 4.786 95.914 ;
               RECT 4.734 97.078 4.786 97.114 ;
               RECT 4.734 98.278 4.786 98.314 ;
               RECT 4.734 99.478 4.786 99.514 ;
               RECT 4.734 100.678 4.786 100.714 ;
               RECT 4.734 101.878 4.786 101.914 ;
               RECT 4.734 103.078 4.786 103.114 ;
               RECT 4.734 104.278 4.786 104.314 ;
               RECT 4.814 0.806 4.866 0.842 ;
               RECT 4.814 2.006 4.866 2.042 ;
               RECT 4.814 3.206 4.866 3.242 ;
               RECT 4.814 4.406 4.866 4.442 ;
               RECT 4.814 5.606 4.866 5.642 ;
               RECT 4.814 6.806 4.866 6.842 ;
               RECT 4.814 8.006 4.866 8.042 ;
               RECT 4.814 9.206 4.866 9.242 ;
               RECT 4.814 10.406 4.866 10.442 ;
               RECT 4.814 11.606 4.866 11.642 ;
               RECT 4.814 12.806 4.866 12.842 ;
               RECT 4.814 14.006 4.866 14.042 ;
               RECT 4.814 15.206 4.866 15.242 ;
               RECT 4.814 16.406 4.866 16.442 ;
               RECT 4.814 17.606 4.866 17.642 ;
               RECT 4.814 18.806 4.866 18.842 ;
               RECT 4.814 20.006 4.866 20.042 ;
               RECT 4.814 21.206 4.866 21.242 ;
               RECT 4.814 22.406 4.866 22.442 ;
               RECT 4.814 23.606 4.866 23.642 ;
               RECT 4.814 24.806 4.866 24.842 ;
               RECT 4.814 26.006 4.866 26.042 ;
               RECT 4.814 27.206 4.866 27.242 ;
               RECT 4.814 28.406 4.866 28.442 ;
               RECT 4.814 29.606 4.866 29.642 ;
               RECT 4.814 30.806 4.866 30.842 ;
               RECT 4.814 32.006 4.866 32.042 ;
               RECT 4.814 33.206 4.866 33.242 ;
               RECT 4.814 34.406 4.866 34.442 ;
               RECT 4.814 35.606 4.866 35.642 ;
               RECT 4.814 36.806 4.866 36.842 ;
               RECT 4.814 38.006 4.866 38.042 ;
               RECT 4.814 39.206 4.866 39.242 ;
               RECT 4.814 40.406 4.866 40.442 ;
               RECT 4.814 41.606 4.866 41.642 ;
               RECT 4.814 42.806 4.866 42.842 ;
               RECT 4.814 44.006 4.866 44.042 ;
               RECT 4.814 45.206 4.866 45.242 ;
               RECT 4.814 46.406 4.866 46.442 ;
               RECT 4.814 47.606 4.866 47.642 ;
               RECT 4.814 49.422 4.866 49.458 ;
               RECT 4.814 49.662 4.866 49.698 ;
               RECT 4.814 55.422 4.866 55.458 ;
               RECT 4.814 55.662 4.866 55.698 ;
               RECT 4.814 56.726 4.866 56.762 ;
               RECT 4.814 57.926 4.866 57.962 ;
               RECT 4.814 59.126 4.866 59.162 ;
               RECT 4.814 60.326 4.866 60.362 ;
               RECT 4.814 61.526 4.866 61.562 ;
               RECT 4.814 62.726 4.866 62.762 ;
               RECT 4.814 63.926 4.866 63.962 ;
               RECT 4.814 65.126 4.866 65.162 ;
               RECT 4.814 66.326 4.866 66.362 ;
               RECT 4.814 67.526 4.866 67.562 ;
               RECT 4.814 68.726 4.866 68.762 ;
               RECT 4.814 69.926 4.866 69.962 ;
               RECT 4.814 71.126 4.866 71.162 ;
               RECT 4.814 72.326 4.866 72.362 ;
               RECT 4.814 73.526 4.866 73.562 ;
               RECT 4.814 74.726 4.866 74.762 ;
               RECT 4.814 75.926 4.866 75.962 ;
               RECT 4.814 77.126 4.866 77.162 ;
               RECT 4.814 78.326 4.866 78.362 ;
               RECT 4.814 79.526 4.866 79.562 ;
               RECT 4.814 80.726 4.866 80.762 ;
               RECT 4.814 81.926 4.866 81.962 ;
               RECT 4.814 83.126 4.866 83.162 ;
               RECT 4.814 84.326 4.866 84.362 ;
               RECT 4.814 85.526 4.866 85.562 ;
               RECT 4.814 86.726 4.866 86.762 ;
               RECT 4.814 87.926 4.866 87.962 ;
               RECT 4.814 89.126 4.866 89.162 ;
               RECT 4.814 90.326 4.866 90.362 ;
               RECT 4.814 91.526 4.866 91.562 ;
               RECT 4.814 92.726 4.866 92.762 ;
               RECT 4.814 93.926 4.866 93.962 ;
               RECT 4.814 95.126 4.866 95.162 ;
               RECT 4.814 96.326 4.866 96.362 ;
               RECT 4.814 97.526 4.866 97.562 ;
               RECT 4.814 98.726 4.866 98.762 ;
               RECT 4.814 99.926 4.866 99.962 ;
               RECT 4.814 101.126 4.866 101.162 ;
               RECT 4.814 102.326 4.866 102.362 ;
               RECT 4.814 103.526 4.866 103.562 ;
               RECT 4.894 1.558 4.946 1.594 ;
               RECT 4.894 2.758 4.946 2.794 ;
               RECT 4.894 3.958 4.946 3.994 ;
               RECT 4.894 5.158 4.946 5.194 ;
               RECT 4.894 6.358 4.946 6.394 ;
               RECT 4.894 7.558 4.946 7.594 ;
               RECT 4.894 8.758 4.946 8.794 ;
               RECT 4.894 9.958 4.946 9.994 ;
               RECT 4.894 11.158 4.946 11.194 ;
               RECT 4.894 12.358 4.946 12.394 ;
               RECT 4.894 13.558 4.946 13.594 ;
               RECT 4.894 14.758 4.946 14.794 ;
               RECT 4.894 15.958 4.946 15.994 ;
               RECT 4.894 17.158 4.946 17.194 ;
               RECT 4.894 18.358 4.946 18.394 ;
               RECT 4.894 19.558 4.946 19.594 ;
               RECT 4.894 20.758 4.946 20.794 ;
               RECT 4.894 21.958 4.946 21.994 ;
               RECT 4.894 23.158 4.946 23.194 ;
               RECT 4.894 24.358 4.946 24.394 ;
               RECT 4.894 25.558 4.946 25.594 ;
               RECT 4.894 26.758 4.946 26.794 ;
               RECT 4.894 27.958 4.946 27.994 ;
               RECT 4.894 29.158 4.946 29.194 ;
               RECT 4.894 30.358 4.946 30.394 ;
               RECT 4.894 31.558 4.946 31.594 ;
               RECT 4.894 32.758 4.946 32.794 ;
               RECT 4.894 33.958 4.946 33.994 ;
               RECT 4.894 35.158 4.946 35.194 ;
               RECT 4.894 36.358 4.946 36.394 ;
               RECT 4.894 37.558 4.946 37.594 ;
               RECT 4.894 38.758 4.946 38.794 ;
               RECT 4.894 39.958 4.946 39.994 ;
               RECT 4.894 41.158 4.946 41.194 ;
               RECT 4.894 42.358 4.946 42.394 ;
               RECT 4.894 43.558 4.946 43.594 ;
               RECT 4.894 44.758 4.946 44.794 ;
               RECT 4.894 45.958 4.946 45.994 ;
               RECT 4.894 47.158 4.946 47.194 ;
               RECT 4.894 48.358 4.946 48.394 ;
               RECT 4.894 50.142 4.946 50.178 ;
               RECT 4.894 50.382 4.946 50.418 ;
               RECT 4.894 54.702 4.946 54.738 ;
               RECT 4.894 54.942 4.946 54.978 ;
               RECT 4.894 57.478 4.946 57.514 ;
               RECT 4.894 58.678 4.946 58.714 ;
               RECT 4.894 59.878 4.946 59.914 ;
               RECT 4.894 61.078 4.946 61.114 ;
               RECT 4.894 62.278 4.946 62.314 ;
               RECT 4.894 63.478 4.946 63.514 ;
               RECT 4.894 64.678 4.946 64.714 ;
               RECT 4.894 65.878 4.946 65.914 ;
               RECT 4.894 67.078 4.946 67.114 ;
               RECT 4.894 68.278 4.946 68.314 ;
               RECT 4.894 69.478 4.946 69.514 ;
               RECT 4.894 70.678 4.946 70.714 ;
               RECT 4.894 71.878 4.946 71.914 ;
               RECT 4.894 73.078 4.946 73.114 ;
               RECT 4.894 74.278 4.946 74.314 ;
               RECT 4.894 75.478 4.946 75.514 ;
               RECT 4.894 76.678 4.946 76.714 ;
               RECT 4.894 77.878 4.946 77.914 ;
               RECT 4.894 79.078 4.946 79.114 ;
               RECT 4.894 80.278 4.946 80.314 ;
               RECT 4.894 81.478 4.946 81.514 ;
               RECT 4.894 82.678 4.946 82.714 ;
               RECT 4.894 83.878 4.946 83.914 ;
               RECT 4.894 85.078 4.946 85.114 ;
               RECT 4.894 86.278 4.946 86.314 ;
               RECT 4.894 87.478 4.946 87.514 ;
               RECT 4.894 88.678 4.946 88.714 ;
               RECT 4.894 89.878 4.946 89.914 ;
               RECT 4.894 91.078 4.946 91.114 ;
               RECT 4.894 92.278 4.946 92.314 ;
               RECT 4.894 93.478 4.946 93.514 ;
               RECT 4.894 94.678 4.946 94.714 ;
               RECT 4.894 95.878 4.946 95.914 ;
               RECT 4.894 97.078 4.946 97.114 ;
               RECT 4.894 98.278 4.946 98.314 ;
               RECT 4.894 99.478 4.946 99.514 ;
               RECT 4.894 100.678 4.946 100.714 ;
               RECT 4.894 101.878 4.946 101.914 ;
               RECT 4.894 103.078 4.946 103.114 ;
               RECT 4.894 104.278 4.946 104.314 ;
               RECT 4.974 0.281 5.026 0.317 ;
               RECT 4.974 104.803 5.026 104.839 ;
               RECT 5.054 0.806 5.106 0.842 ;
               RECT 5.054 2.006 5.106 2.042 ;
               RECT 5.054 3.206 5.106 3.242 ;
               RECT 5.054 4.406 5.106 4.442 ;
               RECT 5.054 5.606 5.106 5.642 ;
               RECT 5.054 6.806 5.106 6.842 ;
               RECT 5.054 8.006 5.106 8.042 ;
               RECT 5.054 9.206 5.106 9.242 ;
               RECT 5.054 10.406 5.106 10.442 ;
               RECT 5.054 11.606 5.106 11.642 ;
               RECT 5.054 12.806 5.106 12.842 ;
               RECT 5.054 14.006 5.106 14.042 ;
               RECT 5.054 15.206 5.106 15.242 ;
               RECT 5.054 16.406 5.106 16.442 ;
               RECT 5.054 17.606 5.106 17.642 ;
               RECT 5.054 18.806 5.106 18.842 ;
               RECT 5.054 20.006 5.106 20.042 ;
               RECT 5.054 21.206 5.106 21.242 ;
               RECT 5.054 22.406 5.106 22.442 ;
               RECT 5.054 23.606 5.106 23.642 ;
               RECT 5.054 24.806 5.106 24.842 ;
               RECT 5.054 26.006 5.106 26.042 ;
               RECT 5.054 27.206 5.106 27.242 ;
               RECT 5.054 28.406 5.106 28.442 ;
               RECT 5.054 29.606 5.106 29.642 ;
               RECT 5.054 30.806 5.106 30.842 ;
               RECT 5.054 32.006 5.106 32.042 ;
               RECT 5.054 33.206 5.106 33.242 ;
               RECT 5.054 34.406 5.106 34.442 ;
               RECT 5.054 35.606 5.106 35.642 ;
               RECT 5.054 36.806 5.106 36.842 ;
               RECT 5.054 38.006 5.106 38.042 ;
               RECT 5.054 39.206 5.106 39.242 ;
               RECT 5.054 40.406 5.106 40.442 ;
               RECT 5.054 41.606 5.106 41.642 ;
               RECT 5.054 42.806 5.106 42.842 ;
               RECT 5.054 44.006 5.106 44.042 ;
               RECT 5.054 45.206 5.106 45.242 ;
               RECT 5.054 46.406 5.106 46.442 ;
               RECT 5.054 47.606 5.106 47.642 ;
               RECT 5.054 49.422 5.106 49.458 ;
               RECT 5.054 49.662 5.106 49.698 ;
               RECT 5.054 51.102 5.106 51.138 ;
               RECT 5.054 51.582 5.106 51.618 ;
               RECT 5.054 53.502 5.106 53.538 ;
               RECT 5.054 53.982 5.106 54.018 ;
               RECT 5.054 55.422 5.106 55.458 ;
               RECT 5.054 55.662 5.106 55.698 ;
               RECT 5.054 56.726 5.106 56.762 ;
               RECT 5.054 57.926 5.106 57.962 ;
               RECT 5.054 59.126 5.106 59.162 ;
               RECT 5.054 60.326 5.106 60.362 ;
               RECT 5.054 61.526 5.106 61.562 ;
               RECT 5.054 62.726 5.106 62.762 ;
               RECT 5.054 63.926 5.106 63.962 ;
               RECT 5.054 65.126 5.106 65.162 ;
               RECT 5.054 66.326 5.106 66.362 ;
               RECT 5.054 67.526 5.106 67.562 ;
               RECT 5.054 68.726 5.106 68.762 ;
               RECT 5.054 69.926 5.106 69.962 ;
               RECT 5.054 71.126 5.106 71.162 ;
               RECT 5.054 72.326 5.106 72.362 ;
               RECT 5.054 73.526 5.106 73.562 ;
               RECT 5.054 74.726 5.106 74.762 ;
               RECT 5.054 75.926 5.106 75.962 ;
               RECT 5.054 77.126 5.106 77.162 ;
               RECT 5.054 78.326 5.106 78.362 ;
               RECT 5.054 79.526 5.106 79.562 ;
               RECT 5.054 80.726 5.106 80.762 ;
               RECT 5.054 81.926 5.106 81.962 ;
               RECT 5.054 83.126 5.106 83.162 ;
               RECT 5.054 84.326 5.106 84.362 ;
               RECT 5.054 85.526 5.106 85.562 ;
               RECT 5.054 86.726 5.106 86.762 ;
               RECT 5.054 87.926 5.106 87.962 ;
               RECT 5.054 89.126 5.106 89.162 ;
               RECT 5.054 90.326 5.106 90.362 ;
               RECT 5.054 91.526 5.106 91.562 ;
               RECT 5.054 92.726 5.106 92.762 ;
               RECT 5.054 93.926 5.106 93.962 ;
               RECT 5.054 95.126 5.106 95.162 ;
               RECT 5.054 96.326 5.106 96.362 ;
               RECT 5.054 97.526 5.106 97.562 ;
               RECT 5.054 98.726 5.106 98.762 ;
               RECT 5.054 99.926 5.106 99.962 ;
               RECT 5.054 101.126 5.106 101.162 ;
               RECT 5.054 102.326 5.106 102.362 ;
               RECT 5.054 103.526 5.106 103.562 ;
               RECT 5.134 1.558 5.186 1.594 ;
               RECT 5.134 2.758 5.186 2.794 ;
               RECT 5.134 3.958 5.186 3.994 ;
               RECT 5.134 5.158 5.186 5.194 ;
               RECT 5.134 6.358 5.186 6.394 ;
               RECT 5.134 7.558 5.186 7.594 ;
               RECT 5.134 8.758 5.186 8.794 ;
               RECT 5.134 9.958 5.186 9.994 ;
               RECT 5.134 11.158 5.186 11.194 ;
               RECT 5.134 12.358 5.186 12.394 ;
               RECT 5.134 13.558 5.186 13.594 ;
               RECT 5.134 14.758 5.186 14.794 ;
               RECT 5.134 15.958 5.186 15.994 ;
               RECT 5.134 17.158 5.186 17.194 ;
               RECT 5.134 18.358 5.186 18.394 ;
               RECT 5.134 19.558 5.186 19.594 ;
               RECT 5.134 20.758 5.186 20.794 ;
               RECT 5.134 21.958 5.186 21.994 ;
               RECT 5.134 23.158 5.186 23.194 ;
               RECT 5.134 24.358 5.186 24.394 ;
               RECT 5.134 25.558 5.186 25.594 ;
               RECT 5.134 26.758 5.186 26.794 ;
               RECT 5.134 27.958 5.186 27.994 ;
               RECT 5.134 29.158 5.186 29.194 ;
               RECT 5.134 30.358 5.186 30.394 ;
               RECT 5.134 31.558 5.186 31.594 ;
               RECT 5.134 32.758 5.186 32.794 ;
               RECT 5.134 33.958 5.186 33.994 ;
               RECT 5.134 35.158 5.186 35.194 ;
               RECT 5.134 36.358 5.186 36.394 ;
               RECT 5.134 37.558 5.186 37.594 ;
               RECT 5.134 38.758 5.186 38.794 ;
               RECT 5.134 39.958 5.186 39.994 ;
               RECT 5.134 41.158 5.186 41.194 ;
               RECT 5.134 42.358 5.186 42.394 ;
               RECT 5.134 43.558 5.186 43.594 ;
               RECT 5.134 44.758 5.186 44.794 ;
               RECT 5.134 45.958 5.186 45.994 ;
               RECT 5.134 47.158 5.186 47.194 ;
               RECT 5.134 48.358 5.186 48.394 ;
               RECT 5.134 50.142 5.186 50.178 ;
               RECT 5.134 50.382 5.186 50.418 ;
               RECT 5.134 54.702 5.186 54.738 ;
               RECT 5.134 54.942 5.186 54.978 ;
               RECT 5.134 57.478 5.186 57.514 ;
               RECT 5.134 58.678 5.186 58.714 ;
               RECT 5.134 59.878 5.186 59.914 ;
               RECT 5.134 61.078 5.186 61.114 ;
               RECT 5.134 62.278 5.186 62.314 ;
               RECT 5.134 63.478 5.186 63.514 ;
               RECT 5.134 64.678 5.186 64.714 ;
               RECT 5.134 65.878 5.186 65.914 ;
               RECT 5.134 67.078 5.186 67.114 ;
               RECT 5.134 68.278 5.186 68.314 ;
               RECT 5.134 69.478 5.186 69.514 ;
               RECT 5.134 70.678 5.186 70.714 ;
               RECT 5.134 71.878 5.186 71.914 ;
               RECT 5.134 73.078 5.186 73.114 ;
               RECT 5.134 74.278 5.186 74.314 ;
               RECT 5.134 75.478 5.186 75.514 ;
               RECT 5.134 76.678 5.186 76.714 ;
               RECT 5.134 77.878 5.186 77.914 ;
               RECT 5.134 79.078 5.186 79.114 ;
               RECT 5.134 80.278 5.186 80.314 ;
               RECT 5.134 81.478 5.186 81.514 ;
               RECT 5.134 82.678 5.186 82.714 ;
               RECT 5.134 83.878 5.186 83.914 ;
               RECT 5.134 85.078 5.186 85.114 ;
               RECT 5.134 86.278 5.186 86.314 ;
               RECT 5.134 87.478 5.186 87.514 ;
               RECT 5.134 88.678 5.186 88.714 ;
               RECT 5.134 89.878 5.186 89.914 ;
               RECT 5.134 91.078 5.186 91.114 ;
               RECT 5.134 92.278 5.186 92.314 ;
               RECT 5.134 93.478 5.186 93.514 ;
               RECT 5.134 94.678 5.186 94.714 ;
               RECT 5.134 95.878 5.186 95.914 ;
               RECT 5.134 97.078 5.186 97.114 ;
               RECT 5.134 98.278 5.186 98.314 ;
               RECT 5.134 99.478 5.186 99.514 ;
               RECT 5.134 100.678 5.186 100.714 ;
               RECT 5.134 101.878 5.186 101.914 ;
               RECT 5.134 103.078 5.186 103.114 ;
               RECT 5.134 104.278 5.186 104.314 ;
               RECT 5.214 0.806 5.266 0.842 ;
               RECT 5.214 2.006 5.266 2.042 ;
               RECT 5.214 3.206 5.266 3.242 ;
               RECT 5.214 4.406 5.266 4.442 ;
               RECT 5.214 5.606 5.266 5.642 ;
               RECT 5.214 6.806 5.266 6.842 ;
               RECT 5.214 8.006 5.266 8.042 ;
               RECT 5.214 9.206 5.266 9.242 ;
               RECT 5.214 10.406 5.266 10.442 ;
               RECT 5.214 11.606 5.266 11.642 ;
               RECT 5.214 12.806 5.266 12.842 ;
               RECT 5.214 14.006 5.266 14.042 ;
               RECT 5.214 15.206 5.266 15.242 ;
               RECT 5.214 16.406 5.266 16.442 ;
               RECT 5.214 17.606 5.266 17.642 ;
               RECT 5.214 18.806 5.266 18.842 ;
               RECT 5.214 20.006 5.266 20.042 ;
               RECT 5.214 21.206 5.266 21.242 ;
               RECT 5.214 22.406 5.266 22.442 ;
               RECT 5.214 23.606 5.266 23.642 ;
               RECT 5.214 24.806 5.266 24.842 ;
               RECT 5.214 26.006 5.266 26.042 ;
               RECT 5.214 27.206 5.266 27.242 ;
               RECT 5.214 28.406 5.266 28.442 ;
               RECT 5.214 29.606 5.266 29.642 ;
               RECT 5.214 30.806 5.266 30.842 ;
               RECT 5.214 32.006 5.266 32.042 ;
               RECT 5.214 33.206 5.266 33.242 ;
               RECT 5.214 34.406 5.266 34.442 ;
               RECT 5.214 35.606 5.266 35.642 ;
               RECT 5.214 36.806 5.266 36.842 ;
               RECT 5.214 38.006 5.266 38.042 ;
               RECT 5.214 39.206 5.266 39.242 ;
               RECT 5.214 40.406 5.266 40.442 ;
               RECT 5.214 41.606 5.266 41.642 ;
               RECT 5.214 42.806 5.266 42.842 ;
               RECT 5.214 44.006 5.266 44.042 ;
               RECT 5.214 45.206 5.266 45.242 ;
               RECT 5.214 46.406 5.266 46.442 ;
               RECT 5.214 47.606 5.266 47.642 ;
               RECT 5.214 49.422 5.266 49.458 ;
               RECT 5.214 49.662 5.266 49.698 ;
               RECT 5.214 55.422 5.266 55.458 ;
               RECT 5.214 55.662 5.266 55.698 ;
               RECT 5.214 56.726 5.266 56.762 ;
               RECT 5.214 57.926 5.266 57.962 ;
               RECT 5.214 59.126 5.266 59.162 ;
               RECT 5.214 60.326 5.266 60.362 ;
               RECT 5.214 61.526 5.266 61.562 ;
               RECT 5.214 62.726 5.266 62.762 ;
               RECT 5.214 63.926 5.266 63.962 ;
               RECT 5.214 65.126 5.266 65.162 ;
               RECT 5.214 66.326 5.266 66.362 ;
               RECT 5.214 67.526 5.266 67.562 ;
               RECT 5.214 68.726 5.266 68.762 ;
               RECT 5.214 69.926 5.266 69.962 ;
               RECT 5.214 71.126 5.266 71.162 ;
               RECT 5.214 72.326 5.266 72.362 ;
               RECT 5.214 73.526 5.266 73.562 ;
               RECT 5.214 74.726 5.266 74.762 ;
               RECT 5.214 75.926 5.266 75.962 ;
               RECT 5.214 77.126 5.266 77.162 ;
               RECT 5.214 78.326 5.266 78.362 ;
               RECT 5.214 79.526 5.266 79.562 ;
               RECT 5.214 80.726 5.266 80.762 ;
               RECT 5.214 81.926 5.266 81.962 ;
               RECT 5.214 83.126 5.266 83.162 ;
               RECT 5.214 84.326 5.266 84.362 ;
               RECT 5.214 85.526 5.266 85.562 ;
               RECT 5.214 86.726 5.266 86.762 ;
               RECT 5.214 87.926 5.266 87.962 ;
               RECT 5.214 89.126 5.266 89.162 ;
               RECT 5.214 90.326 5.266 90.362 ;
               RECT 5.214 91.526 5.266 91.562 ;
               RECT 5.214 92.726 5.266 92.762 ;
               RECT 5.214 93.926 5.266 93.962 ;
               RECT 5.214 95.126 5.266 95.162 ;
               RECT 5.214 96.326 5.266 96.362 ;
               RECT 5.214 97.526 5.266 97.562 ;
               RECT 5.214 98.726 5.266 98.762 ;
               RECT 5.214 99.926 5.266 99.962 ;
               RECT 5.214 101.126 5.266 101.162 ;
               RECT 5.214 102.326 5.266 102.362 ;
               RECT 5.214 103.526 5.266 103.562 ;
               RECT 5.294 1.558 5.346 1.594 ;
               RECT 5.294 2.758 5.346 2.794 ;
               RECT 5.294 3.958 5.346 3.994 ;
               RECT 5.294 5.158 5.346 5.194 ;
               RECT 5.294 6.358 5.346 6.394 ;
               RECT 5.294 7.558 5.346 7.594 ;
               RECT 5.294 8.758 5.346 8.794 ;
               RECT 5.294 9.958 5.346 9.994 ;
               RECT 5.294 11.158 5.346 11.194 ;
               RECT 5.294 12.358 5.346 12.394 ;
               RECT 5.294 13.558 5.346 13.594 ;
               RECT 5.294 14.758 5.346 14.794 ;
               RECT 5.294 15.958 5.346 15.994 ;
               RECT 5.294 17.158 5.346 17.194 ;
               RECT 5.294 18.358 5.346 18.394 ;
               RECT 5.294 19.558 5.346 19.594 ;
               RECT 5.294 20.758 5.346 20.794 ;
               RECT 5.294 21.958 5.346 21.994 ;
               RECT 5.294 23.158 5.346 23.194 ;
               RECT 5.294 24.358 5.346 24.394 ;
               RECT 5.294 25.558 5.346 25.594 ;
               RECT 5.294 26.758 5.346 26.794 ;
               RECT 5.294 27.958 5.346 27.994 ;
               RECT 5.294 29.158 5.346 29.194 ;
               RECT 5.294 30.358 5.346 30.394 ;
               RECT 5.294 31.558 5.346 31.594 ;
               RECT 5.294 32.758 5.346 32.794 ;
               RECT 5.294 33.958 5.346 33.994 ;
               RECT 5.294 35.158 5.346 35.194 ;
               RECT 5.294 36.358 5.346 36.394 ;
               RECT 5.294 37.558 5.346 37.594 ;
               RECT 5.294 38.758 5.346 38.794 ;
               RECT 5.294 39.958 5.346 39.994 ;
               RECT 5.294 41.158 5.346 41.194 ;
               RECT 5.294 42.358 5.346 42.394 ;
               RECT 5.294 43.558 5.346 43.594 ;
               RECT 5.294 44.758 5.346 44.794 ;
               RECT 5.294 45.958 5.346 45.994 ;
               RECT 5.294 47.158 5.346 47.194 ;
               RECT 5.294 48.358 5.346 48.394 ;
               RECT 5.294 50.142 5.346 50.178 ;
               RECT 5.294 50.382 5.346 50.418 ;
               RECT 5.294 54.702 5.346 54.738 ;
               RECT 5.294 54.942 5.346 54.978 ;
               RECT 5.294 57.478 5.346 57.514 ;
               RECT 5.294 58.678 5.346 58.714 ;
               RECT 5.294 59.878 5.346 59.914 ;
               RECT 5.294 61.078 5.346 61.114 ;
               RECT 5.294 62.278 5.346 62.314 ;
               RECT 5.294 63.478 5.346 63.514 ;
               RECT 5.294 64.678 5.346 64.714 ;
               RECT 5.294 65.878 5.346 65.914 ;
               RECT 5.294 67.078 5.346 67.114 ;
               RECT 5.294 68.278 5.346 68.314 ;
               RECT 5.294 69.478 5.346 69.514 ;
               RECT 5.294 70.678 5.346 70.714 ;
               RECT 5.294 71.878 5.346 71.914 ;
               RECT 5.294 73.078 5.346 73.114 ;
               RECT 5.294 74.278 5.346 74.314 ;
               RECT 5.294 75.478 5.346 75.514 ;
               RECT 5.294 76.678 5.346 76.714 ;
               RECT 5.294 77.878 5.346 77.914 ;
               RECT 5.294 79.078 5.346 79.114 ;
               RECT 5.294 80.278 5.346 80.314 ;
               RECT 5.294 81.478 5.346 81.514 ;
               RECT 5.294 82.678 5.346 82.714 ;
               RECT 5.294 83.878 5.346 83.914 ;
               RECT 5.294 85.078 5.346 85.114 ;
               RECT 5.294 86.278 5.346 86.314 ;
               RECT 5.294 87.478 5.346 87.514 ;
               RECT 5.294 88.678 5.346 88.714 ;
               RECT 5.294 89.878 5.346 89.914 ;
               RECT 5.294 91.078 5.346 91.114 ;
               RECT 5.294 92.278 5.346 92.314 ;
               RECT 5.294 93.478 5.346 93.514 ;
               RECT 5.294 94.678 5.346 94.714 ;
               RECT 5.294 95.878 5.346 95.914 ;
               RECT 5.294 97.078 5.346 97.114 ;
               RECT 5.294 98.278 5.346 98.314 ;
               RECT 5.294 99.478 5.346 99.514 ;
               RECT 5.294 100.678 5.346 100.714 ;
               RECT 5.294 101.878 5.346 101.914 ;
               RECT 5.294 103.078 5.346 103.114 ;
               RECT 5.294 104.278 5.346 104.314 ;
               RECT 5.374 0.281 5.426 0.317 ;
               RECT 5.374 104.803 5.426 104.839 ;
               RECT 5.454 0.806 5.506 0.842 ;
               RECT 5.454 2.006 5.506 2.042 ;
               RECT 5.454 3.206 5.506 3.242 ;
               RECT 5.454 4.406 5.506 4.442 ;
               RECT 5.454 5.606 5.506 5.642 ;
               RECT 5.454 6.806 5.506 6.842 ;
               RECT 5.454 8.006 5.506 8.042 ;
               RECT 5.454 9.206 5.506 9.242 ;
               RECT 5.454 10.406 5.506 10.442 ;
               RECT 5.454 11.606 5.506 11.642 ;
               RECT 5.454 12.806 5.506 12.842 ;
               RECT 5.454 14.006 5.506 14.042 ;
               RECT 5.454 15.206 5.506 15.242 ;
               RECT 5.454 16.406 5.506 16.442 ;
               RECT 5.454 17.606 5.506 17.642 ;
               RECT 5.454 18.806 5.506 18.842 ;
               RECT 5.454 20.006 5.506 20.042 ;
               RECT 5.454 21.206 5.506 21.242 ;
               RECT 5.454 22.406 5.506 22.442 ;
               RECT 5.454 23.606 5.506 23.642 ;
               RECT 5.454 24.806 5.506 24.842 ;
               RECT 5.454 26.006 5.506 26.042 ;
               RECT 5.454 27.206 5.506 27.242 ;
               RECT 5.454 28.406 5.506 28.442 ;
               RECT 5.454 29.606 5.506 29.642 ;
               RECT 5.454 30.806 5.506 30.842 ;
               RECT 5.454 32.006 5.506 32.042 ;
               RECT 5.454 33.206 5.506 33.242 ;
               RECT 5.454 34.406 5.506 34.442 ;
               RECT 5.454 35.606 5.506 35.642 ;
               RECT 5.454 36.806 5.506 36.842 ;
               RECT 5.454 38.006 5.506 38.042 ;
               RECT 5.454 39.206 5.506 39.242 ;
               RECT 5.454 40.406 5.506 40.442 ;
               RECT 5.454 41.606 5.506 41.642 ;
               RECT 5.454 42.806 5.506 42.842 ;
               RECT 5.454 44.006 5.506 44.042 ;
               RECT 5.454 45.206 5.506 45.242 ;
               RECT 5.454 46.406 5.506 46.442 ;
               RECT 5.454 47.606 5.506 47.642 ;
               RECT 5.454 49.422 5.506 49.458 ;
               RECT 5.454 49.662 5.506 49.698 ;
               RECT 5.454 55.422 5.506 55.458 ;
               RECT 5.454 55.662 5.506 55.698 ;
               RECT 5.454 56.726 5.506 56.762 ;
               RECT 5.454 57.926 5.506 57.962 ;
               RECT 5.454 59.126 5.506 59.162 ;
               RECT 5.454 60.326 5.506 60.362 ;
               RECT 5.454 61.526 5.506 61.562 ;
               RECT 5.454 62.726 5.506 62.762 ;
               RECT 5.454 63.926 5.506 63.962 ;
               RECT 5.454 65.126 5.506 65.162 ;
               RECT 5.454 66.326 5.506 66.362 ;
               RECT 5.454 67.526 5.506 67.562 ;
               RECT 5.454 68.726 5.506 68.762 ;
               RECT 5.454 69.926 5.506 69.962 ;
               RECT 5.454 71.126 5.506 71.162 ;
               RECT 5.454 72.326 5.506 72.362 ;
               RECT 5.454 73.526 5.506 73.562 ;
               RECT 5.454 74.726 5.506 74.762 ;
               RECT 5.454 75.926 5.506 75.962 ;
               RECT 5.454 77.126 5.506 77.162 ;
               RECT 5.454 78.326 5.506 78.362 ;
               RECT 5.454 79.526 5.506 79.562 ;
               RECT 5.454 80.726 5.506 80.762 ;
               RECT 5.454 81.926 5.506 81.962 ;
               RECT 5.454 83.126 5.506 83.162 ;
               RECT 5.454 84.326 5.506 84.362 ;
               RECT 5.454 85.526 5.506 85.562 ;
               RECT 5.454 86.726 5.506 86.762 ;
               RECT 5.454 87.926 5.506 87.962 ;
               RECT 5.454 89.126 5.506 89.162 ;
               RECT 5.454 90.326 5.506 90.362 ;
               RECT 5.454 91.526 5.506 91.562 ;
               RECT 5.454 92.726 5.506 92.762 ;
               RECT 5.454 93.926 5.506 93.962 ;
               RECT 5.454 95.126 5.506 95.162 ;
               RECT 5.454 96.326 5.506 96.362 ;
               RECT 5.454 97.526 5.506 97.562 ;
               RECT 5.454 98.726 5.506 98.762 ;
               RECT 5.454 99.926 5.506 99.962 ;
               RECT 5.454 101.126 5.506 101.162 ;
               RECT 5.454 102.326 5.506 102.362 ;
               RECT 5.454 103.526 5.506 103.562 ;
               RECT 5.534 1.558 5.586 1.594 ;
               RECT 5.534 2.758 5.586 2.794 ;
               RECT 5.534 3.958 5.586 3.994 ;
               RECT 5.534 5.158 5.586 5.194 ;
               RECT 5.534 6.358 5.586 6.394 ;
               RECT 5.534 7.558 5.586 7.594 ;
               RECT 5.534 8.758 5.586 8.794 ;
               RECT 5.534 9.958 5.586 9.994 ;
               RECT 5.534 11.158 5.586 11.194 ;
               RECT 5.534 12.358 5.586 12.394 ;
               RECT 5.534 13.558 5.586 13.594 ;
               RECT 5.534 14.758 5.586 14.794 ;
               RECT 5.534 15.958 5.586 15.994 ;
               RECT 5.534 17.158 5.586 17.194 ;
               RECT 5.534 18.358 5.586 18.394 ;
               RECT 5.534 19.558 5.586 19.594 ;
               RECT 5.534 20.758 5.586 20.794 ;
               RECT 5.534 21.958 5.586 21.994 ;
               RECT 5.534 23.158 5.586 23.194 ;
               RECT 5.534 24.358 5.586 24.394 ;
               RECT 5.534 25.558 5.586 25.594 ;
               RECT 5.534 26.758 5.586 26.794 ;
               RECT 5.534 27.958 5.586 27.994 ;
               RECT 5.534 29.158 5.586 29.194 ;
               RECT 5.534 30.358 5.586 30.394 ;
               RECT 5.534 31.558 5.586 31.594 ;
               RECT 5.534 32.758 5.586 32.794 ;
               RECT 5.534 33.958 5.586 33.994 ;
               RECT 5.534 35.158 5.586 35.194 ;
               RECT 5.534 36.358 5.586 36.394 ;
               RECT 5.534 37.558 5.586 37.594 ;
               RECT 5.534 38.758 5.586 38.794 ;
               RECT 5.534 39.958 5.586 39.994 ;
               RECT 5.534 41.158 5.586 41.194 ;
               RECT 5.534 42.358 5.586 42.394 ;
               RECT 5.534 43.558 5.586 43.594 ;
               RECT 5.534 44.758 5.586 44.794 ;
               RECT 5.534 45.958 5.586 45.994 ;
               RECT 5.534 47.158 5.586 47.194 ;
               RECT 5.534 48.358 5.586 48.394 ;
               RECT 5.534 50.142 5.586 50.178 ;
               RECT 5.534 50.382 5.586 50.418 ;
               RECT 5.534 54.702 5.586 54.738 ;
               RECT 5.534 54.942 5.586 54.978 ;
               RECT 5.534 57.478 5.586 57.514 ;
               RECT 5.534 58.678 5.586 58.714 ;
               RECT 5.534 59.878 5.586 59.914 ;
               RECT 5.534 61.078 5.586 61.114 ;
               RECT 5.534 62.278 5.586 62.314 ;
               RECT 5.534 63.478 5.586 63.514 ;
               RECT 5.534 64.678 5.586 64.714 ;
               RECT 5.534 65.878 5.586 65.914 ;
               RECT 5.534 67.078 5.586 67.114 ;
               RECT 5.534 68.278 5.586 68.314 ;
               RECT 5.534 69.478 5.586 69.514 ;
               RECT 5.534 70.678 5.586 70.714 ;
               RECT 5.534 71.878 5.586 71.914 ;
               RECT 5.534 73.078 5.586 73.114 ;
               RECT 5.534 74.278 5.586 74.314 ;
               RECT 5.534 75.478 5.586 75.514 ;
               RECT 5.534 76.678 5.586 76.714 ;
               RECT 5.534 77.878 5.586 77.914 ;
               RECT 5.534 79.078 5.586 79.114 ;
               RECT 5.534 80.278 5.586 80.314 ;
               RECT 5.534 81.478 5.586 81.514 ;
               RECT 5.534 82.678 5.586 82.714 ;
               RECT 5.534 83.878 5.586 83.914 ;
               RECT 5.534 85.078 5.586 85.114 ;
               RECT 5.534 86.278 5.586 86.314 ;
               RECT 5.534 87.478 5.586 87.514 ;
               RECT 5.534 88.678 5.586 88.714 ;
               RECT 5.534 89.878 5.586 89.914 ;
               RECT 5.534 91.078 5.586 91.114 ;
               RECT 5.534 92.278 5.586 92.314 ;
               RECT 5.534 93.478 5.586 93.514 ;
               RECT 5.534 94.678 5.586 94.714 ;
               RECT 5.534 95.878 5.586 95.914 ;
               RECT 5.534 97.078 5.586 97.114 ;
               RECT 5.534 98.278 5.586 98.314 ;
               RECT 5.534 99.478 5.586 99.514 ;
               RECT 5.534 100.678 5.586 100.714 ;
               RECT 5.534 101.878 5.586 101.914 ;
               RECT 5.534 103.078 5.586 103.114 ;
               RECT 5.534 104.278 5.586 104.314 ;
               RECT 5.614 0.806 5.666 0.842 ;
               RECT 5.614 2.006 5.666 2.042 ;
               RECT 5.614 3.206 5.666 3.242 ;
               RECT 5.614 4.406 5.666 4.442 ;
               RECT 5.614 5.606 5.666 5.642 ;
               RECT 5.614 6.806 5.666 6.842 ;
               RECT 5.614 8.006 5.666 8.042 ;
               RECT 5.614 9.206 5.666 9.242 ;
               RECT 5.614 10.406 5.666 10.442 ;
               RECT 5.614 11.606 5.666 11.642 ;
               RECT 5.614 12.806 5.666 12.842 ;
               RECT 5.614 14.006 5.666 14.042 ;
               RECT 5.614 15.206 5.666 15.242 ;
               RECT 5.614 16.406 5.666 16.442 ;
               RECT 5.614 17.606 5.666 17.642 ;
               RECT 5.614 18.806 5.666 18.842 ;
               RECT 5.614 20.006 5.666 20.042 ;
               RECT 5.614 21.206 5.666 21.242 ;
               RECT 5.614 22.406 5.666 22.442 ;
               RECT 5.614 23.606 5.666 23.642 ;
               RECT 5.614 24.806 5.666 24.842 ;
               RECT 5.614 26.006 5.666 26.042 ;
               RECT 5.614 27.206 5.666 27.242 ;
               RECT 5.614 28.406 5.666 28.442 ;
               RECT 5.614 29.606 5.666 29.642 ;
               RECT 5.614 30.806 5.666 30.842 ;
               RECT 5.614 32.006 5.666 32.042 ;
               RECT 5.614 33.206 5.666 33.242 ;
               RECT 5.614 34.406 5.666 34.442 ;
               RECT 5.614 35.606 5.666 35.642 ;
               RECT 5.614 36.806 5.666 36.842 ;
               RECT 5.614 38.006 5.666 38.042 ;
               RECT 5.614 39.206 5.666 39.242 ;
               RECT 5.614 40.406 5.666 40.442 ;
               RECT 5.614 41.606 5.666 41.642 ;
               RECT 5.614 42.806 5.666 42.842 ;
               RECT 5.614 44.006 5.666 44.042 ;
               RECT 5.614 45.206 5.666 45.242 ;
               RECT 5.614 46.406 5.666 46.442 ;
               RECT 5.614 47.606 5.666 47.642 ;
               RECT 5.614 49.422 5.666 49.458 ;
               RECT 5.614 49.662 5.666 49.698 ;
               RECT 5.614 55.422 5.666 55.458 ;
               RECT 5.614 55.662 5.666 55.698 ;
               RECT 5.614 56.726 5.666 56.762 ;
               RECT 5.614 57.926 5.666 57.962 ;
               RECT 5.614 59.126 5.666 59.162 ;
               RECT 5.614 60.326 5.666 60.362 ;
               RECT 5.614 61.526 5.666 61.562 ;
               RECT 5.614 62.726 5.666 62.762 ;
               RECT 5.614 63.926 5.666 63.962 ;
               RECT 5.614 65.126 5.666 65.162 ;
               RECT 5.614 66.326 5.666 66.362 ;
               RECT 5.614 67.526 5.666 67.562 ;
               RECT 5.614 68.726 5.666 68.762 ;
               RECT 5.614 69.926 5.666 69.962 ;
               RECT 5.614 71.126 5.666 71.162 ;
               RECT 5.614 72.326 5.666 72.362 ;
               RECT 5.614 73.526 5.666 73.562 ;
               RECT 5.614 74.726 5.666 74.762 ;
               RECT 5.614 75.926 5.666 75.962 ;
               RECT 5.614 77.126 5.666 77.162 ;
               RECT 5.614 78.326 5.666 78.362 ;
               RECT 5.614 79.526 5.666 79.562 ;
               RECT 5.614 80.726 5.666 80.762 ;
               RECT 5.614 81.926 5.666 81.962 ;
               RECT 5.614 83.126 5.666 83.162 ;
               RECT 5.614 84.326 5.666 84.362 ;
               RECT 5.614 85.526 5.666 85.562 ;
               RECT 5.614 86.726 5.666 86.762 ;
               RECT 5.614 87.926 5.666 87.962 ;
               RECT 5.614 89.126 5.666 89.162 ;
               RECT 5.614 90.326 5.666 90.362 ;
               RECT 5.614 91.526 5.666 91.562 ;
               RECT 5.614 92.726 5.666 92.762 ;
               RECT 5.614 93.926 5.666 93.962 ;
               RECT 5.614 95.126 5.666 95.162 ;
               RECT 5.614 96.326 5.666 96.362 ;
               RECT 5.614 97.526 5.666 97.562 ;
               RECT 5.614 98.726 5.666 98.762 ;
               RECT 5.614 99.926 5.666 99.962 ;
               RECT 5.614 101.126 5.666 101.162 ;
               RECT 5.614 102.326 5.666 102.362 ;
               RECT 5.614 103.526 5.666 103.562 ;
               RECT 5.694 1.558 5.746 1.594 ;
               RECT 5.694 2.758 5.746 2.794 ;
               RECT 5.694 3.958 5.746 3.994 ;
               RECT 5.694 5.158 5.746 5.194 ;
               RECT 5.694 6.358 5.746 6.394 ;
               RECT 5.694 7.558 5.746 7.594 ;
               RECT 5.694 8.758 5.746 8.794 ;
               RECT 5.694 9.958 5.746 9.994 ;
               RECT 5.694 11.158 5.746 11.194 ;
               RECT 5.694 12.358 5.746 12.394 ;
               RECT 5.694 13.558 5.746 13.594 ;
               RECT 5.694 14.758 5.746 14.794 ;
               RECT 5.694 15.958 5.746 15.994 ;
               RECT 5.694 17.158 5.746 17.194 ;
               RECT 5.694 18.358 5.746 18.394 ;
               RECT 5.694 19.558 5.746 19.594 ;
               RECT 5.694 20.758 5.746 20.794 ;
               RECT 5.694 21.958 5.746 21.994 ;
               RECT 5.694 23.158 5.746 23.194 ;
               RECT 5.694 24.358 5.746 24.394 ;
               RECT 5.694 25.558 5.746 25.594 ;
               RECT 5.694 26.758 5.746 26.794 ;
               RECT 5.694 27.958 5.746 27.994 ;
               RECT 5.694 29.158 5.746 29.194 ;
               RECT 5.694 30.358 5.746 30.394 ;
               RECT 5.694 31.558 5.746 31.594 ;
               RECT 5.694 32.758 5.746 32.794 ;
               RECT 5.694 33.958 5.746 33.994 ;
               RECT 5.694 35.158 5.746 35.194 ;
               RECT 5.694 36.358 5.746 36.394 ;
               RECT 5.694 37.558 5.746 37.594 ;
               RECT 5.694 38.758 5.746 38.794 ;
               RECT 5.694 39.958 5.746 39.994 ;
               RECT 5.694 41.158 5.746 41.194 ;
               RECT 5.694 42.358 5.746 42.394 ;
               RECT 5.694 43.558 5.746 43.594 ;
               RECT 5.694 44.758 5.746 44.794 ;
               RECT 5.694 45.958 5.746 45.994 ;
               RECT 5.694 47.158 5.746 47.194 ;
               RECT 5.694 48.358 5.746 48.394 ;
               RECT 5.694 50.142 5.746 50.178 ;
               RECT 5.694 50.382 5.746 50.418 ;
               RECT 5.694 54.702 5.746 54.738 ;
               RECT 5.694 54.942 5.746 54.978 ;
               RECT 5.694 57.478 5.746 57.514 ;
               RECT 5.694 58.678 5.746 58.714 ;
               RECT 5.694 59.878 5.746 59.914 ;
               RECT 5.694 61.078 5.746 61.114 ;
               RECT 5.694 62.278 5.746 62.314 ;
               RECT 5.694 63.478 5.746 63.514 ;
               RECT 5.694 64.678 5.746 64.714 ;
               RECT 5.694 65.878 5.746 65.914 ;
               RECT 5.694 67.078 5.746 67.114 ;
               RECT 5.694 68.278 5.746 68.314 ;
               RECT 5.694 69.478 5.746 69.514 ;
               RECT 5.694 70.678 5.746 70.714 ;
               RECT 5.694 71.878 5.746 71.914 ;
               RECT 5.694 73.078 5.746 73.114 ;
               RECT 5.694 74.278 5.746 74.314 ;
               RECT 5.694 75.478 5.746 75.514 ;
               RECT 5.694 76.678 5.746 76.714 ;
               RECT 5.694 77.878 5.746 77.914 ;
               RECT 5.694 79.078 5.746 79.114 ;
               RECT 5.694 80.278 5.746 80.314 ;
               RECT 5.694 81.478 5.746 81.514 ;
               RECT 5.694 82.678 5.746 82.714 ;
               RECT 5.694 83.878 5.746 83.914 ;
               RECT 5.694 85.078 5.746 85.114 ;
               RECT 5.694 86.278 5.746 86.314 ;
               RECT 5.694 87.478 5.746 87.514 ;
               RECT 5.694 88.678 5.746 88.714 ;
               RECT 5.694 89.878 5.746 89.914 ;
               RECT 5.694 91.078 5.746 91.114 ;
               RECT 5.694 92.278 5.746 92.314 ;
               RECT 5.694 93.478 5.746 93.514 ;
               RECT 5.694 94.678 5.746 94.714 ;
               RECT 5.694 95.878 5.746 95.914 ;
               RECT 5.694 97.078 5.746 97.114 ;
               RECT 5.694 98.278 5.746 98.314 ;
               RECT 5.694 99.478 5.746 99.514 ;
               RECT 5.694 100.678 5.746 100.714 ;
               RECT 5.694 101.878 5.746 101.914 ;
               RECT 5.694 103.078 5.746 103.114 ;
               RECT 5.694 104.278 5.746 104.314 ;
               RECT 5.774 0.281 5.826 0.317 ;
               RECT 5.774 104.803 5.826 104.839 ;
               RECT 5.854 0.806 5.906 0.842 ;
               RECT 5.854 2.006 5.906 2.042 ;
               RECT 5.854 3.206 5.906 3.242 ;
               RECT 5.854 4.406 5.906 4.442 ;
               RECT 5.854 5.606 5.906 5.642 ;
               RECT 5.854 6.806 5.906 6.842 ;
               RECT 5.854 8.006 5.906 8.042 ;
               RECT 5.854 9.206 5.906 9.242 ;
               RECT 5.854 10.406 5.906 10.442 ;
               RECT 5.854 11.606 5.906 11.642 ;
               RECT 5.854 12.806 5.906 12.842 ;
               RECT 5.854 14.006 5.906 14.042 ;
               RECT 5.854 15.206 5.906 15.242 ;
               RECT 5.854 16.406 5.906 16.442 ;
               RECT 5.854 17.606 5.906 17.642 ;
               RECT 5.854 18.806 5.906 18.842 ;
               RECT 5.854 20.006 5.906 20.042 ;
               RECT 5.854 21.206 5.906 21.242 ;
               RECT 5.854 22.406 5.906 22.442 ;
               RECT 5.854 23.606 5.906 23.642 ;
               RECT 5.854 24.806 5.906 24.842 ;
               RECT 5.854 26.006 5.906 26.042 ;
               RECT 5.854 27.206 5.906 27.242 ;
               RECT 5.854 28.406 5.906 28.442 ;
               RECT 5.854 29.606 5.906 29.642 ;
               RECT 5.854 30.806 5.906 30.842 ;
               RECT 5.854 32.006 5.906 32.042 ;
               RECT 5.854 33.206 5.906 33.242 ;
               RECT 5.854 34.406 5.906 34.442 ;
               RECT 5.854 35.606 5.906 35.642 ;
               RECT 5.854 36.806 5.906 36.842 ;
               RECT 5.854 38.006 5.906 38.042 ;
               RECT 5.854 39.206 5.906 39.242 ;
               RECT 5.854 40.406 5.906 40.442 ;
               RECT 5.854 41.606 5.906 41.642 ;
               RECT 5.854 42.806 5.906 42.842 ;
               RECT 5.854 44.006 5.906 44.042 ;
               RECT 5.854 45.206 5.906 45.242 ;
               RECT 5.854 46.406 5.906 46.442 ;
               RECT 5.854 47.606 5.906 47.642 ;
               RECT 5.854 49.422 5.906 49.458 ;
               RECT 5.854 49.662 5.906 49.698 ;
               RECT 5.854 51.102 5.906 51.138 ;
               RECT 5.854 51.582 5.906 51.618 ;
               RECT 5.854 53.502 5.906 53.538 ;
               RECT 5.854 53.982 5.906 54.018 ;
               RECT 5.854 55.422 5.906 55.458 ;
               RECT 5.854 55.662 5.906 55.698 ;
               RECT 5.854 56.726 5.906 56.762 ;
               RECT 5.854 57.926 5.906 57.962 ;
               RECT 5.854 59.126 5.906 59.162 ;
               RECT 5.854 60.326 5.906 60.362 ;
               RECT 5.854 61.526 5.906 61.562 ;
               RECT 5.854 62.726 5.906 62.762 ;
               RECT 5.854 63.926 5.906 63.962 ;
               RECT 5.854 65.126 5.906 65.162 ;
               RECT 5.854 66.326 5.906 66.362 ;
               RECT 5.854 67.526 5.906 67.562 ;
               RECT 5.854 68.726 5.906 68.762 ;
               RECT 5.854 69.926 5.906 69.962 ;
               RECT 5.854 71.126 5.906 71.162 ;
               RECT 5.854 72.326 5.906 72.362 ;
               RECT 5.854 73.526 5.906 73.562 ;
               RECT 5.854 74.726 5.906 74.762 ;
               RECT 5.854 75.926 5.906 75.962 ;
               RECT 5.854 77.126 5.906 77.162 ;
               RECT 5.854 78.326 5.906 78.362 ;
               RECT 5.854 79.526 5.906 79.562 ;
               RECT 5.854 80.726 5.906 80.762 ;
               RECT 5.854 81.926 5.906 81.962 ;
               RECT 5.854 83.126 5.906 83.162 ;
               RECT 5.854 84.326 5.906 84.362 ;
               RECT 5.854 85.526 5.906 85.562 ;
               RECT 5.854 86.726 5.906 86.762 ;
               RECT 5.854 87.926 5.906 87.962 ;
               RECT 5.854 89.126 5.906 89.162 ;
               RECT 5.854 90.326 5.906 90.362 ;
               RECT 5.854 91.526 5.906 91.562 ;
               RECT 5.854 92.726 5.906 92.762 ;
               RECT 5.854 93.926 5.906 93.962 ;
               RECT 5.854 95.126 5.906 95.162 ;
               RECT 5.854 96.326 5.906 96.362 ;
               RECT 5.854 97.526 5.906 97.562 ;
               RECT 5.854 98.726 5.906 98.762 ;
               RECT 5.854 99.926 5.906 99.962 ;
               RECT 5.854 101.126 5.906 101.162 ;
               RECT 5.854 102.326 5.906 102.362 ;
               RECT 5.854 103.526 5.906 103.562 ;
               RECT 5.934 1.558 5.986 1.594 ;
               RECT 5.934 2.758 5.986 2.794 ;
               RECT 5.934 3.958 5.986 3.994 ;
               RECT 5.934 5.158 5.986 5.194 ;
               RECT 5.934 6.358 5.986 6.394 ;
               RECT 5.934 7.558 5.986 7.594 ;
               RECT 5.934 8.758 5.986 8.794 ;
               RECT 5.934 9.958 5.986 9.994 ;
               RECT 5.934 11.158 5.986 11.194 ;
               RECT 5.934 12.358 5.986 12.394 ;
               RECT 5.934 13.558 5.986 13.594 ;
               RECT 5.934 14.758 5.986 14.794 ;
               RECT 5.934 15.958 5.986 15.994 ;
               RECT 5.934 17.158 5.986 17.194 ;
               RECT 5.934 18.358 5.986 18.394 ;
               RECT 5.934 19.558 5.986 19.594 ;
               RECT 5.934 20.758 5.986 20.794 ;
               RECT 5.934 21.958 5.986 21.994 ;
               RECT 5.934 23.158 5.986 23.194 ;
               RECT 5.934 24.358 5.986 24.394 ;
               RECT 5.934 25.558 5.986 25.594 ;
               RECT 5.934 26.758 5.986 26.794 ;
               RECT 5.934 27.958 5.986 27.994 ;
               RECT 5.934 29.158 5.986 29.194 ;
               RECT 5.934 30.358 5.986 30.394 ;
               RECT 5.934 31.558 5.986 31.594 ;
               RECT 5.934 32.758 5.986 32.794 ;
               RECT 5.934 33.958 5.986 33.994 ;
               RECT 5.934 35.158 5.986 35.194 ;
               RECT 5.934 36.358 5.986 36.394 ;
               RECT 5.934 37.558 5.986 37.594 ;
               RECT 5.934 38.758 5.986 38.794 ;
               RECT 5.934 39.958 5.986 39.994 ;
               RECT 5.934 41.158 5.986 41.194 ;
               RECT 5.934 42.358 5.986 42.394 ;
               RECT 5.934 43.558 5.986 43.594 ;
               RECT 5.934 44.758 5.986 44.794 ;
               RECT 5.934 45.958 5.986 45.994 ;
               RECT 5.934 47.158 5.986 47.194 ;
               RECT 5.934 48.358 5.986 48.394 ;
               RECT 5.934 50.142 5.986 50.178 ;
               RECT 5.934 50.382 5.986 50.418 ;
               RECT 5.934 54.702 5.986 54.738 ;
               RECT 5.934 54.942 5.986 54.978 ;
               RECT 5.934 57.478 5.986 57.514 ;
               RECT 5.934 58.678 5.986 58.714 ;
               RECT 5.934 59.878 5.986 59.914 ;
               RECT 5.934 61.078 5.986 61.114 ;
               RECT 5.934 62.278 5.986 62.314 ;
               RECT 5.934 63.478 5.986 63.514 ;
               RECT 5.934 64.678 5.986 64.714 ;
               RECT 5.934 65.878 5.986 65.914 ;
               RECT 5.934 67.078 5.986 67.114 ;
               RECT 5.934 68.278 5.986 68.314 ;
               RECT 5.934 69.478 5.986 69.514 ;
               RECT 5.934 70.678 5.986 70.714 ;
               RECT 5.934 71.878 5.986 71.914 ;
               RECT 5.934 73.078 5.986 73.114 ;
               RECT 5.934 74.278 5.986 74.314 ;
               RECT 5.934 75.478 5.986 75.514 ;
               RECT 5.934 76.678 5.986 76.714 ;
               RECT 5.934 77.878 5.986 77.914 ;
               RECT 5.934 79.078 5.986 79.114 ;
               RECT 5.934 80.278 5.986 80.314 ;
               RECT 5.934 81.478 5.986 81.514 ;
               RECT 5.934 82.678 5.986 82.714 ;
               RECT 5.934 83.878 5.986 83.914 ;
               RECT 5.934 85.078 5.986 85.114 ;
               RECT 5.934 86.278 5.986 86.314 ;
               RECT 5.934 87.478 5.986 87.514 ;
               RECT 5.934 88.678 5.986 88.714 ;
               RECT 5.934 89.878 5.986 89.914 ;
               RECT 5.934 91.078 5.986 91.114 ;
               RECT 5.934 92.278 5.986 92.314 ;
               RECT 5.934 93.478 5.986 93.514 ;
               RECT 5.934 94.678 5.986 94.714 ;
               RECT 5.934 95.878 5.986 95.914 ;
               RECT 5.934 97.078 5.986 97.114 ;
               RECT 5.934 98.278 5.986 98.314 ;
               RECT 5.934 99.478 5.986 99.514 ;
               RECT 5.934 100.678 5.986 100.714 ;
               RECT 5.934 101.878 5.986 101.914 ;
               RECT 5.934 103.078 5.986 103.114 ;
               RECT 5.934 104.278 5.986 104.314 ;
               RECT 6.014 0.806 6.066 0.842 ;
               RECT 6.014 2.006 6.066 2.042 ;
               RECT 6.014 3.206 6.066 3.242 ;
               RECT 6.014 4.406 6.066 4.442 ;
               RECT 6.014 5.606 6.066 5.642 ;
               RECT 6.014 6.806 6.066 6.842 ;
               RECT 6.014 8.006 6.066 8.042 ;
               RECT 6.014 9.206 6.066 9.242 ;
               RECT 6.014 10.406 6.066 10.442 ;
               RECT 6.014 11.606 6.066 11.642 ;
               RECT 6.014 12.806 6.066 12.842 ;
               RECT 6.014 14.006 6.066 14.042 ;
               RECT 6.014 15.206 6.066 15.242 ;
               RECT 6.014 16.406 6.066 16.442 ;
               RECT 6.014 17.606 6.066 17.642 ;
               RECT 6.014 18.806 6.066 18.842 ;
               RECT 6.014 20.006 6.066 20.042 ;
               RECT 6.014 21.206 6.066 21.242 ;
               RECT 6.014 22.406 6.066 22.442 ;
               RECT 6.014 23.606 6.066 23.642 ;
               RECT 6.014 24.806 6.066 24.842 ;
               RECT 6.014 26.006 6.066 26.042 ;
               RECT 6.014 27.206 6.066 27.242 ;
               RECT 6.014 28.406 6.066 28.442 ;
               RECT 6.014 29.606 6.066 29.642 ;
               RECT 6.014 30.806 6.066 30.842 ;
               RECT 6.014 32.006 6.066 32.042 ;
               RECT 6.014 33.206 6.066 33.242 ;
               RECT 6.014 34.406 6.066 34.442 ;
               RECT 6.014 35.606 6.066 35.642 ;
               RECT 6.014 36.806 6.066 36.842 ;
               RECT 6.014 38.006 6.066 38.042 ;
               RECT 6.014 39.206 6.066 39.242 ;
               RECT 6.014 40.406 6.066 40.442 ;
               RECT 6.014 41.606 6.066 41.642 ;
               RECT 6.014 42.806 6.066 42.842 ;
               RECT 6.014 44.006 6.066 44.042 ;
               RECT 6.014 45.206 6.066 45.242 ;
               RECT 6.014 46.406 6.066 46.442 ;
               RECT 6.014 47.606 6.066 47.642 ;
               RECT 6.014 49.422 6.066 49.458 ;
               RECT 6.014 49.662 6.066 49.698 ;
               RECT 6.014 55.422 6.066 55.458 ;
               RECT 6.014 55.662 6.066 55.698 ;
               RECT 6.014 56.726 6.066 56.762 ;
               RECT 6.014 57.926 6.066 57.962 ;
               RECT 6.014 59.126 6.066 59.162 ;
               RECT 6.014 60.326 6.066 60.362 ;
               RECT 6.014 61.526 6.066 61.562 ;
               RECT 6.014 62.726 6.066 62.762 ;
               RECT 6.014 63.926 6.066 63.962 ;
               RECT 6.014 65.126 6.066 65.162 ;
               RECT 6.014 66.326 6.066 66.362 ;
               RECT 6.014 67.526 6.066 67.562 ;
               RECT 6.014 68.726 6.066 68.762 ;
               RECT 6.014 69.926 6.066 69.962 ;
               RECT 6.014 71.126 6.066 71.162 ;
               RECT 6.014 72.326 6.066 72.362 ;
               RECT 6.014 73.526 6.066 73.562 ;
               RECT 6.014 74.726 6.066 74.762 ;
               RECT 6.014 75.926 6.066 75.962 ;
               RECT 6.014 77.126 6.066 77.162 ;
               RECT 6.014 78.326 6.066 78.362 ;
               RECT 6.014 79.526 6.066 79.562 ;
               RECT 6.014 80.726 6.066 80.762 ;
               RECT 6.014 81.926 6.066 81.962 ;
               RECT 6.014 83.126 6.066 83.162 ;
               RECT 6.014 84.326 6.066 84.362 ;
               RECT 6.014 85.526 6.066 85.562 ;
               RECT 6.014 86.726 6.066 86.762 ;
               RECT 6.014 87.926 6.066 87.962 ;
               RECT 6.014 89.126 6.066 89.162 ;
               RECT 6.014 90.326 6.066 90.362 ;
               RECT 6.014 91.526 6.066 91.562 ;
               RECT 6.014 92.726 6.066 92.762 ;
               RECT 6.014 93.926 6.066 93.962 ;
               RECT 6.014 95.126 6.066 95.162 ;
               RECT 6.014 96.326 6.066 96.362 ;
               RECT 6.014 97.526 6.066 97.562 ;
               RECT 6.014 98.726 6.066 98.762 ;
               RECT 6.014 99.926 6.066 99.962 ;
               RECT 6.014 101.126 6.066 101.162 ;
               RECT 6.014 102.326 6.066 102.362 ;
               RECT 6.014 103.526 6.066 103.562 ;
               RECT 6.094 1.558 6.146 1.594 ;
               RECT 6.094 2.758 6.146 2.794 ;
               RECT 6.094 3.958 6.146 3.994 ;
               RECT 6.094 5.158 6.146 5.194 ;
               RECT 6.094 6.358 6.146 6.394 ;
               RECT 6.094 7.558 6.146 7.594 ;
               RECT 6.094 8.758 6.146 8.794 ;
               RECT 6.094 9.958 6.146 9.994 ;
               RECT 6.094 11.158 6.146 11.194 ;
               RECT 6.094 12.358 6.146 12.394 ;
               RECT 6.094 13.558 6.146 13.594 ;
               RECT 6.094 14.758 6.146 14.794 ;
               RECT 6.094 15.958 6.146 15.994 ;
               RECT 6.094 17.158 6.146 17.194 ;
               RECT 6.094 18.358 6.146 18.394 ;
               RECT 6.094 19.558 6.146 19.594 ;
               RECT 6.094 20.758 6.146 20.794 ;
               RECT 6.094 21.958 6.146 21.994 ;
               RECT 6.094 23.158 6.146 23.194 ;
               RECT 6.094 24.358 6.146 24.394 ;
               RECT 6.094 25.558 6.146 25.594 ;
               RECT 6.094 26.758 6.146 26.794 ;
               RECT 6.094 27.958 6.146 27.994 ;
               RECT 6.094 29.158 6.146 29.194 ;
               RECT 6.094 30.358 6.146 30.394 ;
               RECT 6.094 31.558 6.146 31.594 ;
               RECT 6.094 32.758 6.146 32.794 ;
               RECT 6.094 33.958 6.146 33.994 ;
               RECT 6.094 35.158 6.146 35.194 ;
               RECT 6.094 36.358 6.146 36.394 ;
               RECT 6.094 37.558 6.146 37.594 ;
               RECT 6.094 38.758 6.146 38.794 ;
               RECT 6.094 39.958 6.146 39.994 ;
               RECT 6.094 41.158 6.146 41.194 ;
               RECT 6.094 42.358 6.146 42.394 ;
               RECT 6.094 43.558 6.146 43.594 ;
               RECT 6.094 44.758 6.146 44.794 ;
               RECT 6.094 45.958 6.146 45.994 ;
               RECT 6.094 47.158 6.146 47.194 ;
               RECT 6.094 48.358 6.146 48.394 ;
               RECT 6.094 50.142 6.146 50.178 ;
               RECT 6.094 50.382 6.146 50.418 ;
               RECT 6.094 54.702 6.146 54.738 ;
               RECT 6.094 54.942 6.146 54.978 ;
               RECT 6.094 57.478 6.146 57.514 ;
               RECT 6.094 58.678 6.146 58.714 ;
               RECT 6.094 59.878 6.146 59.914 ;
               RECT 6.094 61.078 6.146 61.114 ;
               RECT 6.094 62.278 6.146 62.314 ;
               RECT 6.094 63.478 6.146 63.514 ;
               RECT 6.094 64.678 6.146 64.714 ;
               RECT 6.094 65.878 6.146 65.914 ;
               RECT 6.094 67.078 6.146 67.114 ;
               RECT 6.094 68.278 6.146 68.314 ;
               RECT 6.094 69.478 6.146 69.514 ;
               RECT 6.094 70.678 6.146 70.714 ;
               RECT 6.094 71.878 6.146 71.914 ;
               RECT 6.094 73.078 6.146 73.114 ;
               RECT 6.094 74.278 6.146 74.314 ;
               RECT 6.094 75.478 6.146 75.514 ;
               RECT 6.094 76.678 6.146 76.714 ;
               RECT 6.094 77.878 6.146 77.914 ;
               RECT 6.094 79.078 6.146 79.114 ;
               RECT 6.094 80.278 6.146 80.314 ;
               RECT 6.094 81.478 6.146 81.514 ;
               RECT 6.094 82.678 6.146 82.714 ;
               RECT 6.094 83.878 6.146 83.914 ;
               RECT 6.094 85.078 6.146 85.114 ;
               RECT 6.094 86.278 6.146 86.314 ;
               RECT 6.094 87.478 6.146 87.514 ;
               RECT 6.094 88.678 6.146 88.714 ;
               RECT 6.094 89.878 6.146 89.914 ;
               RECT 6.094 91.078 6.146 91.114 ;
               RECT 6.094 92.278 6.146 92.314 ;
               RECT 6.094 93.478 6.146 93.514 ;
               RECT 6.094 94.678 6.146 94.714 ;
               RECT 6.094 95.878 6.146 95.914 ;
               RECT 6.094 97.078 6.146 97.114 ;
               RECT 6.094 98.278 6.146 98.314 ;
               RECT 6.094 99.478 6.146 99.514 ;
               RECT 6.094 100.678 6.146 100.714 ;
               RECT 6.094 101.878 6.146 101.914 ;
               RECT 6.094 103.078 6.146 103.114 ;
               RECT 6.094 104.278 6.146 104.314 ;
               RECT 6.174 0.281 6.226 0.317 ;
               RECT 6.174 104.803 6.226 104.839 ;
               RECT 6.254 0.806 6.306 0.842 ;
               RECT 6.254 2.006 6.306 2.042 ;
               RECT 6.254 3.206 6.306 3.242 ;
               RECT 6.254 4.406 6.306 4.442 ;
               RECT 6.254 5.606 6.306 5.642 ;
               RECT 6.254 6.806 6.306 6.842 ;
               RECT 6.254 8.006 6.306 8.042 ;
               RECT 6.254 9.206 6.306 9.242 ;
               RECT 6.254 10.406 6.306 10.442 ;
               RECT 6.254 11.606 6.306 11.642 ;
               RECT 6.254 12.806 6.306 12.842 ;
               RECT 6.254 14.006 6.306 14.042 ;
               RECT 6.254 15.206 6.306 15.242 ;
               RECT 6.254 16.406 6.306 16.442 ;
               RECT 6.254 17.606 6.306 17.642 ;
               RECT 6.254 18.806 6.306 18.842 ;
               RECT 6.254 20.006 6.306 20.042 ;
               RECT 6.254 21.206 6.306 21.242 ;
               RECT 6.254 22.406 6.306 22.442 ;
               RECT 6.254 23.606 6.306 23.642 ;
               RECT 6.254 24.806 6.306 24.842 ;
               RECT 6.254 26.006 6.306 26.042 ;
               RECT 6.254 27.206 6.306 27.242 ;
               RECT 6.254 28.406 6.306 28.442 ;
               RECT 6.254 29.606 6.306 29.642 ;
               RECT 6.254 30.806 6.306 30.842 ;
               RECT 6.254 32.006 6.306 32.042 ;
               RECT 6.254 33.206 6.306 33.242 ;
               RECT 6.254 34.406 6.306 34.442 ;
               RECT 6.254 35.606 6.306 35.642 ;
               RECT 6.254 36.806 6.306 36.842 ;
               RECT 6.254 38.006 6.306 38.042 ;
               RECT 6.254 39.206 6.306 39.242 ;
               RECT 6.254 40.406 6.306 40.442 ;
               RECT 6.254 41.606 6.306 41.642 ;
               RECT 6.254 42.806 6.306 42.842 ;
               RECT 6.254 44.006 6.306 44.042 ;
               RECT 6.254 45.206 6.306 45.242 ;
               RECT 6.254 46.406 6.306 46.442 ;
               RECT 6.254 47.606 6.306 47.642 ;
               RECT 6.254 49.422 6.306 49.458 ;
               RECT 6.254 49.662 6.306 49.698 ;
               RECT 6.254 55.422 6.306 55.458 ;
               RECT 6.254 55.662 6.306 55.698 ;
               RECT 6.254 56.726 6.306 56.762 ;
               RECT 6.254 57.926 6.306 57.962 ;
               RECT 6.254 59.126 6.306 59.162 ;
               RECT 6.254 60.326 6.306 60.362 ;
               RECT 6.254 61.526 6.306 61.562 ;
               RECT 6.254 62.726 6.306 62.762 ;
               RECT 6.254 63.926 6.306 63.962 ;
               RECT 6.254 65.126 6.306 65.162 ;
               RECT 6.254 66.326 6.306 66.362 ;
               RECT 6.254 67.526 6.306 67.562 ;
               RECT 6.254 68.726 6.306 68.762 ;
               RECT 6.254 69.926 6.306 69.962 ;
               RECT 6.254 71.126 6.306 71.162 ;
               RECT 6.254 72.326 6.306 72.362 ;
               RECT 6.254 73.526 6.306 73.562 ;
               RECT 6.254 74.726 6.306 74.762 ;
               RECT 6.254 75.926 6.306 75.962 ;
               RECT 6.254 77.126 6.306 77.162 ;
               RECT 6.254 78.326 6.306 78.362 ;
               RECT 6.254 79.526 6.306 79.562 ;
               RECT 6.254 80.726 6.306 80.762 ;
               RECT 6.254 81.926 6.306 81.962 ;
               RECT 6.254 83.126 6.306 83.162 ;
               RECT 6.254 84.326 6.306 84.362 ;
               RECT 6.254 85.526 6.306 85.562 ;
               RECT 6.254 86.726 6.306 86.762 ;
               RECT 6.254 87.926 6.306 87.962 ;
               RECT 6.254 89.126 6.306 89.162 ;
               RECT 6.254 90.326 6.306 90.362 ;
               RECT 6.254 91.526 6.306 91.562 ;
               RECT 6.254 92.726 6.306 92.762 ;
               RECT 6.254 93.926 6.306 93.962 ;
               RECT 6.254 95.126 6.306 95.162 ;
               RECT 6.254 96.326 6.306 96.362 ;
               RECT 6.254 97.526 6.306 97.562 ;
               RECT 6.254 98.726 6.306 98.762 ;
               RECT 6.254 99.926 6.306 99.962 ;
               RECT 6.254 101.126 6.306 101.162 ;
               RECT 6.254 102.326 6.306 102.362 ;
               RECT 6.254 103.526 6.306 103.562 ;
               RECT 6.334 1.558 6.386 1.594 ;
               RECT 6.334 2.758 6.386 2.794 ;
               RECT 6.334 3.958 6.386 3.994 ;
               RECT 6.334 5.158 6.386 5.194 ;
               RECT 6.334 6.358 6.386 6.394 ;
               RECT 6.334 7.558 6.386 7.594 ;
               RECT 6.334 8.758 6.386 8.794 ;
               RECT 6.334 9.958 6.386 9.994 ;
               RECT 6.334 11.158 6.386 11.194 ;
               RECT 6.334 12.358 6.386 12.394 ;
               RECT 6.334 13.558 6.386 13.594 ;
               RECT 6.334 14.758 6.386 14.794 ;
               RECT 6.334 15.958 6.386 15.994 ;
               RECT 6.334 17.158 6.386 17.194 ;
               RECT 6.334 18.358 6.386 18.394 ;
               RECT 6.334 19.558 6.386 19.594 ;
               RECT 6.334 20.758 6.386 20.794 ;
               RECT 6.334 21.958 6.386 21.994 ;
               RECT 6.334 23.158 6.386 23.194 ;
               RECT 6.334 24.358 6.386 24.394 ;
               RECT 6.334 25.558 6.386 25.594 ;
               RECT 6.334 26.758 6.386 26.794 ;
               RECT 6.334 27.958 6.386 27.994 ;
               RECT 6.334 29.158 6.386 29.194 ;
               RECT 6.334 30.358 6.386 30.394 ;
               RECT 6.334 31.558 6.386 31.594 ;
               RECT 6.334 32.758 6.386 32.794 ;
               RECT 6.334 33.958 6.386 33.994 ;
               RECT 6.334 35.158 6.386 35.194 ;
               RECT 6.334 36.358 6.386 36.394 ;
               RECT 6.334 37.558 6.386 37.594 ;
               RECT 6.334 38.758 6.386 38.794 ;
               RECT 6.334 39.958 6.386 39.994 ;
               RECT 6.334 41.158 6.386 41.194 ;
               RECT 6.334 42.358 6.386 42.394 ;
               RECT 6.334 43.558 6.386 43.594 ;
               RECT 6.334 44.758 6.386 44.794 ;
               RECT 6.334 45.958 6.386 45.994 ;
               RECT 6.334 47.158 6.386 47.194 ;
               RECT 6.334 48.358 6.386 48.394 ;
               RECT 6.334 50.142 6.386 50.178 ;
               RECT 6.334 50.382 6.386 50.418 ;
               RECT 6.334 54.702 6.386 54.738 ;
               RECT 6.334 54.942 6.386 54.978 ;
               RECT 6.334 57.478 6.386 57.514 ;
               RECT 6.334 58.678 6.386 58.714 ;
               RECT 6.334 59.878 6.386 59.914 ;
               RECT 6.334 61.078 6.386 61.114 ;
               RECT 6.334 62.278 6.386 62.314 ;
               RECT 6.334 63.478 6.386 63.514 ;
               RECT 6.334 64.678 6.386 64.714 ;
               RECT 6.334 65.878 6.386 65.914 ;
               RECT 6.334 67.078 6.386 67.114 ;
               RECT 6.334 68.278 6.386 68.314 ;
               RECT 6.334 69.478 6.386 69.514 ;
               RECT 6.334 70.678 6.386 70.714 ;
               RECT 6.334 71.878 6.386 71.914 ;
               RECT 6.334 73.078 6.386 73.114 ;
               RECT 6.334 74.278 6.386 74.314 ;
               RECT 6.334 75.478 6.386 75.514 ;
               RECT 6.334 76.678 6.386 76.714 ;
               RECT 6.334 77.878 6.386 77.914 ;
               RECT 6.334 79.078 6.386 79.114 ;
               RECT 6.334 80.278 6.386 80.314 ;
               RECT 6.334 81.478 6.386 81.514 ;
               RECT 6.334 82.678 6.386 82.714 ;
               RECT 6.334 83.878 6.386 83.914 ;
               RECT 6.334 85.078 6.386 85.114 ;
               RECT 6.334 86.278 6.386 86.314 ;
               RECT 6.334 87.478 6.386 87.514 ;
               RECT 6.334 88.678 6.386 88.714 ;
               RECT 6.334 89.878 6.386 89.914 ;
               RECT 6.334 91.078 6.386 91.114 ;
               RECT 6.334 92.278 6.386 92.314 ;
               RECT 6.334 93.478 6.386 93.514 ;
               RECT 6.334 94.678 6.386 94.714 ;
               RECT 6.334 95.878 6.386 95.914 ;
               RECT 6.334 97.078 6.386 97.114 ;
               RECT 6.334 98.278 6.386 98.314 ;
               RECT 6.334 99.478 6.386 99.514 ;
               RECT 6.334 100.678 6.386 100.714 ;
               RECT 6.334 101.878 6.386 101.914 ;
               RECT 6.334 103.078 6.386 103.114 ;
               RECT 6.334 104.278 6.386 104.314 ;
               RECT 6.414 0.806 6.466 0.842 ;
               RECT 6.414 2.006 6.466 2.042 ;
               RECT 6.414 3.206 6.466 3.242 ;
               RECT 6.414 4.406 6.466 4.442 ;
               RECT 6.414 5.606 6.466 5.642 ;
               RECT 6.414 6.806 6.466 6.842 ;
               RECT 6.414 8.006 6.466 8.042 ;
               RECT 6.414 9.206 6.466 9.242 ;
               RECT 6.414 10.406 6.466 10.442 ;
               RECT 6.414 11.606 6.466 11.642 ;
               RECT 6.414 12.806 6.466 12.842 ;
               RECT 6.414 14.006 6.466 14.042 ;
               RECT 6.414 15.206 6.466 15.242 ;
               RECT 6.414 16.406 6.466 16.442 ;
               RECT 6.414 17.606 6.466 17.642 ;
               RECT 6.414 18.806 6.466 18.842 ;
               RECT 6.414 20.006 6.466 20.042 ;
               RECT 6.414 21.206 6.466 21.242 ;
               RECT 6.414 22.406 6.466 22.442 ;
               RECT 6.414 23.606 6.466 23.642 ;
               RECT 6.414 24.806 6.466 24.842 ;
               RECT 6.414 26.006 6.466 26.042 ;
               RECT 6.414 27.206 6.466 27.242 ;
               RECT 6.414 28.406 6.466 28.442 ;
               RECT 6.414 29.606 6.466 29.642 ;
               RECT 6.414 30.806 6.466 30.842 ;
               RECT 6.414 32.006 6.466 32.042 ;
               RECT 6.414 33.206 6.466 33.242 ;
               RECT 6.414 34.406 6.466 34.442 ;
               RECT 6.414 35.606 6.466 35.642 ;
               RECT 6.414 36.806 6.466 36.842 ;
               RECT 6.414 38.006 6.466 38.042 ;
               RECT 6.414 39.206 6.466 39.242 ;
               RECT 6.414 40.406 6.466 40.442 ;
               RECT 6.414 41.606 6.466 41.642 ;
               RECT 6.414 42.806 6.466 42.842 ;
               RECT 6.414 44.006 6.466 44.042 ;
               RECT 6.414 45.206 6.466 45.242 ;
               RECT 6.414 46.406 6.466 46.442 ;
               RECT 6.414 47.606 6.466 47.642 ;
               RECT 6.414 49.422 6.466 49.458 ;
               RECT 6.414 49.662 6.466 49.698 ;
               RECT 6.414 55.422 6.466 55.458 ;
               RECT 6.414 55.662 6.466 55.698 ;
               RECT 6.414 56.726 6.466 56.762 ;
               RECT 6.414 57.926 6.466 57.962 ;
               RECT 6.414 59.126 6.466 59.162 ;
               RECT 6.414 60.326 6.466 60.362 ;
               RECT 6.414 61.526 6.466 61.562 ;
               RECT 6.414 62.726 6.466 62.762 ;
               RECT 6.414 63.926 6.466 63.962 ;
               RECT 6.414 65.126 6.466 65.162 ;
               RECT 6.414 66.326 6.466 66.362 ;
               RECT 6.414 67.526 6.466 67.562 ;
               RECT 6.414 68.726 6.466 68.762 ;
               RECT 6.414 69.926 6.466 69.962 ;
               RECT 6.414 71.126 6.466 71.162 ;
               RECT 6.414 72.326 6.466 72.362 ;
               RECT 6.414 73.526 6.466 73.562 ;
               RECT 6.414 74.726 6.466 74.762 ;
               RECT 6.414 75.926 6.466 75.962 ;
               RECT 6.414 77.126 6.466 77.162 ;
               RECT 6.414 78.326 6.466 78.362 ;
               RECT 6.414 79.526 6.466 79.562 ;
               RECT 6.414 80.726 6.466 80.762 ;
               RECT 6.414 81.926 6.466 81.962 ;
               RECT 6.414 83.126 6.466 83.162 ;
               RECT 6.414 84.326 6.466 84.362 ;
               RECT 6.414 85.526 6.466 85.562 ;
               RECT 6.414 86.726 6.466 86.762 ;
               RECT 6.414 87.926 6.466 87.962 ;
               RECT 6.414 89.126 6.466 89.162 ;
               RECT 6.414 90.326 6.466 90.362 ;
               RECT 6.414 91.526 6.466 91.562 ;
               RECT 6.414 92.726 6.466 92.762 ;
               RECT 6.414 93.926 6.466 93.962 ;
               RECT 6.414 95.126 6.466 95.162 ;
               RECT 6.414 96.326 6.466 96.362 ;
               RECT 6.414 97.526 6.466 97.562 ;
               RECT 6.414 98.726 6.466 98.762 ;
               RECT 6.414 99.926 6.466 99.962 ;
               RECT 6.414 101.126 6.466 101.162 ;
               RECT 6.414 102.326 6.466 102.362 ;
               RECT 6.414 103.526 6.466 103.562 ;
               RECT 6.494 1.558 6.546 1.594 ;
               RECT 6.494 2.758 6.546 2.794 ;
               RECT 6.494 3.958 6.546 3.994 ;
               RECT 6.494 5.158 6.546 5.194 ;
               RECT 6.494 6.358 6.546 6.394 ;
               RECT 6.494 7.558 6.546 7.594 ;
               RECT 6.494 8.758 6.546 8.794 ;
               RECT 6.494 9.958 6.546 9.994 ;
               RECT 6.494 11.158 6.546 11.194 ;
               RECT 6.494 12.358 6.546 12.394 ;
               RECT 6.494 13.558 6.546 13.594 ;
               RECT 6.494 14.758 6.546 14.794 ;
               RECT 6.494 15.958 6.546 15.994 ;
               RECT 6.494 17.158 6.546 17.194 ;
               RECT 6.494 18.358 6.546 18.394 ;
               RECT 6.494 19.558 6.546 19.594 ;
               RECT 6.494 20.758 6.546 20.794 ;
               RECT 6.494 21.958 6.546 21.994 ;
               RECT 6.494 23.158 6.546 23.194 ;
               RECT 6.494 24.358 6.546 24.394 ;
               RECT 6.494 25.558 6.546 25.594 ;
               RECT 6.494 26.758 6.546 26.794 ;
               RECT 6.494 27.958 6.546 27.994 ;
               RECT 6.494 29.158 6.546 29.194 ;
               RECT 6.494 30.358 6.546 30.394 ;
               RECT 6.494 31.558 6.546 31.594 ;
               RECT 6.494 32.758 6.546 32.794 ;
               RECT 6.494 33.958 6.546 33.994 ;
               RECT 6.494 35.158 6.546 35.194 ;
               RECT 6.494 36.358 6.546 36.394 ;
               RECT 6.494 37.558 6.546 37.594 ;
               RECT 6.494 38.758 6.546 38.794 ;
               RECT 6.494 39.958 6.546 39.994 ;
               RECT 6.494 41.158 6.546 41.194 ;
               RECT 6.494 42.358 6.546 42.394 ;
               RECT 6.494 43.558 6.546 43.594 ;
               RECT 6.494 44.758 6.546 44.794 ;
               RECT 6.494 45.958 6.546 45.994 ;
               RECT 6.494 47.158 6.546 47.194 ;
               RECT 6.494 48.358 6.546 48.394 ;
               RECT 6.494 50.142 6.546 50.178 ;
               RECT 6.494 50.382 6.546 50.418 ;
               RECT 6.494 54.702 6.546 54.738 ;
               RECT 6.494 54.942 6.546 54.978 ;
               RECT 6.494 57.478 6.546 57.514 ;
               RECT 6.494 58.678 6.546 58.714 ;
               RECT 6.494 59.878 6.546 59.914 ;
               RECT 6.494 61.078 6.546 61.114 ;
               RECT 6.494 62.278 6.546 62.314 ;
               RECT 6.494 63.478 6.546 63.514 ;
               RECT 6.494 64.678 6.546 64.714 ;
               RECT 6.494 65.878 6.546 65.914 ;
               RECT 6.494 67.078 6.546 67.114 ;
               RECT 6.494 68.278 6.546 68.314 ;
               RECT 6.494 69.478 6.546 69.514 ;
               RECT 6.494 70.678 6.546 70.714 ;
               RECT 6.494 71.878 6.546 71.914 ;
               RECT 6.494 73.078 6.546 73.114 ;
               RECT 6.494 74.278 6.546 74.314 ;
               RECT 6.494 75.478 6.546 75.514 ;
               RECT 6.494 76.678 6.546 76.714 ;
               RECT 6.494 77.878 6.546 77.914 ;
               RECT 6.494 79.078 6.546 79.114 ;
               RECT 6.494 80.278 6.546 80.314 ;
               RECT 6.494 81.478 6.546 81.514 ;
               RECT 6.494 82.678 6.546 82.714 ;
               RECT 6.494 83.878 6.546 83.914 ;
               RECT 6.494 85.078 6.546 85.114 ;
               RECT 6.494 86.278 6.546 86.314 ;
               RECT 6.494 87.478 6.546 87.514 ;
               RECT 6.494 88.678 6.546 88.714 ;
               RECT 6.494 89.878 6.546 89.914 ;
               RECT 6.494 91.078 6.546 91.114 ;
               RECT 6.494 92.278 6.546 92.314 ;
               RECT 6.494 93.478 6.546 93.514 ;
               RECT 6.494 94.678 6.546 94.714 ;
               RECT 6.494 95.878 6.546 95.914 ;
               RECT 6.494 97.078 6.546 97.114 ;
               RECT 6.494 98.278 6.546 98.314 ;
               RECT 6.494 99.478 6.546 99.514 ;
               RECT 6.494 100.678 6.546 100.714 ;
               RECT 6.494 101.878 6.546 101.914 ;
               RECT 6.494 103.078 6.546 103.114 ;
               RECT 6.494 104.278 6.546 104.314 ;
               RECT 6.574 0.281 6.626 0.317 ;
               RECT 6.574 104.803 6.626 104.839 ;
               RECT 6.654 0.806 6.706 0.842 ;
               RECT 6.654 2.006 6.706 2.042 ;
               RECT 6.654 3.206 6.706 3.242 ;
               RECT 6.654 4.406 6.706 4.442 ;
               RECT 6.654 5.606 6.706 5.642 ;
               RECT 6.654 6.806 6.706 6.842 ;
               RECT 6.654 8.006 6.706 8.042 ;
               RECT 6.654 9.206 6.706 9.242 ;
               RECT 6.654 10.406 6.706 10.442 ;
               RECT 6.654 11.606 6.706 11.642 ;
               RECT 6.654 12.806 6.706 12.842 ;
               RECT 6.654 14.006 6.706 14.042 ;
               RECT 6.654 15.206 6.706 15.242 ;
               RECT 6.654 16.406 6.706 16.442 ;
               RECT 6.654 17.606 6.706 17.642 ;
               RECT 6.654 18.806 6.706 18.842 ;
               RECT 6.654 20.006 6.706 20.042 ;
               RECT 6.654 21.206 6.706 21.242 ;
               RECT 6.654 22.406 6.706 22.442 ;
               RECT 6.654 23.606 6.706 23.642 ;
               RECT 6.654 24.806 6.706 24.842 ;
               RECT 6.654 26.006 6.706 26.042 ;
               RECT 6.654 27.206 6.706 27.242 ;
               RECT 6.654 28.406 6.706 28.442 ;
               RECT 6.654 29.606 6.706 29.642 ;
               RECT 6.654 30.806 6.706 30.842 ;
               RECT 6.654 32.006 6.706 32.042 ;
               RECT 6.654 33.206 6.706 33.242 ;
               RECT 6.654 34.406 6.706 34.442 ;
               RECT 6.654 35.606 6.706 35.642 ;
               RECT 6.654 36.806 6.706 36.842 ;
               RECT 6.654 38.006 6.706 38.042 ;
               RECT 6.654 39.206 6.706 39.242 ;
               RECT 6.654 40.406 6.706 40.442 ;
               RECT 6.654 41.606 6.706 41.642 ;
               RECT 6.654 42.806 6.706 42.842 ;
               RECT 6.654 44.006 6.706 44.042 ;
               RECT 6.654 45.206 6.706 45.242 ;
               RECT 6.654 46.406 6.706 46.442 ;
               RECT 6.654 47.606 6.706 47.642 ;
               RECT 6.654 49.422 6.706 49.458 ;
               RECT 6.654 49.662 6.706 49.698 ;
               RECT 6.654 51.102 6.706 51.138 ;
               RECT 6.654 51.582 6.706 51.618 ;
               RECT 6.654 53.502 6.706 53.538 ;
               RECT 6.654 53.982 6.706 54.018 ;
               RECT 6.654 55.422 6.706 55.458 ;
               RECT 6.654 55.662 6.706 55.698 ;
               RECT 6.654 56.726 6.706 56.762 ;
               RECT 6.654 57.926 6.706 57.962 ;
               RECT 6.654 59.126 6.706 59.162 ;
               RECT 6.654 60.326 6.706 60.362 ;
               RECT 6.654 61.526 6.706 61.562 ;
               RECT 6.654 62.726 6.706 62.762 ;
               RECT 6.654 63.926 6.706 63.962 ;
               RECT 6.654 65.126 6.706 65.162 ;
               RECT 6.654 66.326 6.706 66.362 ;
               RECT 6.654 67.526 6.706 67.562 ;
               RECT 6.654 68.726 6.706 68.762 ;
               RECT 6.654 69.926 6.706 69.962 ;
               RECT 6.654 71.126 6.706 71.162 ;
               RECT 6.654 72.326 6.706 72.362 ;
               RECT 6.654 73.526 6.706 73.562 ;
               RECT 6.654 74.726 6.706 74.762 ;
               RECT 6.654 75.926 6.706 75.962 ;
               RECT 6.654 77.126 6.706 77.162 ;
               RECT 6.654 78.326 6.706 78.362 ;
               RECT 6.654 79.526 6.706 79.562 ;
               RECT 6.654 80.726 6.706 80.762 ;
               RECT 6.654 81.926 6.706 81.962 ;
               RECT 6.654 83.126 6.706 83.162 ;
               RECT 6.654 84.326 6.706 84.362 ;
               RECT 6.654 85.526 6.706 85.562 ;
               RECT 6.654 86.726 6.706 86.762 ;
               RECT 6.654 87.926 6.706 87.962 ;
               RECT 6.654 89.126 6.706 89.162 ;
               RECT 6.654 90.326 6.706 90.362 ;
               RECT 6.654 91.526 6.706 91.562 ;
               RECT 6.654 92.726 6.706 92.762 ;
               RECT 6.654 93.926 6.706 93.962 ;
               RECT 6.654 95.126 6.706 95.162 ;
               RECT 6.654 96.326 6.706 96.362 ;
               RECT 6.654 97.526 6.706 97.562 ;
               RECT 6.654 98.726 6.706 98.762 ;
               RECT 6.654 99.926 6.706 99.962 ;
               RECT 6.654 101.126 6.706 101.162 ;
               RECT 6.654 102.326 6.706 102.362 ;
               RECT 6.654 103.526 6.706 103.562 ;
               RECT 6.734 1.558 6.786 1.594 ;
               RECT 6.734 2.758 6.786 2.794 ;
               RECT 6.734 3.958 6.786 3.994 ;
               RECT 6.734 5.158 6.786 5.194 ;
               RECT 6.734 6.358 6.786 6.394 ;
               RECT 6.734 7.558 6.786 7.594 ;
               RECT 6.734 8.758 6.786 8.794 ;
               RECT 6.734 9.958 6.786 9.994 ;
               RECT 6.734 11.158 6.786 11.194 ;
               RECT 6.734 12.358 6.786 12.394 ;
               RECT 6.734 13.558 6.786 13.594 ;
               RECT 6.734 14.758 6.786 14.794 ;
               RECT 6.734 15.958 6.786 15.994 ;
               RECT 6.734 17.158 6.786 17.194 ;
               RECT 6.734 18.358 6.786 18.394 ;
               RECT 6.734 19.558 6.786 19.594 ;
               RECT 6.734 20.758 6.786 20.794 ;
               RECT 6.734 21.958 6.786 21.994 ;
               RECT 6.734 23.158 6.786 23.194 ;
               RECT 6.734 24.358 6.786 24.394 ;
               RECT 6.734 25.558 6.786 25.594 ;
               RECT 6.734 26.758 6.786 26.794 ;
               RECT 6.734 27.958 6.786 27.994 ;
               RECT 6.734 29.158 6.786 29.194 ;
               RECT 6.734 30.358 6.786 30.394 ;
               RECT 6.734 31.558 6.786 31.594 ;
               RECT 6.734 32.758 6.786 32.794 ;
               RECT 6.734 33.958 6.786 33.994 ;
               RECT 6.734 35.158 6.786 35.194 ;
               RECT 6.734 36.358 6.786 36.394 ;
               RECT 6.734 37.558 6.786 37.594 ;
               RECT 6.734 38.758 6.786 38.794 ;
               RECT 6.734 39.958 6.786 39.994 ;
               RECT 6.734 41.158 6.786 41.194 ;
               RECT 6.734 42.358 6.786 42.394 ;
               RECT 6.734 43.558 6.786 43.594 ;
               RECT 6.734 44.758 6.786 44.794 ;
               RECT 6.734 45.958 6.786 45.994 ;
               RECT 6.734 47.158 6.786 47.194 ;
               RECT 6.734 48.358 6.786 48.394 ;
               RECT 6.734 50.142 6.786 50.178 ;
               RECT 6.734 50.382 6.786 50.418 ;
               RECT 6.734 54.702 6.786 54.738 ;
               RECT 6.734 54.942 6.786 54.978 ;
               RECT 6.734 57.478 6.786 57.514 ;
               RECT 6.734 58.678 6.786 58.714 ;
               RECT 6.734 59.878 6.786 59.914 ;
               RECT 6.734 61.078 6.786 61.114 ;
               RECT 6.734 62.278 6.786 62.314 ;
               RECT 6.734 63.478 6.786 63.514 ;
               RECT 6.734 64.678 6.786 64.714 ;
               RECT 6.734 65.878 6.786 65.914 ;
               RECT 6.734 67.078 6.786 67.114 ;
               RECT 6.734 68.278 6.786 68.314 ;
               RECT 6.734 69.478 6.786 69.514 ;
               RECT 6.734 70.678 6.786 70.714 ;
               RECT 6.734 71.878 6.786 71.914 ;
               RECT 6.734 73.078 6.786 73.114 ;
               RECT 6.734 74.278 6.786 74.314 ;
               RECT 6.734 75.478 6.786 75.514 ;
               RECT 6.734 76.678 6.786 76.714 ;
               RECT 6.734 77.878 6.786 77.914 ;
               RECT 6.734 79.078 6.786 79.114 ;
               RECT 6.734 80.278 6.786 80.314 ;
               RECT 6.734 81.478 6.786 81.514 ;
               RECT 6.734 82.678 6.786 82.714 ;
               RECT 6.734 83.878 6.786 83.914 ;
               RECT 6.734 85.078 6.786 85.114 ;
               RECT 6.734 86.278 6.786 86.314 ;
               RECT 6.734 87.478 6.786 87.514 ;
               RECT 6.734 88.678 6.786 88.714 ;
               RECT 6.734 89.878 6.786 89.914 ;
               RECT 6.734 91.078 6.786 91.114 ;
               RECT 6.734 92.278 6.786 92.314 ;
               RECT 6.734 93.478 6.786 93.514 ;
               RECT 6.734 94.678 6.786 94.714 ;
               RECT 6.734 95.878 6.786 95.914 ;
               RECT 6.734 97.078 6.786 97.114 ;
               RECT 6.734 98.278 6.786 98.314 ;
               RECT 6.734 99.478 6.786 99.514 ;
               RECT 6.734 100.678 6.786 100.714 ;
               RECT 6.734 101.878 6.786 101.914 ;
               RECT 6.734 103.078 6.786 103.114 ;
               RECT 6.734 104.278 6.786 104.314 ;
               RECT 6.814 0.806 6.866 0.842 ;
               RECT 6.814 2.006 6.866 2.042 ;
               RECT 6.814 3.206 6.866 3.242 ;
               RECT 6.814 4.406 6.866 4.442 ;
               RECT 6.814 5.606 6.866 5.642 ;
               RECT 6.814 6.806 6.866 6.842 ;
               RECT 6.814 8.006 6.866 8.042 ;
               RECT 6.814 9.206 6.866 9.242 ;
               RECT 6.814 10.406 6.866 10.442 ;
               RECT 6.814 11.606 6.866 11.642 ;
               RECT 6.814 12.806 6.866 12.842 ;
               RECT 6.814 14.006 6.866 14.042 ;
               RECT 6.814 15.206 6.866 15.242 ;
               RECT 6.814 16.406 6.866 16.442 ;
               RECT 6.814 17.606 6.866 17.642 ;
               RECT 6.814 18.806 6.866 18.842 ;
               RECT 6.814 20.006 6.866 20.042 ;
               RECT 6.814 21.206 6.866 21.242 ;
               RECT 6.814 22.406 6.866 22.442 ;
               RECT 6.814 23.606 6.866 23.642 ;
               RECT 6.814 24.806 6.866 24.842 ;
               RECT 6.814 26.006 6.866 26.042 ;
               RECT 6.814 27.206 6.866 27.242 ;
               RECT 6.814 28.406 6.866 28.442 ;
               RECT 6.814 29.606 6.866 29.642 ;
               RECT 6.814 30.806 6.866 30.842 ;
               RECT 6.814 32.006 6.866 32.042 ;
               RECT 6.814 33.206 6.866 33.242 ;
               RECT 6.814 34.406 6.866 34.442 ;
               RECT 6.814 35.606 6.866 35.642 ;
               RECT 6.814 36.806 6.866 36.842 ;
               RECT 6.814 38.006 6.866 38.042 ;
               RECT 6.814 39.206 6.866 39.242 ;
               RECT 6.814 40.406 6.866 40.442 ;
               RECT 6.814 41.606 6.866 41.642 ;
               RECT 6.814 42.806 6.866 42.842 ;
               RECT 6.814 44.006 6.866 44.042 ;
               RECT 6.814 45.206 6.866 45.242 ;
               RECT 6.814 46.406 6.866 46.442 ;
               RECT 6.814 47.606 6.866 47.642 ;
               RECT 6.814 49.422 6.866 49.458 ;
               RECT 6.814 49.662 6.866 49.698 ;
               RECT 6.814 55.422 6.866 55.458 ;
               RECT 6.814 55.662 6.866 55.698 ;
               RECT 6.814 56.726 6.866 56.762 ;
               RECT 6.814 57.926 6.866 57.962 ;
               RECT 6.814 59.126 6.866 59.162 ;
               RECT 6.814 60.326 6.866 60.362 ;
               RECT 6.814 61.526 6.866 61.562 ;
               RECT 6.814 62.726 6.866 62.762 ;
               RECT 6.814 63.926 6.866 63.962 ;
               RECT 6.814 65.126 6.866 65.162 ;
               RECT 6.814 66.326 6.866 66.362 ;
               RECT 6.814 67.526 6.866 67.562 ;
               RECT 6.814 68.726 6.866 68.762 ;
               RECT 6.814 69.926 6.866 69.962 ;
               RECT 6.814 71.126 6.866 71.162 ;
               RECT 6.814 72.326 6.866 72.362 ;
               RECT 6.814 73.526 6.866 73.562 ;
               RECT 6.814 74.726 6.866 74.762 ;
               RECT 6.814 75.926 6.866 75.962 ;
               RECT 6.814 77.126 6.866 77.162 ;
               RECT 6.814 78.326 6.866 78.362 ;
               RECT 6.814 79.526 6.866 79.562 ;
               RECT 6.814 80.726 6.866 80.762 ;
               RECT 6.814 81.926 6.866 81.962 ;
               RECT 6.814 83.126 6.866 83.162 ;
               RECT 6.814 84.326 6.866 84.362 ;
               RECT 6.814 85.526 6.866 85.562 ;
               RECT 6.814 86.726 6.866 86.762 ;
               RECT 6.814 87.926 6.866 87.962 ;
               RECT 6.814 89.126 6.866 89.162 ;
               RECT 6.814 90.326 6.866 90.362 ;
               RECT 6.814 91.526 6.866 91.562 ;
               RECT 6.814 92.726 6.866 92.762 ;
               RECT 6.814 93.926 6.866 93.962 ;
               RECT 6.814 95.126 6.866 95.162 ;
               RECT 6.814 96.326 6.866 96.362 ;
               RECT 6.814 97.526 6.866 97.562 ;
               RECT 6.814 98.726 6.866 98.762 ;
               RECT 6.814 99.926 6.866 99.962 ;
               RECT 6.814 101.126 6.866 101.162 ;
               RECT 6.814 102.326 6.866 102.362 ;
               RECT 6.814 103.526 6.866 103.562 ;
               RECT 6.894 1.558 6.946 1.594 ;
               RECT 6.894 2.758 6.946 2.794 ;
               RECT 6.894 3.958 6.946 3.994 ;
               RECT 6.894 5.158 6.946 5.194 ;
               RECT 6.894 6.358 6.946 6.394 ;
               RECT 6.894 7.558 6.946 7.594 ;
               RECT 6.894 8.758 6.946 8.794 ;
               RECT 6.894 9.958 6.946 9.994 ;
               RECT 6.894 11.158 6.946 11.194 ;
               RECT 6.894 12.358 6.946 12.394 ;
               RECT 6.894 13.558 6.946 13.594 ;
               RECT 6.894 14.758 6.946 14.794 ;
               RECT 6.894 15.958 6.946 15.994 ;
               RECT 6.894 17.158 6.946 17.194 ;
               RECT 6.894 18.358 6.946 18.394 ;
               RECT 6.894 19.558 6.946 19.594 ;
               RECT 6.894 20.758 6.946 20.794 ;
               RECT 6.894 21.958 6.946 21.994 ;
               RECT 6.894 23.158 6.946 23.194 ;
               RECT 6.894 24.358 6.946 24.394 ;
               RECT 6.894 25.558 6.946 25.594 ;
               RECT 6.894 26.758 6.946 26.794 ;
               RECT 6.894 27.958 6.946 27.994 ;
               RECT 6.894 29.158 6.946 29.194 ;
               RECT 6.894 30.358 6.946 30.394 ;
               RECT 6.894 31.558 6.946 31.594 ;
               RECT 6.894 32.758 6.946 32.794 ;
               RECT 6.894 33.958 6.946 33.994 ;
               RECT 6.894 35.158 6.946 35.194 ;
               RECT 6.894 36.358 6.946 36.394 ;
               RECT 6.894 37.558 6.946 37.594 ;
               RECT 6.894 38.758 6.946 38.794 ;
               RECT 6.894 39.958 6.946 39.994 ;
               RECT 6.894 41.158 6.946 41.194 ;
               RECT 6.894 42.358 6.946 42.394 ;
               RECT 6.894 43.558 6.946 43.594 ;
               RECT 6.894 44.758 6.946 44.794 ;
               RECT 6.894 45.958 6.946 45.994 ;
               RECT 6.894 47.158 6.946 47.194 ;
               RECT 6.894 48.358 6.946 48.394 ;
               RECT 6.894 50.142 6.946 50.178 ;
               RECT 6.894 50.382 6.946 50.418 ;
               RECT 6.894 54.702 6.946 54.738 ;
               RECT 6.894 54.942 6.946 54.978 ;
               RECT 6.894 57.478 6.946 57.514 ;
               RECT 6.894 58.678 6.946 58.714 ;
               RECT 6.894 59.878 6.946 59.914 ;
               RECT 6.894 61.078 6.946 61.114 ;
               RECT 6.894 62.278 6.946 62.314 ;
               RECT 6.894 63.478 6.946 63.514 ;
               RECT 6.894 64.678 6.946 64.714 ;
               RECT 6.894 65.878 6.946 65.914 ;
               RECT 6.894 67.078 6.946 67.114 ;
               RECT 6.894 68.278 6.946 68.314 ;
               RECT 6.894 69.478 6.946 69.514 ;
               RECT 6.894 70.678 6.946 70.714 ;
               RECT 6.894 71.878 6.946 71.914 ;
               RECT 6.894 73.078 6.946 73.114 ;
               RECT 6.894 74.278 6.946 74.314 ;
               RECT 6.894 75.478 6.946 75.514 ;
               RECT 6.894 76.678 6.946 76.714 ;
               RECT 6.894 77.878 6.946 77.914 ;
               RECT 6.894 79.078 6.946 79.114 ;
               RECT 6.894 80.278 6.946 80.314 ;
               RECT 6.894 81.478 6.946 81.514 ;
               RECT 6.894 82.678 6.946 82.714 ;
               RECT 6.894 83.878 6.946 83.914 ;
               RECT 6.894 85.078 6.946 85.114 ;
               RECT 6.894 86.278 6.946 86.314 ;
               RECT 6.894 87.478 6.946 87.514 ;
               RECT 6.894 88.678 6.946 88.714 ;
               RECT 6.894 89.878 6.946 89.914 ;
               RECT 6.894 91.078 6.946 91.114 ;
               RECT 6.894 92.278 6.946 92.314 ;
               RECT 6.894 93.478 6.946 93.514 ;
               RECT 6.894 94.678 6.946 94.714 ;
               RECT 6.894 95.878 6.946 95.914 ;
               RECT 6.894 97.078 6.946 97.114 ;
               RECT 6.894 98.278 6.946 98.314 ;
               RECT 6.894 99.478 6.946 99.514 ;
               RECT 6.894 100.678 6.946 100.714 ;
               RECT 6.894 101.878 6.946 101.914 ;
               RECT 6.894 103.078 6.946 103.114 ;
               RECT 6.894 104.278 6.946 104.314 ;
               RECT 6.974 0.281 7.026 0.317 ;
               RECT 6.974 104.803 7.026 104.839 ;
               RECT 7.054 0.806 7.106 0.842 ;
               RECT 7.054 2.006 7.106 2.042 ;
               RECT 7.054 3.206 7.106 3.242 ;
               RECT 7.054 4.406 7.106 4.442 ;
               RECT 7.054 5.606 7.106 5.642 ;
               RECT 7.054 6.806 7.106 6.842 ;
               RECT 7.054 8.006 7.106 8.042 ;
               RECT 7.054 9.206 7.106 9.242 ;
               RECT 7.054 10.406 7.106 10.442 ;
               RECT 7.054 11.606 7.106 11.642 ;
               RECT 7.054 12.806 7.106 12.842 ;
               RECT 7.054 14.006 7.106 14.042 ;
               RECT 7.054 15.206 7.106 15.242 ;
               RECT 7.054 16.406 7.106 16.442 ;
               RECT 7.054 17.606 7.106 17.642 ;
               RECT 7.054 18.806 7.106 18.842 ;
               RECT 7.054 20.006 7.106 20.042 ;
               RECT 7.054 21.206 7.106 21.242 ;
               RECT 7.054 22.406 7.106 22.442 ;
               RECT 7.054 23.606 7.106 23.642 ;
               RECT 7.054 24.806 7.106 24.842 ;
               RECT 7.054 26.006 7.106 26.042 ;
               RECT 7.054 27.206 7.106 27.242 ;
               RECT 7.054 28.406 7.106 28.442 ;
               RECT 7.054 29.606 7.106 29.642 ;
               RECT 7.054 30.806 7.106 30.842 ;
               RECT 7.054 32.006 7.106 32.042 ;
               RECT 7.054 33.206 7.106 33.242 ;
               RECT 7.054 34.406 7.106 34.442 ;
               RECT 7.054 35.606 7.106 35.642 ;
               RECT 7.054 36.806 7.106 36.842 ;
               RECT 7.054 38.006 7.106 38.042 ;
               RECT 7.054 39.206 7.106 39.242 ;
               RECT 7.054 40.406 7.106 40.442 ;
               RECT 7.054 41.606 7.106 41.642 ;
               RECT 7.054 42.806 7.106 42.842 ;
               RECT 7.054 44.006 7.106 44.042 ;
               RECT 7.054 45.206 7.106 45.242 ;
               RECT 7.054 46.406 7.106 46.442 ;
               RECT 7.054 47.606 7.106 47.642 ;
               RECT 7.054 49.422 7.106 49.458 ;
               RECT 7.054 49.662 7.106 49.698 ;
               RECT 7.054 55.422 7.106 55.458 ;
               RECT 7.054 55.662 7.106 55.698 ;
               RECT 7.054 56.726 7.106 56.762 ;
               RECT 7.054 57.926 7.106 57.962 ;
               RECT 7.054 59.126 7.106 59.162 ;
               RECT 7.054 60.326 7.106 60.362 ;
               RECT 7.054 61.526 7.106 61.562 ;
               RECT 7.054 62.726 7.106 62.762 ;
               RECT 7.054 63.926 7.106 63.962 ;
               RECT 7.054 65.126 7.106 65.162 ;
               RECT 7.054 66.326 7.106 66.362 ;
               RECT 7.054 67.526 7.106 67.562 ;
               RECT 7.054 68.726 7.106 68.762 ;
               RECT 7.054 69.926 7.106 69.962 ;
               RECT 7.054 71.126 7.106 71.162 ;
               RECT 7.054 72.326 7.106 72.362 ;
               RECT 7.054 73.526 7.106 73.562 ;
               RECT 7.054 74.726 7.106 74.762 ;
               RECT 7.054 75.926 7.106 75.962 ;
               RECT 7.054 77.126 7.106 77.162 ;
               RECT 7.054 78.326 7.106 78.362 ;
               RECT 7.054 79.526 7.106 79.562 ;
               RECT 7.054 80.726 7.106 80.762 ;
               RECT 7.054 81.926 7.106 81.962 ;
               RECT 7.054 83.126 7.106 83.162 ;
               RECT 7.054 84.326 7.106 84.362 ;
               RECT 7.054 85.526 7.106 85.562 ;
               RECT 7.054 86.726 7.106 86.762 ;
               RECT 7.054 87.926 7.106 87.962 ;
               RECT 7.054 89.126 7.106 89.162 ;
               RECT 7.054 90.326 7.106 90.362 ;
               RECT 7.054 91.526 7.106 91.562 ;
               RECT 7.054 92.726 7.106 92.762 ;
               RECT 7.054 93.926 7.106 93.962 ;
               RECT 7.054 95.126 7.106 95.162 ;
               RECT 7.054 96.326 7.106 96.362 ;
               RECT 7.054 97.526 7.106 97.562 ;
               RECT 7.054 98.726 7.106 98.762 ;
               RECT 7.054 99.926 7.106 99.962 ;
               RECT 7.054 101.126 7.106 101.162 ;
               RECT 7.054 102.326 7.106 102.362 ;
               RECT 7.054 103.526 7.106 103.562 ;
               RECT 7.134 1.558 7.186 1.594 ;
               RECT 7.134 2.758 7.186 2.794 ;
               RECT 7.134 3.958 7.186 3.994 ;
               RECT 7.134 5.158 7.186 5.194 ;
               RECT 7.134 6.358 7.186 6.394 ;
               RECT 7.134 7.558 7.186 7.594 ;
               RECT 7.134 8.758 7.186 8.794 ;
               RECT 7.134 9.958 7.186 9.994 ;
               RECT 7.134 11.158 7.186 11.194 ;
               RECT 7.134 12.358 7.186 12.394 ;
               RECT 7.134 13.558 7.186 13.594 ;
               RECT 7.134 14.758 7.186 14.794 ;
               RECT 7.134 15.958 7.186 15.994 ;
               RECT 7.134 17.158 7.186 17.194 ;
               RECT 7.134 18.358 7.186 18.394 ;
               RECT 7.134 19.558 7.186 19.594 ;
               RECT 7.134 20.758 7.186 20.794 ;
               RECT 7.134 21.958 7.186 21.994 ;
               RECT 7.134 23.158 7.186 23.194 ;
               RECT 7.134 24.358 7.186 24.394 ;
               RECT 7.134 25.558 7.186 25.594 ;
               RECT 7.134 26.758 7.186 26.794 ;
               RECT 7.134 27.958 7.186 27.994 ;
               RECT 7.134 29.158 7.186 29.194 ;
               RECT 7.134 30.358 7.186 30.394 ;
               RECT 7.134 31.558 7.186 31.594 ;
               RECT 7.134 32.758 7.186 32.794 ;
               RECT 7.134 33.958 7.186 33.994 ;
               RECT 7.134 35.158 7.186 35.194 ;
               RECT 7.134 36.358 7.186 36.394 ;
               RECT 7.134 37.558 7.186 37.594 ;
               RECT 7.134 38.758 7.186 38.794 ;
               RECT 7.134 39.958 7.186 39.994 ;
               RECT 7.134 41.158 7.186 41.194 ;
               RECT 7.134 42.358 7.186 42.394 ;
               RECT 7.134 43.558 7.186 43.594 ;
               RECT 7.134 44.758 7.186 44.794 ;
               RECT 7.134 45.958 7.186 45.994 ;
               RECT 7.134 47.158 7.186 47.194 ;
               RECT 7.134 48.358 7.186 48.394 ;
               RECT 7.134 50.142 7.186 50.178 ;
               RECT 7.134 50.382 7.186 50.418 ;
               RECT 7.134 54.702 7.186 54.738 ;
               RECT 7.134 54.942 7.186 54.978 ;
               RECT 7.134 57.478 7.186 57.514 ;
               RECT 7.134 58.678 7.186 58.714 ;
               RECT 7.134 59.878 7.186 59.914 ;
               RECT 7.134 61.078 7.186 61.114 ;
               RECT 7.134 62.278 7.186 62.314 ;
               RECT 7.134 63.478 7.186 63.514 ;
               RECT 7.134 64.678 7.186 64.714 ;
               RECT 7.134 65.878 7.186 65.914 ;
               RECT 7.134 67.078 7.186 67.114 ;
               RECT 7.134 68.278 7.186 68.314 ;
               RECT 7.134 69.478 7.186 69.514 ;
               RECT 7.134 70.678 7.186 70.714 ;
               RECT 7.134 71.878 7.186 71.914 ;
               RECT 7.134 73.078 7.186 73.114 ;
               RECT 7.134 74.278 7.186 74.314 ;
               RECT 7.134 75.478 7.186 75.514 ;
               RECT 7.134 76.678 7.186 76.714 ;
               RECT 7.134 77.878 7.186 77.914 ;
               RECT 7.134 79.078 7.186 79.114 ;
               RECT 7.134 80.278 7.186 80.314 ;
               RECT 7.134 81.478 7.186 81.514 ;
               RECT 7.134 82.678 7.186 82.714 ;
               RECT 7.134 83.878 7.186 83.914 ;
               RECT 7.134 85.078 7.186 85.114 ;
               RECT 7.134 86.278 7.186 86.314 ;
               RECT 7.134 87.478 7.186 87.514 ;
               RECT 7.134 88.678 7.186 88.714 ;
               RECT 7.134 89.878 7.186 89.914 ;
               RECT 7.134 91.078 7.186 91.114 ;
               RECT 7.134 92.278 7.186 92.314 ;
               RECT 7.134 93.478 7.186 93.514 ;
               RECT 7.134 94.678 7.186 94.714 ;
               RECT 7.134 95.878 7.186 95.914 ;
               RECT 7.134 97.078 7.186 97.114 ;
               RECT 7.134 98.278 7.186 98.314 ;
               RECT 7.134 99.478 7.186 99.514 ;
               RECT 7.134 100.678 7.186 100.714 ;
               RECT 7.134 101.878 7.186 101.914 ;
               RECT 7.134 103.078 7.186 103.114 ;
               RECT 7.134 104.278 7.186 104.314 ;
               RECT 7.214 0.806 7.266 0.842 ;
               RECT 7.214 2.006 7.266 2.042 ;
               RECT 7.214 3.206 7.266 3.242 ;
               RECT 7.214 4.406 7.266 4.442 ;
               RECT 7.214 5.606 7.266 5.642 ;
               RECT 7.214 6.806 7.266 6.842 ;
               RECT 7.214 8.006 7.266 8.042 ;
               RECT 7.214 9.206 7.266 9.242 ;
               RECT 7.214 10.406 7.266 10.442 ;
               RECT 7.214 11.606 7.266 11.642 ;
               RECT 7.214 12.806 7.266 12.842 ;
               RECT 7.214 14.006 7.266 14.042 ;
               RECT 7.214 15.206 7.266 15.242 ;
               RECT 7.214 16.406 7.266 16.442 ;
               RECT 7.214 17.606 7.266 17.642 ;
               RECT 7.214 18.806 7.266 18.842 ;
               RECT 7.214 20.006 7.266 20.042 ;
               RECT 7.214 21.206 7.266 21.242 ;
               RECT 7.214 22.406 7.266 22.442 ;
               RECT 7.214 23.606 7.266 23.642 ;
               RECT 7.214 24.806 7.266 24.842 ;
               RECT 7.214 26.006 7.266 26.042 ;
               RECT 7.214 27.206 7.266 27.242 ;
               RECT 7.214 28.406 7.266 28.442 ;
               RECT 7.214 29.606 7.266 29.642 ;
               RECT 7.214 30.806 7.266 30.842 ;
               RECT 7.214 32.006 7.266 32.042 ;
               RECT 7.214 33.206 7.266 33.242 ;
               RECT 7.214 34.406 7.266 34.442 ;
               RECT 7.214 35.606 7.266 35.642 ;
               RECT 7.214 36.806 7.266 36.842 ;
               RECT 7.214 38.006 7.266 38.042 ;
               RECT 7.214 39.206 7.266 39.242 ;
               RECT 7.214 40.406 7.266 40.442 ;
               RECT 7.214 41.606 7.266 41.642 ;
               RECT 7.214 42.806 7.266 42.842 ;
               RECT 7.214 44.006 7.266 44.042 ;
               RECT 7.214 45.206 7.266 45.242 ;
               RECT 7.214 46.406 7.266 46.442 ;
               RECT 7.214 47.606 7.266 47.642 ;
               RECT 7.214 49.422 7.266 49.458 ;
               RECT 7.214 49.662 7.266 49.698 ;
               RECT 7.214 55.422 7.266 55.458 ;
               RECT 7.214 55.662 7.266 55.698 ;
               RECT 7.214 56.726 7.266 56.762 ;
               RECT 7.214 57.926 7.266 57.962 ;
               RECT 7.214 59.126 7.266 59.162 ;
               RECT 7.214 60.326 7.266 60.362 ;
               RECT 7.214 61.526 7.266 61.562 ;
               RECT 7.214 62.726 7.266 62.762 ;
               RECT 7.214 63.926 7.266 63.962 ;
               RECT 7.214 65.126 7.266 65.162 ;
               RECT 7.214 66.326 7.266 66.362 ;
               RECT 7.214 67.526 7.266 67.562 ;
               RECT 7.214 68.726 7.266 68.762 ;
               RECT 7.214 69.926 7.266 69.962 ;
               RECT 7.214 71.126 7.266 71.162 ;
               RECT 7.214 72.326 7.266 72.362 ;
               RECT 7.214 73.526 7.266 73.562 ;
               RECT 7.214 74.726 7.266 74.762 ;
               RECT 7.214 75.926 7.266 75.962 ;
               RECT 7.214 77.126 7.266 77.162 ;
               RECT 7.214 78.326 7.266 78.362 ;
               RECT 7.214 79.526 7.266 79.562 ;
               RECT 7.214 80.726 7.266 80.762 ;
               RECT 7.214 81.926 7.266 81.962 ;
               RECT 7.214 83.126 7.266 83.162 ;
               RECT 7.214 84.326 7.266 84.362 ;
               RECT 7.214 85.526 7.266 85.562 ;
               RECT 7.214 86.726 7.266 86.762 ;
               RECT 7.214 87.926 7.266 87.962 ;
               RECT 7.214 89.126 7.266 89.162 ;
               RECT 7.214 90.326 7.266 90.362 ;
               RECT 7.214 91.526 7.266 91.562 ;
               RECT 7.214 92.726 7.266 92.762 ;
               RECT 7.214 93.926 7.266 93.962 ;
               RECT 7.214 95.126 7.266 95.162 ;
               RECT 7.214 96.326 7.266 96.362 ;
               RECT 7.214 97.526 7.266 97.562 ;
               RECT 7.214 98.726 7.266 98.762 ;
               RECT 7.214 99.926 7.266 99.962 ;
               RECT 7.214 101.126 7.266 101.162 ;
               RECT 7.214 102.326 7.266 102.362 ;
               RECT 7.214 103.526 7.266 103.562 ;
               RECT 7.294 1.558 7.346 1.594 ;
               RECT 7.294 2.758 7.346 2.794 ;
               RECT 7.294 3.958 7.346 3.994 ;
               RECT 7.294 5.158 7.346 5.194 ;
               RECT 7.294 6.358 7.346 6.394 ;
               RECT 7.294 7.558 7.346 7.594 ;
               RECT 7.294 8.758 7.346 8.794 ;
               RECT 7.294 9.958 7.346 9.994 ;
               RECT 7.294 11.158 7.346 11.194 ;
               RECT 7.294 12.358 7.346 12.394 ;
               RECT 7.294 13.558 7.346 13.594 ;
               RECT 7.294 14.758 7.346 14.794 ;
               RECT 7.294 15.958 7.346 15.994 ;
               RECT 7.294 17.158 7.346 17.194 ;
               RECT 7.294 18.358 7.346 18.394 ;
               RECT 7.294 19.558 7.346 19.594 ;
               RECT 7.294 20.758 7.346 20.794 ;
               RECT 7.294 21.958 7.346 21.994 ;
               RECT 7.294 23.158 7.346 23.194 ;
               RECT 7.294 24.358 7.346 24.394 ;
               RECT 7.294 25.558 7.346 25.594 ;
               RECT 7.294 26.758 7.346 26.794 ;
               RECT 7.294 27.958 7.346 27.994 ;
               RECT 7.294 29.158 7.346 29.194 ;
               RECT 7.294 30.358 7.346 30.394 ;
               RECT 7.294 31.558 7.346 31.594 ;
               RECT 7.294 32.758 7.346 32.794 ;
               RECT 7.294 33.958 7.346 33.994 ;
               RECT 7.294 35.158 7.346 35.194 ;
               RECT 7.294 36.358 7.346 36.394 ;
               RECT 7.294 37.558 7.346 37.594 ;
               RECT 7.294 38.758 7.346 38.794 ;
               RECT 7.294 39.958 7.346 39.994 ;
               RECT 7.294 41.158 7.346 41.194 ;
               RECT 7.294 42.358 7.346 42.394 ;
               RECT 7.294 43.558 7.346 43.594 ;
               RECT 7.294 44.758 7.346 44.794 ;
               RECT 7.294 45.958 7.346 45.994 ;
               RECT 7.294 47.158 7.346 47.194 ;
               RECT 7.294 48.358 7.346 48.394 ;
               RECT 7.294 50.142 7.346 50.178 ;
               RECT 7.294 50.382 7.346 50.418 ;
               RECT 7.294 54.702 7.346 54.738 ;
               RECT 7.294 54.942 7.346 54.978 ;
               RECT 7.294 57.478 7.346 57.514 ;
               RECT 7.294 58.678 7.346 58.714 ;
               RECT 7.294 59.878 7.346 59.914 ;
               RECT 7.294 61.078 7.346 61.114 ;
               RECT 7.294 62.278 7.346 62.314 ;
               RECT 7.294 63.478 7.346 63.514 ;
               RECT 7.294 64.678 7.346 64.714 ;
               RECT 7.294 65.878 7.346 65.914 ;
               RECT 7.294 67.078 7.346 67.114 ;
               RECT 7.294 68.278 7.346 68.314 ;
               RECT 7.294 69.478 7.346 69.514 ;
               RECT 7.294 70.678 7.346 70.714 ;
               RECT 7.294 71.878 7.346 71.914 ;
               RECT 7.294 73.078 7.346 73.114 ;
               RECT 7.294 74.278 7.346 74.314 ;
               RECT 7.294 75.478 7.346 75.514 ;
               RECT 7.294 76.678 7.346 76.714 ;
               RECT 7.294 77.878 7.346 77.914 ;
               RECT 7.294 79.078 7.346 79.114 ;
               RECT 7.294 80.278 7.346 80.314 ;
               RECT 7.294 81.478 7.346 81.514 ;
               RECT 7.294 82.678 7.346 82.714 ;
               RECT 7.294 83.878 7.346 83.914 ;
               RECT 7.294 85.078 7.346 85.114 ;
               RECT 7.294 86.278 7.346 86.314 ;
               RECT 7.294 87.478 7.346 87.514 ;
               RECT 7.294 88.678 7.346 88.714 ;
               RECT 7.294 89.878 7.346 89.914 ;
               RECT 7.294 91.078 7.346 91.114 ;
               RECT 7.294 92.278 7.346 92.314 ;
               RECT 7.294 93.478 7.346 93.514 ;
               RECT 7.294 94.678 7.346 94.714 ;
               RECT 7.294 95.878 7.346 95.914 ;
               RECT 7.294 97.078 7.346 97.114 ;
               RECT 7.294 98.278 7.346 98.314 ;
               RECT 7.294 99.478 7.346 99.514 ;
               RECT 7.294 100.678 7.346 100.714 ;
               RECT 7.294 101.878 7.346 101.914 ;
               RECT 7.294 103.078 7.346 103.114 ;
               RECT 7.294 104.278 7.346 104.314 ;
               RECT 7.374 0.281 7.426 0.317 ;
               RECT 7.374 104.803 7.426 104.839 ;
               RECT 7.454 0.806 7.506 0.842 ;
               RECT 7.454 2.006 7.506 2.042 ;
               RECT 7.454 3.206 7.506 3.242 ;
               RECT 7.454 4.406 7.506 4.442 ;
               RECT 7.454 5.606 7.506 5.642 ;
               RECT 7.454 6.806 7.506 6.842 ;
               RECT 7.454 8.006 7.506 8.042 ;
               RECT 7.454 9.206 7.506 9.242 ;
               RECT 7.454 10.406 7.506 10.442 ;
               RECT 7.454 11.606 7.506 11.642 ;
               RECT 7.454 12.806 7.506 12.842 ;
               RECT 7.454 14.006 7.506 14.042 ;
               RECT 7.454 15.206 7.506 15.242 ;
               RECT 7.454 16.406 7.506 16.442 ;
               RECT 7.454 17.606 7.506 17.642 ;
               RECT 7.454 18.806 7.506 18.842 ;
               RECT 7.454 20.006 7.506 20.042 ;
               RECT 7.454 21.206 7.506 21.242 ;
               RECT 7.454 22.406 7.506 22.442 ;
               RECT 7.454 23.606 7.506 23.642 ;
               RECT 7.454 24.806 7.506 24.842 ;
               RECT 7.454 26.006 7.506 26.042 ;
               RECT 7.454 27.206 7.506 27.242 ;
               RECT 7.454 28.406 7.506 28.442 ;
               RECT 7.454 29.606 7.506 29.642 ;
               RECT 7.454 30.806 7.506 30.842 ;
               RECT 7.454 32.006 7.506 32.042 ;
               RECT 7.454 33.206 7.506 33.242 ;
               RECT 7.454 34.406 7.506 34.442 ;
               RECT 7.454 35.606 7.506 35.642 ;
               RECT 7.454 36.806 7.506 36.842 ;
               RECT 7.454 38.006 7.506 38.042 ;
               RECT 7.454 39.206 7.506 39.242 ;
               RECT 7.454 40.406 7.506 40.442 ;
               RECT 7.454 41.606 7.506 41.642 ;
               RECT 7.454 42.806 7.506 42.842 ;
               RECT 7.454 44.006 7.506 44.042 ;
               RECT 7.454 45.206 7.506 45.242 ;
               RECT 7.454 46.406 7.506 46.442 ;
               RECT 7.454 47.606 7.506 47.642 ;
               RECT 7.454 49.422 7.506 49.458 ;
               RECT 7.454 49.662 7.506 49.698 ;
               RECT 7.454 51.102 7.506 51.138 ;
               RECT 7.454 51.582 7.506 51.618 ;
               RECT 7.454 53.502 7.506 53.538 ;
               RECT 7.454 53.982 7.506 54.018 ;
               RECT 7.454 55.422 7.506 55.458 ;
               RECT 7.454 55.662 7.506 55.698 ;
               RECT 7.454 56.726 7.506 56.762 ;
               RECT 7.454 57.926 7.506 57.962 ;
               RECT 7.454 59.126 7.506 59.162 ;
               RECT 7.454 60.326 7.506 60.362 ;
               RECT 7.454 61.526 7.506 61.562 ;
               RECT 7.454 62.726 7.506 62.762 ;
               RECT 7.454 63.926 7.506 63.962 ;
               RECT 7.454 65.126 7.506 65.162 ;
               RECT 7.454 66.326 7.506 66.362 ;
               RECT 7.454 67.526 7.506 67.562 ;
               RECT 7.454 68.726 7.506 68.762 ;
               RECT 7.454 69.926 7.506 69.962 ;
               RECT 7.454 71.126 7.506 71.162 ;
               RECT 7.454 72.326 7.506 72.362 ;
               RECT 7.454 73.526 7.506 73.562 ;
               RECT 7.454 74.726 7.506 74.762 ;
               RECT 7.454 75.926 7.506 75.962 ;
               RECT 7.454 77.126 7.506 77.162 ;
               RECT 7.454 78.326 7.506 78.362 ;
               RECT 7.454 79.526 7.506 79.562 ;
               RECT 7.454 80.726 7.506 80.762 ;
               RECT 7.454 81.926 7.506 81.962 ;
               RECT 7.454 83.126 7.506 83.162 ;
               RECT 7.454 84.326 7.506 84.362 ;
               RECT 7.454 85.526 7.506 85.562 ;
               RECT 7.454 86.726 7.506 86.762 ;
               RECT 7.454 87.926 7.506 87.962 ;
               RECT 7.454 89.126 7.506 89.162 ;
               RECT 7.454 90.326 7.506 90.362 ;
               RECT 7.454 91.526 7.506 91.562 ;
               RECT 7.454 92.726 7.506 92.762 ;
               RECT 7.454 93.926 7.506 93.962 ;
               RECT 7.454 95.126 7.506 95.162 ;
               RECT 7.454 96.326 7.506 96.362 ;
               RECT 7.454 97.526 7.506 97.562 ;
               RECT 7.454 98.726 7.506 98.762 ;
               RECT 7.454 99.926 7.506 99.962 ;
               RECT 7.454 101.126 7.506 101.162 ;
               RECT 7.454 102.326 7.506 102.362 ;
               RECT 7.454 103.526 7.506 103.562 ;
               RECT 7.534 1.558 7.586 1.594 ;
               RECT 7.534 2.758 7.586 2.794 ;
               RECT 7.534 3.958 7.586 3.994 ;
               RECT 7.534 5.158 7.586 5.194 ;
               RECT 7.534 6.358 7.586 6.394 ;
               RECT 7.534 7.558 7.586 7.594 ;
               RECT 7.534 8.758 7.586 8.794 ;
               RECT 7.534 9.958 7.586 9.994 ;
               RECT 7.534 11.158 7.586 11.194 ;
               RECT 7.534 12.358 7.586 12.394 ;
               RECT 7.534 13.558 7.586 13.594 ;
               RECT 7.534 14.758 7.586 14.794 ;
               RECT 7.534 15.958 7.586 15.994 ;
               RECT 7.534 17.158 7.586 17.194 ;
               RECT 7.534 18.358 7.586 18.394 ;
               RECT 7.534 19.558 7.586 19.594 ;
               RECT 7.534 20.758 7.586 20.794 ;
               RECT 7.534 21.958 7.586 21.994 ;
               RECT 7.534 23.158 7.586 23.194 ;
               RECT 7.534 24.358 7.586 24.394 ;
               RECT 7.534 25.558 7.586 25.594 ;
               RECT 7.534 26.758 7.586 26.794 ;
               RECT 7.534 27.958 7.586 27.994 ;
               RECT 7.534 29.158 7.586 29.194 ;
               RECT 7.534 30.358 7.586 30.394 ;
               RECT 7.534 31.558 7.586 31.594 ;
               RECT 7.534 32.758 7.586 32.794 ;
               RECT 7.534 33.958 7.586 33.994 ;
               RECT 7.534 35.158 7.586 35.194 ;
               RECT 7.534 36.358 7.586 36.394 ;
               RECT 7.534 37.558 7.586 37.594 ;
               RECT 7.534 38.758 7.586 38.794 ;
               RECT 7.534 39.958 7.586 39.994 ;
               RECT 7.534 41.158 7.586 41.194 ;
               RECT 7.534 42.358 7.586 42.394 ;
               RECT 7.534 43.558 7.586 43.594 ;
               RECT 7.534 44.758 7.586 44.794 ;
               RECT 7.534 45.958 7.586 45.994 ;
               RECT 7.534 47.158 7.586 47.194 ;
               RECT 7.534 48.358 7.586 48.394 ;
               RECT 7.534 50.142 7.586 50.178 ;
               RECT 7.534 50.382 7.586 50.418 ;
               RECT 7.534 54.702 7.586 54.738 ;
               RECT 7.534 54.942 7.586 54.978 ;
               RECT 7.534 57.478 7.586 57.514 ;
               RECT 7.534 58.678 7.586 58.714 ;
               RECT 7.534 59.878 7.586 59.914 ;
               RECT 7.534 61.078 7.586 61.114 ;
               RECT 7.534 62.278 7.586 62.314 ;
               RECT 7.534 63.478 7.586 63.514 ;
               RECT 7.534 64.678 7.586 64.714 ;
               RECT 7.534 65.878 7.586 65.914 ;
               RECT 7.534 67.078 7.586 67.114 ;
               RECT 7.534 68.278 7.586 68.314 ;
               RECT 7.534 69.478 7.586 69.514 ;
               RECT 7.534 70.678 7.586 70.714 ;
               RECT 7.534 71.878 7.586 71.914 ;
               RECT 7.534 73.078 7.586 73.114 ;
               RECT 7.534 74.278 7.586 74.314 ;
               RECT 7.534 75.478 7.586 75.514 ;
               RECT 7.534 76.678 7.586 76.714 ;
               RECT 7.534 77.878 7.586 77.914 ;
               RECT 7.534 79.078 7.586 79.114 ;
               RECT 7.534 80.278 7.586 80.314 ;
               RECT 7.534 81.478 7.586 81.514 ;
               RECT 7.534 82.678 7.586 82.714 ;
               RECT 7.534 83.878 7.586 83.914 ;
               RECT 7.534 85.078 7.586 85.114 ;
               RECT 7.534 86.278 7.586 86.314 ;
               RECT 7.534 87.478 7.586 87.514 ;
               RECT 7.534 88.678 7.586 88.714 ;
               RECT 7.534 89.878 7.586 89.914 ;
               RECT 7.534 91.078 7.586 91.114 ;
               RECT 7.534 92.278 7.586 92.314 ;
               RECT 7.534 93.478 7.586 93.514 ;
               RECT 7.534 94.678 7.586 94.714 ;
               RECT 7.534 95.878 7.586 95.914 ;
               RECT 7.534 97.078 7.586 97.114 ;
               RECT 7.534 98.278 7.586 98.314 ;
               RECT 7.534 99.478 7.586 99.514 ;
               RECT 7.534 100.678 7.586 100.714 ;
               RECT 7.534 101.878 7.586 101.914 ;
               RECT 7.534 103.078 7.586 103.114 ;
               RECT 7.534 104.278 7.586 104.314 ;
               RECT 7.614 0.806 7.666 0.842 ;
               RECT 7.614 2.006 7.666 2.042 ;
               RECT 7.614 3.206 7.666 3.242 ;
               RECT 7.614 4.406 7.666 4.442 ;
               RECT 7.614 5.606 7.666 5.642 ;
               RECT 7.614 6.806 7.666 6.842 ;
               RECT 7.614 8.006 7.666 8.042 ;
               RECT 7.614 9.206 7.666 9.242 ;
               RECT 7.614 10.406 7.666 10.442 ;
               RECT 7.614 11.606 7.666 11.642 ;
               RECT 7.614 12.806 7.666 12.842 ;
               RECT 7.614 14.006 7.666 14.042 ;
               RECT 7.614 15.206 7.666 15.242 ;
               RECT 7.614 16.406 7.666 16.442 ;
               RECT 7.614 17.606 7.666 17.642 ;
               RECT 7.614 18.806 7.666 18.842 ;
               RECT 7.614 20.006 7.666 20.042 ;
               RECT 7.614 21.206 7.666 21.242 ;
               RECT 7.614 22.406 7.666 22.442 ;
               RECT 7.614 23.606 7.666 23.642 ;
               RECT 7.614 24.806 7.666 24.842 ;
               RECT 7.614 26.006 7.666 26.042 ;
               RECT 7.614 27.206 7.666 27.242 ;
               RECT 7.614 28.406 7.666 28.442 ;
               RECT 7.614 29.606 7.666 29.642 ;
               RECT 7.614 30.806 7.666 30.842 ;
               RECT 7.614 32.006 7.666 32.042 ;
               RECT 7.614 33.206 7.666 33.242 ;
               RECT 7.614 34.406 7.666 34.442 ;
               RECT 7.614 35.606 7.666 35.642 ;
               RECT 7.614 36.806 7.666 36.842 ;
               RECT 7.614 38.006 7.666 38.042 ;
               RECT 7.614 39.206 7.666 39.242 ;
               RECT 7.614 40.406 7.666 40.442 ;
               RECT 7.614 41.606 7.666 41.642 ;
               RECT 7.614 42.806 7.666 42.842 ;
               RECT 7.614 44.006 7.666 44.042 ;
               RECT 7.614 45.206 7.666 45.242 ;
               RECT 7.614 46.406 7.666 46.442 ;
               RECT 7.614 47.606 7.666 47.642 ;
               RECT 7.614 49.422 7.666 49.458 ;
               RECT 7.614 49.662 7.666 49.698 ;
               RECT 7.614 55.422 7.666 55.458 ;
               RECT 7.614 55.662 7.666 55.698 ;
               RECT 7.614 56.726 7.666 56.762 ;
               RECT 7.614 57.926 7.666 57.962 ;
               RECT 7.614 59.126 7.666 59.162 ;
               RECT 7.614 60.326 7.666 60.362 ;
               RECT 7.614 61.526 7.666 61.562 ;
               RECT 7.614 62.726 7.666 62.762 ;
               RECT 7.614 63.926 7.666 63.962 ;
               RECT 7.614 65.126 7.666 65.162 ;
               RECT 7.614 66.326 7.666 66.362 ;
               RECT 7.614 67.526 7.666 67.562 ;
               RECT 7.614 68.726 7.666 68.762 ;
               RECT 7.614 69.926 7.666 69.962 ;
               RECT 7.614 71.126 7.666 71.162 ;
               RECT 7.614 72.326 7.666 72.362 ;
               RECT 7.614 73.526 7.666 73.562 ;
               RECT 7.614 74.726 7.666 74.762 ;
               RECT 7.614 75.926 7.666 75.962 ;
               RECT 7.614 77.126 7.666 77.162 ;
               RECT 7.614 78.326 7.666 78.362 ;
               RECT 7.614 79.526 7.666 79.562 ;
               RECT 7.614 80.726 7.666 80.762 ;
               RECT 7.614 81.926 7.666 81.962 ;
               RECT 7.614 83.126 7.666 83.162 ;
               RECT 7.614 84.326 7.666 84.362 ;
               RECT 7.614 85.526 7.666 85.562 ;
               RECT 7.614 86.726 7.666 86.762 ;
               RECT 7.614 87.926 7.666 87.962 ;
               RECT 7.614 89.126 7.666 89.162 ;
               RECT 7.614 90.326 7.666 90.362 ;
               RECT 7.614 91.526 7.666 91.562 ;
               RECT 7.614 92.726 7.666 92.762 ;
               RECT 7.614 93.926 7.666 93.962 ;
               RECT 7.614 95.126 7.666 95.162 ;
               RECT 7.614 96.326 7.666 96.362 ;
               RECT 7.614 97.526 7.666 97.562 ;
               RECT 7.614 98.726 7.666 98.762 ;
               RECT 7.614 99.926 7.666 99.962 ;
               RECT 7.614 101.126 7.666 101.162 ;
               RECT 7.614 102.326 7.666 102.362 ;
               RECT 7.614 103.526 7.666 103.562 ;
               RECT 7.694 1.558 7.746 1.594 ;
               RECT 7.694 2.758 7.746 2.794 ;
               RECT 7.694 3.958 7.746 3.994 ;
               RECT 7.694 5.158 7.746 5.194 ;
               RECT 7.694 6.358 7.746 6.394 ;
               RECT 7.694 7.558 7.746 7.594 ;
               RECT 7.694 8.758 7.746 8.794 ;
               RECT 7.694 9.958 7.746 9.994 ;
               RECT 7.694 11.158 7.746 11.194 ;
               RECT 7.694 12.358 7.746 12.394 ;
               RECT 7.694 13.558 7.746 13.594 ;
               RECT 7.694 14.758 7.746 14.794 ;
               RECT 7.694 15.958 7.746 15.994 ;
               RECT 7.694 17.158 7.746 17.194 ;
               RECT 7.694 18.358 7.746 18.394 ;
               RECT 7.694 19.558 7.746 19.594 ;
               RECT 7.694 20.758 7.746 20.794 ;
               RECT 7.694 21.958 7.746 21.994 ;
               RECT 7.694 23.158 7.746 23.194 ;
               RECT 7.694 24.358 7.746 24.394 ;
               RECT 7.694 25.558 7.746 25.594 ;
               RECT 7.694 26.758 7.746 26.794 ;
               RECT 7.694 27.958 7.746 27.994 ;
               RECT 7.694 29.158 7.746 29.194 ;
               RECT 7.694 30.358 7.746 30.394 ;
               RECT 7.694 31.558 7.746 31.594 ;
               RECT 7.694 32.758 7.746 32.794 ;
               RECT 7.694 33.958 7.746 33.994 ;
               RECT 7.694 35.158 7.746 35.194 ;
               RECT 7.694 36.358 7.746 36.394 ;
               RECT 7.694 37.558 7.746 37.594 ;
               RECT 7.694 38.758 7.746 38.794 ;
               RECT 7.694 39.958 7.746 39.994 ;
               RECT 7.694 41.158 7.746 41.194 ;
               RECT 7.694 42.358 7.746 42.394 ;
               RECT 7.694 43.558 7.746 43.594 ;
               RECT 7.694 44.758 7.746 44.794 ;
               RECT 7.694 45.958 7.746 45.994 ;
               RECT 7.694 47.158 7.746 47.194 ;
               RECT 7.694 48.358 7.746 48.394 ;
               RECT 7.694 50.142 7.746 50.178 ;
               RECT 7.694 50.382 7.746 50.418 ;
               RECT 7.694 54.702 7.746 54.738 ;
               RECT 7.694 54.942 7.746 54.978 ;
               RECT 7.694 57.478 7.746 57.514 ;
               RECT 7.694 58.678 7.746 58.714 ;
               RECT 7.694 59.878 7.746 59.914 ;
               RECT 7.694 61.078 7.746 61.114 ;
               RECT 7.694 62.278 7.746 62.314 ;
               RECT 7.694 63.478 7.746 63.514 ;
               RECT 7.694 64.678 7.746 64.714 ;
               RECT 7.694 65.878 7.746 65.914 ;
               RECT 7.694 67.078 7.746 67.114 ;
               RECT 7.694 68.278 7.746 68.314 ;
               RECT 7.694 69.478 7.746 69.514 ;
               RECT 7.694 70.678 7.746 70.714 ;
               RECT 7.694 71.878 7.746 71.914 ;
               RECT 7.694 73.078 7.746 73.114 ;
               RECT 7.694 74.278 7.746 74.314 ;
               RECT 7.694 75.478 7.746 75.514 ;
               RECT 7.694 76.678 7.746 76.714 ;
               RECT 7.694 77.878 7.746 77.914 ;
               RECT 7.694 79.078 7.746 79.114 ;
               RECT 7.694 80.278 7.746 80.314 ;
               RECT 7.694 81.478 7.746 81.514 ;
               RECT 7.694 82.678 7.746 82.714 ;
               RECT 7.694 83.878 7.746 83.914 ;
               RECT 7.694 85.078 7.746 85.114 ;
               RECT 7.694 86.278 7.746 86.314 ;
               RECT 7.694 87.478 7.746 87.514 ;
               RECT 7.694 88.678 7.746 88.714 ;
               RECT 7.694 89.878 7.746 89.914 ;
               RECT 7.694 91.078 7.746 91.114 ;
               RECT 7.694 92.278 7.746 92.314 ;
               RECT 7.694 93.478 7.746 93.514 ;
               RECT 7.694 94.678 7.746 94.714 ;
               RECT 7.694 95.878 7.746 95.914 ;
               RECT 7.694 97.078 7.746 97.114 ;
               RECT 7.694 98.278 7.746 98.314 ;
               RECT 7.694 99.478 7.746 99.514 ;
               RECT 7.694 100.678 7.746 100.714 ;
               RECT 7.694 101.878 7.746 101.914 ;
               RECT 7.694 103.078 7.746 103.114 ;
               RECT 7.694 104.278 7.746 104.314 ;
               RECT 7.774 0.281 7.826 0.317 ;
               RECT 7.774 104.803 7.826 104.839 ;
               RECT 7.854 0.806 7.906 0.842 ;
               RECT 7.854 2.006 7.906 2.042 ;
               RECT 7.854 3.206 7.906 3.242 ;
               RECT 7.854 4.406 7.906 4.442 ;
               RECT 7.854 5.606 7.906 5.642 ;
               RECT 7.854 6.806 7.906 6.842 ;
               RECT 7.854 8.006 7.906 8.042 ;
               RECT 7.854 9.206 7.906 9.242 ;
               RECT 7.854 10.406 7.906 10.442 ;
               RECT 7.854 11.606 7.906 11.642 ;
               RECT 7.854 12.806 7.906 12.842 ;
               RECT 7.854 14.006 7.906 14.042 ;
               RECT 7.854 15.206 7.906 15.242 ;
               RECT 7.854 16.406 7.906 16.442 ;
               RECT 7.854 17.606 7.906 17.642 ;
               RECT 7.854 18.806 7.906 18.842 ;
               RECT 7.854 20.006 7.906 20.042 ;
               RECT 7.854 21.206 7.906 21.242 ;
               RECT 7.854 22.406 7.906 22.442 ;
               RECT 7.854 23.606 7.906 23.642 ;
               RECT 7.854 24.806 7.906 24.842 ;
               RECT 7.854 26.006 7.906 26.042 ;
               RECT 7.854 27.206 7.906 27.242 ;
               RECT 7.854 28.406 7.906 28.442 ;
               RECT 7.854 29.606 7.906 29.642 ;
               RECT 7.854 30.806 7.906 30.842 ;
               RECT 7.854 32.006 7.906 32.042 ;
               RECT 7.854 33.206 7.906 33.242 ;
               RECT 7.854 34.406 7.906 34.442 ;
               RECT 7.854 35.606 7.906 35.642 ;
               RECT 7.854 36.806 7.906 36.842 ;
               RECT 7.854 38.006 7.906 38.042 ;
               RECT 7.854 39.206 7.906 39.242 ;
               RECT 7.854 40.406 7.906 40.442 ;
               RECT 7.854 41.606 7.906 41.642 ;
               RECT 7.854 42.806 7.906 42.842 ;
               RECT 7.854 44.006 7.906 44.042 ;
               RECT 7.854 45.206 7.906 45.242 ;
               RECT 7.854 46.406 7.906 46.442 ;
               RECT 7.854 47.606 7.906 47.642 ;
               RECT 7.854 49.422 7.906 49.458 ;
               RECT 7.854 49.662 7.906 49.698 ;
               RECT 7.854 55.422 7.906 55.458 ;
               RECT 7.854 55.662 7.906 55.698 ;
               RECT 7.854 56.726 7.906 56.762 ;
               RECT 7.854 57.926 7.906 57.962 ;
               RECT 7.854 59.126 7.906 59.162 ;
               RECT 7.854 60.326 7.906 60.362 ;
               RECT 7.854 61.526 7.906 61.562 ;
               RECT 7.854 62.726 7.906 62.762 ;
               RECT 7.854 63.926 7.906 63.962 ;
               RECT 7.854 65.126 7.906 65.162 ;
               RECT 7.854 66.326 7.906 66.362 ;
               RECT 7.854 67.526 7.906 67.562 ;
               RECT 7.854 68.726 7.906 68.762 ;
               RECT 7.854 69.926 7.906 69.962 ;
               RECT 7.854 71.126 7.906 71.162 ;
               RECT 7.854 72.326 7.906 72.362 ;
               RECT 7.854 73.526 7.906 73.562 ;
               RECT 7.854 74.726 7.906 74.762 ;
               RECT 7.854 75.926 7.906 75.962 ;
               RECT 7.854 77.126 7.906 77.162 ;
               RECT 7.854 78.326 7.906 78.362 ;
               RECT 7.854 79.526 7.906 79.562 ;
               RECT 7.854 80.726 7.906 80.762 ;
               RECT 7.854 81.926 7.906 81.962 ;
               RECT 7.854 83.126 7.906 83.162 ;
               RECT 7.854 84.326 7.906 84.362 ;
               RECT 7.854 85.526 7.906 85.562 ;
               RECT 7.854 86.726 7.906 86.762 ;
               RECT 7.854 87.926 7.906 87.962 ;
               RECT 7.854 89.126 7.906 89.162 ;
               RECT 7.854 90.326 7.906 90.362 ;
               RECT 7.854 91.526 7.906 91.562 ;
               RECT 7.854 92.726 7.906 92.762 ;
               RECT 7.854 93.926 7.906 93.962 ;
               RECT 7.854 95.126 7.906 95.162 ;
               RECT 7.854 96.326 7.906 96.362 ;
               RECT 7.854 97.526 7.906 97.562 ;
               RECT 7.854 98.726 7.906 98.762 ;
               RECT 7.854 99.926 7.906 99.962 ;
               RECT 7.854 101.126 7.906 101.162 ;
               RECT 7.854 102.326 7.906 102.362 ;
               RECT 7.854 103.526 7.906 103.562 ;
               RECT 7.934 1.558 7.986 1.594 ;
               RECT 7.934 2.758 7.986 2.794 ;
               RECT 7.934 3.958 7.986 3.994 ;
               RECT 7.934 5.158 7.986 5.194 ;
               RECT 7.934 6.358 7.986 6.394 ;
               RECT 7.934 7.558 7.986 7.594 ;
               RECT 7.934 8.758 7.986 8.794 ;
               RECT 7.934 9.958 7.986 9.994 ;
               RECT 7.934 11.158 7.986 11.194 ;
               RECT 7.934 12.358 7.986 12.394 ;
               RECT 7.934 13.558 7.986 13.594 ;
               RECT 7.934 14.758 7.986 14.794 ;
               RECT 7.934 15.958 7.986 15.994 ;
               RECT 7.934 17.158 7.986 17.194 ;
               RECT 7.934 18.358 7.986 18.394 ;
               RECT 7.934 19.558 7.986 19.594 ;
               RECT 7.934 20.758 7.986 20.794 ;
               RECT 7.934 21.958 7.986 21.994 ;
               RECT 7.934 23.158 7.986 23.194 ;
               RECT 7.934 24.358 7.986 24.394 ;
               RECT 7.934 25.558 7.986 25.594 ;
               RECT 7.934 26.758 7.986 26.794 ;
               RECT 7.934 27.958 7.986 27.994 ;
               RECT 7.934 29.158 7.986 29.194 ;
               RECT 7.934 30.358 7.986 30.394 ;
               RECT 7.934 31.558 7.986 31.594 ;
               RECT 7.934 32.758 7.986 32.794 ;
               RECT 7.934 33.958 7.986 33.994 ;
               RECT 7.934 35.158 7.986 35.194 ;
               RECT 7.934 36.358 7.986 36.394 ;
               RECT 7.934 37.558 7.986 37.594 ;
               RECT 7.934 38.758 7.986 38.794 ;
               RECT 7.934 39.958 7.986 39.994 ;
               RECT 7.934 41.158 7.986 41.194 ;
               RECT 7.934 42.358 7.986 42.394 ;
               RECT 7.934 43.558 7.986 43.594 ;
               RECT 7.934 44.758 7.986 44.794 ;
               RECT 7.934 45.958 7.986 45.994 ;
               RECT 7.934 47.158 7.986 47.194 ;
               RECT 7.934 48.358 7.986 48.394 ;
               RECT 7.934 50.142 7.986 50.178 ;
               RECT 7.934 50.382 7.986 50.418 ;
               RECT 7.934 54.702 7.986 54.738 ;
               RECT 7.934 54.942 7.986 54.978 ;
               RECT 7.934 57.478 7.986 57.514 ;
               RECT 7.934 58.678 7.986 58.714 ;
               RECT 7.934 59.878 7.986 59.914 ;
               RECT 7.934 61.078 7.986 61.114 ;
               RECT 7.934 62.278 7.986 62.314 ;
               RECT 7.934 63.478 7.986 63.514 ;
               RECT 7.934 64.678 7.986 64.714 ;
               RECT 7.934 65.878 7.986 65.914 ;
               RECT 7.934 67.078 7.986 67.114 ;
               RECT 7.934 68.278 7.986 68.314 ;
               RECT 7.934 69.478 7.986 69.514 ;
               RECT 7.934 70.678 7.986 70.714 ;
               RECT 7.934 71.878 7.986 71.914 ;
               RECT 7.934 73.078 7.986 73.114 ;
               RECT 7.934 74.278 7.986 74.314 ;
               RECT 7.934 75.478 7.986 75.514 ;
               RECT 7.934 76.678 7.986 76.714 ;
               RECT 7.934 77.878 7.986 77.914 ;
               RECT 7.934 79.078 7.986 79.114 ;
               RECT 7.934 80.278 7.986 80.314 ;
               RECT 7.934 81.478 7.986 81.514 ;
               RECT 7.934 82.678 7.986 82.714 ;
               RECT 7.934 83.878 7.986 83.914 ;
               RECT 7.934 85.078 7.986 85.114 ;
               RECT 7.934 86.278 7.986 86.314 ;
               RECT 7.934 87.478 7.986 87.514 ;
               RECT 7.934 88.678 7.986 88.714 ;
               RECT 7.934 89.878 7.986 89.914 ;
               RECT 7.934 91.078 7.986 91.114 ;
               RECT 7.934 92.278 7.986 92.314 ;
               RECT 7.934 93.478 7.986 93.514 ;
               RECT 7.934 94.678 7.986 94.714 ;
               RECT 7.934 95.878 7.986 95.914 ;
               RECT 7.934 97.078 7.986 97.114 ;
               RECT 7.934 98.278 7.986 98.314 ;
               RECT 7.934 99.478 7.986 99.514 ;
               RECT 7.934 100.678 7.986 100.714 ;
               RECT 7.934 101.878 7.986 101.914 ;
               RECT 7.934 103.078 7.986 103.114 ;
               RECT 7.934 104.278 7.986 104.314 ;
               RECT 8.014 0.806 8.066 0.842 ;
               RECT 8.014 2.006 8.066 2.042 ;
               RECT 8.014 3.206 8.066 3.242 ;
               RECT 8.014 4.406 8.066 4.442 ;
               RECT 8.014 5.606 8.066 5.642 ;
               RECT 8.014 6.806 8.066 6.842 ;
               RECT 8.014 8.006 8.066 8.042 ;
               RECT 8.014 9.206 8.066 9.242 ;
               RECT 8.014 10.406 8.066 10.442 ;
               RECT 8.014 11.606 8.066 11.642 ;
               RECT 8.014 12.806 8.066 12.842 ;
               RECT 8.014 14.006 8.066 14.042 ;
               RECT 8.014 15.206 8.066 15.242 ;
               RECT 8.014 16.406 8.066 16.442 ;
               RECT 8.014 17.606 8.066 17.642 ;
               RECT 8.014 18.806 8.066 18.842 ;
               RECT 8.014 20.006 8.066 20.042 ;
               RECT 8.014 21.206 8.066 21.242 ;
               RECT 8.014 22.406 8.066 22.442 ;
               RECT 8.014 23.606 8.066 23.642 ;
               RECT 8.014 24.806 8.066 24.842 ;
               RECT 8.014 26.006 8.066 26.042 ;
               RECT 8.014 27.206 8.066 27.242 ;
               RECT 8.014 28.406 8.066 28.442 ;
               RECT 8.014 29.606 8.066 29.642 ;
               RECT 8.014 30.806 8.066 30.842 ;
               RECT 8.014 32.006 8.066 32.042 ;
               RECT 8.014 33.206 8.066 33.242 ;
               RECT 8.014 34.406 8.066 34.442 ;
               RECT 8.014 35.606 8.066 35.642 ;
               RECT 8.014 36.806 8.066 36.842 ;
               RECT 8.014 38.006 8.066 38.042 ;
               RECT 8.014 39.206 8.066 39.242 ;
               RECT 8.014 40.406 8.066 40.442 ;
               RECT 8.014 41.606 8.066 41.642 ;
               RECT 8.014 42.806 8.066 42.842 ;
               RECT 8.014 44.006 8.066 44.042 ;
               RECT 8.014 45.206 8.066 45.242 ;
               RECT 8.014 46.406 8.066 46.442 ;
               RECT 8.014 47.606 8.066 47.642 ;
               RECT 8.014 49.422 8.066 49.458 ;
               RECT 8.014 49.662 8.066 49.698 ;
               RECT 8.014 55.422 8.066 55.458 ;
               RECT 8.014 55.662 8.066 55.698 ;
               RECT 8.014 56.726 8.066 56.762 ;
               RECT 8.014 57.926 8.066 57.962 ;
               RECT 8.014 59.126 8.066 59.162 ;
               RECT 8.014 60.326 8.066 60.362 ;
               RECT 8.014 61.526 8.066 61.562 ;
               RECT 8.014 62.726 8.066 62.762 ;
               RECT 8.014 63.926 8.066 63.962 ;
               RECT 8.014 65.126 8.066 65.162 ;
               RECT 8.014 66.326 8.066 66.362 ;
               RECT 8.014 67.526 8.066 67.562 ;
               RECT 8.014 68.726 8.066 68.762 ;
               RECT 8.014 69.926 8.066 69.962 ;
               RECT 8.014 71.126 8.066 71.162 ;
               RECT 8.014 72.326 8.066 72.362 ;
               RECT 8.014 73.526 8.066 73.562 ;
               RECT 8.014 74.726 8.066 74.762 ;
               RECT 8.014 75.926 8.066 75.962 ;
               RECT 8.014 77.126 8.066 77.162 ;
               RECT 8.014 78.326 8.066 78.362 ;
               RECT 8.014 79.526 8.066 79.562 ;
               RECT 8.014 80.726 8.066 80.762 ;
               RECT 8.014 81.926 8.066 81.962 ;
               RECT 8.014 83.126 8.066 83.162 ;
               RECT 8.014 84.326 8.066 84.362 ;
               RECT 8.014 85.526 8.066 85.562 ;
               RECT 8.014 86.726 8.066 86.762 ;
               RECT 8.014 87.926 8.066 87.962 ;
               RECT 8.014 89.126 8.066 89.162 ;
               RECT 8.014 90.326 8.066 90.362 ;
               RECT 8.014 91.526 8.066 91.562 ;
               RECT 8.014 92.726 8.066 92.762 ;
               RECT 8.014 93.926 8.066 93.962 ;
               RECT 8.014 95.126 8.066 95.162 ;
               RECT 8.014 96.326 8.066 96.362 ;
               RECT 8.014 97.526 8.066 97.562 ;
               RECT 8.014 98.726 8.066 98.762 ;
               RECT 8.014 99.926 8.066 99.962 ;
               RECT 8.014 101.126 8.066 101.162 ;
               RECT 8.014 102.326 8.066 102.362 ;
               RECT 8.014 103.526 8.066 103.562 ;
               RECT 8.094 1.558 8.146 1.594 ;
               RECT 8.094 2.758 8.146 2.794 ;
               RECT 8.094 3.958 8.146 3.994 ;
               RECT 8.094 5.158 8.146 5.194 ;
               RECT 8.094 6.358 8.146 6.394 ;
               RECT 8.094 7.558 8.146 7.594 ;
               RECT 8.094 8.758 8.146 8.794 ;
               RECT 8.094 9.958 8.146 9.994 ;
               RECT 8.094 11.158 8.146 11.194 ;
               RECT 8.094 12.358 8.146 12.394 ;
               RECT 8.094 13.558 8.146 13.594 ;
               RECT 8.094 14.758 8.146 14.794 ;
               RECT 8.094 15.958 8.146 15.994 ;
               RECT 8.094 17.158 8.146 17.194 ;
               RECT 8.094 18.358 8.146 18.394 ;
               RECT 8.094 19.558 8.146 19.594 ;
               RECT 8.094 20.758 8.146 20.794 ;
               RECT 8.094 21.958 8.146 21.994 ;
               RECT 8.094 23.158 8.146 23.194 ;
               RECT 8.094 24.358 8.146 24.394 ;
               RECT 8.094 25.558 8.146 25.594 ;
               RECT 8.094 26.758 8.146 26.794 ;
               RECT 8.094 27.958 8.146 27.994 ;
               RECT 8.094 29.158 8.146 29.194 ;
               RECT 8.094 30.358 8.146 30.394 ;
               RECT 8.094 31.558 8.146 31.594 ;
               RECT 8.094 32.758 8.146 32.794 ;
               RECT 8.094 33.958 8.146 33.994 ;
               RECT 8.094 35.158 8.146 35.194 ;
               RECT 8.094 36.358 8.146 36.394 ;
               RECT 8.094 37.558 8.146 37.594 ;
               RECT 8.094 38.758 8.146 38.794 ;
               RECT 8.094 39.958 8.146 39.994 ;
               RECT 8.094 41.158 8.146 41.194 ;
               RECT 8.094 42.358 8.146 42.394 ;
               RECT 8.094 43.558 8.146 43.594 ;
               RECT 8.094 44.758 8.146 44.794 ;
               RECT 8.094 45.958 8.146 45.994 ;
               RECT 8.094 47.158 8.146 47.194 ;
               RECT 8.094 48.358 8.146 48.394 ;
               RECT 8.094 50.142 8.146 50.178 ;
               RECT 8.094 50.382 8.146 50.418 ;
               RECT 8.094 54.702 8.146 54.738 ;
               RECT 8.094 54.942 8.146 54.978 ;
               RECT 8.094 57.478 8.146 57.514 ;
               RECT 8.094 58.678 8.146 58.714 ;
               RECT 8.094 59.878 8.146 59.914 ;
               RECT 8.094 61.078 8.146 61.114 ;
               RECT 8.094 62.278 8.146 62.314 ;
               RECT 8.094 63.478 8.146 63.514 ;
               RECT 8.094 64.678 8.146 64.714 ;
               RECT 8.094 65.878 8.146 65.914 ;
               RECT 8.094 67.078 8.146 67.114 ;
               RECT 8.094 68.278 8.146 68.314 ;
               RECT 8.094 69.478 8.146 69.514 ;
               RECT 8.094 70.678 8.146 70.714 ;
               RECT 8.094 71.878 8.146 71.914 ;
               RECT 8.094 73.078 8.146 73.114 ;
               RECT 8.094 74.278 8.146 74.314 ;
               RECT 8.094 75.478 8.146 75.514 ;
               RECT 8.094 76.678 8.146 76.714 ;
               RECT 8.094 77.878 8.146 77.914 ;
               RECT 8.094 79.078 8.146 79.114 ;
               RECT 8.094 80.278 8.146 80.314 ;
               RECT 8.094 81.478 8.146 81.514 ;
               RECT 8.094 82.678 8.146 82.714 ;
               RECT 8.094 83.878 8.146 83.914 ;
               RECT 8.094 85.078 8.146 85.114 ;
               RECT 8.094 86.278 8.146 86.314 ;
               RECT 8.094 87.478 8.146 87.514 ;
               RECT 8.094 88.678 8.146 88.714 ;
               RECT 8.094 89.878 8.146 89.914 ;
               RECT 8.094 91.078 8.146 91.114 ;
               RECT 8.094 92.278 8.146 92.314 ;
               RECT 8.094 93.478 8.146 93.514 ;
               RECT 8.094 94.678 8.146 94.714 ;
               RECT 8.094 95.878 8.146 95.914 ;
               RECT 8.094 97.078 8.146 97.114 ;
               RECT 8.094 98.278 8.146 98.314 ;
               RECT 8.094 99.478 8.146 99.514 ;
               RECT 8.094 100.678 8.146 100.714 ;
               RECT 8.094 101.878 8.146 101.914 ;
               RECT 8.094 103.078 8.146 103.114 ;
               RECT 8.094 104.278 8.146 104.314 ;
               RECT 8.174 0.281 8.226 0.317 ;
               RECT 8.174 104.803 8.226 104.839 ;
               RECT 8.254 0.806 8.306 0.842 ;
               RECT 8.254 2.006 8.306 2.042 ;
               RECT 8.254 3.206 8.306 3.242 ;
               RECT 8.254 4.406 8.306 4.442 ;
               RECT 8.254 5.606 8.306 5.642 ;
               RECT 8.254 6.806 8.306 6.842 ;
               RECT 8.254 8.006 8.306 8.042 ;
               RECT 8.254 9.206 8.306 9.242 ;
               RECT 8.254 10.406 8.306 10.442 ;
               RECT 8.254 11.606 8.306 11.642 ;
               RECT 8.254 12.806 8.306 12.842 ;
               RECT 8.254 14.006 8.306 14.042 ;
               RECT 8.254 15.206 8.306 15.242 ;
               RECT 8.254 16.406 8.306 16.442 ;
               RECT 8.254 17.606 8.306 17.642 ;
               RECT 8.254 18.806 8.306 18.842 ;
               RECT 8.254 20.006 8.306 20.042 ;
               RECT 8.254 21.206 8.306 21.242 ;
               RECT 8.254 22.406 8.306 22.442 ;
               RECT 8.254 23.606 8.306 23.642 ;
               RECT 8.254 24.806 8.306 24.842 ;
               RECT 8.254 26.006 8.306 26.042 ;
               RECT 8.254 27.206 8.306 27.242 ;
               RECT 8.254 28.406 8.306 28.442 ;
               RECT 8.254 29.606 8.306 29.642 ;
               RECT 8.254 30.806 8.306 30.842 ;
               RECT 8.254 32.006 8.306 32.042 ;
               RECT 8.254 33.206 8.306 33.242 ;
               RECT 8.254 34.406 8.306 34.442 ;
               RECT 8.254 35.606 8.306 35.642 ;
               RECT 8.254 36.806 8.306 36.842 ;
               RECT 8.254 38.006 8.306 38.042 ;
               RECT 8.254 39.206 8.306 39.242 ;
               RECT 8.254 40.406 8.306 40.442 ;
               RECT 8.254 41.606 8.306 41.642 ;
               RECT 8.254 42.806 8.306 42.842 ;
               RECT 8.254 44.006 8.306 44.042 ;
               RECT 8.254 45.206 8.306 45.242 ;
               RECT 8.254 46.406 8.306 46.442 ;
               RECT 8.254 47.606 8.306 47.642 ;
               RECT 8.254 49.422 8.306 49.458 ;
               RECT 8.254 49.662 8.306 49.698 ;
               RECT 8.254 51.102 8.306 51.138 ;
               RECT 8.254 51.582 8.306 51.618 ;
               RECT 8.254 53.502 8.306 53.538 ;
               RECT 8.254 53.982 8.306 54.018 ;
               RECT 8.254 55.422 8.306 55.458 ;
               RECT 8.254 55.662 8.306 55.698 ;
               RECT 8.254 56.726 8.306 56.762 ;
               RECT 8.254 57.926 8.306 57.962 ;
               RECT 8.254 59.126 8.306 59.162 ;
               RECT 8.254 60.326 8.306 60.362 ;
               RECT 8.254 61.526 8.306 61.562 ;
               RECT 8.254 62.726 8.306 62.762 ;
               RECT 8.254 63.926 8.306 63.962 ;
               RECT 8.254 65.126 8.306 65.162 ;
               RECT 8.254 66.326 8.306 66.362 ;
               RECT 8.254 67.526 8.306 67.562 ;
               RECT 8.254 68.726 8.306 68.762 ;
               RECT 8.254 69.926 8.306 69.962 ;
               RECT 8.254 71.126 8.306 71.162 ;
               RECT 8.254 72.326 8.306 72.362 ;
               RECT 8.254 73.526 8.306 73.562 ;
               RECT 8.254 74.726 8.306 74.762 ;
               RECT 8.254 75.926 8.306 75.962 ;
               RECT 8.254 77.126 8.306 77.162 ;
               RECT 8.254 78.326 8.306 78.362 ;
               RECT 8.254 79.526 8.306 79.562 ;
               RECT 8.254 80.726 8.306 80.762 ;
               RECT 8.254 81.926 8.306 81.962 ;
               RECT 8.254 83.126 8.306 83.162 ;
               RECT 8.254 84.326 8.306 84.362 ;
               RECT 8.254 85.526 8.306 85.562 ;
               RECT 8.254 86.726 8.306 86.762 ;
               RECT 8.254 87.926 8.306 87.962 ;
               RECT 8.254 89.126 8.306 89.162 ;
               RECT 8.254 90.326 8.306 90.362 ;
               RECT 8.254 91.526 8.306 91.562 ;
               RECT 8.254 92.726 8.306 92.762 ;
               RECT 8.254 93.926 8.306 93.962 ;
               RECT 8.254 95.126 8.306 95.162 ;
               RECT 8.254 96.326 8.306 96.362 ;
               RECT 8.254 97.526 8.306 97.562 ;
               RECT 8.254 98.726 8.306 98.762 ;
               RECT 8.254 99.926 8.306 99.962 ;
               RECT 8.254 101.126 8.306 101.162 ;
               RECT 8.254 102.326 8.306 102.362 ;
               RECT 8.254 103.526 8.306 103.562 ;
               RECT 8.334 1.558 8.386 1.594 ;
               RECT 8.334 2.758 8.386 2.794 ;
               RECT 8.334 3.958 8.386 3.994 ;
               RECT 8.334 5.158 8.386 5.194 ;
               RECT 8.334 6.358 8.386 6.394 ;
               RECT 8.334 7.558 8.386 7.594 ;
               RECT 8.334 8.758 8.386 8.794 ;
               RECT 8.334 9.958 8.386 9.994 ;
               RECT 8.334 11.158 8.386 11.194 ;
               RECT 8.334 12.358 8.386 12.394 ;
               RECT 8.334 13.558 8.386 13.594 ;
               RECT 8.334 14.758 8.386 14.794 ;
               RECT 8.334 15.958 8.386 15.994 ;
               RECT 8.334 17.158 8.386 17.194 ;
               RECT 8.334 18.358 8.386 18.394 ;
               RECT 8.334 19.558 8.386 19.594 ;
               RECT 8.334 20.758 8.386 20.794 ;
               RECT 8.334 21.958 8.386 21.994 ;
               RECT 8.334 23.158 8.386 23.194 ;
               RECT 8.334 24.358 8.386 24.394 ;
               RECT 8.334 25.558 8.386 25.594 ;
               RECT 8.334 26.758 8.386 26.794 ;
               RECT 8.334 27.958 8.386 27.994 ;
               RECT 8.334 29.158 8.386 29.194 ;
               RECT 8.334 30.358 8.386 30.394 ;
               RECT 8.334 31.558 8.386 31.594 ;
               RECT 8.334 32.758 8.386 32.794 ;
               RECT 8.334 33.958 8.386 33.994 ;
               RECT 8.334 35.158 8.386 35.194 ;
               RECT 8.334 36.358 8.386 36.394 ;
               RECT 8.334 37.558 8.386 37.594 ;
               RECT 8.334 38.758 8.386 38.794 ;
               RECT 8.334 39.958 8.386 39.994 ;
               RECT 8.334 41.158 8.386 41.194 ;
               RECT 8.334 42.358 8.386 42.394 ;
               RECT 8.334 43.558 8.386 43.594 ;
               RECT 8.334 44.758 8.386 44.794 ;
               RECT 8.334 45.958 8.386 45.994 ;
               RECT 8.334 47.158 8.386 47.194 ;
               RECT 8.334 48.358 8.386 48.394 ;
               RECT 8.334 50.142 8.386 50.178 ;
               RECT 8.334 50.382 8.386 50.418 ;
               RECT 8.334 54.702 8.386 54.738 ;
               RECT 8.334 54.942 8.386 54.978 ;
               RECT 8.334 57.478 8.386 57.514 ;
               RECT 8.334 58.678 8.386 58.714 ;
               RECT 8.334 59.878 8.386 59.914 ;
               RECT 8.334 61.078 8.386 61.114 ;
               RECT 8.334 62.278 8.386 62.314 ;
               RECT 8.334 63.478 8.386 63.514 ;
               RECT 8.334 64.678 8.386 64.714 ;
               RECT 8.334 65.878 8.386 65.914 ;
               RECT 8.334 67.078 8.386 67.114 ;
               RECT 8.334 68.278 8.386 68.314 ;
               RECT 8.334 69.478 8.386 69.514 ;
               RECT 8.334 70.678 8.386 70.714 ;
               RECT 8.334 71.878 8.386 71.914 ;
               RECT 8.334 73.078 8.386 73.114 ;
               RECT 8.334 74.278 8.386 74.314 ;
               RECT 8.334 75.478 8.386 75.514 ;
               RECT 8.334 76.678 8.386 76.714 ;
               RECT 8.334 77.878 8.386 77.914 ;
               RECT 8.334 79.078 8.386 79.114 ;
               RECT 8.334 80.278 8.386 80.314 ;
               RECT 8.334 81.478 8.386 81.514 ;
               RECT 8.334 82.678 8.386 82.714 ;
               RECT 8.334 83.878 8.386 83.914 ;
               RECT 8.334 85.078 8.386 85.114 ;
               RECT 8.334 86.278 8.386 86.314 ;
               RECT 8.334 87.478 8.386 87.514 ;
               RECT 8.334 88.678 8.386 88.714 ;
               RECT 8.334 89.878 8.386 89.914 ;
               RECT 8.334 91.078 8.386 91.114 ;
               RECT 8.334 92.278 8.386 92.314 ;
               RECT 8.334 93.478 8.386 93.514 ;
               RECT 8.334 94.678 8.386 94.714 ;
               RECT 8.334 95.878 8.386 95.914 ;
               RECT 8.334 97.078 8.386 97.114 ;
               RECT 8.334 98.278 8.386 98.314 ;
               RECT 8.334 99.478 8.386 99.514 ;
               RECT 8.334 100.678 8.386 100.714 ;
               RECT 8.334 101.878 8.386 101.914 ;
               RECT 8.334 103.078 8.386 103.114 ;
               RECT 8.334 104.278 8.386 104.314 ;
               RECT 8.414 0.806 8.466 0.842 ;
               RECT 8.414 2.006 8.466 2.042 ;
               RECT 8.414 3.206 8.466 3.242 ;
               RECT 8.414 4.406 8.466 4.442 ;
               RECT 8.414 5.606 8.466 5.642 ;
               RECT 8.414 6.806 8.466 6.842 ;
               RECT 8.414 8.006 8.466 8.042 ;
               RECT 8.414 9.206 8.466 9.242 ;
               RECT 8.414 10.406 8.466 10.442 ;
               RECT 8.414 11.606 8.466 11.642 ;
               RECT 8.414 12.806 8.466 12.842 ;
               RECT 8.414 14.006 8.466 14.042 ;
               RECT 8.414 15.206 8.466 15.242 ;
               RECT 8.414 16.406 8.466 16.442 ;
               RECT 8.414 17.606 8.466 17.642 ;
               RECT 8.414 18.806 8.466 18.842 ;
               RECT 8.414 20.006 8.466 20.042 ;
               RECT 8.414 21.206 8.466 21.242 ;
               RECT 8.414 22.406 8.466 22.442 ;
               RECT 8.414 23.606 8.466 23.642 ;
               RECT 8.414 24.806 8.466 24.842 ;
               RECT 8.414 26.006 8.466 26.042 ;
               RECT 8.414 27.206 8.466 27.242 ;
               RECT 8.414 28.406 8.466 28.442 ;
               RECT 8.414 29.606 8.466 29.642 ;
               RECT 8.414 30.806 8.466 30.842 ;
               RECT 8.414 32.006 8.466 32.042 ;
               RECT 8.414 33.206 8.466 33.242 ;
               RECT 8.414 34.406 8.466 34.442 ;
               RECT 8.414 35.606 8.466 35.642 ;
               RECT 8.414 36.806 8.466 36.842 ;
               RECT 8.414 38.006 8.466 38.042 ;
               RECT 8.414 39.206 8.466 39.242 ;
               RECT 8.414 40.406 8.466 40.442 ;
               RECT 8.414 41.606 8.466 41.642 ;
               RECT 8.414 42.806 8.466 42.842 ;
               RECT 8.414 44.006 8.466 44.042 ;
               RECT 8.414 45.206 8.466 45.242 ;
               RECT 8.414 46.406 8.466 46.442 ;
               RECT 8.414 47.606 8.466 47.642 ;
               RECT 8.414 49.422 8.466 49.458 ;
               RECT 8.414 49.662 8.466 49.698 ;
               RECT 8.414 55.422 8.466 55.458 ;
               RECT 8.414 55.662 8.466 55.698 ;
               RECT 8.414 56.726 8.466 56.762 ;
               RECT 8.414 57.926 8.466 57.962 ;
               RECT 8.414 59.126 8.466 59.162 ;
               RECT 8.414 60.326 8.466 60.362 ;
               RECT 8.414 61.526 8.466 61.562 ;
               RECT 8.414 62.726 8.466 62.762 ;
               RECT 8.414 63.926 8.466 63.962 ;
               RECT 8.414 65.126 8.466 65.162 ;
               RECT 8.414 66.326 8.466 66.362 ;
               RECT 8.414 67.526 8.466 67.562 ;
               RECT 8.414 68.726 8.466 68.762 ;
               RECT 8.414 69.926 8.466 69.962 ;
               RECT 8.414 71.126 8.466 71.162 ;
               RECT 8.414 72.326 8.466 72.362 ;
               RECT 8.414 73.526 8.466 73.562 ;
               RECT 8.414 74.726 8.466 74.762 ;
               RECT 8.414 75.926 8.466 75.962 ;
               RECT 8.414 77.126 8.466 77.162 ;
               RECT 8.414 78.326 8.466 78.362 ;
               RECT 8.414 79.526 8.466 79.562 ;
               RECT 8.414 80.726 8.466 80.762 ;
               RECT 8.414 81.926 8.466 81.962 ;
               RECT 8.414 83.126 8.466 83.162 ;
               RECT 8.414 84.326 8.466 84.362 ;
               RECT 8.414 85.526 8.466 85.562 ;
               RECT 8.414 86.726 8.466 86.762 ;
               RECT 8.414 87.926 8.466 87.962 ;
               RECT 8.414 89.126 8.466 89.162 ;
               RECT 8.414 90.326 8.466 90.362 ;
               RECT 8.414 91.526 8.466 91.562 ;
               RECT 8.414 92.726 8.466 92.762 ;
               RECT 8.414 93.926 8.466 93.962 ;
               RECT 8.414 95.126 8.466 95.162 ;
               RECT 8.414 96.326 8.466 96.362 ;
               RECT 8.414 97.526 8.466 97.562 ;
               RECT 8.414 98.726 8.466 98.762 ;
               RECT 8.414 99.926 8.466 99.962 ;
               RECT 8.414 101.126 8.466 101.162 ;
               RECT 8.414 102.326 8.466 102.362 ;
               RECT 8.414 103.526 8.466 103.562 ;
               RECT 8.494 1.558 8.546 1.594 ;
               RECT 8.494 2.758 8.546 2.794 ;
               RECT 8.494 3.958 8.546 3.994 ;
               RECT 8.494 5.158 8.546 5.194 ;
               RECT 8.494 6.358 8.546 6.394 ;
               RECT 8.494 7.558 8.546 7.594 ;
               RECT 8.494 8.758 8.546 8.794 ;
               RECT 8.494 9.958 8.546 9.994 ;
               RECT 8.494 11.158 8.546 11.194 ;
               RECT 8.494 12.358 8.546 12.394 ;
               RECT 8.494 13.558 8.546 13.594 ;
               RECT 8.494 14.758 8.546 14.794 ;
               RECT 8.494 15.958 8.546 15.994 ;
               RECT 8.494 17.158 8.546 17.194 ;
               RECT 8.494 18.358 8.546 18.394 ;
               RECT 8.494 19.558 8.546 19.594 ;
               RECT 8.494 20.758 8.546 20.794 ;
               RECT 8.494 21.958 8.546 21.994 ;
               RECT 8.494 23.158 8.546 23.194 ;
               RECT 8.494 24.358 8.546 24.394 ;
               RECT 8.494 25.558 8.546 25.594 ;
               RECT 8.494 26.758 8.546 26.794 ;
               RECT 8.494 27.958 8.546 27.994 ;
               RECT 8.494 29.158 8.546 29.194 ;
               RECT 8.494 30.358 8.546 30.394 ;
               RECT 8.494 31.558 8.546 31.594 ;
               RECT 8.494 32.758 8.546 32.794 ;
               RECT 8.494 33.958 8.546 33.994 ;
               RECT 8.494 35.158 8.546 35.194 ;
               RECT 8.494 36.358 8.546 36.394 ;
               RECT 8.494 37.558 8.546 37.594 ;
               RECT 8.494 38.758 8.546 38.794 ;
               RECT 8.494 39.958 8.546 39.994 ;
               RECT 8.494 41.158 8.546 41.194 ;
               RECT 8.494 42.358 8.546 42.394 ;
               RECT 8.494 43.558 8.546 43.594 ;
               RECT 8.494 44.758 8.546 44.794 ;
               RECT 8.494 45.958 8.546 45.994 ;
               RECT 8.494 47.158 8.546 47.194 ;
               RECT 8.494 48.358 8.546 48.394 ;
               RECT 8.494 50.142 8.546 50.178 ;
               RECT 8.494 50.382 8.546 50.418 ;
               RECT 8.494 54.702 8.546 54.738 ;
               RECT 8.494 54.942 8.546 54.978 ;
               RECT 8.494 57.478 8.546 57.514 ;
               RECT 8.494 58.678 8.546 58.714 ;
               RECT 8.494 59.878 8.546 59.914 ;
               RECT 8.494 61.078 8.546 61.114 ;
               RECT 8.494 62.278 8.546 62.314 ;
               RECT 8.494 63.478 8.546 63.514 ;
               RECT 8.494 64.678 8.546 64.714 ;
               RECT 8.494 65.878 8.546 65.914 ;
               RECT 8.494 67.078 8.546 67.114 ;
               RECT 8.494 68.278 8.546 68.314 ;
               RECT 8.494 69.478 8.546 69.514 ;
               RECT 8.494 70.678 8.546 70.714 ;
               RECT 8.494 71.878 8.546 71.914 ;
               RECT 8.494 73.078 8.546 73.114 ;
               RECT 8.494 74.278 8.546 74.314 ;
               RECT 8.494 75.478 8.546 75.514 ;
               RECT 8.494 76.678 8.546 76.714 ;
               RECT 8.494 77.878 8.546 77.914 ;
               RECT 8.494 79.078 8.546 79.114 ;
               RECT 8.494 80.278 8.546 80.314 ;
               RECT 8.494 81.478 8.546 81.514 ;
               RECT 8.494 82.678 8.546 82.714 ;
               RECT 8.494 83.878 8.546 83.914 ;
               RECT 8.494 85.078 8.546 85.114 ;
               RECT 8.494 86.278 8.546 86.314 ;
               RECT 8.494 87.478 8.546 87.514 ;
               RECT 8.494 88.678 8.546 88.714 ;
               RECT 8.494 89.878 8.546 89.914 ;
               RECT 8.494 91.078 8.546 91.114 ;
               RECT 8.494 92.278 8.546 92.314 ;
               RECT 8.494 93.478 8.546 93.514 ;
               RECT 8.494 94.678 8.546 94.714 ;
               RECT 8.494 95.878 8.546 95.914 ;
               RECT 8.494 97.078 8.546 97.114 ;
               RECT 8.494 98.278 8.546 98.314 ;
               RECT 8.494 99.478 8.546 99.514 ;
               RECT 8.494 100.678 8.546 100.714 ;
               RECT 8.494 101.878 8.546 101.914 ;
               RECT 8.494 103.078 8.546 103.114 ;
               RECT 8.494 104.278 8.546 104.314 ;
               RECT 8.574 0.281 8.626 0.317 ;
               RECT 8.574 104.803 8.626 104.839 ;
               RECT 8.654 0.806 8.706 0.842 ;
               RECT 8.654 2.006 8.706 2.042 ;
               RECT 8.654 3.206 8.706 3.242 ;
               RECT 8.654 4.406 8.706 4.442 ;
               RECT 8.654 5.606 8.706 5.642 ;
               RECT 8.654 6.806 8.706 6.842 ;
               RECT 8.654 8.006 8.706 8.042 ;
               RECT 8.654 9.206 8.706 9.242 ;
               RECT 8.654 10.406 8.706 10.442 ;
               RECT 8.654 11.606 8.706 11.642 ;
               RECT 8.654 12.806 8.706 12.842 ;
               RECT 8.654 14.006 8.706 14.042 ;
               RECT 8.654 15.206 8.706 15.242 ;
               RECT 8.654 16.406 8.706 16.442 ;
               RECT 8.654 17.606 8.706 17.642 ;
               RECT 8.654 18.806 8.706 18.842 ;
               RECT 8.654 20.006 8.706 20.042 ;
               RECT 8.654 21.206 8.706 21.242 ;
               RECT 8.654 22.406 8.706 22.442 ;
               RECT 8.654 23.606 8.706 23.642 ;
               RECT 8.654 24.806 8.706 24.842 ;
               RECT 8.654 26.006 8.706 26.042 ;
               RECT 8.654 27.206 8.706 27.242 ;
               RECT 8.654 28.406 8.706 28.442 ;
               RECT 8.654 29.606 8.706 29.642 ;
               RECT 8.654 30.806 8.706 30.842 ;
               RECT 8.654 32.006 8.706 32.042 ;
               RECT 8.654 33.206 8.706 33.242 ;
               RECT 8.654 34.406 8.706 34.442 ;
               RECT 8.654 35.606 8.706 35.642 ;
               RECT 8.654 36.806 8.706 36.842 ;
               RECT 8.654 38.006 8.706 38.042 ;
               RECT 8.654 39.206 8.706 39.242 ;
               RECT 8.654 40.406 8.706 40.442 ;
               RECT 8.654 41.606 8.706 41.642 ;
               RECT 8.654 42.806 8.706 42.842 ;
               RECT 8.654 44.006 8.706 44.042 ;
               RECT 8.654 45.206 8.706 45.242 ;
               RECT 8.654 46.406 8.706 46.442 ;
               RECT 8.654 47.606 8.706 47.642 ;
               RECT 8.654 49.422 8.706 49.458 ;
               RECT 8.654 49.662 8.706 49.698 ;
               RECT 8.654 55.422 8.706 55.458 ;
               RECT 8.654 55.662 8.706 55.698 ;
               RECT 8.654 56.726 8.706 56.762 ;
               RECT 8.654 57.926 8.706 57.962 ;
               RECT 8.654 59.126 8.706 59.162 ;
               RECT 8.654 60.326 8.706 60.362 ;
               RECT 8.654 61.526 8.706 61.562 ;
               RECT 8.654 62.726 8.706 62.762 ;
               RECT 8.654 63.926 8.706 63.962 ;
               RECT 8.654 65.126 8.706 65.162 ;
               RECT 8.654 66.326 8.706 66.362 ;
               RECT 8.654 67.526 8.706 67.562 ;
               RECT 8.654 68.726 8.706 68.762 ;
               RECT 8.654 69.926 8.706 69.962 ;
               RECT 8.654 71.126 8.706 71.162 ;
               RECT 8.654 72.326 8.706 72.362 ;
               RECT 8.654 73.526 8.706 73.562 ;
               RECT 8.654 74.726 8.706 74.762 ;
               RECT 8.654 75.926 8.706 75.962 ;
               RECT 8.654 77.126 8.706 77.162 ;
               RECT 8.654 78.326 8.706 78.362 ;
               RECT 8.654 79.526 8.706 79.562 ;
               RECT 8.654 80.726 8.706 80.762 ;
               RECT 8.654 81.926 8.706 81.962 ;
               RECT 8.654 83.126 8.706 83.162 ;
               RECT 8.654 84.326 8.706 84.362 ;
               RECT 8.654 85.526 8.706 85.562 ;
               RECT 8.654 86.726 8.706 86.762 ;
               RECT 8.654 87.926 8.706 87.962 ;
               RECT 8.654 89.126 8.706 89.162 ;
               RECT 8.654 90.326 8.706 90.362 ;
               RECT 8.654 91.526 8.706 91.562 ;
               RECT 8.654 92.726 8.706 92.762 ;
               RECT 8.654 93.926 8.706 93.962 ;
               RECT 8.654 95.126 8.706 95.162 ;
               RECT 8.654 96.326 8.706 96.362 ;
               RECT 8.654 97.526 8.706 97.562 ;
               RECT 8.654 98.726 8.706 98.762 ;
               RECT 8.654 99.926 8.706 99.962 ;
               RECT 8.654 101.126 8.706 101.162 ;
               RECT 8.654 102.326 8.706 102.362 ;
               RECT 8.654 103.526 8.706 103.562 ;
               RECT 8.734 1.558 8.786 1.594 ;
               RECT 8.734 2.758 8.786 2.794 ;
               RECT 8.734 3.958 8.786 3.994 ;
               RECT 8.734 5.158 8.786 5.194 ;
               RECT 8.734 6.358 8.786 6.394 ;
               RECT 8.734 7.558 8.786 7.594 ;
               RECT 8.734 8.758 8.786 8.794 ;
               RECT 8.734 9.958 8.786 9.994 ;
               RECT 8.734 11.158 8.786 11.194 ;
               RECT 8.734 12.358 8.786 12.394 ;
               RECT 8.734 13.558 8.786 13.594 ;
               RECT 8.734 14.758 8.786 14.794 ;
               RECT 8.734 15.958 8.786 15.994 ;
               RECT 8.734 17.158 8.786 17.194 ;
               RECT 8.734 18.358 8.786 18.394 ;
               RECT 8.734 19.558 8.786 19.594 ;
               RECT 8.734 20.758 8.786 20.794 ;
               RECT 8.734 21.958 8.786 21.994 ;
               RECT 8.734 23.158 8.786 23.194 ;
               RECT 8.734 24.358 8.786 24.394 ;
               RECT 8.734 25.558 8.786 25.594 ;
               RECT 8.734 26.758 8.786 26.794 ;
               RECT 8.734 27.958 8.786 27.994 ;
               RECT 8.734 29.158 8.786 29.194 ;
               RECT 8.734 30.358 8.786 30.394 ;
               RECT 8.734 31.558 8.786 31.594 ;
               RECT 8.734 32.758 8.786 32.794 ;
               RECT 8.734 33.958 8.786 33.994 ;
               RECT 8.734 35.158 8.786 35.194 ;
               RECT 8.734 36.358 8.786 36.394 ;
               RECT 8.734 37.558 8.786 37.594 ;
               RECT 8.734 38.758 8.786 38.794 ;
               RECT 8.734 39.958 8.786 39.994 ;
               RECT 8.734 41.158 8.786 41.194 ;
               RECT 8.734 42.358 8.786 42.394 ;
               RECT 8.734 43.558 8.786 43.594 ;
               RECT 8.734 44.758 8.786 44.794 ;
               RECT 8.734 45.958 8.786 45.994 ;
               RECT 8.734 47.158 8.786 47.194 ;
               RECT 8.734 48.358 8.786 48.394 ;
               RECT 8.734 50.142 8.786 50.178 ;
               RECT 8.734 50.382 8.786 50.418 ;
               RECT 8.734 54.702 8.786 54.738 ;
               RECT 8.734 54.942 8.786 54.978 ;
               RECT 8.734 57.478 8.786 57.514 ;
               RECT 8.734 58.678 8.786 58.714 ;
               RECT 8.734 59.878 8.786 59.914 ;
               RECT 8.734 61.078 8.786 61.114 ;
               RECT 8.734 62.278 8.786 62.314 ;
               RECT 8.734 63.478 8.786 63.514 ;
               RECT 8.734 64.678 8.786 64.714 ;
               RECT 8.734 65.878 8.786 65.914 ;
               RECT 8.734 67.078 8.786 67.114 ;
               RECT 8.734 68.278 8.786 68.314 ;
               RECT 8.734 69.478 8.786 69.514 ;
               RECT 8.734 70.678 8.786 70.714 ;
               RECT 8.734 71.878 8.786 71.914 ;
               RECT 8.734 73.078 8.786 73.114 ;
               RECT 8.734 74.278 8.786 74.314 ;
               RECT 8.734 75.478 8.786 75.514 ;
               RECT 8.734 76.678 8.786 76.714 ;
               RECT 8.734 77.878 8.786 77.914 ;
               RECT 8.734 79.078 8.786 79.114 ;
               RECT 8.734 80.278 8.786 80.314 ;
               RECT 8.734 81.478 8.786 81.514 ;
               RECT 8.734 82.678 8.786 82.714 ;
               RECT 8.734 83.878 8.786 83.914 ;
               RECT 8.734 85.078 8.786 85.114 ;
               RECT 8.734 86.278 8.786 86.314 ;
               RECT 8.734 87.478 8.786 87.514 ;
               RECT 8.734 88.678 8.786 88.714 ;
               RECT 8.734 89.878 8.786 89.914 ;
               RECT 8.734 91.078 8.786 91.114 ;
               RECT 8.734 92.278 8.786 92.314 ;
               RECT 8.734 93.478 8.786 93.514 ;
               RECT 8.734 94.678 8.786 94.714 ;
               RECT 8.734 95.878 8.786 95.914 ;
               RECT 8.734 97.078 8.786 97.114 ;
               RECT 8.734 98.278 8.786 98.314 ;
               RECT 8.734 99.478 8.786 99.514 ;
               RECT 8.734 100.678 8.786 100.714 ;
               RECT 8.734 101.878 8.786 101.914 ;
               RECT 8.734 103.078 8.786 103.114 ;
               RECT 8.734 104.278 8.786 104.314 ;
               RECT 8.814 0.806 8.866 0.842 ;
               RECT 8.814 2.006 8.866 2.042 ;
               RECT 8.814 3.206 8.866 3.242 ;
               RECT 8.814 4.406 8.866 4.442 ;
               RECT 8.814 5.606 8.866 5.642 ;
               RECT 8.814 6.806 8.866 6.842 ;
               RECT 8.814 8.006 8.866 8.042 ;
               RECT 8.814 9.206 8.866 9.242 ;
               RECT 8.814 10.406 8.866 10.442 ;
               RECT 8.814 11.606 8.866 11.642 ;
               RECT 8.814 12.806 8.866 12.842 ;
               RECT 8.814 14.006 8.866 14.042 ;
               RECT 8.814 15.206 8.866 15.242 ;
               RECT 8.814 16.406 8.866 16.442 ;
               RECT 8.814 17.606 8.866 17.642 ;
               RECT 8.814 18.806 8.866 18.842 ;
               RECT 8.814 20.006 8.866 20.042 ;
               RECT 8.814 21.206 8.866 21.242 ;
               RECT 8.814 22.406 8.866 22.442 ;
               RECT 8.814 23.606 8.866 23.642 ;
               RECT 8.814 24.806 8.866 24.842 ;
               RECT 8.814 26.006 8.866 26.042 ;
               RECT 8.814 27.206 8.866 27.242 ;
               RECT 8.814 28.406 8.866 28.442 ;
               RECT 8.814 29.606 8.866 29.642 ;
               RECT 8.814 30.806 8.866 30.842 ;
               RECT 8.814 32.006 8.866 32.042 ;
               RECT 8.814 33.206 8.866 33.242 ;
               RECT 8.814 34.406 8.866 34.442 ;
               RECT 8.814 35.606 8.866 35.642 ;
               RECT 8.814 36.806 8.866 36.842 ;
               RECT 8.814 38.006 8.866 38.042 ;
               RECT 8.814 39.206 8.866 39.242 ;
               RECT 8.814 40.406 8.866 40.442 ;
               RECT 8.814 41.606 8.866 41.642 ;
               RECT 8.814 42.806 8.866 42.842 ;
               RECT 8.814 44.006 8.866 44.042 ;
               RECT 8.814 45.206 8.866 45.242 ;
               RECT 8.814 46.406 8.866 46.442 ;
               RECT 8.814 47.606 8.866 47.642 ;
               RECT 8.814 49.422 8.866 49.458 ;
               RECT 8.814 49.662 8.866 49.698 ;
               RECT 8.814 55.422 8.866 55.458 ;
               RECT 8.814 55.662 8.866 55.698 ;
               RECT 8.814 56.726 8.866 56.762 ;
               RECT 8.814 57.926 8.866 57.962 ;
               RECT 8.814 59.126 8.866 59.162 ;
               RECT 8.814 60.326 8.866 60.362 ;
               RECT 8.814 61.526 8.866 61.562 ;
               RECT 8.814 62.726 8.866 62.762 ;
               RECT 8.814 63.926 8.866 63.962 ;
               RECT 8.814 65.126 8.866 65.162 ;
               RECT 8.814 66.326 8.866 66.362 ;
               RECT 8.814 67.526 8.866 67.562 ;
               RECT 8.814 68.726 8.866 68.762 ;
               RECT 8.814 69.926 8.866 69.962 ;
               RECT 8.814 71.126 8.866 71.162 ;
               RECT 8.814 72.326 8.866 72.362 ;
               RECT 8.814 73.526 8.866 73.562 ;
               RECT 8.814 74.726 8.866 74.762 ;
               RECT 8.814 75.926 8.866 75.962 ;
               RECT 8.814 77.126 8.866 77.162 ;
               RECT 8.814 78.326 8.866 78.362 ;
               RECT 8.814 79.526 8.866 79.562 ;
               RECT 8.814 80.726 8.866 80.762 ;
               RECT 8.814 81.926 8.866 81.962 ;
               RECT 8.814 83.126 8.866 83.162 ;
               RECT 8.814 84.326 8.866 84.362 ;
               RECT 8.814 85.526 8.866 85.562 ;
               RECT 8.814 86.726 8.866 86.762 ;
               RECT 8.814 87.926 8.866 87.962 ;
               RECT 8.814 89.126 8.866 89.162 ;
               RECT 8.814 90.326 8.866 90.362 ;
               RECT 8.814 91.526 8.866 91.562 ;
               RECT 8.814 92.726 8.866 92.762 ;
               RECT 8.814 93.926 8.866 93.962 ;
               RECT 8.814 95.126 8.866 95.162 ;
               RECT 8.814 96.326 8.866 96.362 ;
               RECT 8.814 97.526 8.866 97.562 ;
               RECT 8.814 98.726 8.866 98.762 ;
               RECT 8.814 99.926 8.866 99.962 ;
               RECT 8.814 101.126 8.866 101.162 ;
               RECT 8.814 102.326 8.866 102.362 ;
               RECT 8.814 103.526 8.866 103.562 ;
               RECT 8.894 1.558 8.946 1.594 ;
               RECT 8.894 2.758 8.946 2.794 ;
               RECT 8.894 3.958 8.946 3.994 ;
               RECT 8.894 5.158 8.946 5.194 ;
               RECT 8.894 6.358 8.946 6.394 ;
               RECT 8.894 7.558 8.946 7.594 ;
               RECT 8.894 8.758 8.946 8.794 ;
               RECT 8.894 9.958 8.946 9.994 ;
               RECT 8.894 11.158 8.946 11.194 ;
               RECT 8.894 12.358 8.946 12.394 ;
               RECT 8.894 13.558 8.946 13.594 ;
               RECT 8.894 14.758 8.946 14.794 ;
               RECT 8.894 15.958 8.946 15.994 ;
               RECT 8.894 17.158 8.946 17.194 ;
               RECT 8.894 18.358 8.946 18.394 ;
               RECT 8.894 19.558 8.946 19.594 ;
               RECT 8.894 20.758 8.946 20.794 ;
               RECT 8.894 21.958 8.946 21.994 ;
               RECT 8.894 23.158 8.946 23.194 ;
               RECT 8.894 24.358 8.946 24.394 ;
               RECT 8.894 25.558 8.946 25.594 ;
               RECT 8.894 26.758 8.946 26.794 ;
               RECT 8.894 27.958 8.946 27.994 ;
               RECT 8.894 29.158 8.946 29.194 ;
               RECT 8.894 30.358 8.946 30.394 ;
               RECT 8.894 31.558 8.946 31.594 ;
               RECT 8.894 32.758 8.946 32.794 ;
               RECT 8.894 33.958 8.946 33.994 ;
               RECT 8.894 35.158 8.946 35.194 ;
               RECT 8.894 36.358 8.946 36.394 ;
               RECT 8.894 37.558 8.946 37.594 ;
               RECT 8.894 38.758 8.946 38.794 ;
               RECT 8.894 39.958 8.946 39.994 ;
               RECT 8.894 41.158 8.946 41.194 ;
               RECT 8.894 42.358 8.946 42.394 ;
               RECT 8.894 43.558 8.946 43.594 ;
               RECT 8.894 44.758 8.946 44.794 ;
               RECT 8.894 45.958 8.946 45.994 ;
               RECT 8.894 47.158 8.946 47.194 ;
               RECT 8.894 48.358 8.946 48.394 ;
               RECT 8.894 50.142 8.946 50.178 ;
               RECT 8.894 50.382 8.946 50.418 ;
               RECT 8.894 54.702 8.946 54.738 ;
               RECT 8.894 54.942 8.946 54.978 ;
               RECT 8.894 57.478 8.946 57.514 ;
               RECT 8.894 58.678 8.946 58.714 ;
               RECT 8.894 59.878 8.946 59.914 ;
               RECT 8.894 61.078 8.946 61.114 ;
               RECT 8.894 62.278 8.946 62.314 ;
               RECT 8.894 63.478 8.946 63.514 ;
               RECT 8.894 64.678 8.946 64.714 ;
               RECT 8.894 65.878 8.946 65.914 ;
               RECT 8.894 67.078 8.946 67.114 ;
               RECT 8.894 68.278 8.946 68.314 ;
               RECT 8.894 69.478 8.946 69.514 ;
               RECT 8.894 70.678 8.946 70.714 ;
               RECT 8.894 71.878 8.946 71.914 ;
               RECT 8.894 73.078 8.946 73.114 ;
               RECT 8.894 74.278 8.946 74.314 ;
               RECT 8.894 75.478 8.946 75.514 ;
               RECT 8.894 76.678 8.946 76.714 ;
               RECT 8.894 77.878 8.946 77.914 ;
               RECT 8.894 79.078 8.946 79.114 ;
               RECT 8.894 80.278 8.946 80.314 ;
               RECT 8.894 81.478 8.946 81.514 ;
               RECT 8.894 82.678 8.946 82.714 ;
               RECT 8.894 83.878 8.946 83.914 ;
               RECT 8.894 85.078 8.946 85.114 ;
               RECT 8.894 86.278 8.946 86.314 ;
               RECT 8.894 87.478 8.946 87.514 ;
               RECT 8.894 88.678 8.946 88.714 ;
               RECT 8.894 89.878 8.946 89.914 ;
               RECT 8.894 91.078 8.946 91.114 ;
               RECT 8.894 92.278 8.946 92.314 ;
               RECT 8.894 93.478 8.946 93.514 ;
               RECT 8.894 94.678 8.946 94.714 ;
               RECT 8.894 95.878 8.946 95.914 ;
               RECT 8.894 97.078 8.946 97.114 ;
               RECT 8.894 98.278 8.946 98.314 ;
               RECT 8.894 99.478 8.946 99.514 ;
               RECT 8.894 100.678 8.946 100.714 ;
               RECT 8.894 101.878 8.946 101.914 ;
               RECT 8.894 103.078 8.946 103.114 ;
               RECT 8.894 104.278 8.946 104.314 ;
               RECT 8.974 0.281 9.026 0.317 ;
               RECT 8.974 104.803 9.026 104.839 ;
               RECT 9.054 0.806 9.106 0.842 ;
               RECT 9.054 2.006 9.106 2.042 ;
               RECT 9.054 3.206 9.106 3.242 ;
               RECT 9.054 4.406 9.106 4.442 ;
               RECT 9.054 5.606 9.106 5.642 ;
               RECT 9.054 6.806 9.106 6.842 ;
               RECT 9.054 8.006 9.106 8.042 ;
               RECT 9.054 9.206 9.106 9.242 ;
               RECT 9.054 10.406 9.106 10.442 ;
               RECT 9.054 11.606 9.106 11.642 ;
               RECT 9.054 12.806 9.106 12.842 ;
               RECT 9.054 14.006 9.106 14.042 ;
               RECT 9.054 15.206 9.106 15.242 ;
               RECT 9.054 16.406 9.106 16.442 ;
               RECT 9.054 17.606 9.106 17.642 ;
               RECT 9.054 18.806 9.106 18.842 ;
               RECT 9.054 20.006 9.106 20.042 ;
               RECT 9.054 21.206 9.106 21.242 ;
               RECT 9.054 22.406 9.106 22.442 ;
               RECT 9.054 23.606 9.106 23.642 ;
               RECT 9.054 24.806 9.106 24.842 ;
               RECT 9.054 26.006 9.106 26.042 ;
               RECT 9.054 27.206 9.106 27.242 ;
               RECT 9.054 28.406 9.106 28.442 ;
               RECT 9.054 29.606 9.106 29.642 ;
               RECT 9.054 30.806 9.106 30.842 ;
               RECT 9.054 32.006 9.106 32.042 ;
               RECT 9.054 33.206 9.106 33.242 ;
               RECT 9.054 34.406 9.106 34.442 ;
               RECT 9.054 35.606 9.106 35.642 ;
               RECT 9.054 36.806 9.106 36.842 ;
               RECT 9.054 38.006 9.106 38.042 ;
               RECT 9.054 39.206 9.106 39.242 ;
               RECT 9.054 40.406 9.106 40.442 ;
               RECT 9.054 41.606 9.106 41.642 ;
               RECT 9.054 42.806 9.106 42.842 ;
               RECT 9.054 44.006 9.106 44.042 ;
               RECT 9.054 45.206 9.106 45.242 ;
               RECT 9.054 46.406 9.106 46.442 ;
               RECT 9.054 47.606 9.106 47.642 ;
               RECT 9.054 49.422 9.106 49.458 ;
               RECT 9.054 49.662 9.106 49.698 ;
               RECT 9.054 51.102 9.106 51.138 ;
               RECT 9.054 51.582 9.106 51.618 ;
               RECT 9.054 53.502 9.106 53.538 ;
               RECT 9.054 53.982 9.106 54.018 ;
               RECT 9.054 55.422 9.106 55.458 ;
               RECT 9.054 55.662 9.106 55.698 ;
               RECT 9.054 56.726 9.106 56.762 ;
               RECT 9.054 57.926 9.106 57.962 ;
               RECT 9.054 59.126 9.106 59.162 ;
               RECT 9.054 60.326 9.106 60.362 ;
               RECT 9.054 61.526 9.106 61.562 ;
               RECT 9.054 62.726 9.106 62.762 ;
               RECT 9.054 63.926 9.106 63.962 ;
               RECT 9.054 65.126 9.106 65.162 ;
               RECT 9.054 66.326 9.106 66.362 ;
               RECT 9.054 67.526 9.106 67.562 ;
               RECT 9.054 68.726 9.106 68.762 ;
               RECT 9.054 69.926 9.106 69.962 ;
               RECT 9.054 71.126 9.106 71.162 ;
               RECT 9.054 72.326 9.106 72.362 ;
               RECT 9.054 73.526 9.106 73.562 ;
               RECT 9.054 74.726 9.106 74.762 ;
               RECT 9.054 75.926 9.106 75.962 ;
               RECT 9.054 77.126 9.106 77.162 ;
               RECT 9.054 78.326 9.106 78.362 ;
               RECT 9.054 79.526 9.106 79.562 ;
               RECT 9.054 80.726 9.106 80.762 ;
               RECT 9.054 81.926 9.106 81.962 ;
               RECT 9.054 83.126 9.106 83.162 ;
               RECT 9.054 84.326 9.106 84.362 ;
               RECT 9.054 85.526 9.106 85.562 ;
               RECT 9.054 86.726 9.106 86.762 ;
               RECT 9.054 87.926 9.106 87.962 ;
               RECT 9.054 89.126 9.106 89.162 ;
               RECT 9.054 90.326 9.106 90.362 ;
               RECT 9.054 91.526 9.106 91.562 ;
               RECT 9.054 92.726 9.106 92.762 ;
               RECT 9.054 93.926 9.106 93.962 ;
               RECT 9.054 95.126 9.106 95.162 ;
               RECT 9.054 96.326 9.106 96.362 ;
               RECT 9.054 97.526 9.106 97.562 ;
               RECT 9.054 98.726 9.106 98.762 ;
               RECT 9.054 99.926 9.106 99.962 ;
               RECT 9.054 101.126 9.106 101.162 ;
               RECT 9.054 102.326 9.106 102.362 ;
               RECT 9.054 103.526 9.106 103.562 ;
               RECT 9.134 1.558 9.186 1.594 ;
               RECT 9.134 2.758 9.186 2.794 ;
               RECT 9.134 3.958 9.186 3.994 ;
               RECT 9.134 5.158 9.186 5.194 ;
               RECT 9.134 6.358 9.186 6.394 ;
               RECT 9.134 7.558 9.186 7.594 ;
               RECT 9.134 8.758 9.186 8.794 ;
               RECT 9.134 9.958 9.186 9.994 ;
               RECT 9.134 11.158 9.186 11.194 ;
               RECT 9.134 12.358 9.186 12.394 ;
               RECT 9.134 13.558 9.186 13.594 ;
               RECT 9.134 14.758 9.186 14.794 ;
               RECT 9.134 15.958 9.186 15.994 ;
               RECT 9.134 17.158 9.186 17.194 ;
               RECT 9.134 18.358 9.186 18.394 ;
               RECT 9.134 19.558 9.186 19.594 ;
               RECT 9.134 20.758 9.186 20.794 ;
               RECT 9.134 21.958 9.186 21.994 ;
               RECT 9.134 23.158 9.186 23.194 ;
               RECT 9.134 24.358 9.186 24.394 ;
               RECT 9.134 25.558 9.186 25.594 ;
               RECT 9.134 26.758 9.186 26.794 ;
               RECT 9.134 27.958 9.186 27.994 ;
               RECT 9.134 29.158 9.186 29.194 ;
               RECT 9.134 30.358 9.186 30.394 ;
               RECT 9.134 31.558 9.186 31.594 ;
               RECT 9.134 32.758 9.186 32.794 ;
               RECT 9.134 33.958 9.186 33.994 ;
               RECT 9.134 35.158 9.186 35.194 ;
               RECT 9.134 36.358 9.186 36.394 ;
               RECT 9.134 37.558 9.186 37.594 ;
               RECT 9.134 38.758 9.186 38.794 ;
               RECT 9.134 39.958 9.186 39.994 ;
               RECT 9.134 41.158 9.186 41.194 ;
               RECT 9.134 42.358 9.186 42.394 ;
               RECT 9.134 43.558 9.186 43.594 ;
               RECT 9.134 44.758 9.186 44.794 ;
               RECT 9.134 45.958 9.186 45.994 ;
               RECT 9.134 47.158 9.186 47.194 ;
               RECT 9.134 48.358 9.186 48.394 ;
               RECT 9.134 50.142 9.186 50.178 ;
               RECT 9.134 50.382 9.186 50.418 ;
               RECT 9.134 54.702 9.186 54.738 ;
               RECT 9.134 54.942 9.186 54.978 ;
               RECT 9.134 57.478 9.186 57.514 ;
               RECT 9.134 58.678 9.186 58.714 ;
               RECT 9.134 59.878 9.186 59.914 ;
               RECT 9.134 61.078 9.186 61.114 ;
               RECT 9.134 62.278 9.186 62.314 ;
               RECT 9.134 63.478 9.186 63.514 ;
               RECT 9.134 64.678 9.186 64.714 ;
               RECT 9.134 65.878 9.186 65.914 ;
               RECT 9.134 67.078 9.186 67.114 ;
               RECT 9.134 68.278 9.186 68.314 ;
               RECT 9.134 69.478 9.186 69.514 ;
               RECT 9.134 70.678 9.186 70.714 ;
               RECT 9.134 71.878 9.186 71.914 ;
               RECT 9.134 73.078 9.186 73.114 ;
               RECT 9.134 74.278 9.186 74.314 ;
               RECT 9.134 75.478 9.186 75.514 ;
               RECT 9.134 76.678 9.186 76.714 ;
               RECT 9.134 77.878 9.186 77.914 ;
               RECT 9.134 79.078 9.186 79.114 ;
               RECT 9.134 80.278 9.186 80.314 ;
               RECT 9.134 81.478 9.186 81.514 ;
               RECT 9.134 82.678 9.186 82.714 ;
               RECT 9.134 83.878 9.186 83.914 ;
               RECT 9.134 85.078 9.186 85.114 ;
               RECT 9.134 86.278 9.186 86.314 ;
               RECT 9.134 87.478 9.186 87.514 ;
               RECT 9.134 88.678 9.186 88.714 ;
               RECT 9.134 89.878 9.186 89.914 ;
               RECT 9.134 91.078 9.186 91.114 ;
               RECT 9.134 92.278 9.186 92.314 ;
               RECT 9.134 93.478 9.186 93.514 ;
               RECT 9.134 94.678 9.186 94.714 ;
               RECT 9.134 95.878 9.186 95.914 ;
               RECT 9.134 97.078 9.186 97.114 ;
               RECT 9.134 98.278 9.186 98.314 ;
               RECT 9.134 99.478 9.186 99.514 ;
               RECT 9.134 100.678 9.186 100.714 ;
               RECT 9.134 101.878 9.186 101.914 ;
               RECT 9.134 103.078 9.186 103.114 ;
               RECT 9.134 104.278 9.186 104.314 ;
               RECT 9.214 0.806 9.266 0.842 ;
               RECT 9.214 2.006 9.266 2.042 ;
               RECT 9.214 3.206 9.266 3.242 ;
               RECT 9.214 4.406 9.266 4.442 ;
               RECT 9.214 5.606 9.266 5.642 ;
               RECT 9.214 6.806 9.266 6.842 ;
               RECT 9.214 8.006 9.266 8.042 ;
               RECT 9.214 9.206 9.266 9.242 ;
               RECT 9.214 10.406 9.266 10.442 ;
               RECT 9.214 11.606 9.266 11.642 ;
               RECT 9.214 12.806 9.266 12.842 ;
               RECT 9.214 14.006 9.266 14.042 ;
               RECT 9.214 15.206 9.266 15.242 ;
               RECT 9.214 16.406 9.266 16.442 ;
               RECT 9.214 17.606 9.266 17.642 ;
               RECT 9.214 18.806 9.266 18.842 ;
               RECT 9.214 20.006 9.266 20.042 ;
               RECT 9.214 21.206 9.266 21.242 ;
               RECT 9.214 22.406 9.266 22.442 ;
               RECT 9.214 23.606 9.266 23.642 ;
               RECT 9.214 24.806 9.266 24.842 ;
               RECT 9.214 26.006 9.266 26.042 ;
               RECT 9.214 27.206 9.266 27.242 ;
               RECT 9.214 28.406 9.266 28.442 ;
               RECT 9.214 29.606 9.266 29.642 ;
               RECT 9.214 30.806 9.266 30.842 ;
               RECT 9.214 32.006 9.266 32.042 ;
               RECT 9.214 33.206 9.266 33.242 ;
               RECT 9.214 34.406 9.266 34.442 ;
               RECT 9.214 35.606 9.266 35.642 ;
               RECT 9.214 36.806 9.266 36.842 ;
               RECT 9.214 38.006 9.266 38.042 ;
               RECT 9.214 39.206 9.266 39.242 ;
               RECT 9.214 40.406 9.266 40.442 ;
               RECT 9.214 41.606 9.266 41.642 ;
               RECT 9.214 42.806 9.266 42.842 ;
               RECT 9.214 44.006 9.266 44.042 ;
               RECT 9.214 45.206 9.266 45.242 ;
               RECT 9.214 46.406 9.266 46.442 ;
               RECT 9.214 47.606 9.266 47.642 ;
               RECT 9.214 49.422 9.266 49.458 ;
               RECT 9.214 49.662 9.266 49.698 ;
               RECT 9.214 55.422 9.266 55.458 ;
               RECT 9.214 55.662 9.266 55.698 ;
               RECT 9.214 56.726 9.266 56.762 ;
               RECT 9.214 57.926 9.266 57.962 ;
               RECT 9.214 59.126 9.266 59.162 ;
               RECT 9.214 60.326 9.266 60.362 ;
               RECT 9.214 61.526 9.266 61.562 ;
               RECT 9.214 62.726 9.266 62.762 ;
               RECT 9.214 63.926 9.266 63.962 ;
               RECT 9.214 65.126 9.266 65.162 ;
               RECT 9.214 66.326 9.266 66.362 ;
               RECT 9.214 67.526 9.266 67.562 ;
               RECT 9.214 68.726 9.266 68.762 ;
               RECT 9.214 69.926 9.266 69.962 ;
               RECT 9.214 71.126 9.266 71.162 ;
               RECT 9.214 72.326 9.266 72.362 ;
               RECT 9.214 73.526 9.266 73.562 ;
               RECT 9.214 74.726 9.266 74.762 ;
               RECT 9.214 75.926 9.266 75.962 ;
               RECT 9.214 77.126 9.266 77.162 ;
               RECT 9.214 78.326 9.266 78.362 ;
               RECT 9.214 79.526 9.266 79.562 ;
               RECT 9.214 80.726 9.266 80.762 ;
               RECT 9.214 81.926 9.266 81.962 ;
               RECT 9.214 83.126 9.266 83.162 ;
               RECT 9.214 84.326 9.266 84.362 ;
               RECT 9.214 85.526 9.266 85.562 ;
               RECT 9.214 86.726 9.266 86.762 ;
               RECT 9.214 87.926 9.266 87.962 ;
               RECT 9.214 89.126 9.266 89.162 ;
               RECT 9.214 90.326 9.266 90.362 ;
               RECT 9.214 91.526 9.266 91.562 ;
               RECT 9.214 92.726 9.266 92.762 ;
               RECT 9.214 93.926 9.266 93.962 ;
               RECT 9.214 95.126 9.266 95.162 ;
               RECT 9.214 96.326 9.266 96.362 ;
               RECT 9.214 97.526 9.266 97.562 ;
               RECT 9.214 98.726 9.266 98.762 ;
               RECT 9.214 99.926 9.266 99.962 ;
               RECT 9.214 101.126 9.266 101.162 ;
               RECT 9.214 102.326 9.266 102.362 ;
               RECT 9.214 103.526 9.266 103.562 ;
               RECT 9.294 1.558 9.346 1.594 ;
               RECT 9.294 2.758 9.346 2.794 ;
               RECT 9.294 3.958 9.346 3.994 ;
               RECT 9.294 5.158 9.346 5.194 ;
               RECT 9.294 6.358 9.346 6.394 ;
               RECT 9.294 7.558 9.346 7.594 ;
               RECT 9.294 8.758 9.346 8.794 ;
               RECT 9.294 9.958 9.346 9.994 ;
               RECT 9.294 11.158 9.346 11.194 ;
               RECT 9.294 12.358 9.346 12.394 ;
               RECT 9.294 13.558 9.346 13.594 ;
               RECT 9.294 14.758 9.346 14.794 ;
               RECT 9.294 15.958 9.346 15.994 ;
               RECT 9.294 17.158 9.346 17.194 ;
               RECT 9.294 18.358 9.346 18.394 ;
               RECT 9.294 19.558 9.346 19.594 ;
               RECT 9.294 20.758 9.346 20.794 ;
               RECT 9.294 21.958 9.346 21.994 ;
               RECT 9.294 23.158 9.346 23.194 ;
               RECT 9.294 24.358 9.346 24.394 ;
               RECT 9.294 25.558 9.346 25.594 ;
               RECT 9.294 26.758 9.346 26.794 ;
               RECT 9.294 27.958 9.346 27.994 ;
               RECT 9.294 29.158 9.346 29.194 ;
               RECT 9.294 30.358 9.346 30.394 ;
               RECT 9.294 31.558 9.346 31.594 ;
               RECT 9.294 32.758 9.346 32.794 ;
               RECT 9.294 33.958 9.346 33.994 ;
               RECT 9.294 35.158 9.346 35.194 ;
               RECT 9.294 36.358 9.346 36.394 ;
               RECT 9.294 37.558 9.346 37.594 ;
               RECT 9.294 38.758 9.346 38.794 ;
               RECT 9.294 39.958 9.346 39.994 ;
               RECT 9.294 41.158 9.346 41.194 ;
               RECT 9.294 42.358 9.346 42.394 ;
               RECT 9.294 43.558 9.346 43.594 ;
               RECT 9.294 44.758 9.346 44.794 ;
               RECT 9.294 45.958 9.346 45.994 ;
               RECT 9.294 47.158 9.346 47.194 ;
               RECT 9.294 48.358 9.346 48.394 ;
               RECT 9.294 50.142 9.346 50.178 ;
               RECT 9.294 50.382 9.346 50.418 ;
               RECT 9.294 54.702 9.346 54.738 ;
               RECT 9.294 54.942 9.346 54.978 ;
               RECT 9.294 57.478 9.346 57.514 ;
               RECT 9.294 58.678 9.346 58.714 ;
               RECT 9.294 59.878 9.346 59.914 ;
               RECT 9.294 61.078 9.346 61.114 ;
               RECT 9.294 62.278 9.346 62.314 ;
               RECT 9.294 63.478 9.346 63.514 ;
               RECT 9.294 64.678 9.346 64.714 ;
               RECT 9.294 65.878 9.346 65.914 ;
               RECT 9.294 67.078 9.346 67.114 ;
               RECT 9.294 68.278 9.346 68.314 ;
               RECT 9.294 69.478 9.346 69.514 ;
               RECT 9.294 70.678 9.346 70.714 ;
               RECT 9.294 71.878 9.346 71.914 ;
               RECT 9.294 73.078 9.346 73.114 ;
               RECT 9.294 74.278 9.346 74.314 ;
               RECT 9.294 75.478 9.346 75.514 ;
               RECT 9.294 76.678 9.346 76.714 ;
               RECT 9.294 77.878 9.346 77.914 ;
               RECT 9.294 79.078 9.346 79.114 ;
               RECT 9.294 80.278 9.346 80.314 ;
               RECT 9.294 81.478 9.346 81.514 ;
               RECT 9.294 82.678 9.346 82.714 ;
               RECT 9.294 83.878 9.346 83.914 ;
               RECT 9.294 85.078 9.346 85.114 ;
               RECT 9.294 86.278 9.346 86.314 ;
               RECT 9.294 87.478 9.346 87.514 ;
               RECT 9.294 88.678 9.346 88.714 ;
               RECT 9.294 89.878 9.346 89.914 ;
               RECT 9.294 91.078 9.346 91.114 ;
               RECT 9.294 92.278 9.346 92.314 ;
               RECT 9.294 93.478 9.346 93.514 ;
               RECT 9.294 94.678 9.346 94.714 ;
               RECT 9.294 95.878 9.346 95.914 ;
               RECT 9.294 97.078 9.346 97.114 ;
               RECT 9.294 98.278 9.346 98.314 ;
               RECT 9.294 99.478 9.346 99.514 ;
               RECT 9.294 100.678 9.346 100.714 ;
               RECT 9.294 101.878 9.346 101.914 ;
               RECT 9.294 103.078 9.346 103.114 ;
               RECT 9.294 104.278 9.346 104.314 ;
               RECT 9.374 0.281 9.426 0.317 ;
               RECT 9.374 104.803 9.426 104.839 ;
               RECT 9.454 0.806 9.506 0.842 ;
               RECT 9.454 2.006 9.506 2.042 ;
               RECT 9.454 3.206 9.506 3.242 ;
               RECT 9.454 4.406 9.506 4.442 ;
               RECT 9.454 5.606 9.506 5.642 ;
               RECT 9.454 6.806 9.506 6.842 ;
               RECT 9.454 8.006 9.506 8.042 ;
               RECT 9.454 9.206 9.506 9.242 ;
               RECT 9.454 10.406 9.506 10.442 ;
               RECT 9.454 11.606 9.506 11.642 ;
               RECT 9.454 12.806 9.506 12.842 ;
               RECT 9.454 14.006 9.506 14.042 ;
               RECT 9.454 15.206 9.506 15.242 ;
               RECT 9.454 16.406 9.506 16.442 ;
               RECT 9.454 17.606 9.506 17.642 ;
               RECT 9.454 18.806 9.506 18.842 ;
               RECT 9.454 20.006 9.506 20.042 ;
               RECT 9.454 21.206 9.506 21.242 ;
               RECT 9.454 22.406 9.506 22.442 ;
               RECT 9.454 23.606 9.506 23.642 ;
               RECT 9.454 24.806 9.506 24.842 ;
               RECT 9.454 26.006 9.506 26.042 ;
               RECT 9.454 27.206 9.506 27.242 ;
               RECT 9.454 28.406 9.506 28.442 ;
               RECT 9.454 29.606 9.506 29.642 ;
               RECT 9.454 30.806 9.506 30.842 ;
               RECT 9.454 32.006 9.506 32.042 ;
               RECT 9.454 33.206 9.506 33.242 ;
               RECT 9.454 34.406 9.506 34.442 ;
               RECT 9.454 35.606 9.506 35.642 ;
               RECT 9.454 36.806 9.506 36.842 ;
               RECT 9.454 38.006 9.506 38.042 ;
               RECT 9.454 39.206 9.506 39.242 ;
               RECT 9.454 40.406 9.506 40.442 ;
               RECT 9.454 41.606 9.506 41.642 ;
               RECT 9.454 42.806 9.506 42.842 ;
               RECT 9.454 44.006 9.506 44.042 ;
               RECT 9.454 45.206 9.506 45.242 ;
               RECT 9.454 46.406 9.506 46.442 ;
               RECT 9.454 47.606 9.506 47.642 ;
               RECT 9.454 49.422 9.506 49.458 ;
               RECT 9.454 49.662 9.506 49.698 ;
               RECT 9.454 55.422 9.506 55.458 ;
               RECT 9.454 55.662 9.506 55.698 ;
               RECT 9.454 56.726 9.506 56.762 ;
               RECT 9.454 57.926 9.506 57.962 ;
               RECT 9.454 59.126 9.506 59.162 ;
               RECT 9.454 60.326 9.506 60.362 ;
               RECT 9.454 61.526 9.506 61.562 ;
               RECT 9.454 62.726 9.506 62.762 ;
               RECT 9.454 63.926 9.506 63.962 ;
               RECT 9.454 65.126 9.506 65.162 ;
               RECT 9.454 66.326 9.506 66.362 ;
               RECT 9.454 67.526 9.506 67.562 ;
               RECT 9.454 68.726 9.506 68.762 ;
               RECT 9.454 69.926 9.506 69.962 ;
               RECT 9.454 71.126 9.506 71.162 ;
               RECT 9.454 72.326 9.506 72.362 ;
               RECT 9.454 73.526 9.506 73.562 ;
               RECT 9.454 74.726 9.506 74.762 ;
               RECT 9.454 75.926 9.506 75.962 ;
               RECT 9.454 77.126 9.506 77.162 ;
               RECT 9.454 78.326 9.506 78.362 ;
               RECT 9.454 79.526 9.506 79.562 ;
               RECT 9.454 80.726 9.506 80.762 ;
               RECT 9.454 81.926 9.506 81.962 ;
               RECT 9.454 83.126 9.506 83.162 ;
               RECT 9.454 84.326 9.506 84.362 ;
               RECT 9.454 85.526 9.506 85.562 ;
               RECT 9.454 86.726 9.506 86.762 ;
               RECT 9.454 87.926 9.506 87.962 ;
               RECT 9.454 89.126 9.506 89.162 ;
               RECT 9.454 90.326 9.506 90.362 ;
               RECT 9.454 91.526 9.506 91.562 ;
               RECT 9.454 92.726 9.506 92.762 ;
               RECT 9.454 93.926 9.506 93.962 ;
               RECT 9.454 95.126 9.506 95.162 ;
               RECT 9.454 96.326 9.506 96.362 ;
               RECT 9.454 97.526 9.506 97.562 ;
               RECT 9.454 98.726 9.506 98.762 ;
               RECT 9.454 99.926 9.506 99.962 ;
               RECT 9.454 101.126 9.506 101.162 ;
               RECT 9.454 102.326 9.506 102.362 ;
               RECT 9.454 103.526 9.506 103.562 ;
               RECT 9.534 1.558 9.586 1.594 ;
               RECT 9.534 2.758 9.586 2.794 ;
               RECT 9.534 3.958 9.586 3.994 ;
               RECT 9.534 5.158 9.586 5.194 ;
               RECT 9.534 6.358 9.586 6.394 ;
               RECT 9.534 7.558 9.586 7.594 ;
               RECT 9.534 8.758 9.586 8.794 ;
               RECT 9.534 9.958 9.586 9.994 ;
               RECT 9.534 11.158 9.586 11.194 ;
               RECT 9.534 12.358 9.586 12.394 ;
               RECT 9.534 13.558 9.586 13.594 ;
               RECT 9.534 14.758 9.586 14.794 ;
               RECT 9.534 15.958 9.586 15.994 ;
               RECT 9.534 17.158 9.586 17.194 ;
               RECT 9.534 18.358 9.586 18.394 ;
               RECT 9.534 19.558 9.586 19.594 ;
               RECT 9.534 20.758 9.586 20.794 ;
               RECT 9.534 21.958 9.586 21.994 ;
               RECT 9.534 23.158 9.586 23.194 ;
               RECT 9.534 24.358 9.586 24.394 ;
               RECT 9.534 25.558 9.586 25.594 ;
               RECT 9.534 26.758 9.586 26.794 ;
               RECT 9.534 27.958 9.586 27.994 ;
               RECT 9.534 29.158 9.586 29.194 ;
               RECT 9.534 30.358 9.586 30.394 ;
               RECT 9.534 31.558 9.586 31.594 ;
               RECT 9.534 32.758 9.586 32.794 ;
               RECT 9.534 33.958 9.586 33.994 ;
               RECT 9.534 35.158 9.586 35.194 ;
               RECT 9.534 36.358 9.586 36.394 ;
               RECT 9.534 37.558 9.586 37.594 ;
               RECT 9.534 38.758 9.586 38.794 ;
               RECT 9.534 39.958 9.586 39.994 ;
               RECT 9.534 41.158 9.586 41.194 ;
               RECT 9.534 42.358 9.586 42.394 ;
               RECT 9.534 43.558 9.586 43.594 ;
               RECT 9.534 44.758 9.586 44.794 ;
               RECT 9.534 45.958 9.586 45.994 ;
               RECT 9.534 47.158 9.586 47.194 ;
               RECT 9.534 48.358 9.586 48.394 ;
               RECT 9.534 50.142 9.586 50.178 ;
               RECT 9.534 50.382 9.586 50.418 ;
               RECT 9.534 54.702 9.586 54.738 ;
               RECT 9.534 54.942 9.586 54.978 ;
               RECT 9.534 57.478 9.586 57.514 ;
               RECT 9.534 58.678 9.586 58.714 ;
               RECT 9.534 59.878 9.586 59.914 ;
               RECT 9.534 61.078 9.586 61.114 ;
               RECT 9.534 62.278 9.586 62.314 ;
               RECT 9.534 63.478 9.586 63.514 ;
               RECT 9.534 64.678 9.586 64.714 ;
               RECT 9.534 65.878 9.586 65.914 ;
               RECT 9.534 67.078 9.586 67.114 ;
               RECT 9.534 68.278 9.586 68.314 ;
               RECT 9.534 69.478 9.586 69.514 ;
               RECT 9.534 70.678 9.586 70.714 ;
               RECT 9.534 71.878 9.586 71.914 ;
               RECT 9.534 73.078 9.586 73.114 ;
               RECT 9.534 74.278 9.586 74.314 ;
               RECT 9.534 75.478 9.586 75.514 ;
               RECT 9.534 76.678 9.586 76.714 ;
               RECT 9.534 77.878 9.586 77.914 ;
               RECT 9.534 79.078 9.586 79.114 ;
               RECT 9.534 80.278 9.586 80.314 ;
               RECT 9.534 81.478 9.586 81.514 ;
               RECT 9.534 82.678 9.586 82.714 ;
               RECT 9.534 83.878 9.586 83.914 ;
               RECT 9.534 85.078 9.586 85.114 ;
               RECT 9.534 86.278 9.586 86.314 ;
               RECT 9.534 87.478 9.586 87.514 ;
               RECT 9.534 88.678 9.586 88.714 ;
               RECT 9.534 89.878 9.586 89.914 ;
               RECT 9.534 91.078 9.586 91.114 ;
               RECT 9.534 92.278 9.586 92.314 ;
               RECT 9.534 93.478 9.586 93.514 ;
               RECT 9.534 94.678 9.586 94.714 ;
               RECT 9.534 95.878 9.586 95.914 ;
               RECT 9.534 97.078 9.586 97.114 ;
               RECT 9.534 98.278 9.586 98.314 ;
               RECT 9.534 99.478 9.586 99.514 ;
               RECT 9.534 100.678 9.586 100.714 ;
               RECT 9.534 101.878 9.586 101.914 ;
               RECT 9.534 103.078 9.586 103.114 ;
               RECT 9.534 104.278 9.586 104.314 ;
               RECT 9.614 0.806 9.666 0.842 ;
               RECT 9.614 2.006 9.666 2.042 ;
               RECT 9.614 3.206 9.666 3.242 ;
               RECT 9.614 4.406 9.666 4.442 ;
               RECT 9.614 5.606 9.666 5.642 ;
               RECT 9.614 6.806 9.666 6.842 ;
               RECT 9.614 8.006 9.666 8.042 ;
               RECT 9.614 9.206 9.666 9.242 ;
               RECT 9.614 10.406 9.666 10.442 ;
               RECT 9.614 11.606 9.666 11.642 ;
               RECT 9.614 12.806 9.666 12.842 ;
               RECT 9.614 14.006 9.666 14.042 ;
               RECT 9.614 15.206 9.666 15.242 ;
               RECT 9.614 16.406 9.666 16.442 ;
               RECT 9.614 17.606 9.666 17.642 ;
               RECT 9.614 18.806 9.666 18.842 ;
               RECT 9.614 20.006 9.666 20.042 ;
               RECT 9.614 21.206 9.666 21.242 ;
               RECT 9.614 22.406 9.666 22.442 ;
               RECT 9.614 23.606 9.666 23.642 ;
               RECT 9.614 24.806 9.666 24.842 ;
               RECT 9.614 26.006 9.666 26.042 ;
               RECT 9.614 27.206 9.666 27.242 ;
               RECT 9.614 28.406 9.666 28.442 ;
               RECT 9.614 29.606 9.666 29.642 ;
               RECT 9.614 30.806 9.666 30.842 ;
               RECT 9.614 32.006 9.666 32.042 ;
               RECT 9.614 33.206 9.666 33.242 ;
               RECT 9.614 34.406 9.666 34.442 ;
               RECT 9.614 35.606 9.666 35.642 ;
               RECT 9.614 36.806 9.666 36.842 ;
               RECT 9.614 38.006 9.666 38.042 ;
               RECT 9.614 39.206 9.666 39.242 ;
               RECT 9.614 40.406 9.666 40.442 ;
               RECT 9.614 41.606 9.666 41.642 ;
               RECT 9.614 42.806 9.666 42.842 ;
               RECT 9.614 44.006 9.666 44.042 ;
               RECT 9.614 45.206 9.666 45.242 ;
               RECT 9.614 46.406 9.666 46.442 ;
               RECT 9.614 47.606 9.666 47.642 ;
               RECT 9.614 49.422 9.666 49.458 ;
               RECT 9.614 49.662 9.666 49.698 ;
               RECT 9.614 55.422 9.666 55.458 ;
               RECT 9.614 55.662 9.666 55.698 ;
               RECT 9.614 56.726 9.666 56.762 ;
               RECT 9.614 57.926 9.666 57.962 ;
               RECT 9.614 59.126 9.666 59.162 ;
               RECT 9.614 60.326 9.666 60.362 ;
               RECT 9.614 61.526 9.666 61.562 ;
               RECT 9.614 62.726 9.666 62.762 ;
               RECT 9.614 63.926 9.666 63.962 ;
               RECT 9.614 65.126 9.666 65.162 ;
               RECT 9.614 66.326 9.666 66.362 ;
               RECT 9.614 67.526 9.666 67.562 ;
               RECT 9.614 68.726 9.666 68.762 ;
               RECT 9.614 69.926 9.666 69.962 ;
               RECT 9.614 71.126 9.666 71.162 ;
               RECT 9.614 72.326 9.666 72.362 ;
               RECT 9.614 73.526 9.666 73.562 ;
               RECT 9.614 74.726 9.666 74.762 ;
               RECT 9.614 75.926 9.666 75.962 ;
               RECT 9.614 77.126 9.666 77.162 ;
               RECT 9.614 78.326 9.666 78.362 ;
               RECT 9.614 79.526 9.666 79.562 ;
               RECT 9.614 80.726 9.666 80.762 ;
               RECT 9.614 81.926 9.666 81.962 ;
               RECT 9.614 83.126 9.666 83.162 ;
               RECT 9.614 84.326 9.666 84.362 ;
               RECT 9.614 85.526 9.666 85.562 ;
               RECT 9.614 86.726 9.666 86.762 ;
               RECT 9.614 87.926 9.666 87.962 ;
               RECT 9.614 89.126 9.666 89.162 ;
               RECT 9.614 90.326 9.666 90.362 ;
               RECT 9.614 91.526 9.666 91.562 ;
               RECT 9.614 92.726 9.666 92.762 ;
               RECT 9.614 93.926 9.666 93.962 ;
               RECT 9.614 95.126 9.666 95.162 ;
               RECT 9.614 96.326 9.666 96.362 ;
               RECT 9.614 97.526 9.666 97.562 ;
               RECT 9.614 98.726 9.666 98.762 ;
               RECT 9.614 99.926 9.666 99.962 ;
               RECT 9.614 101.126 9.666 101.162 ;
               RECT 9.614 102.326 9.666 102.362 ;
               RECT 9.614 103.526 9.666 103.562 ;
               RECT 9.694 1.558 9.746 1.594 ;
               RECT 9.694 2.758 9.746 2.794 ;
               RECT 9.694 3.958 9.746 3.994 ;
               RECT 9.694 5.158 9.746 5.194 ;
               RECT 9.694 6.358 9.746 6.394 ;
               RECT 9.694 7.558 9.746 7.594 ;
               RECT 9.694 8.758 9.746 8.794 ;
               RECT 9.694 9.958 9.746 9.994 ;
               RECT 9.694 11.158 9.746 11.194 ;
               RECT 9.694 12.358 9.746 12.394 ;
               RECT 9.694 13.558 9.746 13.594 ;
               RECT 9.694 14.758 9.746 14.794 ;
               RECT 9.694 15.958 9.746 15.994 ;
               RECT 9.694 17.158 9.746 17.194 ;
               RECT 9.694 18.358 9.746 18.394 ;
               RECT 9.694 19.558 9.746 19.594 ;
               RECT 9.694 20.758 9.746 20.794 ;
               RECT 9.694 21.958 9.746 21.994 ;
               RECT 9.694 23.158 9.746 23.194 ;
               RECT 9.694 24.358 9.746 24.394 ;
               RECT 9.694 25.558 9.746 25.594 ;
               RECT 9.694 26.758 9.746 26.794 ;
               RECT 9.694 27.958 9.746 27.994 ;
               RECT 9.694 29.158 9.746 29.194 ;
               RECT 9.694 30.358 9.746 30.394 ;
               RECT 9.694 31.558 9.746 31.594 ;
               RECT 9.694 32.758 9.746 32.794 ;
               RECT 9.694 33.958 9.746 33.994 ;
               RECT 9.694 35.158 9.746 35.194 ;
               RECT 9.694 36.358 9.746 36.394 ;
               RECT 9.694 37.558 9.746 37.594 ;
               RECT 9.694 38.758 9.746 38.794 ;
               RECT 9.694 39.958 9.746 39.994 ;
               RECT 9.694 41.158 9.746 41.194 ;
               RECT 9.694 42.358 9.746 42.394 ;
               RECT 9.694 43.558 9.746 43.594 ;
               RECT 9.694 44.758 9.746 44.794 ;
               RECT 9.694 45.958 9.746 45.994 ;
               RECT 9.694 47.158 9.746 47.194 ;
               RECT 9.694 48.358 9.746 48.394 ;
               RECT 9.694 50.142 9.746 50.178 ;
               RECT 9.694 50.382 9.746 50.418 ;
               RECT 9.694 54.702 9.746 54.738 ;
               RECT 9.694 54.942 9.746 54.978 ;
               RECT 9.694 57.478 9.746 57.514 ;
               RECT 9.694 58.678 9.746 58.714 ;
               RECT 9.694 59.878 9.746 59.914 ;
               RECT 9.694 61.078 9.746 61.114 ;
               RECT 9.694 62.278 9.746 62.314 ;
               RECT 9.694 63.478 9.746 63.514 ;
               RECT 9.694 64.678 9.746 64.714 ;
               RECT 9.694 65.878 9.746 65.914 ;
               RECT 9.694 67.078 9.746 67.114 ;
               RECT 9.694 68.278 9.746 68.314 ;
               RECT 9.694 69.478 9.746 69.514 ;
               RECT 9.694 70.678 9.746 70.714 ;
               RECT 9.694 71.878 9.746 71.914 ;
               RECT 9.694 73.078 9.746 73.114 ;
               RECT 9.694 74.278 9.746 74.314 ;
               RECT 9.694 75.478 9.746 75.514 ;
               RECT 9.694 76.678 9.746 76.714 ;
               RECT 9.694 77.878 9.746 77.914 ;
               RECT 9.694 79.078 9.746 79.114 ;
               RECT 9.694 80.278 9.746 80.314 ;
               RECT 9.694 81.478 9.746 81.514 ;
               RECT 9.694 82.678 9.746 82.714 ;
               RECT 9.694 83.878 9.746 83.914 ;
               RECT 9.694 85.078 9.746 85.114 ;
               RECT 9.694 86.278 9.746 86.314 ;
               RECT 9.694 87.478 9.746 87.514 ;
               RECT 9.694 88.678 9.746 88.714 ;
               RECT 9.694 89.878 9.746 89.914 ;
               RECT 9.694 91.078 9.746 91.114 ;
               RECT 9.694 92.278 9.746 92.314 ;
               RECT 9.694 93.478 9.746 93.514 ;
               RECT 9.694 94.678 9.746 94.714 ;
               RECT 9.694 95.878 9.746 95.914 ;
               RECT 9.694 97.078 9.746 97.114 ;
               RECT 9.694 98.278 9.746 98.314 ;
               RECT 9.694 99.478 9.746 99.514 ;
               RECT 9.694 100.678 9.746 100.714 ;
               RECT 9.694 101.878 9.746 101.914 ;
               RECT 9.694 103.078 9.746 103.114 ;
               RECT 9.694 104.278 9.746 104.314 ;
               RECT 9.774 0.281 9.826 0.317 ;
               RECT 9.774 104.803 9.826 104.839 ;
               RECT 9.854 0.806 9.906 0.842 ;
               RECT 9.854 2.006 9.906 2.042 ;
               RECT 9.854 3.206 9.906 3.242 ;
               RECT 9.854 4.406 9.906 4.442 ;
               RECT 9.854 5.606 9.906 5.642 ;
               RECT 9.854 6.806 9.906 6.842 ;
               RECT 9.854 8.006 9.906 8.042 ;
               RECT 9.854 9.206 9.906 9.242 ;
               RECT 9.854 10.406 9.906 10.442 ;
               RECT 9.854 11.606 9.906 11.642 ;
               RECT 9.854 12.806 9.906 12.842 ;
               RECT 9.854 14.006 9.906 14.042 ;
               RECT 9.854 15.206 9.906 15.242 ;
               RECT 9.854 16.406 9.906 16.442 ;
               RECT 9.854 17.606 9.906 17.642 ;
               RECT 9.854 18.806 9.906 18.842 ;
               RECT 9.854 20.006 9.906 20.042 ;
               RECT 9.854 21.206 9.906 21.242 ;
               RECT 9.854 22.406 9.906 22.442 ;
               RECT 9.854 23.606 9.906 23.642 ;
               RECT 9.854 24.806 9.906 24.842 ;
               RECT 9.854 26.006 9.906 26.042 ;
               RECT 9.854 27.206 9.906 27.242 ;
               RECT 9.854 28.406 9.906 28.442 ;
               RECT 9.854 29.606 9.906 29.642 ;
               RECT 9.854 30.806 9.906 30.842 ;
               RECT 9.854 32.006 9.906 32.042 ;
               RECT 9.854 33.206 9.906 33.242 ;
               RECT 9.854 34.406 9.906 34.442 ;
               RECT 9.854 35.606 9.906 35.642 ;
               RECT 9.854 36.806 9.906 36.842 ;
               RECT 9.854 38.006 9.906 38.042 ;
               RECT 9.854 39.206 9.906 39.242 ;
               RECT 9.854 40.406 9.906 40.442 ;
               RECT 9.854 41.606 9.906 41.642 ;
               RECT 9.854 42.806 9.906 42.842 ;
               RECT 9.854 44.006 9.906 44.042 ;
               RECT 9.854 45.206 9.906 45.242 ;
               RECT 9.854 46.406 9.906 46.442 ;
               RECT 9.854 47.606 9.906 47.642 ;
               RECT 9.854 49.422 9.906 49.458 ;
               RECT 9.854 49.662 9.906 49.698 ;
               RECT 9.854 51.102 9.906 51.138 ;
               RECT 9.854 51.582 9.906 51.618 ;
               RECT 9.854 53.502 9.906 53.538 ;
               RECT 9.854 53.982 9.906 54.018 ;
               RECT 9.854 55.422 9.906 55.458 ;
               RECT 9.854 55.662 9.906 55.698 ;
               RECT 9.854 56.726 9.906 56.762 ;
               RECT 9.854 57.926 9.906 57.962 ;
               RECT 9.854 59.126 9.906 59.162 ;
               RECT 9.854 60.326 9.906 60.362 ;
               RECT 9.854 61.526 9.906 61.562 ;
               RECT 9.854 62.726 9.906 62.762 ;
               RECT 9.854 63.926 9.906 63.962 ;
               RECT 9.854 65.126 9.906 65.162 ;
               RECT 9.854 66.326 9.906 66.362 ;
               RECT 9.854 67.526 9.906 67.562 ;
               RECT 9.854 68.726 9.906 68.762 ;
               RECT 9.854 69.926 9.906 69.962 ;
               RECT 9.854 71.126 9.906 71.162 ;
               RECT 9.854 72.326 9.906 72.362 ;
               RECT 9.854 73.526 9.906 73.562 ;
               RECT 9.854 74.726 9.906 74.762 ;
               RECT 9.854 75.926 9.906 75.962 ;
               RECT 9.854 77.126 9.906 77.162 ;
               RECT 9.854 78.326 9.906 78.362 ;
               RECT 9.854 79.526 9.906 79.562 ;
               RECT 9.854 80.726 9.906 80.762 ;
               RECT 9.854 81.926 9.906 81.962 ;
               RECT 9.854 83.126 9.906 83.162 ;
               RECT 9.854 84.326 9.906 84.362 ;
               RECT 9.854 85.526 9.906 85.562 ;
               RECT 9.854 86.726 9.906 86.762 ;
               RECT 9.854 87.926 9.906 87.962 ;
               RECT 9.854 89.126 9.906 89.162 ;
               RECT 9.854 90.326 9.906 90.362 ;
               RECT 9.854 91.526 9.906 91.562 ;
               RECT 9.854 92.726 9.906 92.762 ;
               RECT 9.854 93.926 9.906 93.962 ;
               RECT 9.854 95.126 9.906 95.162 ;
               RECT 9.854 96.326 9.906 96.362 ;
               RECT 9.854 97.526 9.906 97.562 ;
               RECT 9.854 98.726 9.906 98.762 ;
               RECT 9.854 99.926 9.906 99.962 ;
               RECT 9.854 101.126 9.906 101.162 ;
               RECT 9.854 102.326 9.906 102.362 ;
               RECT 9.854 103.526 9.906 103.562 ;
               RECT 9.934 1.558 9.986 1.594 ;
               RECT 9.934 2.758 9.986 2.794 ;
               RECT 9.934 3.958 9.986 3.994 ;
               RECT 9.934 5.158 9.986 5.194 ;
               RECT 9.934 6.358 9.986 6.394 ;
               RECT 9.934 7.558 9.986 7.594 ;
               RECT 9.934 8.758 9.986 8.794 ;
               RECT 9.934 9.958 9.986 9.994 ;
               RECT 9.934 11.158 9.986 11.194 ;
               RECT 9.934 12.358 9.986 12.394 ;
               RECT 9.934 13.558 9.986 13.594 ;
               RECT 9.934 14.758 9.986 14.794 ;
               RECT 9.934 15.958 9.986 15.994 ;
               RECT 9.934 17.158 9.986 17.194 ;
               RECT 9.934 18.358 9.986 18.394 ;
               RECT 9.934 19.558 9.986 19.594 ;
               RECT 9.934 20.758 9.986 20.794 ;
               RECT 9.934 21.958 9.986 21.994 ;
               RECT 9.934 23.158 9.986 23.194 ;
               RECT 9.934 24.358 9.986 24.394 ;
               RECT 9.934 25.558 9.986 25.594 ;
               RECT 9.934 26.758 9.986 26.794 ;
               RECT 9.934 27.958 9.986 27.994 ;
               RECT 9.934 29.158 9.986 29.194 ;
               RECT 9.934 30.358 9.986 30.394 ;
               RECT 9.934 31.558 9.986 31.594 ;
               RECT 9.934 32.758 9.986 32.794 ;
               RECT 9.934 33.958 9.986 33.994 ;
               RECT 9.934 35.158 9.986 35.194 ;
               RECT 9.934 36.358 9.986 36.394 ;
               RECT 9.934 37.558 9.986 37.594 ;
               RECT 9.934 38.758 9.986 38.794 ;
               RECT 9.934 39.958 9.986 39.994 ;
               RECT 9.934 41.158 9.986 41.194 ;
               RECT 9.934 42.358 9.986 42.394 ;
               RECT 9.934 43.558 9.986 43.594 ;
               RECT 9.934 44.758 9.986 44.794 ;
               RECT 9.934 45.958 9.986 45.994 ;
               RECT 9.934 47.158 9.986 47.194 ;
               RECT 9.934 48.358 9.986 48.394 ;
               RECT 9.934 50.142 9.986 50.178 ;
               RECT 9.934 50.382 9.986 50.418 ;
               RECT 9.934 54.702 9.986 54.738 ;
               RECT 9.934 54.942 9.986 54.978 ;
               RECT 9.934 57.478 9.986 57.514 ;
               RECT 9.934 58.678 9.986 58.714 ;
               RECT 9.934 59.878 9.986 59.914 ;
               RECT 9.934 61.078 9.986 61.114 ;
               RECT 9.934 62.278 9.986 62.314 ;
               RECT 9.934 63.478 9.986 63.514 ;
               RECT 9.934 64.678 9.986 64.714 ;
               RECT 9.934 65.878 9.986 65.914 ;
               RECT 9.934 67.078 9.986 67.114 ;
               RECT 9.934 68.278 9.986 68.314 ;
               RECT 9.934 69.478 9.986 69.514 ;
               RECT 9.934 70.678 9.986 70.714 ;
               RECT 9.934 71.878 9.986 71.914 ;
               RECT 9.934 73.078 9.986 73.114 ;
               RECT 9.934 74.278 9.986 74.314 ;
               RECT 9.934 75.478 9.986 75.514 ;
               RECT 9.934 76.678 9.986 76.714 ;
               RECT 9.934 77.878 9.986 77.914 ;
               RECT 9.934 79.078 9.986 79.114 ;
               RECT 9.934 80.278 9.986 80.314 ;
               RECT 9.934 81.478 9.986 81.514 ;
               RECT 9.934 82.678 9.986 82.714 ;
               RECT 9.934 83.878 9.986 83.914 ;
               RECT 9.934 85.078 9.986 85.114 ;
               RECT 9.934 86.278 9.986 86.314 ;
               RECT 9.934 87.478 9.986 87.514 ;
               RECT 9.934 88.678 9.986 88.714 ;
               RECT 9.934 89.878 9.986 89.914 ;
               RECT 9.934 91.078 9.986 91.114 ;
               RECT 9.934 92.278 9.986 92.314 ;
               RECT 9.934 93.478 9.986 93.514 ;
               RECT 9.934 94.678 9.986 94.714 ;
               RECT 9.934 95.878 9.986 95.914 ;
               RECT 9.934 97.078 9.986 97.114 ;
               RECT 9.934 98.278 9.986 98.314 ;
               RECT 9.934 99.478 9.986 99.514 ;
               RECT 9.934 100.678 9.986 100.714 ;
               RECT 9.934 101.878 9.986 101.914 ;
               RECT 9.934 103.078 9.986 103.114 ;
               RECT 9.934 104.278 9.986 104.314 ;
               RECT 10.014 0.806 10.066 0.842 ;
               RECT 10.014 2.006 10.066 2.042 ;
               RECT 10.014 3.206 10.066 3.242 ;
               RECT 10.014 4.406 10.066 4.442 ;
               RECT 10.014 5.606 10.066 5.642 ;
               RECT 10.014 6.806 10.066 6.842 ;
               RECT 10.014 8.006 10.066 8.042 ;
               RECT 10.014 9.206 10.066 9.242 ;
               RECT 10.014 10.406 10.066 10.442 ;
               RECT 10.014 11.606 10.066 11.642 ;
               RECT 10.014 12.806 10.066 12.842 ;
               RECT 10.014 14.006 10.066 14.042 ;
               RECT 10.014 15.206 10.066 15.242 ;
               RECT 10.014 16.406 10.066 16.442 ;
               RECT 10.014 17.606 10.066 17.642 ;
               RECT 10.014 18.806 10.066 18.842 ;
               RECT 10.014 20.006 10.066 20.042 ;
               RECT 10.014 21.206 10.066 21.242 ;
               RECT 10.014 22.406 10.066 22.442 ;
               RECT 10.014 23.606 10.066 23.642 ;
               RECT 10.014 24.806 10.066 24.842 ;
               RECT 10.014 26.006 10.066 26.042 ;
               RECT 10.014 27.206 10.066 27.242 ;
               RECT 10.014 28.406 10.066 28.442 ;
               RECT 10.014 29.606 10.066 29.642 ;
               RECT 10.014 30.806 10.066 30.842 ;
               RECT 10.014 32.006 10.066 32.042 ;
               RECT 10.014 33.206 10.066 33.242 ;
               RECT 10.014 34.406 10.066 34.442 ;
               RECT 10.014 35.606 10.066 35.642 ;
               RECT 10.014 36.806 10.066 36.842 ;
               RECT 10.014 38.006 10.066 38.042 ;
               RECT 10.014 39.206 10.066 39.242 ;
               RECT 10.014 40.406 10.066 40.442 ;
               RECT 10.014 41.606 10.066 41.642 ;
               RECT 10.014 42.806 10.066 42.842 ;
               RECT 10.014 44.006 10.066 44.042 ;
               RECT 10.014 45.206 10.066 45.242 ;
               RECT 10.014 46.406 10.066 46.442 ;
               RECT 10.014 47.606 10.066 47.642 ;
               RECT 10.014 49.422 10.066 49.458 ;
               RECT 10.014 49.662 10.066 49.698 ;
               RECT 10.014 55.422 10.066 55.458 ;
               RECT 10.014 55.662 10.066 55.698 ;
               RECT 10.014 56.726 10.066 56.762 ;
               RECT 10.014 57.926 10.066 57.962 ;
               RECT 10.014 59.126 10.066 59.162 ;
               RECT 10.014 60.326 10.066 60.362 ;
               RECT 10.014 61.526 10.066 61.562 ;
               RECT 10.014 62.726 10.066 62.762 ;
               RECT 10.014 63.926 10.066 63.962 ;
               RECT 10.014 65.126 10.066 65.162 ;
               RECT 10.014 66.326 10.066 66.362 ;
               RECT 10.014 67.526 10.066 67.562 ;
               RECT 10.014 68.726 10.066 68.762 ;
               RECT 10.014 69.926 10.066 69.962 ;
               RECT 10.014 71.126 10.066 71.162 ;
               RECT 10.014 72.326 10.066 72.362 ;
               RECT 10.014 73.526 10.066 73.562 ;
               RECT 10.014 74.726 10.066 74.762 ;
               RECT 10.014 75.926 10.066 75.962 ;
               RECT 10.014 77.126 10.066 77.162 ;
               RECT 10.014 78.326 10.066 78.362 ;
               RECT 10.014 79.526 10.066 79.562 ;
               RECT 10.014 80.726 10.066 80.762 ;
               RECT 10.014 81.926 10.066 81.962 ;
               RECT 10.014 83.126 10.066 83.162 ;
               RECT 10.014 84.326 10.066 84.362 ;
               RECT 10.014 85.526 10.066 85.562 ;
               RECT 10.014 86.726 10.066 86.762 ;
               RECT 10.014 87.926 10.066 87.962 ;
               RECT 10.014 89.126 10.066 89.162 ;
               RECT 10.014 90.326 10.066 90.362 ;
               RECT 10.014 91.526 10.066 91.562 ;
               RECT 10.014 92.726 10.066 92.762 ;
               RECT 10.014 93.926 10.066 93.962 ;
               RECT 10.014 95.126 10.066 95.162 ;
               RECT 10.014 96.326 10.066 96.362 ;
               RECT 10.014 97.526 10.066 97.562 ;
               RECT 10.014 98.726 10.066 98.762 ;
               RECT 10.014 99.926 10.066 99.962 ;
               RECT 10.014 101.126 10.066 101.162 ;
               RECT 10.014 102.326 10.066 102.362 ;
               RECT 10.014 103.526 10.066 103.562 ;
               RECT 10.094 1.558 10.146 1.594 ;
               RECT 10.094 2.758 10.146 2.794 ;
               RECT 10.094 3.958 10.146 3.994 ;
               RECT 10.094 5.158 10.146 5.194 ;
               RECT 10.094 6.358 10.146 6.394 ;
               RECT 10.094 7.558 10.146 7.594 ;
               RECT 10.094 8.758 10.146 8.794 ;
               RECT 10.094 9.958 10.146 9.994 ;
               RECT 10.094 11.158 10.146 11.194 ;
               RECT 10.094 12.358 10.146 12.394 ;
               RECT 10.094 13.558 10.146 13.594 ;
               RECT 10.094 14.758 10.146 14.794 ;
               RECT 10.094 15.958 10.146 15.994 ;
               RECT 10.094 17.158 10.146 17.194 ;
               RECT 10.094 18.358 10.146 18.394 ;
               RECT 10.094 19.558 10.146 19.594 ;
               RECT 10.094 20.758 10.146 20.794 ;
               RECT 10.094 21.958 10.146 21.994 ;
               RECT 10.094 23.158 10.146 23.194 ;
               RECT 10.094 24.358 10.146 24.394 ;
               RECT 10.094 25.558 10.146 25.594 ;
               RECT 10.094 26.758 10.146 26.794 ;
               RECT 10.094 27.958 10.146 27.994 ;
               RECT 10.094 29.158 10.146 29.194 ;
               RECT 10.094 30.358 10.146 30.394 ;
               RECT 10.094 31.558 10.146 31.594 ;
               RECT 10.094 32.758 10.146 32.794 ;
               RECT 10.094 33.958 10.146 33.994 ;
               RECT 10.094 35.158 10.146 35.194 ;
               RECT 10.094 36.358 10.146 36.394 ;
               RECT 10.094 37.558 10.146 37.594 ;
               RECT 10.094 38.758 10.146 38.794 ;
               RECT 10.094 39.958 10.146 39.994 ;
               RECT 10.094 41.158 10.146 41.194 ;
               RECT 10.094 42.358 10.146 42.394 ;
               RECT 10.094 43.558 10.146 43.594 ;
               RECT 10.094 44.758 10.146 44.794 ;
               RECT 10.094 45.958 10.146 45.994 ;
               RECT 10.094 47.158 10.146 47.194 ;
               RECT 10.094 48.358 10.146 48.394 ;
               RECT 10.094 50.142 10.146 50.178 ;
               RECT 10.094 50.382 10.146 50.418 ;
               RECT 10.094 54.702 10.146 54.738 ;
               RECT 10.094 54.942 10.146 54.978 ;
               RECT 10.094 57.478 10.146 57.514 ;
               RECT 10.094 58.678 10.146 58.714 ;
               RECT 10.094 59.878 10.146 59.914 ;
               RECT 10.094 61.078 10.146 61.114 ;
               RECT 10.094 62.278 10.146 62.314 ;
               RECT 10.094 63.478 10.146 63.514 ;
               RECT 10.094 64.678 10.146 64.714 ;
               RECT 10.094 65.878 10.146 65.914 ;
               RECT 10.094 67.078 10.146 67.114 ;
               RECT 10.094 68.278 10.146 68.314 ;
               RECT 10.094 69.478 10.146 69.514 ;
               RECT 10.094 70.678 10.146 70.714 ;
               RECT 10.094 71.878 10.146 71.914 ;
               RECT 10.094 73.078 10.146 73.114 ;
               RECT 10.094 74.278 10.146 74.314 ;
               RECT 10.094 75.478 10.146 75.514 ;
               RECT 10.094 76.678 10.146 76.714 ;
               RECT 10.094 77.878 10.146 77.914 ;
               RECT 10.094 79.078 10.146 79.114 ;
               RECT 10.094 80.278 10.146 80.314 ;
               RECT 10.094 81.478 10.146 81.514 ;
               RECT 10.094 82.678 10.146 82.714 ;
               RECT 10.094 83.878 10.146 83.914 ;
               RECT 10.094 85.078 10.146 85.114 ;
               RECT 10.094 86.278 10.146 86.314 ;
               RECT 10.094 87.478 10.146 87.514 ;
               RECT 10.094 88.678 10.146 88.714 ;
               RECT 10.094 89.878 10.146 89.914 ;
               RECT 10.094 91.078 10.146 91.114 ;
               RECT 10.094 92.278 10.146 92.314 ;
               RECT 10.094 93.478 10.146 93.514 ;
               RECT 10.094 94.678 10.146 94.714 ;
               RECT 10.094 95.878 10.146 95.914 ;
               RECT 10.094 97.078 10.146 97.114 ;
               RECT 10.094 98.278 10.146 98.314 ;
               RECT 10.094 99.478 10.146 99.514 ;
               RECT 10.094 100.678 10.146 100.714 ;
               RECT 10.094 101.878 10.146 101.914 ;
               RECT 10.094 103.078 10.146 103.114 ;
               RECT 10.094 104.278 10.146 104.314 ;
               RECT 10.174 0.281 10.226 0.317 ;
               RECT 10.174 104.803 10.226 104.839 ;
               RECT 10.254 0.806 10.306 0.842 ;
               RECT 10.254 2.006 10.306 2.042 ;
               RECT 10.254 3.206 10.306 3.242 ;
               RECT 10.254 4.406 10.306 4.442 ;
               RECT 10.254 5.606 10.306 5.642 ;
               RECT 10.254 6.806 10.306 6.842 ;
               RECT 10.254 8.006 10.306 8.042 ;
               RECT 10.254 9.206 10.306 9.242 ;
               RECT 10.254 10.406 10.306 10.442 ;
               RECT 10.254 11.606 10.306 11.642 ;
               RECT 10.254 12.806 10.306 12.842 ;
               RECT 10.254 14.006 10.306 14.042 ;
               RECT 10.254 15.206 10.306 15.242 ;
               RECT 10.254 16.406 10.306 16.442 ;
               RECT 10.254 17.606 10.306 17.642 ;
               RECT 10.254 18.806 10.306 18.842 ;
               RECT 10.254 20.006 10.306 20.042 ;
               RECT 10.254 21.206 10.306 21.242 ;
               RECT 10.254 22.406 10.306 22.442 ;
               RECT 10.254 23.606 10.306 23.642 ;
               RECT 10.254 24.806 10.306 24.842 ;
               RECT 10.254 26.006 10.306 26.042 ;
               RECT 10.254 27.206 10.306 27.242 ;
               RECT 10.254 28.406 10.306 28.442 ;
               RECT 10.254 29.606 10.306 29.642 ;
               RECT 10.254 30.806 10.306 30.842 ;
               RECT 10.254 32.006 10.306 32.042 ;
               RECT 10.254 33.206 10.306 33.242 ;
               RECT 10.254 34.406 10.306 34.442 ;
               RECT 10.254 35.606 10.306 35.642 ;
               RECT 10.254 36.806 10.306 36.842 ;
               RECT 10.254 38.006 10.306 38.042 ;
               RECT 10.254 39.206 10.306 39.242 ;
               RECT 10.254 40.406 10.306 40.442 ;
               RECT 10.254 41.606 10.306 41.642 ;
               RECT 10.254 42.806 10.306 42.842 ;
               RECT 10.254 44.006 10.306 44.042 ;
               RECT 10.254 45.206 10.306 45.242 ;
               RECT 10.254 46.406 10.306 46.442 ;
               RECT 10.254 47.606 10.306 47.642 ;
               RECT 10.254 49.422 10.306 49.458 ;
               RECT 10.254 49.662 10.306 49.698 ;
               RECT 10.254 55.422 10.306 55.458 ;
               RECT 10.254 55.662 10.306 55.698 ;
               RECT 10.254 56.726 10.306 56.762 ;
               RECT 10.254 57.926 10.306 57.962 ;
               RECT 10.254 59.126 10.306 59.162 ;
               RECT 10.254 60.326 10.306 60.362 ;
               RECT 10.254 61.526 10.306 61.562 ;
               RECT 10.254 62.726 10.306 62.762 ;
               RECT 10.254 63.926 10.306 63.962 ;
               RECT 10.254 65.126 10.306 65.162 ;
               RECT 10.254 66.326 10.306 66.362 ;
               RECT 10.254 67.526 10.306 67.562 ;
               RECT 10.254 68.726 10.306 68.762 ;
               RECT 10.254 69.926 10.306 69.962 ;
               RECT 10.254 71.126 10.306 71.162 ;
               RECT 10.254 72.326 10.306 72.362 ;
               RECT 10.254 73.526 10.306 73.562 ;
               RECT 10.254 74.726 10.306 74.762 ;
               RECT 10.254 75.926 10.306 75.962 ;
               RECT 10.254 77.126 10.306 77.162 ;
               RECT 10.254 78.326 10.306 78.362 ;
               RECT 10.254 79.526 10.306 79.562 ;
               RECT 10.254 80.726 10.306 80.762 ;
               RECT 10.254 81.926 10.306 81.962 ;
               RECT 10.254 83.126 10.306 83.162 ;
               RECT 10.254 84.326 10.306 84.362 ;
               RECT 10.254 85.526 10.306 85.562 ;
               RECT 10.254 86.726 10.306 86.762 ;
               RECT 10.254 87.926 10.306 87.962 ;
               RECT 10.254 89.126 10.306 89.162 ;
               RECT 10.254 90.326 10.306 90.362 ;
               RECT 10.254 91.526 10.306 91.562 ;
               RECT 10.254 92.726 10.306 92.762 ;
               RECT 10.254 93.926 10.306 93.962 ;
               RECT 10.254 95.126 10.306 95.162 ;
               RECT 10.254 96.326 10.306 96.362 ;
               RECT 10.254 97.526 10.306 97.562 ;
               RECT 10.254 98.726 10.306 98.762 ;
               RECT 10.254 99.926 10.306 99.962 ;
               RECT 10.254 101.126 10.306 101.162 ;
               RECT 10.254 102.326 10.306 102.362 ;
               RECT 10.254 103.526 10.306 103.562 ;
               RECT 10.334 1.558 10.386 1.594 ;
               RECT 10.334 2.758 10.386 2.794 ;
               RECT 10.334 3.958 10.386 3.994 ;
               RECT 10.334 5.158 10.386 5.194 ;
               RECT 10.334 6.358 10.386 6.394 ;
               RECT 10.334 7.558 10.386 7.594 ;
               RECT 10.334 8.758 10.386 8.794 ;
               RECT 10.334 9.958 10.386 9.994 ;
               RECT 10.334 11.158 10.386 11.194 ;
               RECT 10.334 12.358 10.386 12.394 ;
               RECT 10.334 13.558 10.386 13.594 ;
               RECT 10.334 14.758 10.386 14.794 ;
               RECT 10.334 15.958 10.386 15.994 ;
               RECT 10.334 17.158 10.386 17.194 ;
               RECT 10.334 18.358 10.386 18.394 ;
               RECT 10.334 19.558 10.386 19.594 ;
               RECT 10.334 20.758 10.386 20.794 ;
               RECT 10.334 21.958 10.386 21.994 ;
               RECT 10.334 23.158 10.386 23.194 ;
               RECT 10.334 24.358 10.386 24.394 ;
               RECT 10.334 25.558 10.386 25.594 ;
               RECT 10.334 26.758 10.386 26.794 ;
               RECT 10.334 27.958 10.386 27.994 ;
               RECT 10.334 29.158 10.386 29.194 ;
               RECT 10.334 30.358 10.386 30.394 ;
               RECT 10.334 31.558 10.386 31.594 ;
               RECT 10.334 32.758 10.386 32.794 ;
               RECT 10.334 33.958 10.386 33.994 ;
               RECT 10.334 35.158 10.386 35.194 ;
               RECT 10.334 36.358 10.386 36.394 ;
               RECT 10.334 37.558 10.386 37.594 ;
               RECT 10.334 38.758 10.386 38.794 ;
               RECT 10.334 39.958 10.386 39.994 ;
               RECT 10.334 41.158 10.386 41.194 ;
               RECT 10.334 42.358 10.386 42.394 ;
               RECT 10.334 43.558 10.386 43.594 ;
               RECT 10.334 44.758 10.386 44.794 ;
               RECT 10.334 45.958 10.386 45.994 ;
               RECT 10.334 47.158 10.386 47.194 ;
               RECT 10.334 48.358 10.386 48.394 ;
               RECT 10.334 50.142 10.386 50.178 ;
               RECT 10.334 50.382 10.386 50.418 ;
               RECT 10.334 54.702 10.386 54.738 ;
               RECT 10.334 54.942 10.386 54.978 ;
               RECT 10.334 57.478 10.386 57.514 ;
               RECT 10.334 58.678 10.386 58.714 ;
               RECT 10.334 59.878 10.386 59.914 ;
               RECT 10.334 61.078 10.386 61.114 ;
               RECT 10.334 62.278 10.386 62.314 ;
               RECT 10.334 63.478 10.386 63.514 ;
               RECT 10.334 64.678 10.386 64.714 ;
               RECT 10.334 65.878 10.386 65.914 ;
               RECT 10.334 67.078 10.386 67.114 ;
               RECT 10.334 68.278 10.386 68.314 ;
               RECT 10.334 69.478 10.386 69.514 ;
               RECT 10.334 70.678 10.386 70.714 ;
               RECT 10.334 71.878 10.386 71.914 ;
               RECT 10.334 73.078 10.386 73.114 ;
               RECT 10.334 74.278 10.386 74.314 ;
               RECT 10.334 75.478 10.386 75.514 ;
               RECT 10.334 76.678 10.386 76.714 ;
               RECT 10.334 77.878 10.386 77.914 ;
               RECT 10.334 79.078 10.386 79.114 ;
               RECT 10.334 80.278 10.386 80.314 ;
               RECT 10.334 81.478 10.386 81.514 ;
               RECT 10.334 82.678 10.386 82.714 ;
               RECT 10.334 83.878 10.386 83.914 ;
               RECT 10.334 85.078 10.386 85.114 ;
               RECT 10.334 86.278 10.386 86.314 ;
               RECT 10.334 87.478 10.386 87.514 ;
               RECT 10.334 88.678 10.386 88.714 ;
               RECT 10.334 89.878 10.386 89.914 ;
               RECT 10.334 91.078 10.386 91.114 ;
               RECT 10.334 92.278 10.386 92.314 ;
               RECT 10.334 93.478 10.386 93.514 ;
               RECT 10.334 94.678 10.386 94.714 ;
               RECT 10.334 95.878 10.386 95.914 ;
               RECT 10.334 97.078 10.386 97.114 ;
               RECT 10.334 98.278 10.386 98.314 ;
               RECT 10.334 99.478 10.386 99.514 ;
               RECT 10.334 100.678 10.386 100.714 ;
               RECT 10.334 101.878 10.386 101.914 ;
               RECT 10.334 103.078 10.386 103.114 ;
               RECT 10.334 104.278 10.386 104.314 ;
               RECT 10.414 0.806 10.466 0.842 ;
               RECT 10.414 2.006 10.466 2.042 ;
               RECT 10.414 3.206 10.466 3.242 ;
               RECT 10.414 4.406 10.466 4.442 ;
               RECT 10.414 5.606 10.466 5.642 ;
               RECT 10.414 6.806 10.466 6.842 ;
               RECT 10.414 8.006 10.466 8.042 ;
               RECT 10.414 9.206 10.466 9.242 ;
               RECT 10.414 10.406 10.466 10.442 ;
               RECT 10.414 11.606 10.466 11.642 ;
               RECT 10.414 12.806 10.466 12.842 ;
               RECT 10.414 14.006 10.466 14.042 ;
               RECT 10.414 15.206 10.466 15.242 ;
               RECT 10.414 16.406 10.466 16.442 ;
               RECT 10.414 17.606 10.466 17.642 ;
               RECT 10.414 18.806 10.466 18.842 ;
               RECT 10.414 20.006 10.466 20.042 ;
               RECT 10.414 21.206 10.466 21.242 ;
               RECT 10.414 22.406 10.466 22.442 ;
               RECT 10.414 23.606 10.466 23.642 ;
               RECT 10.414 24.806 10.466 24.842 ;
               RECT 10.414 26.006 10.466 26.042 ;
               RECT 10.414 27.206 10.466 27.242 ;
               RECT 10.414 28.406 10.466 28.442 ;
               RECT 10.414 29.606 10.466 29.642 ;
               RECT 10.414 30.806 10.466 30.842 ;
               RECT 10.414 32.006 10.466 32.042 ;
               RECT 10.414 33.206 10.466 33.242 ;
               RECT 10.414 34.406 10.466 34.442 ;
               RECT 10.414 35.606 10.466 35.642 ;
               RECT 10.414 36.806 10.466 36.842 ;
               RECT 10.414 38.006 10.466 38.042 ;
               RECT 10.414 39.206 10.466 39.242 ;
               RECT 10.414 40.406 10.466 40.442 ;
               RECT 10.414 41.606 10.466 41.642 ;
               RECT 10.414 42.806 10.466 42.842 ;
               RECT 10.414 44.006 10.466 44.042 ;
               RECT 10.414 45.206 10.466 45.242 ;
               RECT 10.414 46.406 10.466 46.442 ;
               RECT 10.414 47.606 10.466 47.642 ;
               RECT 10.414 49.422 10.466 49.458 ;
               RECT 10.414 49.662 10.466 49.698 ;
               RECT 10.414 55.422 10.466 55.458 ;
               RECT 10.414 55.662 10.466 55.698 ;
               RECT 10.414 56.726 10.466 56.762 ;
               RECT 10.414 57.926 10.466 57.962 ;
               RECT 10.414 59.126 10.466 59.162 ;
               RECT 10.414 60.326 10.466 60.362 ;
               RECT 10.414 61.526 10.466 61.562 ;
               RECT 10.414 62.726 10.466 62.762 ;
               RECT 10.414 63.926 10.466 63.962 ;
               RECT 10.414 65.126 10.466 65.162 ;
               RECT 10.414 66.326 10.466 66.362 ;
               RECT 10.414 67.526 10.466 67.562 ;
               RECT 10.414 68.726 10.466 68.762 ;
               RECT 10.414 69.926 10.466 69.962 ;
               RECT 10.414 71.126 10.466 71.162 ;
               RECT 10.414 72.326 10.466 72.362 ;
               RECT 10.414 73.526 10.466 73.562 ;
               RECT 10.414 74.726 10.466 74.762 ;
               RECT 10.414 75.926 10.466 75.962 ;
               RECT 10.414 77.126 10.466 77.162 ;
               RECT 10.414 78.326 10.466 78.362 ;
               RECT 10.414 79.526 10.466 79.562 ;
               RECT 10.414 80.726 10.466 80.762 ;
               RECT 10.414 81.926 10.466 81.962 ;
               RECT 10.414 83.126 10.466 83.162 ;
               RECT 10.414 84.326 10.466 84.362 ;
               RECT 10.414 85.526 10.466 85.562 ;
               RECT 10.414 86.726 10.466 86.762 ;
               RECT 10.414 87.926 10.466 87.962 ;
               RECT 10.414 89.126 10.466 89.162 ;
               RECT 10.414 90.326 10.466 90.362 ;
               RECT 10.414 91.526 10.466 91.562 ;
               RECT 10.414 92.726 10.466 92.762 ;
               RECT 10.414 93.926 10.466 93.962 ;
               RECT 10.414 95.126 10.466 95.162 ;
               RECT 10.414 96.326 10.466 96.362 ;
               RECT 10.414 97.526 10.466 97.562 ;
               RECT 10.414 98.726 10.466 98.762 ;
               RECT 10.414 99.926 10.466 99.962 ;
               RECT 10.414 101.126 10.466 101.162 ;
               RECT 10.414 102.326 10.466 102.362 ;
               RECT 10.414 103.526 10.466 103.562 ;
               RECT 10.494 1.558 10.546 1.594 ;
               RECT 10.494 2.758 10.546 2.794 ;
               RECT 10.494 3.958 10.546 3.994 ;
               RECT 10.494 5.158 10.546 5.194 ;
               RECT 10.494 6.358 10.546 6.394 ;
               RECT 10.494 7.558 10.546 7.594 ;
               RECT 10.494 8.758 10.546 8.794 ;
               RECT 10.494 9.958 10.546 9.994 ;
               RECT 10.494 11.158 10.546 11.194 ;
               RECT 10.494 12.358 10.546 12.394 ;
               RECT 10.494 13.558 10.546 13.594 ;
               RECT 10.494 14.758 10.546 14.794 ;
               RECT 10.494 15.958 10.546 15.994 ;
               RECT 10.494 17.158 10.546 17.194 ;
               RECT 10.494 18.358 10.546 18.394 ;
               RECT 10.494 19.558 10.546 19.594 ;
               RECT 10.494 20.758 10.546 20.794 ;
               RECT 10.494 21.958 10.546 21.994 ;
               RECT 10.494 23.158 10.546 23.194 ;
               RECT 10.494 24.358 10.546 24.394 ;
               RECT 10.494 25.558 10.546 25.594 ;
               RECT 10.494 26.758 10.546 26.794 ;
               RECT 10.494 27.958 10.546 27.994 ;
               RECT 10.494 29.158 10.546 29.194 ;
               RECT 10.494 30.358 10.546 30.394 ;
               RECT 10.494 31.558 10.546 31.594 ;
               RECT 10.494 32.758 10.546 32.794 ;
               RECT 10.494 33.958 10.546 33.994 ;
               RECT 10.494 35.158 10.546 35.194 ;
               RECT 10.494 36.358 10.546 36.394 ;
               RECT 10.494 37.558 10.546 37.594 ;
               RECT 10.494 38.758 10.546 38.794 ;
               RECT 10.494 39.958 10.546 39.994 ;
               RECT 10.494 41.158 10.546 41.194 ;
               RECT 10.494 42.358 10.546 42.394 ;
               RECT 10.494 43.558 10.546 43.594 ;
               RECT 10.494 44.758 10.546 44.794 ;
               RECT 10.494 45.958 10.546 45.994 ;
               RECT 10.494 47.158 10.546 47.194 ;
               RECT 10.494 48.358 10.546 48.394 ;
               RECT 10.494 50.142 10.546 50.178 ;
               RECT 10.494 50.382 10.546 50.418 ;
               RECT 10.494 54.702 10.546 54.738 ;
               RECT 10.494 54.942 10.546 54.978 ;
               RECT 10.494 57.478 10.546 57.514 ;
               RECT 10.494 58.678 10.546 58.714 ;
               RECT 10.494 59.878 10.546 59.914 ;
               RECT 10.494 61.078 10.546 61.114 ;
               RECT 10.494 62.278 10.546 62.314 ;
               RECT 10.494 63.478 10.546 63.514 ;
               RECT 10.494 64.678 10.546 64.714 ;
               RECT 10.494 65.878 10.546 65.914 ;
               RECT 10.494 67.078 10.546 67.114 ;
               RECT 10.494 68.278 10.546 68.314 ;
               RECT 10.494 69.478 10.546 69.514 ;
               RECT 10.494 70.678 10.546 70.714 ;
               RECT 10.494 71.878 10.546 71.914 ;
               RECT 10.494 73.078 10.546 73.114 ;
               RECT 10.494 74.278 10.546 74.314 ;
               RECT 10.494 75.478 10.546 75.514 ;
               RECT 10.494 76.678 10.546 76.714 ;
               RECT 10.494 77.878 10.546 77.914 ;
               RECT 10.494 79.078 10.546 79.114 ;
               RECT 10.494 80.278 10.546 80.314 ;
               RECT 10.494 81.478 10.546 81.514 ;
               RECT 10.494 82.678 10.546 82.714 ;
               RECT 10.494 83.878 10.546 83.914 ;
               RECT 10.494 85.078 10.546 85.114 ;
               RECT 10.494 86.278 10.546 86.314 ;
               RECT 10.494 87.478 10.546 87.514 ;
               RECT 10.494 88.678 10.546 88.714 ;
               RECT 10.494 89.878 10.546 89.914 ;
               RECT 10.494 91.078 10.546 91.114 ;
               RECT 10.494 92.278 10.546 92.314 ;
               RECT 10.494 93.478 10.546 93.514 ;
               RECT 10.494 94.678 10.546 94.714 ;
               RECT 10.494 95.878 10.546 95.914 ;
               RECT 10.494 97.078 10.546 97.114 ;
               RECT 10.494 98.278 10.546 98.314 ;
               RECT 10.494 99.478 10.546 99.514 ;
               RECT 10.494 100.678 10.546 100.714 ;
               RECT 10.494 101.878 10.546 101.914 ;
               RECT 10.494 103.078 10.546 103.114 ;
               RECT 10.494 104.278 10.546 104.314 ;
               RECT 10.574 0.281 10.626 0.317 ;
               RECT 10.574 104.803 10.626 104.839 ;
               RECT 10.654 0.806 10.706 0.842 ;
               RECT 10.654 2.006 10.706 2.042 ;
               RECT 10.654 3.206 10.706 3.242 ;
               RECT 10.654 4.406 10.706 4.442 ;
               RECT 10.654 5.606 10.706 5.642 ;
               RECT 10.654 6.806 10.706 6.842 ;
               RECT 10.654 8.006 10.706 8.042 ;
               RECT 10.654 9.206 10.706 9.242 ;
               RECT 10.654 10.406 10.706 10.442 ;
               RECT 10.654 11.606 10.706 11.642 ;
               RECT 10.654 12.806 10.706 12.842 ;
               RECT 10.654 14.006 10.706 14.042 ;
               RECT 10.654 15.206 10.706 15.242 ;
               RECT 10.654 16.406 10.706 16.442 ;
               RECT 10.654 17.606 10.706 17.642 ;
               RECT 10.654 18.806 10.706 18.842 ;
               RECT 10.654 20.006 10.706 20.042 ;
               RECT 10.654 21.206 10.706 21.242 ;
               RECT 10.654 22.406 10.706 22.442 ;
               RECT 10.654 23.606 10.706 23.642 ;
               RECT 10.654 24.806 10.706 24.842 ;
               RECT 10.654 26.006 10.706 26.042 ;
               RECT 10.654 27.206 10.706 27.242 ;
               RECT 10.654 28.406 10.706 28.442 ;
               RECT 10.654 29.606 10.706 29.642 ;
               RECT 10.654 30.806 10.706 30.842 ;
               RECT 10.654 32.006 10.706 32.042 ;
               RECT 10.654 33.206 10.706 33.242 ;
               RECT 10.654 34.406 10.706 34.442 ;
               RECT 10.654 35.606 10.706 35.642 ;
               RECT 10.654 36.806 10.706 36.842 ;
               RECT 10.654 38.006 10.706 38.042 ;
               RECT 10.654 39.206 10.706 39.242 ;
               RECT 10.654 40.406 10.706 40.442 ;
               RECT 10.654 41.606 10.706 41.642 ;
               RECT 10.654 42.806 10.706 42.842 ;
               RECT 10.654 44.006 10.706 44.042 ;
               RECT 10.654 45.206 10.706 45.242 ;
               RECT 10.654 46.406 10.706 46.442 ;
               RECT 10.654 47.606 10.706 47.642 ;
               RECT 10.654 49.422 10.706 49.458 ;
               RECT 10.654 49.662 10.706 49.698 ;
               RECT 10.654 51.102 10.706 51.138 ;
               RECT 10.654 51.582 10.706 51.618 ;
               RECT 10.654 53.502 10.706 53.538 ;
               RECT 10.654 53.982 10.706 54.018 ;
               RECT 10.654 55.422 10.706 55.458 ;
               RECT 10.654 55.662 10.706 55.698 ;
               RECT 10.654 56.726 10.706 56.762 ;
               RECT 10.654 57.926 10.706 57.962 ;
               RECT 10.654 59.126 10.706 59.162 ;
               RECT 10.654 60.326 10.706 60.362 ;
               RECT 10.654 61.526 10.706 61.562 ;
               RECT 10.654 62.726 10.706 62.762 ;
               RECT 10.654 63.926 10.706 63.962 ;
               RECT 10.654 65.126 10.706 65.162 ;
               RECT 10.654 66.326 10.706 66.362 ;
               RECT 10.654 67.526 10.706 67.562 ;
               RECT 10.654 68.726 10.706 68.762 ;
               RECT 10.654 69.926 10.706 69.962 ;
               RECT 10.654 71.126 10.706 71.162 ;
               RECT 10.654 72.326 10.706 72.362 ;
               RECT 10.654 73.526 10.706 73.562 ;
               RECT 10.654 74.726 10.706 74.762 ;
               RECT 10.654 75.926 10.706 75.962 ;
               RECT 10.654 77.126 10.706 77.162 ;
               RECT 10.654 78.326 10.706 78.362 ;
               RECT 10.654 79.526 10.706 79.562 ;
               RECT 10.654 80.726 10.706 80.762 ;
               RECT 10.654 81.926 10.706 81.962 ;
               RECT 10.654 83.126 10.706 83.162 ;
               RECT 10.654 84.326 10.706 84.362 ;
               RECT 10.654 85.526 10.706 85.562 ;
               RECT 10.654 86.726 10.706 86.762 ;
               RECT 10.654 87.926 10.706 87.962 ;
               RECT 10.654 89.126 10.706 89.162 ;
               RECT 10.654 90.326 10.706 90.362 ;
               RECT 10.654 91.526 10.706 91.562 ;
               RECT 10.654 92.726 10.706 92.762 ;
               RECT 10.654 93.926 10.706 93.962 ;
               RECT 10.654 95.126 10.706 95.162 ;
               RECT 10.654 96.326 10.706 96.362 ;
               RECT 10.654 97.526 10.706 97.562 ;
               RECT 10.654 98.726 10.706 98.762 ;
               RECT 10.654 99.926 10.706 99.962 ;
               RECT 10.654 101.126 10.706 101.162 ;
               RECT 10.654 102.326 10.706 102.362 ;
               RECT 10.654 103.526 10.706 103.562 ;
               RECT 10.734 1.558 10.786 1.594 ;
               RECT 10.734 2.758 10.786 2.794 ;
               RECT 10.734 3.958 10.786 3.994 ;
               RECT 10.734 5.158 10.786 5.194 ;
               RECT 10.734 6.358 10.786 6.394 ;
               RECT 10.734 7.558 10.786 7.594 ;
               RECT 10.734 8.758 10.786 8.794 ;
               RECT 10.734 9.958 10.786 9.994 ;
               RECT 10.734 11.158 10.786 11.194 ;
               RECT 10.734 12.358 10.786 12.394 ;
               RECT 10.734 13.558 10.786 13.594 ;
               RECT 10.734 14.758 10.786 14.794 ;
               RECT 10.734 15.958 10.786 15.994 ;
               RECT 10.734 17.158 10.786 17.194 ;
               RECT 10.734 18.358 10.786 18.394 ;
               RECT 10.734 19.558 10.786 19.594 ;
               RECT 10.734 20.758 10.786 20.794 ;
               RECT 10.734 21.958 10.786 21.994 ;
               RECT 10.734 23.158 10.786 23.194 ;
               RECT 10.734 24.358 10.786 24.394 ;
               RECT 10.734 25.558 10.786 25.594 ;
               RECT 10.734 26.758 10.786 26.794 ;
               RECT 10.734 27.958 10.786 27.994 ;
               RECT 10.734 29.158 10.786 29.194 ;
               RECT 10.734 30.358 10.786 30.394 ;
               RECT 10.734 31.558 10.786 31.594 ;
               RECT 10.734 32.758 10.786 32.794 ;
               RECT 10.734 33.958 10.786 33.994 ;
               RECT 10.734 35.158 10.786 35.194 ;
               RECT 10.734 36.358 10.786 36.394 ;
               RECT 10.734 37.558 10.786 37.594 ;
               RECT 10.734 38.758 10.786 38.794 ;
               RECT 10.734 39.958 10.786 39.994 ;
               RECT 10.734 41.158 10.786 41.194 ;
               RECT 10.734 42.358 10.786 42.394 ;
               RECT 10.734 43.558 10.786 43.594 ;
               RECT 10.734 44.758 10.786 44.794 ;
               RECT 10.734 45.958 10.786 45.994 ;
               RECT 10.734 47.158 10.786 47.194 ;
               RECT 10.734 48.358 10.786 48.394 ;
               RECT 10.734 50.142 10.786 50.178 ;
               RECT 10.734 50.382 10.786 50.418 ;
               RECT 10.734 54.702 10.786 54.738 ;
               RECT 10.734 54.942 10.786 54.978 ;
               RECT 10.734 57.478 10.786 57.514 ;
               RECT 10.734 58.678 10.786 58.714 ;
               RECT 10.734 59.878 10.786 59.914 ;
               RECT 10.734 61.078 10.786 61.114 ;
               RECT 10.734 62.278 10.786 62.314 ;
               RECT 10.734 63.478 10.786 63.514 ;
               RECT 10.734 64.678 10.786 64.714 ;
               RECT 10.734 65.878 10.786 65.914 ;
               RECT 10.734 67.078 10.786 67.114 ;
               RECT 10.734 68.278 10.786 68.314 ;
               RECT 10.734 69.478 10.786 69.514 ;
               RECT 10.734 70.678 10.786 70.714 ;
               RECT 10.734 71.878 10.786 71.914 ;
               RECT 10.734 73.078 10.786 73.114 ;
               RECT 10.734 74.278 10.786 74.314 ;
               RECT 10.734 75.478 10.786 75.514 ;
               RECT 10.734 76.678 10.786 76.714 ;
               RECT 10.734 77.878 10.786 77.914 ;
               RECT 10.734 79.078 10.786 79.114 ;
               RECT 10.734 80.278 10.786 80.314 ;
               RECT 10.734 81.478 10.786 81.514 ;
               RECT 10.734 82.678 10.786 82.714 ;
               RECT 10.734 83.878 10.786 83.914 ;
               RECT 10.734 85.078 10.786 85.114 ;
               RECT 10.734 86.278 10.786 86.314 ;
               RECT 10.734 87.478 10.786 87.514 ;
               RECT 10.734 88.678 10.786 88.714 ;
               RECT 10.734 89.878 10.786 89.914 ;
               RECT 10.734 91.078 10.786 91.114 ;
               RECT 10.734 92.278 10.786 92.314 ;
               RECT 10.734 93.478 10.786 93.514 ;
               RECT 10.734 94.678 10.786 94.714 ;
               RECT 10.734 95.878 10.786 95.914 ;
               RECT 10.734 97.078 10.786 97.114 ;
               RECT 10.734 98.278 10.786 98.314 ;
               RECT 10.734 99.478 10.786 99.514 ;
               RECT 10.734 100.678 10.786 100.714 ;
               RECT 10.734 101.878 10.786 101.914 ;
               RECT 10.734 103.078 10.786 103.114 ;
               RECT 10.734 104.278 10.786 104.314 ;
               RECT 10.814 0.806 10.866 0.842 ;
               RECT 10.814 2.006 10.866 2.042 ;
               RECT 10.814 3.206 10.866 3.242 ;
               RECT 10.814 4.406 10.866 4.442 ;
               RECT 10.814 5.606 10.866 5.642 ;
               RECT 10.814 6.806 10.866 6.842 ;
               RECT 10.814 8.006 10.866 8.042 ;
               RECT 10.814 9.206 10.866 9.242 ;
               RECT 10.814 10.406 10.866 10.442 ;
               RECT 10.814 11.606 10.866 11.642 ;
               RECT 10.814 12.806 10.866 12.842 ;
               RECT 10.814 14.006 10.866 14.042 ;
               RECT 10.814 15.206 10.866 15.242 ;
               RECT 10.814 16.406 10.866 16.442 ;
               RECT 10.814 17.606 10.866 17.642 ;
               RECT 10.814 18.806 10.866 18.842 ;
               RECT 10.814 20.006 10.866 20.042 ;
               RECT 10.814 21.206 10.866 21.242 ;
               RECT 10.814 22.406 10.866 22.442 ;
               RECT 10.814 23.606 10.866 23.642 ;
               RECT 10.814 24.806 10.866 24.842 ;
               RECT 10.814 26.006 10.866 26.042 ;
               RECT 10.814 27.206 10.866 27.242 ;
               RECT 10.814 28.406 10.866 28.442 ;
               RECT 10.814 29.606 10.866 29.642 ;
               RECT 10.814 30.806 10.866 30.842 ;
               RECT 10.814 32.006 10.866 32.042 ;
               RECT 10.814 33.206 10.866 33.242 ;
               RECT 10.814 34.406 10.866 34.442 ;
               RECT 10.814 35.606 10.866 35.642 ;
               RECT 10.814 36.806 10.866 36.842 ;
               RECT 10.814 38.006 10.866 38.042 ;
               RECT 10.814 39.206 10.866 39.242 ;
               RECT 10.814 40.406 10.866 40.442 ;
               RECT 10.814 41.606 10.866 41.642 ;
               RECT 10.814 42.806 10.866 42.842 ;
               RECT 10.814 44.006 10.866 44.042 ;
               RECT 10.814 45.206 10.866 45.242 ;
               RECT 10.814 46.406 10.866 46.442 ;
               RECT 10.814 47.606 10.866 47.642 ;
               RECT 10.814 49.422 10.866 49.458 ;
               RECT 10.814 49.662 10.866 49.698 ;
               RECT 10.814 55.422 10.866 55.458 ;
               RECT 10.814 55.662 10.866 55.698 ;
               RECT 10.814 56.726 10.866 56.762 ;
               RECT 10.814 57.926 10.866 57.962 ;
               RECT 10.814 59.126 10.866 59.162 ;
               RECT 10.814 60.326 10.866 60.362 ;
               RECT 10.814 61.526 10.866 61.562 ;
               RECT 10.814 62.726 10.866 62.762 ;
               RECT 10.814 63.926 10.866 63.962 ;
               RECT 10.814 65.126 10.866 65.162 ;
               RECT 10.814 66.326 10.866 66.362 ;
               RECT 10.814 67.526 10.866 67.562 ;
               RECT 10.814 68.726 10.866 68.762 ;
               RECT 10.814 69.926 10.866 69.962 ;
               RECT 10.814 71.126 10.866 71.162 ;
               RECT 10.814 72.326 10.866 72.362 ;
               RECT 10.814 73.526 10.866 73.562 ;
               RECT 10.814 74.726 10.866 74.762 ;
               RECT 10.814 75.926 10.866 75.962 ;
               RECT 10.814 77.126 10.866 77.162 ;
               RECT 10.814 78.326 10.866 78.362 ;
               RECT 10.814 79.526 10.866 79.562 ;
               RECT 10.814 80.726 10.866 80.762 ;
               RECT 10.814 81.926 10.866 81.962 ;
               RECT 10.814 83.126 10.866 83.162 ;
               RECT 10.814 84.326 10.866 84.362 ;
               RECT 10.814 85.526 10.866 85.562 ;
               RECT 10.814 86.726 10.866 86.762 ;
               RECT 10.814 87.926 10.866 87.962 ;
               RECT 10.814 89.126 10.866 89.162 ;
               RECT 10.814 90.326 10.866 90.362 ;
               RECT 10.814 91.526 10.866 91.562 ;
               RECT 10.814 92.726 10.866 92.762 ;
               RECT 10.814 93.926 10.866 93.962 ;
               RECT 10.814 95.126 10.866 95.162 ;
               RECT 10.814 96.326 10.866 96.362 ;
               RECT 10.814 97.526 10.866 97.562 ;
               RECT 10.814 98.726 10.866 98.762 ;
               RECT 10.814 99.926 10.866 99.962 ;
               RECT 10.814 101.126 10.866 101.162 ;
               RECT 10.814 102.326 10.866 102.362 ;
               RECT 10.814 103.526 10.866 103.562 ;
               RECT 10.894 1.558 10.946 1.594 ;
               RECT 10.894 2.758 10.946 2.794 ;
               RECT 10.894 3.958 10.946 3.994 ;
               RECT 10.894 5.158 10.946 5.194 ;
               RECT 10.894 6.358 10.946 6.394 ;
               RECT 10.894 7.558 10.946 7.594 ;
               RECT 10.894 8.758 10.946 8.794 ;
               RECT 10.894 9.958 10.946 9.994 ;
               RECT 10.894 11.158 10.946 11.194 ;
               RECT 10.894 12.358 10.946 12.394 ;
               RECT 10.894 13.558 10.946 13.594 ;
               RECT 10.894 14.758 10.946 14.794 ;
               RECT 10.894 15.958 10.946 15.994 ;
               RECT 10.894 17.158 10.946 17.194 ;
               RECT 10.894 18.358 10.946 18.394 ;
               RECT 10.894 19.558 10.946 19.594 ;
               RECT 10.894 20.758 10.946 20.794 ;
               RECT 10.894 21.958 10.946 21.994 ;
               RECT 10.894 23.158 10.946 23.194 ;
               RECT 10.894 24.358 10.946 24.394 ;
               RECT 10.894 25.558 10.946 25.594 ;
               RECT 10.894 26.758 10.946 26.794 ;
               RECT 10.894 27.958 10.946 27.994 ;
               RECT 10.894 29.158 10.946 29.194 ;
               RECT 10.894 30.358 10.946 30.394 ;
               RECT 10.894 31.558 10.946 31.594 ;
               RECT 10.894 32.758 10.946 32.794 ;
               RECT 10.894 33.958 10.946 33.994 ;
               RECT 10.894 35.158 10.946 35.194 ;
               RECT 10.894 36.358 10.946 36.394 ;
               RECT 10.894 37.558 10.946 37.594 ;
               RECT 10.894 38.758 10.946 38.794 ;
               RECT 10.894 39.958 10.946 39.994 ;
               RECT 10.894 41.158 10.946 41.194 ;
               RECT 10.894 42.358 10.946 42.394 ;
               RECT 10.894 43.558 10.946 43.594 ;
               RECT 10.894 44.758 10.946 44.794 ;
               RECT 10.894 45.958 10.946 45.994 ;
               RECT 10.894 47.158 10.946 47.194 ;
               RECT 10.894 48.358 10.946 48.394 ;
               RECT 10.894 50.142 10.946 50.178 ;
               RECT 10.894 50.382 10.946 50.418 ;
               RECT 10.894 54.702 10.946 54.738 ;
               RECT 10.894 54.942 10.946 54.978 ;
               RECT 10.894 57.478 10.946 57.514 ;
               RECT 10.894 58.678 10.946 58.714 ;
               RECT 10.894 59.878 10.946 59.914 ;
               RECT 10.894 61.078 10.946 61.114 ;
               RECT 10.894 62.278 10.946 62.314 ;
               RECT 10.894 63.478 10.946 63.514 ;
               RECT 10.894 64.678 10.946 64.714 ;
               RECT 10.894 65.878 10.946 65.914 ;
               RECT 10.894 67.078 10.946 67.114 ;
               RECT 10.894 68.278 10.946 68.314 ;
               RECT 10.894 69.478 10.946 69.514 ;
               RECT 10.894 70.678 10.946 70.714 ;
               RECT 10.894 71.878 10.946 71.914 ;
               RECT 10.894 73.078 10.946 73.114 ;
               RECT 10.894 74.278 10.946 74.314 ;
               RECT 10.894 75.478 10.946 75.514 ;
               RECT 10.894 76.678 10.946 76.714 ;
               RECT 10.894 77.878 10.946 77.914 ;
               RECT 10.894 79.078 10.946 79.114 ;
               RECT 10.894 80.278 10.946 80.314 ;
               RECT 10.894 81.478 10.946 81.514 ;
               RECT 10.894 82.678 10.946 82.714 ;
               RECT 10.894 83.878 10.946 83.914 ;
               RECT 10.894 85.078 10.946 85.114 ;
               RECT 10.894 86.278 10.946 86.314 ;
               RECT 10.894 87.478 10.946 87.514 ;
               RECT 10.894 88.678 10.946 88.714 ;
               RECT 10.894 89.878 10.946 89.914 ;
               RECT 10.894 91.078 10.946 91.114 ;
               RECT 10.894 92.278 10.946 92.314 ;
               RECT 10.894 93.478 10.946 93.514 ;
               RECT 10.894 94.678 10.946 94.714 ;
               RECT 10.894 95.878 10.946 95.914 ;
               RECT 10.894 97.078 10.946 97.114 ;
               RECT 10.894 98.278 10.946 98.314 ;
               RECT 10.894 99.478 10.946 99.514 ;
               RECT 10.894 100.678 10.946 100.714 ;
               RECT 10.894 101.878 10.946 101.914 ;
               RECT 10.894 103.078 10.946 103.114 ;
               RECT 10.894 104.278 10.946 104.314 ;
               RECT 10.974 0.281 11.026 0.317 ;
               RECT 10.974 104.803 11.026 104.839 ;
               RECT 11.054 0.806 11.106 0.842 ;
               RECT 11.054 2.006 11.106 2.042 ;
               RECT 11.054 3.206 11.106 3.242 ;
               RECT 11.054 4.406 11.106 4.442 ;
               RECT 11.054 5.606 11.106 5.642 ;
               RECT 11.054 6.806 11.106 6.842 ;
               RECT 11.054 8.006 11.106 8.042 ;
               RECT 11.054 9.206 11.106 9.242 ;
               RECT 11.054 10.406 11.106 10.442 ;
               RECT 11.054 11.606 11.106 11.642 ;
               RECT 11.054 12.806 11.106 12.842 ;
               RECT 11.054 14.006 11.106 14.042 ;
               RECT 11.054 15.206 11.106 15.242 ;
               RECT 11.054 16.406 11.106 16.442 ;
               RECT 11.054 17.606 11.106 17.642 ;
               RECT 11.054 18.806 11.106 18.842 ;
               RECT 11.054 20.006 11.106 20.042 ;
               RECT 11.054 21.206 11.106 21.242 ;
               RECT 11.054 22.406 11.106 22.442 ;
               RECT 11.054 23.606 11.106 23.642 ;
               RECT 11.054 24.806 11.106 24.842 ;
               RECT 11.054 26.006 11.106 26.042 ;
               RECT 11.054 27.206 11.106 27.242 ;
               RECT 11.054 28.406 11.106 28.442 ;
               RECT 11.054 29.606 11.106 29.642 ;
               RECT 11.054 30.806 11.106 30.842 ;
               RECT 11.054 32.006 11.106 32.042 ;
               RECT 11.054 33.206 11.106 33.242 ;
               RECT 11.054 34.406 11.106 34.442 ;
               RECT 11.054 35.606 11.106 35.642 ;
               RECT 11.054 36.806 11.106 36.842 ;
               RECT 11.054 38.006 11.106 38.042 ;
               RECT 11.054 39.206 11.106 39.242 ;
               RECT 11.054 40.406 11.106 40.442 ;
               RECT 11.054 41.606 11.106 41.642 ;
               RECT 11.054 42.806 11.106 42.842 ;
               RECT 11.054 44.006 11.106 44.042 ;
               RECT 11.054 45.206 11.106 45.242 ;
               RECT 11.054 46.406 11.106 46.442 ;
               RECT 11.054 47.606 11.106 47.642 ;
               RECT 11.054 49.422 11.106 49.458 ;
               RECT 11.054 49.662 11.106 49.698 ;
               RECT 11.054 55.422 11.106 55.458 ;
               RECT 11.054 55.662 11.106 55.698 ;
               RECT 11.054 56.726 11.106 56.762 ;
               RECT 11.054 57.926 11.106 57.962 ;
               RECT 11.054 59.126 11.106 59.162 ;
               RECT 11.054 60.326 11.106 60.362 ;
               RECT 11.054 61.526 11.106 61.562 ;
               RECT 11.054 62.726 11.106 62.762 ;
               RECT 11.054 63.926 11.106 63.962 ;
               RECT 11.054 65.126 11.106 65.162 ;
               RECT 11.054 66.326 11.106 66.362 ;
               RECT 11.054 67.526 11.106 67.562 ;
               RECT 11.054 68.726 11.106 68.762 ;
               RECT 11.054 69.926 11.106 69.962 ;
               RECT 11.054 71.126 11.106 71.162 ;
               RECT 11.054 72.326 11.106 72.362 ;
               RECT 11.054 73.526 11.106 73.562 ;
               RECT 11.054 74.726 11.106 74.762 ;
               RECT 11.054 75.926 11.106 75.962 ;
               RECT 11.054 77.126 11.106 77.162 ;
               RECT 11.054 78.326 11.106 78.362 ;
               RECT 11.054 79.526 11.106 79.562 ;
               RECT 11.054 80.726 11.106 80.762 ;
               RECT 11.054 81.926 11.106 81.962 ;
               RECT 11.054 83.126 11.106 83.162 ;
               RECT 11.054 84.326 11.106 84.362 ;
               RECT 11.054 85.526 11.106 85.562 ;
               RECT 11.054 86.726 11.106 86.762 ;
               RECT 11.054 87.926 11.106 87.962 ;
               RECT 11.054 89.126 11.106 89.162 ;
               RECT 11.054 90.326 11.106 90.362 ;
               RECT 11.054 91.526 11.106 91.562 ;
               RECT 11.054 92.726 11.106 92.762 ;
               RECT 11.054 93.926 11.106 93.962 ;
               RECT 11.054 95.126 11.106 95.162 ;
               RECT 11.054 96.326 11.106 96.362 ;
               RECT 11.054 97.526 11.106 97.562 ;
               RECT 11.054 98.726 11.106 98.762 ;
               RECT 11.054 99.926 11.106 99.962 ;
               RECT 11.054 101.126 11.106 101.162 ;
               RECT 11.054 102.326 11.106 102.362 ;
               RECT 11.054 103.526 11.106 103.562 ;
               RECT 11.134 1.558 11.186 1.594 ;
               RECT 11.134 2.758 11.186 2.794 ;
               RECT 11.134 3.958 11.186 3.994 ;
               RECT 11.134 5.158 11.186 5.194 ;
               RECT 11.134 6.358 11.186 6.394 ;
               RECT 11.134 7.558 11.186 7.594 ;
               RECT 11.134 8.758 11.186 8.794 ;
               RECT 11.134 9.958 11.186 9.994 ;
               RECT 11.134 11.158 11.186 11.194 ;
               RECT 11.134 12.358 11.186 12.394 ;
               RECT 11.134 13.558 11.186 13.594 ;
               RECT 11.134 14.758 11.186 14.794 ;
               RECT 11.134 15.958 11.186 15.994 ;
               RECT 11.134 17.158 11.186 17.194 ;
               RECT 11.134 18.358 11.186 18.394 ;
               RECT 11.134 19.558 11.186 19.594 ;
               RECT 11.134 20.758 11.186 20.794 ;
               RECT 11.134 21.958 11.186 21.994 ;
               RECT 11.134 23.158 11.186 23.194 ;
               RECT 11.134 24.358 11.186 24.394 ;
               RECT 11.134 25.558 11.186 25.594 ;
               RECT 11.134 26.758 11.186 26.794 ;
               RECT 11.134 27.958 11.186 27.994 ;
               RECT 11.134 29.158 11.186 29.194 ;
               RECT 11.134 30.358 11.186 30.394 ;
               RECT 11.134 31.558 11.186 31.594 ;
               RECT 11.134 32.758 11.186 32.794 ;
               RECT 11.134 33.958 11.186 33.994 ;
               RECT 11.134 35.158 11.186 35.194 ;
               RECT 11.134 36.358 11.186 36.394 ;
               RECT 11.134 37.558 11.186 37.594 ;
               RECT 11.134 38.758 11.186 38.794 ;
               RECT 11.134 39.958 11.186 39.994 ;
               RECT 11.134 41.158 11.186 41.194 ;
               RECT 11.134 42.358 11.186 42.394 ;
               RECT 11.134 43.558 11.186 43.594 ;
               RECT 11.134 44.758 11.186 44.794 ;
               RECT 11.134 45.958 11.186 45.994 ;
               RECT 11.134 47.158 11.186 47.194 ;
               RECT 11.134 48.358 11.186 48.394 ;
               RECT 11.134 50.142 11.186 50.178 ;
               RECT 11.134 50.382 11.186 50.418 ;
               RECT 11.134 54.702 11.186 54.738 ;
               RECT 11.134 54.942 11.186 54.978 ;
               RECT 11.134 57.478 11.186 57.514 ;
               RECT 11.134 58.678 11.186 58.714 ;
               RECT 11.134 59.878 11.186 59.914 ;
               RECT 11.134 61.078 11.186 61.114 ;
               RECT 11.134 62.278 11.186 62.314 ;
               RECT 11.134 63.478 11.186 63.514 ;
               RECT 11.134 64.678 11.186 64.714 ;
               RECT 11.134 65.878 11.186 65.914 ;
               RECT 11.134 67.078 11.186 67.114 ;
               RECT 11.134 68.278 11.186 68.314 ;
               RECT 11.134 69.478 11.186 69.514 ;
               RECT 11.134 70.678 11.186 70.714 ;
               RECT 11.134 71.878 11.186 71.914 ;
               RECT 11.134 73.078 11.186 73.114 ;
               RECT 11.134 74.278 11.186 74.314 ;
               RECT 11.134 75.478 11.186 75.514 ;
               RECT 11.134 76.678 11.186 76.714 ;
               RECT 11.134 77.878 11.186 77.914 ;
               RECT 11.134 79.078 11.186 79.114 ;
               RECT 11.134 80.278 11.186 80.314 ;
               RECT 11.134 81.478 11.186 81.514 ;
               RECT 11.134 82.678 11.186 82.714 ;
               RECT 11.134 83.878 11.186 83.914 ;
               RECT 11.134 85.078 11.186 85.114 ;
               RECT 11.134 86.278 11.186 86.314 ;
               RECT 11.134 87.478 11.186 87.514 ;
               RECT 11.134 88.678 11.186 88.714 ;
               RECT 11.134 89.878 11.186 89.914 ;
               RECT 11.134 91.078 11.186 91.114 ;
               RECT 11.134 92.278 11.186 92.314 ;
               RECT 11.134 93.478 11.186 93.514 ;
               RECT 11.134 94.678 11.186 94.714 ;
               RECT 11.134 95.878 11.186 95.914 ;
               RECT 11.134 97.078 11.186 97.114 ;
               RECT 11.134 98.278 11.186 98.314 ;
               RECT 11.134 99.478 11.186 99.514 ;
               RECT 11.134 100.678 11.186 100.714 ;
               RECT 11.134 101.878 11.186 101.914 ;
               RECT 11.134 103.078 11.186 103.114 ;
               RECT 11.134 104.278 11.186 104.314 ;
               RECT 11.214 0.806 11.266 0.842 ;
               RECT 11.214 2.006 11.266 2.042 ;
               RECT 11.214 3.206 11.266 3.242 ;
               RECT 11.214 4.406 11.266 4.442 ;
               RECT 11.214 5.606 11.266 5.642 ;
               RECT 11.214 6.806 11.266 6.842 ;
               RECT 11.214 8.006 11.266 8.042 ;
               RECT 11.214 9.206 11.266 9.242 ;
               RECT 11.214 10.406 11.266 10.442 ;
               RECT 11.214 11.606 11.266 11.642 ;
               RECT 11.214 12.806 11.266 12.842 ;
               RECT 11.214 14.006 11.266 14.042 ;
               RECT 11.214 15.206 11.266 15.242 ;
               RECT 11.214 16.406 11.266 16.442 ;
               RECT 11.214 17.606 11.266 17.642 ;
               RECT 11.214 18.806 11.266 18.842 ;
               RECT 11.214 20.006 11.266 20.042 ;
               RECT 11.214 21.206 11.266 21.242 ;
               RECT 11.214 22.406 11.266 22.442 ;
               RECT 11.214 23.606 11.266 23.642 ;
               RECT 11.214 24.806 11.266 24.842 ;
               RECT 11.214 26.006 11.266 26.042 ;
               RECT 11.214 27.206 11.266 27.242 ;
               RECT 11.214 28.406 11.266 28.442 ;
               RECT 11.214 29.606 11.266 29.642 ;
               RECT 11.214 30.806 11.266 30.842 ;
               RECT 11.214 32.006 11.266 32.042 ;
               RECT 11.214 33.206 11.266 33.242 ;
               RECT 11.214 34.406 11.266 34.442 ;
               RECT 11.214 35.606 11.266 35.642 ;
               RECT 11.214 36.806 11.266 36.842 ;
               RECT 11.214 38.006 11.266 38.042 ;
               RECT 11.214 39.206 11.266 39.242 ;
               RECT 11.214 40.406 11.266 40.442 ;
               RECT 11.214 41.606 11.266 41.642 ;
               RECT 11.214 42.806 11.266 42.842 ;
               RECT 11.214 44.006 11.266 44.042 ;
               RECT 11.214 45.206 11.266 45.242 ;
               RECT 11.214 46.406 11.266 46.442 ;
               RECT 11.214 47.606 11.266 47.642 ;
               RECT 11.214 49.422 11.266 49.458 ;
               RECT 11.214 49.662 11.266 49.698 ;
               RECT 11.214 55.422 11.266 55.458 ;
               RECT 11.214 55.662 11.266 55.698 ;
               RECT 11.214 56.726 11.266 56.762 ;
               RECT 11.214 57.926 11.266 57.962 ;
               RECT 11.214 59.126 11.266 59.162 ;
               RECT 11.214 60.326 11.266 60.362 ;
               RECT 11.214 61.526 11.266 61.562 ;
               RECT 11.214 62.726 11.266 62.762 ;
               RECT 11.214 63.926 11.266 63.962 ;
               RECT 11.214 65.126 11.266 65.162 ;
               RECT 11.214 66.326 11.266 66.362 ;
               RECT 11.214 67.526 11.266 67.562 ;
               RECT 11.214 68.726 11.266 68.762 ;
               RECT 11.214 69.926 11.266 69.962 ;
               RECT 11.214 71.126 11.266 71.162 ;
               RECT 11.214 72.326 11.266 72.362 ;
               RECT 11.214 73.526 11.266 73.562 ;
               RECT 11.214 74.726 11.266 74.762 ;
               RECT 11.214 75.926 11.266 75.962 ;
               RECT 11.214 77.126 11.266 77.162 ;
               RECT 11.214 78.326 11.266 78.362 ;
               RECT 11.214 79.526 11.266 79.562 ;
               RECT 11.214 80.726 11.266 80.762 ;
               RECT 11.214 81.926 11.266 81.962 ;
               RECT 11.214 83.126 11.266 83.162 ;
               RECT 11.214 84.326 11.266 84.362 ;
               RECT 11.214 85.526 11.266 85.562 ;
               RECT 11.214 86.726 11.266 86.762 ;
               RECT 11.214 87.926 11.266 87.962 ;
               RECT 11.214 89.126 11.266 89.162 ;
               RECT 11.214 90.326 11.266 90.362 ;
               RECT 11.214 91.526 11.266 91.562 ;
               RECT 11.214 92.726 11.266 92.762 ;
               RECT 11.214 93.926 11.266 93.962 ;
               RECT 11.214 95.126 11.266 95.162 ;
               RECT 11.214 96.326 11.266 96.362 ;
               RECT 11.214 97.526 11.266 97.562 ;
               RECT 11.214 98.726 11.266 98.762 ;
               RECT 11.214 99.926 11.266 99.962 ;
               RECT 11.214 101.126 11.266 101.162 ;
               RECT 11.214 102.326 11.266 102.362 ;
               RECT 11.214 103.526 11.266 103.562 ;
               RECT 11.294 1.558 11.346 1.594 ;
               RECT 11.294 2.758 11.346 2.794 ;
               RECT 11.294 3.958 11.346 3.994 ;
               RECT 11.294 5.158 11.346 5.194 ;
               RECT 11.294 6.358 11.346 6.394 ;
               RECT 11.294 7.558 11.346 7.594 ;
               RECT 11.294 8.758 11.346 8.794 ;
               RECT 11.294 9.958 11.346 9.994 ;
               RECT 11.294 11.158 11.346 11.194 ;
               RECT 11.294 12.358 11.346 12.394 ;
               RECT 11.294 13.558 11.346 13.594 ;
               RECT 11.294 14.758 11.346 14.794 ;
               RECT 11.294 15.958 11.346 15.994 ;
               RECT 11.294 17.158 11.346 17.194 ;
               RECT 11.294 18.358 11.346 18.394 ;
               RECT 11.294 19.558 11.346 19.594 ;
               RECT 11.294 20.758 11.346 20.794 ;
               RECT 11.294 21.958 11.346 21.994 ;
               RECT 11.294 23.158 11.346 23.194 ;
               RECT 11.294 24.358 11.346 24.394 ;
               RECT 11.294 25.558 11.346 25.594 ;
               RECT 11.294 26.758 11.346 26.794 ;
               RECT 11.294 27.958 11.346 27.994 ;
               RECT 11.294 29.158 11.346 29.194 ;
               RECT 11.294 30.358 11.346 30.394 ;
               RECT 11.294 31.558 11.346 31.594 ;
               RECT 11.294 32.758 11.346 32.794 ;
               RECT 11.294 33.958 11.346 33.994 ;
               RECT 11.294 35.158 11.346 35.194 ;
               RECT 11.294 36.358 11.346 36.394 ;
               RECT 11.294 37.558 11.346 37.594 ;
               RECT 11.294 38.758 11.346 38.794 ;
               RECT 11.294 39.958 11.346 39.994 ;
               RECT 11.294 41.158 11.346 41.194 ;
               RECT 11.294 42.358 11.346 42.394 ;
               RECT 11.294 43.558 11.346 43.594 ;
               RECT 11.294 44.758 11.346 44.794 ;
               RECT 11.294 45.958 11.346 45.994 ;
               RECT 11.294 47.158 11.346 47.194 ;
               RECT 11.294 48.358 11.346 48.394 ;
               RECT 11.294 50.142 11.346 50.178 ;
               RECT 11.294 50.382 11.346 50.418 ;
               RECT 11.294 54.702 11.346 54.738 ;
               RECT 11.294 54.942 11.346 54.978 ;
               RECT 11.294 57.478 11.346 57.514 ;
               RECT 11.294 58.678 11.346 58.714 ;
               RECT 11.294 59.878 11.346 59.914 ;
               RECT 11.294 61.078 11.346 61.114 ;
               RECT 11.294 62.278 11.346 62.314 ;
               RECT 11.294 63.478 11.346 63.514 ;
               RECT 11.294 64.678 11.346 64.714 ;
               RECT 11.294 65.878 11.346 65.914 ;
               RECT 11.294 67.078 11.346 67.114 ;
               RECT 11.294 68.278 11.346 68.314 ;
               RECT 11.294 69.478 11.346 69.514 ;
               RECT 11.294 70.678 11.346 70.714 ;
               RECT 11.294 71.878 11.346 71.914 ;
               RECT 11.294 73.078 11.346 73.114 ;
               RECT 11.294 74.278 11.346 74.314 ;
               RECT 11.294 75.478 11.346 75.514 ;
               RECT 11.294 76.678 11.346 76.714 ;
               RECT 11.294 77.878 11.346 77.914 ;
               RECT 11.294 79.078 11.346 79.114 ;
               RECT 11.294 80.278 11.346 80.314 ;
               RECT 11.294 81.478 11.346 81.514 ;
               RECT 11.294 82.678 11.346 82.714 ;
               RECT 11.294 83.878 11.346 83.914 ;
               RECT 11.294 85.078 11.346 85.114 ;
               RECT 11.294 86.278 11.346 86.314 ;
               RECT 11.294 87.478 11.346 87.514 ;
               RECT 11.294 88.678 11.346 88.714 ;
               RECT 11.294 89.878 11.346 89.914 ;
               RECT 11.294 91.078 11.346 91.114 ;
               RECT 11.294 92.278 11.346 92.314 ;
               RECT 11.294 93.478 11.346 93.514 ;
               RECT 11.294 94.678 11.346 94.714 ;
               RECT 11.294 95.878 11.346 95.914 ;
               RECT 11.294 97.078 11.346 97.114 ;
               RECT 11.294 98.278 11.346 98.314 ;
               RECT 11.294 99.478 11.346 99.514 ;
               RECT 11.294 100.678 11.346 100.714 ;
               RECT 11.294 101.878 11.346 101.914 ;
               RECT 11.294 103.078 11.346 103.114 ;
               RECT 11.294 104.278 11.346 104.314 ;
               RECT 11.374 0.281 11.426 0.317 ;
               RECT 11.374 104.803 11.426 104.839 ;
               RECT 11.454 0.806 11.506 0.842 ;
               RECT 11.454 2.006 11.506 2.042 ;
               RECT 11.454 3.206 11.506 3.242 ;
               RECT 11.454 4.406 11.506 4.442 ;
               RECT 11.454 5.606 11.506 5.642 ;
               RECT 11.454 6.806 11.506 6.842 ;
               RECT 11.454 8.006 11.506 8.042 ;
               RECT 11.454 9.206 11.506 9.242 ;
               RECT 11.454 10.406 11.506 10.442 ;
               RECT 11.454 11.606 11.506 11.642 ;
               RECT 11.454 12.806 11.506 12.842 ;
               RECT 11.454 14.006 11.506 14.042 ;
               RECT 11.454 15.206 11.506 15.242 ;
               RECT 11.454 16.406 11.506 16.442 ;
               RECT 11.454 17.606 11.506 17.642 ;
               RECT 11.454 18.806 11.506 18.842 ;
               RECT 11.454 20.006 11.506 20.042 ;
               RECT 11.454 21.206 11.506 21.242 ;
               RECT 11.454 22.406 11.506 22.442 ;
               RECT 11.454 23.606 11.506 23.642 ;
               RECT 11.454 24.806 11.506 24.842 ;
               RECT 11.454 26.006 11.506 26.042 ;
               RECT 11.454 27.206 11.506 27.242 ;
               RECT 11.454 28.406 11.506 28.442 ;
               RECT 11.454 29.606 11.506 29.642 ;
               RECT 11.454 30.806 11.506 30.842 ;
               RECT 11.454 32.006 11.506 32.042 ;
               RECT 11.454 33.206 11.506 33.242 ;
               RECT 11.454 34.406 11.506 34.442 ;
               RECT 11.454 35.606 11.506 35.642 ;
               RECT 11.454 36.806 11.506 36.842 ;
               RECT 11.454 38.006 11.506 38.042 ;
               RECT 11.454 39.206 11.506 39.242 ;
               RECT 11.454 40.406 11.506 40.442 ;
               RECT 11.454 41.606 11.506 41.642 ;
               RECT 11.454 42.806 11.506 42.842 ;
               RECT 11.454 44.006 11.506 44.042 ;
               RECT 11.454 45.206 11.506 45.242 ;
               RECT 11.454 46.406 11.506 46.442 ;
               RECT 11.454 47.606 11.506 47.642 ;
               RECT 11.454 49.422 11.506 49.458 ;
               RECT 11.454 49.662 11.506 49.698 ;
               RECT 11.454 51.102 11.506 51.138 ;
               RECT 11.454 51.582 11.506 51.618 ;
               RECT 11.454 53.502 11.506 53.538 ;
               RECT 11.454 53.982 11.506 54.018 ;
               RECT 11.454 55.422 11.506 55.458 ;
               RECT 11.454 55.662 11.506 55.698 ;
               RECT 11.454 56.726 11.506 56.762 ;
               RECT 11.454 57.926 11.506 57.962 ;
               RECT 11.454 59.126 11.506 59.162 ;
               RECT 11.454 60.326 11.506 60.362 ;
               RECT 11.454 61.526 11.506 61.562 ;
               RECT 11.454 62.726 11.506 62.762 ;
               RECT 11.454 63.926 11.506 63.962 ;
               RECT 11.454 65.126 11.506 65.162 ;
               RECT 11.454 66.326 11.506 66.362 ;
               RECT 11.454 67.526 11.506 67.562 ;
               RECT 11.454 68.726 11.506 68.762 ;
               RECT 11.454 69.926 11.506 69.962 ;
               RECT 11.454 71.126 11.506 71.162 ;
               RECT 11.454 72.326 11.506 72.362 ;
               RECT 11.454 73.526 11.506 73.562 ;
               RECT 11.454 74.726 11.506 74.762 ;
               RECT 11.454 75.926 11.506 75.962 ;
               RECT 11.454 77.126 11.506 77.162 ;
               RECT 11.454 78.326 11.506 78.362 ;
               RECT 11.454 79.526 11.506 79.562 ;
               RECT 11.454 80.726 11.506 80.762 ;
               RECT 11.454 81.926 11.506 81.962 ;
               RECT 11.454 83.126 11.506 83.162 ;
               RECT 11.454 84.326 11.506 84.362 ;
               RECT 11.454 85.526 11.506 85.562 ;
               RECT 11.454 86.726 11.506 86.762 ;
               RECT 11.454 87.926 11.506 87.962 ;
               RECT 11.454 89.126 11.506 89.162 ;
               RECT 11.454 90.326 11.506 90.362 ;
               RECT 11.454 91.526 11.506 91.562 ;
               RECT 11.454 92.726 11.506 92.762 ;
               RECT 11.454 93.926 11.506 93.962 ;
               RECT 11.454 95.126 11.506 95.162 ;
               RECT 11.454 96.326 11.506 96.362 ;
               RECT 11.454 97.526 11.506 97.562 ;
               RECT 11.454 98.726 11.506 98.762 ;
               RECT 11.454 99.926 11.506 99.962 ;
               RECT 11.454 101.126 11.506 101.162 ;
               RECT 11.454 102.326 11.506 102.362 ;
               RECT 11.454 103.526 11.506 103.562 ;
               RECT 11.534 1.558 11.586 1.594 ;
               RECT 11.534 2.758 11.586 2.794 ;
               RECT 11.534 3.958 11.586 3.994 ;
               RECT 11.534 5.158 11.586 5.194 ;
               RECT 11.534 6.358 11.586 6.394 ;
               RECT 11.534 7.558 11.586 7.594 ;
               RECT 11.534 8.758 11.586 8.794 ;
               RECT 11.534 9.958 11.586 9.994 ;
               RECT 11.534 11.158 11.586 11.194 ;
               RECT 11.534 12.358 11.586 12.394 ;
               RECT 11.534 13.558 11.586 13.594 ;
               RECT 11.534 14.758 11.586 14.794 ;
               RECT 11.534 15.958 11.586 15.994 ;
               RECT 11.534 17.158 11.586 17.194 ;
               RECT 11.534 18.358 11.586 18.394 ;
               RECT 11.534 19.558 11.586 19.594 ;
               RECT 11.534 20.758 11.586 20.794 ;
               RECT 11.534 21.958 11.586 21.994 ;
               RECT 11.534 23.158 11.586 23.194 ;
               RECT 11.534 24.358 11.586 24.394 ;
               RECT 11.534 25.558 11.586 25.594 ;
               RECT 11.534 26.758 11.586 26.794 ;
               RECT 11.534 27.958 11.586 27.994 ;
               RECT 11.534 29.158 11.586 29.194 ;
               RECT 11.534 30.358 11.586 30.394 ;
               RECT 11.534 31.558 11.586 31.594 ;
               RECT 11.534 32.758 11.586 32.794 ;
               RECT 11.534 33.958 11.586 33.994 ;
               RECT 11.534 35.158 11.586 35.194 ;
               RECT 11.534 36.358 11.586 36.394 ;
               RECT 11.534 37.558 11.586 37.594 ;
               RECT 11.534 38.758 11.586 38.794 ;
               RECT 11.534 39.958 11.586 39.994 ;
               RECT 11.534 41.158 11.586 41.194 ;
               RECT 11.534 42.358 11.586 42.394 ;
               RECT 11.534 43.558 11.586 43.594 ;
               RECT 11.534 44.758 11.586 44.794 ;
               RECT 11.534 45.958 11.586 45.994 ;
               RECT 11.534 47.158 11.586 47.194 ;
               RECT 11.534 48.358 11.586 48.394 ;
               RECT 11.534 50.142 11.586 50.178 ;
               RECT 11.534 50.382 11.586 50.418 ;
               RECT 11.534 54.702 11.586 54.738 ;
               RECT 11.534 54.942 11.586 54.978 ;
               RECT 11.534 57.478 11.586 57.514 ;
               RECT 11.534 58.678 11.586 58.714 ;
               RECT 11.534 59.878 11.586 59.914 ;
               RECT 11.534 61.078 11.586 61.114 ;
               RECT 11.534 62.278 11.586 62.314 ;
               RECT 11.534 63.478 11.586 63.514 ;
               RECT 11.534 64.678 11.586 64.714 ;
               RECT 11.534 65.878 11.586 65.914 ;
               RECT 11.534 67.078 11.586 67.114 ;
               RECT 11.534 68.278 11.586 68.314 ;
               RECT 11.534 69.478 11.586 69.514 ;
               RECT 11.534 70.678 11.586 70.714 ;
               RECT 11.534 71.878 11.586 71.914 ;
               RECT 11.534 73.078 11.586 73.114 ;
               RECT 11.534 74.278 11.586 74.314 ;
               RECT 11.534 75.478 11.586 75.514 ;
               RECT 11.534 76.678 11.586 76.714 ;
               RECT 11.534 77.878 11.586 77.914 ;
               RECT 11.534 79.078 11.586 79.114 ;
               RECT 11.534 80.278 11.586 80.314 ;
               RECT 11.534 81.478 11.586 81.514 ;
               RECT 11.534 82.678 11.586 82.714 ;
               RECT 11.534 83.878 11.586 83.914 ;
               RECT 11.534 85.078 11.586 85.114 ;
               RECT 11.534 86.278 11.586 86.314 ;
               RECT 11.534 87.478 11.586 87.514 ;
               RECT 11.534 88.678 11.586 88.714 ;
               RECT 11.534 89.878 11.586 89.914 ;
               RECT 11.534 91.078 11.586 91.114 ;
               RECT 11.534 92.278 11.586 92.314 ;
               RECT 11.534 93.478 11.586 93.514 ;
               RECT 11.534 94.678 11.586 94.714 ;
               RECT 11.534 95.878 11.586 95.914 ;
               RECT 11.534 97.078 11.586 97.114 ;
               RECT 11.534 98.278 11.586 98.314 ;
               RECT 11.534 99.478 11.586 99.514 ;
               RECT 11.534 100.678 11.586 100.714 ;
               RECT 11.534 101.878 11.586 101.914 ;
               RECT 11.534 103.078 11.586 103.114 ;
               RECT 11.534 104.278 11.586 104.314 ;
               RECT 11.614 0.806 11.666 0.842 ;
               RECT 11.614 2.006 11.666 2.042 ;
               RECT 11.614 3.206 11.666 3.242 ;
               RECT 11.614 4.406 11.666 4.442 ;
               RECT 11.614 5.606 11.666 5.642 ;
               RECT 11.614 6.806 11.666 6.842 ;
               RECT 11.614 8.006 11.666 8.042 ;
               RECT 11.614 9.206 11.666 9.242 ;
               RECT 11.614 10.406 11.666 10.442 ;
               RECT 11.614 11.606 11.666 11.642 ;
               RECT 11.614 12.806 11.666 12.842 ;
               RECT 11.614 14.006 11.666 14.042 ;
               RECT 11.614 15.206 11.666 15.242 ;
               RECT 11.614 16.406 11.666 16.442 ;
               RECT 11.614 17.606 11.666 17.642 ;
               RECT 11.614 18.806 11.666 18.842 ;
               RECT 11.614 20.006 11.666 20.042 ;
               RECT 11.614 21.206 11.666 21.242 ;
               RECT 11.614 22.406 11.666 22.442 ;
               RECT 11.614 23.606 11.666 23.642 ;
               RECT 11.614 24.806 11.666 24.842 ;
               RECT 11.614 26.006 11.666 26.042 ;
               RECT 11.614 27.206 11.666 27.242 ;
               RECT 11.614 28.406 11.666 28.442 ;
               RECT 11.614 29.606 11.666 29.642 ;
               RECT 11.614 30.806 11.666 30.842 ;
               RECT 11.614 32.006 11.666 32.042 ;
               RECT 11.614 33.206 11.666 33.242 ;
               RECT 11.614 34.406 11.666 34.442 ;
               RECT 11.614 35.606 11.666 35.642 ;
               RECT 11.614 36.806 11.666 36.842 ;
               RECT 11.614 38.006 11.666 38.042 ;
               RECT 11.614 39.206 11.666 39.242 ;
               RECT 11.614 40.406 11.666 40.442 ;
               RECT 11.614 41.606 11.666 41.642 ;
               RECT 11.614 42.806 11.666 42.842 ;
               RECT 11.614 44.006 11.666 44.042 ;
               RECT 11.614 45.206 11.666 45.242 ;
               RECT 11.614 46.406 11.666 46.442 ;
               RECT 11.614 47.606 11.666 47.642 ;
               RECT 11.614 49.422 11.666 49.458 ;
               RECT 11.614 49.662 11.666 49.698 ;
               RECT 11.614 55.422 11.666 55.458 ;
               RECT 11.614 55.662 11.666 55.698 ;
               RECT 11.614 56.726 11.666 56.762 ;
               RECT 11.614 57.926 11.666 57.962 ;
               RECT 11.614 59.126 11.666 59.162 ;
               RECT 11.614 60.326 11.666 60.362 ;
               RECT 11.614 61.526 11.666 61.562 ;
               RECT 11.614 62.726 11.666 62.762 ;
               RECT 11.614 63.926 11.666 63.962 ;
               RECT 11.614 65.126 11.666 65.162 ;
               RECT 11.614 66.326 11.666 66.362 ;
               RECT 11.614 67.526 11.666 67.562 ;
               RECT 11.614 68.726 11.666 68.762 ;
               RECT 11.614 69.926 11.666 69.962 ;
               RECT 11.614 71.126 11.666 71.162 ;
               RECT 11.614 72.326 11.666 72.362 ;
               RECT 11.614 73.526 11.666 73.562 ;
               RECT 11.614 74.726 11.666 74.762 ;
               RECT 11.614 75.926 11.666 75.962 ;
               RECT 11.614 77.126 11.666 77.162 ;
               RECT 11.614 78.326 11.666 78.362 ;
               RECT 11.614 79.526 11.666 79.562 ;
               RECT 11.614 80.726 11.666 80.762 ;
               RECT 11.614 81.926 11.666 81.962 ;
               RECT 11.614 83.126 11.666 83.162 ;
               RECT 11.614 84.326 11.666 84.362 ;
               RECT 11.614 85.526 11.666 85.562 ;
               RECT 11.614 86.726 11.666 86.762 ;
               RECT 11.614 87.926 11.666 87.962 ;
               RECT 11.614 89.126 11.666 89.162 ;
               RECT 11.614 90.326 11.666 90.362 ;
               RECT 11.614 91.526 11.666 91.562 ;
               RECT 11.614 92.726 11.666 92.762 ;
               RECT 11.614 93.926 11.666 93.962 ;
               RECT 11.614 95.126 11.666 95.162 ;
               RECT 11.614 96.326 11.666 96.362 ;
               RECT 11.614 97.526 11.666 97.562 ;
               RECT 11.614 98.726 11.666 98.762 ;
               RECT 11.614 99.926 11.666 99.962 ;
               RECT 11.614 101.126 11.666 101.162 ;
               RECT 11.614 102.326 11.666 102.362 ;
               RECT 11.614 103.526 11.666 103.562 ;
               RECT 11.694 1.558 11.746 1.594 ;
               RECT 11.694 2.758 11.746 2.794 ;
               RECT 11.694 3.958 11.746 3.994 ;
               RECT 11.694 5.158 11.746 5.194 ;
               RECT 11.694 6.358 11.746 6.394 ;
               RECT 11.694 7.558 11.746 7.594 ;
               RECT 11.694 8.758 11.746 8.794 ;
               RECT 11.694 9.958 11.746 9.994 ;
               RECT 11.694 11.158 11.746 11.194 ;
               RECT 11.694 12.358 11.746 12.394 ;
               RECT 11.694 13.558 11.746 13.594 ;
               RECT 11.694 14.758 11.746 14.794 ;
               RECT 11.694 15.958 11.746 15.994 ;
               RECT 11.694 17.158 11.746 17.194 ;
               RECT 11.694 18.358 11.746 18.394 ;
               RECT 11.694 19.558 11.746 19.594 ;
               RECT 11.694 20.758 11.746 20.794 ;
               RECT 11.694 21.958 11.746 21.994 ;
               RECT 11.694 23.158 11.746 23.194 ;
               RECT 11.694 24.358 11.746 24.394 ;
               RECT 11.694 25.558 11.746 25.594 ;
               RECT 11.694 26.758 11.746 26.794 ;
               RECT 11.694 27.958 11.746 27.994 ;
               RECT 11.694 29.158 11.746 29.194 ;
               RECT 11.694 30.358 11.746 30.394 ;
               RECT 11.694 31.558 11.746 31.594 ;
               RECT 11.694 32.758 11.746 32.794 ;
               RECT 11.694 33.958 11.746 33.994 ;
               RECT 11.694 35.158 11.746 35.194 ;
               RECT 11.694 36.358 11.746 36.394 ;
               RECT 11.694 37.558 11.746 37.594 ;
               RECT 11.694 38.758 11.746 38.794 ;
               RECT 11.694 39.958 11.746 39.994 ;
               RECT 11.694 41.158 11.746 41.194 ;
               RECT 11.694 42.358 11.746 42.394 ;
               RECT 11.694 43.558 11.746 43.594 ;
               RECT 11.694 44.758 11.746 44.794 ;
               RECT 11.694 45.958 11.746 45.994 ;
               RECT 11.694 47.158 11.746 47.194 ;
               RECT 11.694 48.358 11.746 48.394 ;
               RECT 11.694 50.142 11.746 50.178 ;
               RECT 11.694 50.382 11.746 50.418 ;
               RECT 11.694 54.702 11.746 54.738 ;
               RECT 11.694 54.942 11.746 54.978 ;
               RECT 11.694 57.478 11.746 57.514 ;
               RECT 11.694 58.678 11.746 58.714 ;
               RECT 11.694 59.878 11.746 59.914 ;
               RECT 11.694 61.078 11.746 61.114 ;
               RECT 11.694 62.278 11.746 62.314 ;
               RECT 11.694 63.478 11.746 63.514 ;
               RECT 11.694 64.678 11.746 64.714 ;
               RECT 11.694 65.878 11.746 65.914 ;
               RECT 11.694 67.078 11.746 67.114 ;
               RECT 11.694 68.278 11.746 68.314 ;
               RECT 11.694 69.478 11.746 69.514 ;
               RECT 11.694 70.678 11.746 70.714 ;
               RECT 11.694 71.878 11.746 71.914 ;
               RECT 11.694 73.078 11.746 73.114 ;
               RECT 11.694 74.278 11.746 74.314 ;
               RECT 11.694 75.478 11.746 75.514 ;
               RECT 11.694 76.678 11.746 76.714 ;
               RECT 11.694 77.878 11.746 77.914 ;
               RECT 11.694 79.078 11.746 79.114 ;
               RECT 11.694 80.278 11.746 80.314 ;
               RECT 11.694 81.478 11.746 81.514 ;
               RECT 11.694 82.678 11.746 82.714 ;
               RECT 11.694 83.878 11.746 83.914 ;
               RECT 11.694 85.078 11.746 85.114 ;
               RECT 11.694 86.278 11.746 86.314 ;
               RECT 11.694 87.478 11.746 87.514 ;
               RECT 11.694 88.678 11.746 88.714 ;
               RECT 11.694 89.878 11.746 89.914 ;
               RECT 11.694 91.078 11.746 91.114 ;
               RECT 11.694 92.278 11.746 92.314 ;
               RECT 11.694 93.478 11.746 93.514 ;
               RECT 11.694 94.678 11.746 94.714 ;
               RECT 11.694 95.878 11.746 95.914 ;
               RECT 11.694 97.078 11.746 97.114 ;
               RECT 11.694 98.278 11.746 98.314 ;
               RECT 11.694 99.478 11.746 99.514 ;
               RECT 11.694 100.678 11.746 100.714 ;
               RECT 11.694 101.878 11.746 101.914 ;
               RECT 11.694 103.078 11.746 103.114 ;
               RECT 11.694 104.278 11.746 104.314 ;
               RECT 11.774 0.281 11.826 0.317 ;
               RECT 11.774 104.803 11.826 104.839 ;
               RECT 11.854 0.806 11.906 0.842 ;
               RECT 11.854 2.006 11.906 2.042 ;
               RECT 11.854 3.206 11.906 3.242 ;
               RECT 11.854 4.406 11.906 4.442 ;
               RECT 11.854 5.606 11.906 5.642 ;
               RECT 11.854 6.806 11.906 6.842 ;
               RECT 11.854 8.006 11.906 8.042 ;
               RECT 11.854 9.206 11.906 9.242 ;
               RECT 11.854 10.406 11.906 10.442 ;
               RECT 11.854 11.606 11.906 11.642 ;
               RECT 11.854 12.806 11.906 12.842 ;
               RECT 11.854 14.006 11.906 14.042 ;
               RECT 11.854 15.206 11.906 15.242 ;
               RECT 11.854 16.406 11.906 16.442 ;
               RECT 11.854 17.606 11.906 17.642 ;
               RECT 11.854 18.806 11.906 18.842 ;
               RECT 11.854 20.006 11.906 20.042 ;
               RECT 11.854 21.206 11.906 21.242 ;
               RECT 11.854 22.406 11.906 22.442 ;
               RECT 11.854 23.606 11.906 23.642 ;
               RECT 11.854 24.806 11.906 24.842 ;
               RECT 11.854 26.006 11.906 26.042 ;
               RECT 11.854 27.206 11.906 27.242 ;
               RECT 11.854 28.406 11.906 28.442 ;
               RECT 11.854 29.606 11.906 29.642 ;
               RECT 11.854 30.806 11.906 30.842 ;
               RECT 11.854 32.006 11.906 32.042 ;
               RECT 11.854 33.206 11.906 33.242 ;
               RECT 11.854 34.406 11.906 34.442 ;
               RECT 11.854 35.606 11.906 35.642 ;
               RECT 11.854 36.806 11.906 36.842 ;
               RECT 11.854 38.006 11.906 38.042 ;
               RECT 11.854 39.206 11.906 39.242 ;
               RECT 11.854 40.406 11.906 40.442 ;
               RECT 11.854 41.606 11.906 41.642 ;
               RECT 11.854 42.806 11.906 42.842 ;
               RECT 11.854 44.006 11.906 44.042 ;
               RECT 11.854 45.206 11.906 45.242 ;
               RECT 11.854 46.406 11.906 46.442 ;
               RECT 11.854 47.606 11.906 47.642 ;
               RECT 11.854 49.422 11.906 49.458 ;
               RECT 11.854 49.662 11.906 49.698 ;
               RECT 11.854 55.422 11.906 55.458 ;
               RECT 11.854 55.662 11.906 55.698 ;
               RECT 11.854 56.726 11.906 56.762 ;
               RECT 11.854 57.926 11.906 57.962 ;
               RECT 11.854 59.126 11.906 59.162 ;
               RECT 11.854 60.326 11.906 60.362 ;
               RECT 11.854 61.526 11.906 61.562 ;
               RECT 11.854 62.726 11.906 62.762 ;
               RECT 11.854 63.926 11.906 63.962 ;
               RECT 11.854 65.126 11.906 65.162 ;
               RECT 11.854 66.326 11.906 66.362 ;
               RECT 11.854 67.526 11.906 67.562 ;
               RECT 11.854 68.726 11.906 68.762 ;
               RECT 11.854 69.926 11.906 69.962 ;
               RECT 11.854 71.126 11.906 71.162 ;
               RECT 11.854 72.326 11.906 72.362 ;
               RECT 11.854 73.526 11.906 73.562 ;
               RECT 11.854 74.726 11.906 74.762 ;
               RECT 11.854 75.926 11.906 75.962 ;
               RECT 11.854 77.126 11.906 77.162 ;
               RECT 11.854 78.326 11.906 78.362 ;
               RECT 11.854 79.526 11.906 79.562 ;
               RECT 11.854 80.726 11.906 80.762 ;
               RECT 11.854 81.926 11.906 81.962 ;
               RECT 11.854 83.126 11.906 83.162 ;
               RECT 11.854 84.326 11.906 84.362 ;
               RECT 11.854 85.526 11.906 85.562 ;
               RECT 11.854 86.726 11.906 86.762 ;
               RECT 11.854 87.926 11.906 87.962 ;
               RECT 11.854 89.126 11.906 89.162 ;
               RECT 11.854 90.326 11.906 90.362 ;
               RECT 11.854 91.526 11.906 91.562 ;
               RECT 11.854 92.726 11.906 92.762 ;
               RECT 11.854 93.926 11.906 93.962 ;
               RECT 11.854 95.126 11.906 95.162 ;
               RECT 11.854 96.326 11.906 96.362 ;
               RECT 11.854 97.526 11.906 97.562 ;
               RECT 11.854 98.726 11.906 98.762 ;
               RECT 11.854 99.926 11.906 99.962 ;
               RECT 11.854 101.126 11.906 101.162 ;
               RECT 11.854 102.326 11.906 102.362 ;
               RECT 11.854 103.526 11.906 103.562 ;
               RECT 11.934 1.558 11.986 1.594 ;
               RECT 11.934 2.758 11.986 2.794 ;
               RECT 11.934 3.958 11.986 3.994 ;
               RECT 11.934 5.158 11.986 5.194 ;
               RECT 11.934 6.358 11.986 6.394 ;
               RECT 11.934 7.558 11.986 7.594 ;
               RECT 11.934 8.758 11.986 8.794 ;
               RECT 11.934 9.958 11.986 9.994 ;
               RECT 11.934 11.158 11.986 11.194 ;
               RECT 11.934 12.358 11.986 12.394 ;
               RECT 11.934 13.558 11.986 13.594 ;
               RECT 11.934 14.758 11.986 14.794 ;
               RECT 11.934 15.958 11.986 15.994 ;
               RECT 11.934 17.158 11.986 17.194 ;
               RECT 11.934 18.358 11.986 18.394 ;
               RECT 11.934 19.558 11.986 19.594 ;
               RECT 11.934 20.758 11.986 20.794 ;
               RECT 11.934 21.958 11.986 21.994 ;
               RECT 11.934 23.158 11.986 23.194 ;
               RECT 11.934 24.358 11.986 24.394 ;
               RECT 11.934 25.558 11.986 25.594 ;
               RECT 11.934 26.758 11.986 26.794 ;
               RECT 11.934 27.958 11.986 27.994 ;
               RECT 11.934 29.158 11.986 29.194 ;
               RECT 11.934 30.358 11.986 30.394 ;
               RECT 11.934 31.558 11.986 31.594 ;
               RECT 11.934 32.758 11.986 32.794 ;
               RECT 11.934 33.958 11.986 33.994 ;
               RECT 11.934 35.158 11.986 35.194 ;
               RECT 11.934 36.358 11.986 36.394 ;
               RECT 11.934 37.558 11.986 37.594 ;
               RECT 11.934 38.758 11.986 38.794 ;
               RECT 11.934 39.958 11.986 39.994 ;
               RECT 11.934 41.158 11.986 41.194 ;
               RECT 11.934 42.358 11.986 42.394 ;
               RECT 11.934 43.558 11.986 43.594 ;
               RECT 11.934 44.758 11.986 44.794 ;
               RECT 11.934 45.958 11.986 45.994 ;
               RECT 11.934 47.158 11.986 47.194 ;
               RECT 11.934 48.358 11.986 48.394 ;
               RECT 11.934 50.142 11.986 50.178 ;
               RECT 11.934 50.382 11.986 50.418 ;
               RECT 11.934 54.702 11.986 54.738 ;
               RECT 11.934 54.942 11.986 54.978 ;
               RECT 11.934 57.478 11.986 57.514 ;
               RECT 11.934 58.678 11.986 58.714 ;
               RECT 11.934 59.878 11.986 59.914 ;
               RECT 11.934 61.078 11.986 61.114 ;
               RECT 11.934 62.278 11.986 62.314 ;
               RECT 11.934 63.478 11.986 63.514 ;
               RECT 11.934 64.678 11.986 64.714 ;
               RECT 11.934 65.878 11.986 65.914 ;
               RECT 11.934 67.078 11.986 67.114 ;
               RECT 11.934 68.278 11.986 68.314 ;
               RECT 11.934 69.478 11.986 69.514 ;
               RECT 11.934 70.678 11.986 70.714 ;
               RECT 11.934 71.878 11.986 71.914 ;
               RECT 11.934 73.078 11.986 73.114 ;
               RECT 11.934 74.278 11.986 74.314 ;
               RECT 11.934 75.478 11.986 75.514 ;
               RECT 11.934 76.678 11.986 76.714 ;
               RECT 11.934 77.878 11.986 77.914 ;
               RECT 11.934 79.078 11.986 79.114 ;
               RECT 11.934 80.278 11.986 80.314 ;
               RECT 11.934 81.478 11.986 81.514 ;
               RECT 11.934 82.678 11.986 82.714 ;
               RECT 11.934 83.878 11.986 83.914 ;
               RECT 11.934 85.078 11.986 85.114 ;
               RECT 11.934 86.278 11.986 86.314 ;
               RECT 11.934 87.478 11.986 87.514 ;
               RECT 11.934 88.678 11.986 88.714 ;
               RECT 11.934 89.878 11.986 89.914 ;
               RECT 11.934 91.078 11.986 91.114 ;
               RECT 11.934 92.278 11.986 92.314 ;
               RECT 11.934 93.478 11.986 93.514 ;
               RECT 11.934 94.678 11.986 94.714 ;
               RECT 11.934 95.878 11.986 95.914 ;
               RECT 11.934 97.078 11.986 97.114 ;
               RECT 11.934 98.278 11.986 98.314 ;
               RECT 11.934 99.478 11.986 99.514 ;
               RECT 11.934 100.678 11.986 100.714 ;
               RECT 11.934 101.878 11.986 101.914 ;
               RECT 11.934 103.078 11.986 103.114 ;
               RECT 11.934 104.278 11.986 104.314 ;
               RECT 12.014 0.806 12.066 0.842 ;
               RECT 12.014 2.006 12.066 2.042 ;
               RECT 12.014 3.206 12.066 3.242 ;
               RECT 12.014 4.406 12.066 4.442 ;
               RECT 12.014 5.606 12.066 5.642 ;
               RECT 12.014 6.806 12.066 6.842 ;
               RECT 12.014 8.006 12.066 8.042 ;
               RECT 12.014 9.206 12.066 9.242 ;
               RECT 12.014 10.406 12.066 10.442 ;
               RECT 12.014 11.606 12.066 11.642 ;
               RECT 12.014 12.806 12.066 12.842 ;
               RECT 12.014 14.006 12.066 14.042 ;
               RECT 12.014 15.206 12.066 15.242 ;
               RECT 12.014 16.406 12.066 16.442 ;
               RECT 12.014 17.606 12.066 17.642 ;
               RECT 12.014 18.806 12.066 18.842 ;
               RECT 12.014 20.006 12.066 20.042 ;
               RECT 12.014 21.206 12.066 21.242 ;
               RECT 12.014 22.406 12.066 22.442 ;
               RECT 12.014 23.606 12.066 23.642 ;
               RECT 12.014 24.806 12.066 24.842 ;
               RECT 12.014 26.006 12.066 26.042 ;
               RECT 12.014 27.206 12.066 27.242 ;
               RECT 12.014 28.406 12.066 28.442 ;
               RECT 12.014 29.606 12.066 29.642 ;
               RECT 12.014 30.806 12.066 30.842 ;
               RECT 12.014 32.006 12.066 32.042 ;
               RECT 12.014 33.206 12.066 33.242 ;
               RECT 12.014 34.406 12.066 34.442 ;
               RECT 12.014 35.606 12.066 35.642 ;
               RECT 12.014 36.806 12.066 36.842 ;
               RECT 12.014 38.006 12.066 38.042 ;
               RECT 12.014 39.206 12.066 39.242 ;
               RECT 12.014 40.406 12.066 40.442 ;
               RECT 12.014 41.606 12.066 41.642 ;
               RECT 12.014 42.806 12.066 42.842 ;
               RECT 12.014 44.006 12.066 44.042 ;
               RECT 12.014 45.206 12.066 45.242 ;
               RECT 12.014 46.406 12.066 46.442 ;
               RECT 12.014 47.606 12.066 47.642 ;
               RECT 12.014 49.422 12.066 49.458 ;
               RECT 12.014 49.662 12.066 49.698 ;
               RECT 12.014 55.422 12.066 55.458 ;
               RECT 12.014 55.662 12.066 55.698 ;
               RECT 12.014 56.726 12.066 56.762 ;
               RECT 12.014 57.926 12.066 57.962 ;
               RECT 12.014 59.126 12.066 59.162 ;
               RECT 12.014 60.326 12.066 60.362 ;
               RECT 12.014 61.526 12.066 61.562 ;
               RECT 12.014 62.726 12.066 62.762 ;
               RECT 12.014 63.926 12.066 63.962 ;
               RECT 12.014 65.126 12.066 65.162 ;
               RECT 12.014 66.326 12.066 66.362 ;
               RECT 12.014 67.526 12.066 67.562 ;
               RECT 12.014 68.726 12.066 68.762 ;
               RECT 12.014 69.926 12.066 69.962 ;
               RECT 12.014 71.126 12.066 71.162 ;
               RECT 12.014 72.326 12.066 72.362 ;
               RECT 12.014 73.526 12.066 73.562 ;
               RECT 12.014 74.726 12.066 74.762 ;
               RECT 12.014 75.926 12.066 75.962 ;
               RECT 12.014 77.126 12.066 77.162 ;
               RECT 12.014 78.326 12.066 78.362 ;
               RECT 12.014 79.526 12.066 79.562 ;
               RECT 12.014 80.726 12.066 80.762 ;
               RECT 12.014 81.926 12.066 81.962 ;
               RECT 12.014 83.126 12.066 83.162 ;
               RECT 12.014 84.326 12.066 84.362 ;
               RECT 12.014 85.526 12.066 85.562 ;
               RECT 12.014 86.726 12.066 86.762 ;
               RECT 12.014 87.926 12.066 87.962 ;
               RECT 12.014 89.126 12.066 89.162 ;
               RECT 12.014 90.326 12.066 90.362 ;
               RECT 12.014 91.526 12.066 91.562 ;
               RECT 12.014 92.726 12.066 92.762 ;
               RECT 12.014 93.926 12.066 93.962 ;
               RECT 12.014 95.126 12.066 95.162 ;
               RECT 12.014 96.326 12.066 96.362 ;
               RECT 12.014 97.526 12.066 97.562 ;
               RECT 12.014 98.726 12.066 98.762 ;
               RECT 12.014 99.926 12.066 99.962 ;
               RECT 12.014 101.126 12.066 101.162 ;
               RECT 12.014 102.326 12.066 102.362 ;
               RECT 12.014 103.526 12.066 103.562 ;
               RECT 12.094 1.558 12.146 1.594 ;
               RECT 12.094 2.758 12.146 2.794 ;
               RECT 12.094 3.958 12.146 3.994 ;
               RECT 12.094 5.158 12.146 5.194 ;
               RECT 12.094 6.358 12.146 6.394 ;
               RECT 12.094 7.558 12.146 7.594 ;
               RECT 12.094 8.758 12.146 8.794 ;
               RECT 12.094 9.958 12.146 9.994 ;
               RECT 12.094 11.158 12.146 11.194 ;
               RECT 12.094 12.358 12.146 12.394 ;
               RECT 12.094 13.558 12.146 13.594 ;
               RECT 12.094 14.758 12.146 14.794 ;
               RECT 12.094 15.958 12.146 15.994 ;
               RECT 12.094 17.158 12.146 17.194 ;
               RECT 12.094 18.358 12.146 18.394 ;
               RECT 12.094 19.558 12.146 19.594 ;
               RECT 12.094 20.758 12.146 20.794 ;
               RECT 12.094 21.958 12.146 21.994 ;
               RECT 12.094 23.158 12.146 23.194 ;
               RECT 12.094 24.358 12.146 24.394 ;
               RECT 12.094 25.558 12.146 25.594 ;
               RECT 12.094 26.758 12.146 26.794 ;
               RECT 12.094 27.958 12.146 27.994 ;
               RECT 12.094 29.158 12.146 29.194 ;
               RECT 12.094 30.358 12.146 30.394 ;
               RECT 12.094 31.558 12.146 31.594 ;
               RECT 12.094 32.758 12.146 32.794 ;
               RECT 12.094 33.958 12.146 33.994 ;
               RECT 12.094 35.158 12.146 35.194 ;
               RECT 12.094 36.358 12.146 36.394 ;
               RECT 12.094 37.558 12.146 37.594 ;
               RECT 12.094 38.758 12.146 38.794 ;
               RECT 12.094 39.958 12.146 39.994 ;
               RECT 12.094 41.158 12.146 41.194 ;
               RECT 12.094 42.358 12.146 42.394 ;
               RECT 12.094 43.558 12.146 43.594 ;
               RECT 12.094 44.758 12.146 44.794 ;
               RECT 12.094 45.958 12.146 45.994 ;
               RECT 12.094 47.158 12.146 47.194 ;
               RECT 12.094 48.358 12.146 48.394 ;
               RECT 12.094 50.142 12.146 50.178 ;
               RECT 12.094 50.382 12.146 50.418 ;
               RECT 12.094 54.702 12.146 54.738 ;
               RECT 12.094 54.942 12.146 54.978 ;
               RECT 12.094 57.478 12.146 57.514 ;
               RECT 12.094 58.678 12.146 58.714 ;
               RECT 12.094 59.878 12.146 59.914 ;
               RECT 12.094 61.078 12.146 61.114 ;
               RECT 12.094 62.278 12.146 62.314 ;
               RECT 12.094 63.478 12.146 63.514 ;
               RECT 12.094 64.678 12.146 64.714 ;
               RECT 12.094 65.878 12.146 65.914 ;
               RECT 12.094 67.078 12.146 67.114 ;
               RECT 12.094 68.278 12.146 68.314 ;
               RECT 12.094 69.478 12.146 69.514 ;
               RECT 12.094 70.678 12.146 70.714 ;
               RECT 12.094 71.878 12.146 71.914 ;
               RECT 12.094 73.078 12.146 73.114 ;
               RECT 12.094 74.278 12.146 74.314 ;
               RECT 12.094 75.478 12.146 75.514 ;
               RECT 12.094 76.678 12.146 76.714 ;
               RECT 12.094 77.878 12.146 77.914 ;
               RECT 12.094 79.078 12.146 79.114 ;
               RECT 12.094 80.278 12.146 80.314 ;
               RECT 12.094 81.478 12.146 81.514 ;
               RECT 12.094 82.678 12.146 82.714 ;
               RECT 12.094 83.878 12.146 83.914 ;
               RECT 12.094 85.078 12.146 85.114 ;
               RECT 12.094 86.278 12.146 86.314 ;
               RECT 12.094 87.478 12.146 87.514 ;
               RECT 12.094 88.678 12.146 88.714 ;
               RECT 12.094 89.878 12.146 89.914 ;
               RECT 12.094 91.078 12.146 91.114 ;
               RECT 12.094 92.278 12.146 92.314 ;
               RECT 12.094 93.478 12.146 93.514 ;
               RECT 12.094 94.678 12.146 94.714 ;
               RECT 12.094 95.878 12.146 95.914 ;
               RECT 12.094 97.078 12.146 97.114 ;
               RECT 12.094 98.278 12.146 98.314 ;
               RECT 12.094 99.478 12.146 99.514 ;
               RECT 12.094 100.678 12.146 100.714 ;
               RECT 12.094 101.878 12.146 101.914 ;
               RECT 12.094 103.078 12.146 103.114 ;
               RECT 12.094 104.278 12.146 104.314 ;
               RECT 12.174 0.281 12.226 0.317 ;
               RECT 12.174 104.803 12.226 104.839 ;
               RECT 12.254 0.806 12.306 0.842 ;
               RECT 12.254 2.006 12.306 2.042 ;
               RECT 12.254 3.206 12.306 3.242 ;
               RECT 12.254 4.406 12.306 4.442 ;
               RECT 12.254 5.606 12.306 5.642 ;
               RECT 12.254 6.806 12.306 6.842 ;
               RECT 12.254 8.006 12.306 8.042 ;
               RECT 12.254 9.206 12.306 9.242 ;
               RECT 12.254 10.406 12.306 10.442 ;
               RECT 12.254 11.606 12.306 11.642 ;
               RECT 12.254 12.806 12.306 12.842 ;
               RECT 12.254 14.006 12.306 14.042 ;
               RECT 12.254 15.206 12.306 15.242 ;
               RECT 12.254 16.406 12.306 16.442 ;
               RECT 12.254 17.606 12.306 17.642 ;
               RECT 12.254 18.806 12.306 18.842 ;
               RECT 12.254 20.006 12.306 20.042 ;
               RECT 12.254 21.206 12.306 21.242 ;
               RECT 12.254 22.406 12.306 22.442 ;
               RECT 12.254 23.606 12.306 23.642 ;
               RECT 12.254 24.806 12.306 24.842 ;
               RECT 12.254 26.006 12.306 26.042 ;
               RECT 12.254 27.206 12.306 27.242 ;
               RECT 12.254 28.406 12.306 28.442 ;
               RECT 12.254 29.606 12.306 29.642 ;
               RECT 12.254 30.806 12.306 30.842 ;
               RECT 12.254 32.006 12.306 32.042 ;
               RECT 12.254 33.206 12.306 33.242 ;
               RECT 12.254 34.406 12.306 34.442 ;
               RECT 12.254 35.606 12.306 35.642 ;
               RECT 12.254 36.806 12.306 36.842 ;
               RECT 12.254 38.006 12.306 38.042 ;
               RECT 12.254 39.206 12.306 39.242 ;
               RECT 12.254 40.406 12.306 40.442 ;
               RECT 12.254 41.606 12.306 41.642 ;
               RECT 12.254 42.806 12.306 42.842 ;
               RECT 12.254 44.006 12.306 44.042 ;
               RECT 12.254 45.206 12.306 45.242 ;
               RECT 12.254 46.406 12.306 46.442 ;
               RECT 12.254 47.606 12.306 47.642 ;
               RECT 12.254 49.422 12.306 49.458 ;
               RECT 12.254 49.662 12.306 49.698 ;
               RECT 12.254 51.102 12.306 51.138 ;
               RECT 12.254 51.582 12.306 51.618 ;
               RECT 12.254 53.502 12.306 53.538 ;
               RECT 12.254 53.982 12.306 54.018 ;
               RECT 12.254 55.422 12.306 55.458 ;
               RECT 12.254 55.662 12.306 55.698 ;
               RECT 12.254 56.726 12.306 56.762 ;
               RECT 12.254 57.926 12.306 57.962 ;
               RECT 12.254 59.126 12.306 59.162 ;
               RECT 12.254 60.326 12.306 60.362 ;
               RECT 12.254 61.526 12.306 61.562 ;
               RECT 12.254 62.726 12.306 62.762 ;
               RECT 12.254 63.926 12.306 63.962 ;
               RECT 12.254 65.126 12.306 65.162 ;
               RECT 12.254 66.326 12.306 66.362 ;
               RECT 12.254 67.526 12.306 67.562 ;
               RECT 12.254 68.726 12.306 68.762 ;
               RECT 12.254 69.926 12.306 69.962 ;
               RECT 12.254 71.126 12.306 71.162 ;
               RECT 12.254 72.326 12.306 72.362 ;
               RECT 12.254 73.526 12.306 73.562 ;
               RECT 12.254 74.726 12.306 74.762 ;
               RECT 12.254 75.926 12.306 75.962 ;
               RECT 12.254 77.126 12.306 77.162 ;
               RECT 12.254 78.326 12.306 78.362 ;
               RECT 12.254 79.526 12.306 79.562 ;
               RECT 12.254 80.726 12.306 80.762 ;
               RECT 12.254 81.926 12.306 81.962 ;
               RECT 12.254 83.126 12.306 83.162 ;
               RECT 12.254 84.326 12.306 84.362 ;
               RECT 12.254 85.526 12.306 85.562 ;
               RECT 12.254 86.726 12.306 86.762 ;
               RECT 12.254 87.926 12.306 87.962 ;
               RECT 12.254 89.126 12.306 89.162 ;
               RECT 12.254 90.326 12.306 90.362 ;
               RECT 12.254 91.526 12.306 91.562 ;
               RECT 12.254 92.726 12.306 92.762 ;
               RECT 12.254 93.926 12.306 93.962 ;
               RECT 12.254 95.126 12.306 95.162 ;
               RECT 12.254 96.326 12.306 96.362 ;
               RECT 12.254 97.526 12.306 97.562 ;
               RECT 12.254 98.726 12.306 98.762 ;
               RECT 12.254 99.926 12.306 99.962 ;
               RECT 12.254 101.126 12.306 101.162 ;
               RECT 12.254 102.326 12.306 102.362 ;
               RECT 12.254 103.526 12.306 103.562 ;
               RECT 12.334 1.558 12.386 1.594 ;
               RECT 12.334 2.758 12.386 2.794 ;
               RECT 12.334 3.958 12.386 3.994 ;
               RECT 12.334 5.158 12.386 5.194 ;
               RECT 12.334 6.358 12.386 6.394 ;
               RECT 12.334 7.558 12.386 7.594 ;
               RECT 12.334 8.758 12.386 8.794 ;
               RECT 12.334 9.958 12.386 9.994 ;
               RECT 12.334 11.158 12.386 11.194 ;
               RECT 12.334 12.358 12.386 12.394 ;
               RECT 12.334 13.558 12.386 13.594 ;
               RECT 12.334 14.758 12.386 14.794 ;
               RECT 12.334 15.958 12.386 15.994 ;
               RECT 12.334 17.158 12.386 17.194 ;
               RECT 12.334 18.358 12.386 18.394 ;
               RECT 12.334 19.558 12.386 19.594 ;
               RECT 12.334 20.758 12.386 20.794 ;
               RECT 12.334 21.958 12.386 21.994 ;
               RECT 12.334 23.158 12.386 23.194 ;
               RECT 12.334 24.358 12.386 24.394 ;
               RECT 12.334 25.558 12.386 25.594 ;
               RECT 12.334 26.758 12.386 26.794 ;
               RECT 12.334 27.958 12.386 27.994 ;
               RECT 12.334 29.158 12.386 29.194 ;
               RECT 12.334 30.358 12.386 30.394 ;
               RECT 12.334 31.558 12.386 31.594 ;
               RECT 12.334 32.758 12.386 32.794 ;
               RECT 12.334 33.958 12.386 33.994 ;
               RECT 12.334 35.158 12.386 35.194 ;
               RECT 12.334 36.358 12.386 36.394 ;
               RECT 12.334 37.558 12.386 37.594 ;
               RECT 12.334 38.758 12.386 38.794 ;
               RECT 12.334 39.958 12.386 39.994 ;
               RECT 12.334 41.158 12.386 41.194 ;
               RECT 12.334 42.358 12.386 42.394 ;
               RECT 12.334 43.558 12.386 43.594 ;
               RECT 12.334 44.758 12.386 44.794 ;
               RECT 12.334 45.958 12.386 45.994 ;
               RECT 12.334 47.158 12.386 47.194 ;
               RECT 12.334 48.358 12.386 48.394 ;
               RECT 12.334 50.142 12.386 50.178 ;
               RECT 12.334 50.382 12.386 50.418 ;
               RECT 12.334 54.702 12.386 54.738 ;
               RECT 12.334 54.942 12.386 54.978 ;
               RECT 12.334 57.478 12.386 57.514 ;
               RECT 12.334 58.678 12.386 58.714 ;
               RECT 12.334 59.878 12.386 59.914 ;
               RECT 12.334 61.078 12.386 61.114 ;
               RECT 12.334 62.278 12.386 62.314 ;
               RECT 12.334 63.478 12.386 63.514 ;
               RECT 12.334 64.678 12.386 64.714 ;
               RECT 12.334 65.878 12.386 65.914 ;
               RECT 12.334 67.078 12.386 67.114 ;
               RECT 12.334 68.278 12.386 68.314 ;
               RECT 12.334 69.478 12.386 69.514 ;
               RECT 12.334 70.678 12.386 70.714 ;
               RECT 12.334 71.878 12.386 71.914 ;
               RECT 12.334 73.078 12.386 73.114 ;
               RECT 12.334 74.278 12.386 74.314 ;
               RECT 12.334 75.478 12.386 75.514 ;
               RECT 12.334 76.678 12.386 76.714 ;
               RECT 12.334 77.878 12.386 77.914 ;
               RECT 12.334 79.078 12.386 79.114 ;
               RECT 12.334 80.278 12.386 80.314 ;
               RECT 12.334 81.478 12.386 81.514 ;
               RECT 12.334 82.678 12.386 82.714 ;
               RECT 12.334 83.878 12.386 83.914 ;
               RECT 12.334 85.078 12.386 85.114 ;
               RECT 12.334 86.278 12.386 86.314 ;
               RECT 12.334 87.478 12.386 87.514 ;
               RECT 12.334 88.678 12.386 88.714 ;
               RECT 12.334 89.878 12.386 89.914 ;
               RECT 12.334 91.078 12.386 91.114 ;
               RECT 12.334 92.278 12.386 92.314 ;
               RECT 12.334 93.478 12.386 93.514 ;
               RECT 12.334 94.678 12.386 94.714 ;
               RECT 12.334 95.878 12.386 95.914 ;
               RECT 12.334 97.078 12.386 97.114 ;
               RECT 12.334 98.278 12.386 98.314 ;
               RECT 12.334 99.478 12.386 99.514 ;
               RECT 12.334 100.678 12.386 100.714 ;
               RECT 12.334 101.878 12.386 101.914 ;
               RECT 12.334 103.078 12.386 103.114 ;
               RECT 12.334 104.278 12.386 104.314 ;
               RECT 12.414 0.806 12.466 0.842 ;
               RECT 12.414 2.006 12.466 2.042 ;
               RECT 12.414 3.206 12.466 3.242 ;
               RECT 12.414 4.406 12.466 4.442 ;
               RECT 12.414 5.606 12.466 5.642 ;
               RECT 12.414 6.806 12.466 6.842 ;
               RECT 12.414 8.006 12.466 8.042 ;
               RECT 12.414 9.206 12.466 9.242 ;
               RECT 12.414 10.406 12.466 10.442 ;
               RECT 12.414 11.606 12.466 11.642 ;
               RECT 12.414 12.806 12.466 12.842 ;
               RECT 12.414 14.006 12.466 14.042 ;
               RECT 12.414 15.206 12.466 15.242 ;
               RECT 12.414 16.406 12.466 16.442 ;
               RECT 12.414 17.606 12.466 17.642 ;
               RECT 12.414 18.806 12.466 18.842 ;
               RECT 12.414 20.006 12.466 20.042 ;
               RECT 12.414 21.206 12.466 21.242 ;
               RECT 12.414 22.406 12.466 22.442 ;
               RECT 12.414 23.606 12.466 23.642 ;
               RECT 12.414 24.806 12.466 24.842 ;
               RECT 12.414 26.006 12.466 26.042 ;
               RECT 12.414 27.206 12.466 27.242 ;
               RECT 12.414 28.406 12.466 28.442 ;
               RECT 12.414 29.606 12.466 29.642 ;
               RECT 12.414 30.806 12.466 30.842 ;
               RECT 12.414 32.006 12.466 32.042 ;
               RECT 12.414 33.206 12.466 33.242 ;
               RECT 12.414 34.406 12.466 34.442 ;
               RECT 12.414 35.606 12.466 35.642 ;
               RECT 12.414 36.806 12.466 36.842 ;
               RECT 12.414 38.006 12.466 38.042 ;
               RECT 12.414 39.206 12.466 39.242 ;
               RECT 12.414 40.406 12.466 40.442 ;
               RECT 12.414 41.606 12.466 41.642 ;
               RECT 12.414 42.806 12.466 42.842 ;
               RECT 12.414 44.006 12.466 44.042 ;
               RECT 12.414 45.206 12.466 45.242 ;
               RECT 12.414 46.406 12.466 46.442 ;
               RECT 12.414 47.606 12.466 47.642 ;
               RECT 12.414 49.422 12.466 49.458 ;
               RECT 12.414 49.662 12.466 49.698 ;
               RECT 12.414 55.422 12.466 55.458 ;
               RECT 12.414 55.662 12.466 55.698 ;
               RECT 12.414 56.726 12.466 56.762 ;
               RECT 12.414 57.926 12.466 57.962 ;
               RECT 12.414 59.126 12.466 59.162 ;
               RECT 12.414 60.326 12.466 60.362 ;
               RECT 12.414 61.526 12.466 61.562 ;
               RECT 12.414 62.726 12.466 62.762 ;
               RECT 12.414 63.926 12.466 63.962 ;
               RECT 12.414 65.126 12.466 65.162 ;
               RECT 12.414 66.326 12.466 66.362 ;
               RECT 12.414 67.526 12.466 67.562 ;
               RECT 12.414 68.726 12.466 68.762 ;
               RECT 12.414 69.926 12.466 69.962 ;
               RECT 12.414 71.126 12.466 71.162 ;
               RECT 12.414 72.326 12.466 72.362 ;
               RECT 12.414 73.526 12.466 73.562 ;
               RECT 12.414 74.726 12.466 74.762 ;
               RECT 12.414 75.926 12.466 75.962 ;
               RECT 12.414 77.126 12.466 77.162 ;
               RECT 12.414 78.326 12.466 78.362 ;
               RECT 12.414 79.526 12.466 79.562 ;
               RECT 12.414 80.726 12.466 80.762 ;
               RECT 12.414 81.926 12.466 81.962 ;
               RECT 12.414 83.126 12.466 83.162 ;
               RECT 12.414 84.326 12.466 84.362 ;
               RECT 12.414 85.526 12.466 85.562 ;
               RECT 12.414 86.726 12.466 86.762 ;
               RECT 12.414 87.926 12.466 87.962 ;
               RECT 12.414 89.126 12.466 89.162 ;
               RECT 12.414 90.326 12.466 90.362 ;
               RECT 12.414 91.526 12.466 91.562 ;
               RECT 12.414 92.726 12.466 92.762 ;
               RECT 12.414 93.926 12.466 93.962 ;
               RECT 12.414 95.126 12.466 95.162 ;
               RECT 12.414 96.326 12.466 96.362 ;
               RECT 12.414 97.526 12.466 97.562 ;
               RECT 12.414 98.726 12.466 98.762 ;
               RECT 12.414 99.926 12.466 99.962 ;
               RECT 12.414 101.126 12.466 101.162 ;
               RECT 12.414 102.326 12.466 102.362 ;
               RECT 12.414 103.526 12.466 103.562 ;
               RECT 12.494 1.558 12.546 1.594 ;
               RECT 12.494 2.758 12.546 2.794 ;
               RECT 12.494 3.958 12.546 3.994 ;
               RECT 12.494 5.158 12.546 5.194 ;
               RECT 12.494 6.358 12.546 6.394 ;
               RECT 12.494 7.558 12.546 7.594 ;
               RECT 12.494 8.758 12.546 8.794 ;
               RECT 12.494 9.958 12.546 9.994 ;
               RECT 12.494 11.158 12.546 11.194 ;
               RECT 12.494 12.358 12.546 12.394 ;
               RECT 12.494 13.558 12.546 13.594 ;
               RECT 12.494 14.758 12.546 14.794 ;
               RECT 12.494 15.958 12.546 15.994 ;
               RECT 12.494 17.158 12.546 17.194 ;
               RECT 12.494 18.358 12.546 18.394 ;
               RECT 12.494 19.558 12.546 19.594 ;
               RECT 12.494 20.758 12.546 20.794 ;
               RECT 12.494 21.958 12.546 21.994 ;
               RECT 12.494 23.158 12.546 23.194 ;
               RECT 12.494 24.358 12.546 24.394 ;
               RECT 12.494 25.558 12.546 25.594 ;
               RECT 12.494 26.758 12.546 26.794 ;
               RECT 12.494 27.958 12.546 27.994 ;
               RECT 12.494 29.158 12.546 29.194 ;
               RECT 12.494 30.358 12.546 30.394 ;
               RECT 12.494 31.558 12.546 31.594 ;
               RECT 12.494 32.758 12.546 32.794 ;
               RECT 12.494 33.958 12.546 33.994 ;
               RECT 12.494 35.158 12.546 35.194 ;
               RECT 12.494 36.358 12.546 36.394 ;
               RECT 12.494 37.558 12.546 37.594 ;
               RECT 12.494 38.758 12.546 38.794 ;
               RECT 12.494 39.958 12.546 39.994 ;
               RECT 12.494 41.158 12.546 41.194 ;
               RECT 12.494 42.358 12.546 42.394 ;
               RECT 12.494 43.558 12.546 43.594 ;
               RECT 12.494 44.758 12.546 44.794 ;
               RECT 12.494 45.958 12.546 45.994 ;
               RECT 12.494 47.158 12.546 47.194 ;
               RECT 12.494 48.358 12.546 48.394 ;
               RECT 12.494 50.142 12.546 50.178 ;
               RECT 12.494 50.382 12.546 50.418 ;
               RECT 12.494 54.702 12.546 54.738 ;
               RECT 12.494 54.942 12.546 54.978 ;
               RECT 12.494 57.478 12.546 57.514 ;
               RECT 12.494 58.678 12.546 58.714 ;
               RECT 12.494 59.878 12.546 59.914 ;
               RECT 12.494 61.078 12.546 61.114 ;
               RECT 12.494 62.278 12.546 62.314 ;
               RECT 12.494 63.478 12.546 63.514 ;
               RECT 12.494 64.678 12.546 64.714 ;
               RECT 12.494 65.878 12.546 65.914 ;
               RECT 12.494 67.078 12.546 67.114 ;
               RECT 12.494 68.278 12.546 68.314 ;
               RECT 12.494 69.478 12.546 69.514 ;
               RECT 12.494 70.678 12.546 70.714 ;
               RECT 12.494 71.878 12.546 71.914 ;
               RECT 12.494 73.078 12.546 73.114 ;
               RECT 12.494 74.278 12.546 74.314 ;
               RECT 12.494 75.478 12.546 75.514 ;
               RECT 12.494 76.678 12.546 76.714 ;
               RECT 12.494 77.878 12.546 77.914 ;
               RECT 12.494 79.078 12.546 79.114 ;
               RECT 12.494 80.278 12.546 80.314 ;
               RECT 12.494 81.478 12.546 81.514 ;
               RECT 12.494 82.678 12.546 82.714 ;
               RECT 12.494 83.878 12.546 83.914 ;
               RECT 12.494 85.078 12.546 85.114 ;
               RECT 12.494 86.278 12.546 86.314 ;
               RECT 12.494 87.478 12.546 87.514 ;
               RECT 12.494 88.678 12.546 88.714 ;
               RECT 12.494 89.878 12.546 89.914 ;
               RECT 12.494 91.078 12.546 91.114 ;
               RECT 12.494 92.278 12.546 92.314 ;
               RECT 12.494 93.478 12.546 93.514 ;
               RECT 12.494 94.678 12.546 94.714 ;
               RECT 12.494 95.878 12.546 95.914 ;
               RECT 12.494 97.078 12.546 97.114 ;
               RECT 12.494 98.278 12.546 98.314 ;
               RECT 12.494 99.478 12.546 99.514 ;
               RECT 12.494 100.678 12.546 100.714 ;
               RECT 12.494 101.878 12.546 101.914 ;
               RECT 12.494 103.078 12.546 103.114 ;
               RECT 12.494 104.278 12.546 104.314 ;
               RECT 12.574 0.281 12.626 0.317 ;
               RECT 12.574 104.803 12.626 104.839 ;
               RECT 12.654 0.806 12.706 0.842 ;
               RECT 12.654 2.006 12.706 2.042 ;
               RECT 12.654 3.206 12.706 3.242 ;
               RECT 12.654 4.406 12.706 4.442 ;
               RECT 12.654 5.606 12.706 5.642 ;
               RECT 12.654 6.806 12.706 6.842 ;
               RECT 12.654 8.006 12.706 8.042 ;
               RECT 12.654 9.206 12.706 9.242 ;
               RECT 12.654 10.406 12.706 10.442 ;
               RECT 12.654 11.606 12.706 11.642 ;
               RECT 12.654 12.806 12.706 12.842 ;
               RECT 12.654 14.006 12.706 14.042 ;
               RECT 12.654 15.206 12.706 15.242 ;
               RECT 12.654 16.406 12.706 16.442 ;
               RECT 12.654 17.606 12.706 17.642 ;
               RECT 12.654 18.806 12.706 18.842 ;
               RECT 12.654 20.006 12.706 20.042 ;
               RECT 12.654 21.206 12.706 21.242 ;
               RECT 12.654 22.406 12.706 22.442 ;
               RECT 12.654 23.606 12.706 23.642 ;
               RECT 12.654 24.806 12.706 24.842 ;
               RECT 12.654 26.006 12.706 26.042 ;
               RECT 12.654 27.206 12.706 27.242 ;
               RECT 12.654 28.406 12.706 28.442 ;
               RECT 12.654 29.606 12.706 29.642 ;
               RECT 12.654 30.806 12.706 30.842 ;
               RECT 12.654 32.006 12.706 32.042 ;
               RECT 12.654 33.206 12.706 33.242 ;
               RECT 12.654 34.406 12.706 34.442 ;
               RECT 12.654 35.606 12.706 35.642 ;
               RECT 12.654 36.806 12.706 36.842 ;
               RECT 12.654 38.006 12.706 38.042 ;
               RECT 12.654 39.206 12.706 39.242 ;
               RECT 12.654 40.406 12.706 40.442 ;
               RECT 12.654 41.606 12.706 41.642 ;
               RECT 12.654 42.806 12.706 42.842 ;
               RECT 12.654 44.006 12.706 44.042 ;
               RECT 12.654 45.206 12.706 45.242 ;
               RECT 12.654 46.406 12.706 46.442 ;
               RECT 12.654 47.606 12.706 47.642 ;
               RECT 12.654 49.422 12.706 49.458 ;
               RECT 12.654 49.662 12.706 49.698 ;
               RECT 12.654 55.422 12.706 55.458 ;
               RECT 12.654 55.662 12.706 55.698 ;
               RECT 12.654 56.726 12.706 56.762 ;
               RECT 12.654 57.926 12.706 57.962 ;
               RECT 12.654 59.126 12.706 59.162 ;
               RECT 12.654 60.326 12.706 60.362 ;
               RECT 12.654 61.526 12.706 61.562 ;
               RECT 12.654 62.726 12.706 62.762 ;
               RECT 12.654 63.926 12.706 63.962 ;
               RECT 12.654 65.126 12.706 65.162 ;
               RECT 12.654 66.326 12.706 66.362 ;
               RECT 12.654 67.526 12.706 67.562 ;
               RECT 12.654 68.726 12.706 68.762 ;
               RECT 12.654 69.926 12.706 69.962 ;
               RECT 12.654 71.126 12.706 71.162 ;
               RECT 12.654 72.326 12.706 72.362 ;
               RECT 12.654 73.526 12.706 73.562 ;
               RECT 12.654 74.726 12.706 74.762 ;
               RECT 12.654 75.926 12.706 75.962 ;
               RECT 12.654 77.126 12.706 77.162 ;
               RECT 12.654 78.326 12.706 78.362 ;
               RECT 12.654 79.526 12.706 79.562 ;
               RECT 12.654 80.726 12.706 80.762 ;
               RECT 12.654 81.926 12.706 81.962 ;
               RECT 12.654 83.126 12.706 83.162 ;
               RECT 12.654 84.326 12.706 84.362 ;
               RECT 12.654 85.526 12.706 85.562 ;
               RECT 12.654 86.726 12.706 86.762 ;
               RECT 12.654 87.926 12.706 87.962 ;
               RECT 12.654 89.126 12.706 89.162 ;
               RECT 12.654 90.326 12.706 90.362 ;
               RECT 12.654 91.526 12.706 91.562 ;
               RECT 12.654 92.726 12.706 92.762 ;
               RECT 12.654 93.926 12.706 93.962 ;
               RECT 12.654 95.126 12.706 95.162 ;
               RECT 12.654 96.326 12.706 96.362 ;
               RECT 12.654 97.526 12.706 97.562 ;
               RECT 12.654 98.726 12.706 98.762 ;
               RECT 12.654 99.926 12.706 99.962 ;
               RECT 12.654 101.126 12.706 101.162 ;
               RECT 12.654 102.326 12.706 102.362 ;
               RECT 12.654 103.526 12.706 103.562 ;
               RECT 12.734 1.558 12.786 1.594 ;
               RECT 12.734 2.758 12.786 2.794 ;
               RECT 12.734 3.958 12.786 3.994 ;
               RECT 12.734 5.158 12.786 5.194 ;
               RECT 12.734 6.358 12.786 6.394 ;
               RECT 12.734 7.558 12.786 7.594 ;
               RECT 12.734 8.758 12.786 8.794 ;
               RECT 12.734 9.958 12.786 9.994 ;
               RECT 12.734 11.158 12.786 11.194 ;
               RECT 12.734 12.358 12.786 12.394 ;
               RECT 12.734 13.558 12.786 13.594 ;
               RECT 12.734 14.758 12.786 14.794 ;
               RECT 12.734 15.958 12.786 15.994 ;
               RECT 12.734 17.158 12.786 17.194 ;
               RECT 12.734 18.358 12.786 18.394 ;
               RECT 12.734 19.558 12.786 19.594 ;
               RECT 12.734 20.758 12.786 20.794 ;
               RECT 12.734 21.958 12.786 21.994 ;
               RECT 12.734 23.158 12.786 23.194 ;
               RECT 12.734 24.358 12.786 24.394 ;
               RECT 12.734 25.558 12.786 25.594 ;
               RECT 12.734 26.758 12.786 26.794 ;
               RECT 12.734 27.958 12.786 27.994 ;
               RECT 12.734 29.158 12.786 29.194 ;
               RECT 12.734 30.358 12.786 30.394 ;
               RECT 12.734 31.558 12.786 31.594 ;
               RECT 12.734 32.758 12.786 32.794 ;
               RECT 12.734 33.958 12.786 33.994 ;
               RECT 12.734 35.158 12.786 35.194 ;
               RECT 12.734 36.358 12.786 36.394 ;
               RECT 12.734 37.558 12.786 37.594 ;
               RECT 12.734 38.758 12.786 38.794 ;
               RECT 12.734 39.958 12.786 39.994 ;
               RECT 12.734 41.158 12.786 41.194 ;
               RECT 12.734 42.358 12.786 42.394 ;
               RECT 12.734 43.558 12.786 43.594 ;
               RECT 12.734 44.758 12.786 44.794 ;
               RECT 12.734 45.958 12.786 45.994 ;
               RECT 12.734 47.158 12.786 47.194 ;
               RECT 12.734 48.358 12.786 48.394 ;
               RECT 12.734 50.142 12.786 50.178 ;
               RECT 12.734 50.382 12.786 50.418 ;
               RECT 12.734 54.702 12.786 54.738 ;
               RECT 12.734 54.942 12.786 54.978 ;
               RECT 12.734 57.478 12.786 57.514 ;
               RECT 12.734 58.678 12.786 58.714 ;
               RECT 12.734 59.878 12.786 59.914 ;
               RECT 12.734 61.078 12.786 61.114 ;
               RECT 12.734 62.278 12.786 62.314 ;
               RECT 12.734 63.478 12.786 63.514 ;
               RECT 12.734 64.678 12.786 64.714 ;
               RECT 12.734 65.878 12.786 65.914 ;
               RECT 12.734 67.078 12.786 67.114 ;
               RECT 12.734 68.278 12.786 68.314 ;
               RECT 12.734 69.478 12.786 69.514 ;
               RECT 12.734 70.678 12.786 70.714 ;
               RECT 12.734 71.878 12.786 71.914 ;
               RECT 12.734 73.078 12.786 73.114 ;
               RECT 12.734 74.278 12.786 74.314 ;
               RECT 12.734 75.478 12.786 75.514 ;
               RECT 12.734 76.678 12.786 76.714 ;
               RECT 12.734 77.878 12.786 77.914 ;
               RECT 12.734 79.078 12.786 79.114 ;
               RECT 12.734 80.278 12.786 80.314 ;
               RECT 12.734 81.478 12.786 81.514 ;
               RECT 12.734 82.678 12.786 82.714 ;
               RECT 12.734 83.878 12.786 83.914 ;
               RECT 12.734 85.078 12.786 85.114 ;
               RECT 12.734 86.278 12.786 86.314 ;
               RECT 12.734 87.478 12.786 87.514 ;
               RECT 12.734 88.678 12.786 88.714 ;
               RECT 12.734 89.878 12.786 89.914 ;
               RECT 12.734 91.078 12.786 91.114 ;
               RECT 12.734 92.278 12.786 92.314 ;
               RECT 12.734 93.478 12.786 93.514 ;
               RECT 12.734 94.678 12.786 94.714 ;
               RECT 12.734 95.878 12.786 95.914 ;
               RECT 12.734 97.078 12.786 97.114 ;
               RECT 12.734 98.278 12.786 98.314 ;
               RECT 12.734 99.478 12.786 99.514 ;
               RECT 12.734 100.678 12.786 100.714 ;
               RECT 12.734 101.878 12.786 101.914 ;
               RECT 12.734 103.078 12.786 103.114 ;
               RECT 12.734 104.278 12.786 104.314 ;
               RECT 12.814 0.806 12.866 0.842 ;
               RECT 12.814 2.006 12.866 2.042 ;
               RECT 12.814 3.206 12.866 3.242 ;
               RECT 12.814 4.406 12.866 4.442 ;
               RECT 12.814 5.606 12.866 5.642 ;
               RECT 12.814 6.806 12.866 6.842 ;
               RECT 12.814 8.006 12.866 8.042 ;
               RECT 12.814 9.206 12.866 9.242 ;
               RECT 12.814 10.406 12.866 10.442 ;
               RECT 12.814 11.606 12.866 11.642 ;
               RECT 12.814 12.806 12.866 12.842 ;
               RECT 12.814 14.006 12.866 14.042 ;
               RECT 12.814 15.206 12.866 15.242 ;
               RECT 12.814 16.406 12.866 16.442 ;
               RECT 12.814 17.606 12.866 17.642 ;
               RECT 12.814 18.806 12.866 18.842 ;
               RECT 12.814 20.006 12.866 20.042 ;
               RECT 12.814 21.206 12.866 21.242 ;
               RECT 12.814 22.406 12.866 22.442 ;
               RECT 12.814 23.606 12.866 23.642 ;
               RECT 12.814 24.806 12.866 24.842 ;
               RECT 12.814 26.006 12.866 26.042 ;
               RECT 12.814 27.206 12.866 27.242 ;
               RECT 12.814 28.406 12.866 28.442 ;
               RECT 12.814 29.606 12.866 29.642 ;
               RECT 12.814 30.806 12.866 30.842 ;
               RECT 12.814 32.006 12.866 32.042 ;
               RECT 12.814 33.206 12.866 33.242 ;
               RECT 12.814 34.406 12.866 34.442 ;
               RECT 12.814 35.606 12.866 35.642 ;
               RECT 12.814 36.806 12.866 36.842 ;
               RECT 12.814 38.006 12.866 38.042 ;
               RECT 12.814 39.206 12.866 39.242 ;
               RECT 12.814 40.406 12.866 40.442 ;
               RECT 12.814 41.606 12.866 41.642 ;
               RECT 12.814 42.806 12.866 42.842 ;
               RECT 12.814 44.006 12.866 44.042 ;
               RECT 12.814 45.206 12.866 45.242 ;
               RECT 12.814 46.406 12.866 46.442 ;
               RECT 12.814 47.606 12.866 47.642 ;
               RECT 12.814 49.422 12.866 49.458 ;
               RECT 12.814 49.662 12.866 49.698 ;
               RECT 12.814 55.422 12.866 55.458 ;
               RECT 12.814 55.662 12.866 55.698 ;
               RECT 12.814 56.726 12.866 56.762 ;
               RECT 12.814 57.926 12.866 57.962 ;
               RECT 12.814 59.126 12.866 59.162 ;
               RECT 12.814 60.326 12.866 60.362 ;
               RECT 12.814 61.526 12.866 61.562 ;
               RECT 12.814 62.726 12.866 62.762 ;
               RECT 12.814 63.926 12.866 63.962 ;
               RECT 12.814 65.126 12.866 65.162 ;
               RECT 12.814 66.326 12.866 66.362 ;
               RECT 12.814 67.526 12.866 67.562 ;
               RECT 12.814 68.726 12.866 68.762 ;
               RECT 12.814 69.926 12.866 69.962 ;
               RECT 12.814 71.126 12.866 71.162 ;
               RECT 12.814 72.326 12.866 72.362 ;
               RECT 12.814 73.526 12.866 73.562 ;
               RECT 12.814 74.726 12.866 74.762 ;
               RECT 12.814 75.926 12.866 75.962 ;
               RECT 12.814 77.126 12.866 77.162 ;
               RECT 12.814 78.326 12.866 78.362 ;
               RECT 12.814 79.526 12.866 79.562 ;
               RECT 12.814 80.726 12.866 80.762 ;
               RECT 12.814 81.926 12.866 81.962 ;
               RECT 12.814 83.126 12.866 83.162 ;
               RECT 12.814 84.326 12.866 84.362 ;
               RECT 12.814 85.526 12.866 85.562 ;
               RECT 12.814 86.726 12.866 86.762 ;
               RECT 12.814 87.926 12.866 87.962 ;
               RECT 12.814 89.126 12.866 89.162 ;
               RECT 12.814 90.326 12.866 90.362 ;
               RECT 12.814 91.526 12.866 91.562 ;
               RECT 12.814 92.726 12.866 92.762 ;
               RECT 12.814 93.926 12.866 93.962 ;
               RECT 12.814 95.126 12.866 95.162 ;
               RECT 12.814 96.326 12.866 96.362 ;
               RECT 12.814 97.526 12.866 97.562 ;
               RECT 12.814 98.726 12.866 98.762 ;
               RECT 12.814 99.926 12.866 99.962 ;
               RECT 12.814 101.126 12.866 101.162 ;
               RECT 12.814 102.326 12.866 102.362 ;
               RECT 12.814 103.526 12.866 103.562 ;
               RECT 12.894 1.558 12.946 1.594 ;
               RECT 12.894 2.758 12.946 2.794 ;
               RECT 12.894 3.958 12.946 3.994 ;
               RECT 12.894 5.158 12.946 5.194 ;
               RECT 12.894 6.358 12.946 6.394 ;
               RECT 12.894 7.558 12.946 7.594 ;
               RECT 12.894 8.758 12.946 8.794 ;
               RECT 12.894 9.958 12.946 9.994 ;
               RECT 12.894 11.158 12.946 11.194 ;
               RECT 12.894 12.358 12.946 12.394 ;
               RECT 12.894 13.558 12.946 13.594 ;
               RECT 12.894 14.758 12.946 14.794 ;
               RECT 12.894 15.958 12.946 15.994 ;
               RECT 12.894 17.158 12.946 17.194 ;
               RECT 12.894 18.358 12.946 18.394 ;
               RECT 12.894 19.558 12.946 19.594 ;
               RECT 12.894 20.758 12.946 20.794 ;
               RECT 12.894 21.958 12.946 21.994 ;
               RECT 12.894 23.158 12.946 23.194 ;
               RECT 12.894 24.358 12.946 24.394 ;
               RECT 12.894 25.558 12.946 25.594 ;
               RECT 12.894 26.758 12.946 26.794 ;
               RECT 12.894 27.958 12.946 27.994 ;
               RECT 12.894 29.158 12.946 29.194 ;
               RECT 12.894 30.358 12.946 30.394 ;
               RECT 12.894 31.558 12.946 31.594 ;
               RECT 12.894 32.758 12.946 32.794 ;
               RECT 12.894 33.958 12.946 33.994 ;
               RECT 12.894 35.158 12.946 35.194 ;
               RECT 12.894 36.358 12.946 36.394 ;
               RECT 12.894 37.558 12.946 37.594 ;
               RECT 12.894 38.758 12.946 38.794 ;
               RECT 12.894 39.958 12.946 39.994 ;
               RECT 12.894 41.158 12.946 41.194 ;
               RECT 12.894 42.358 12.946 42.394 ;
               RECT 12.894 43.558 12.946 43.594 ;
               RECT 12.894 44.758 12.946 44.794 ;
               RECT 12.894 45.958 12.946 45.994 ;
               RECT 12.894 47.158 12.946 47.194 ;
               RECT 12.894 48.358 12.946 48.394 ;
               RECT 12.894 50.142 12.946 50.178 ;
               RECT 12.894 50.382 12.946 50.418 ;
               RECT 12.894 54.702 12.946 54.738 ;
               RECT 12.894 54.942 12.946 54.978 ;
               RECT 12.894 57.478 12.946 57.514 ;
               RECT 12.894 58.678 12.946 58.714 ;
               RECT 12.894 59.878 12.946 59.914 ;
               RECT 12.894 61.078 12.946 61.114 ;
               RECT 12.894 62.278 12.946 62.314 ;
               RECT 12.894 63.478 12.946 63.514 ;
               RECT 12.894 64.678 12.946 64.714 ;
               RECT 12.894 65.878 12.946 65.914 ;
               RECT 12.894 67.078 12.946 67.114 ;
               RECT 12.894 68.278 12.946 68.314 ;
               RECT 12.894 69.478 12.946 69.514 ;
               RECT 12.894 70.678 12.946 70.714 ;
               RECT 12.894 71.878 12.946 71.914 ;
               RECT 12.894 73.078 12.946 73.114 ;
               RECT 12.894 74.278 12.946 74.314 ;
               RECT 12.894 75.478 12.946 75.514 ;
               RECT 12.894 76.678 12.946 76.714 ;
               RECT 12.894 77.878 12.946 77.914 ;
               RECT 12.894 79.078 12.946 79.114 ;
               RECT 12.894 80.278 12.946 80.314 ;
               RECT 12.894 81.478 12.946 81.514 ;
               RECT 12.894 82.678 12.946 82.714 ;
               RECT 12.894 83.878 12.946 83.914 ;
               RECT 12.894 85.078 12.946 85.114 ;
               RECT 12.894 86.278 12.946 86.314 ;
               RECT 12.894 87.478 12.946 87.514 ;
               RECT 12.894 88.678 12.946 88.714 ;
               RECT 12.894 89.878 12.946 89.914 ;
               RECT 12.894 91.078 12.946 91.114 ;
               RECT 12.894 92.278 12.946 92.314 ;
               RECT 12.894 93.478 12.946 93.514 ;
               RECT 12.894 94.678 12.946 94.714 ;
               RECT 12.894 95.878 12.946 95.914 ;
               RECT 12.894 97.078 12.946 97.114 ;
               RECT 12.894 98.278 12.946 98.314 ;
               RECT 12.894 99.478 12.946 99.514 ;
               RECT 12.894 100.678 12.946 100.714 ;
               RECT 12.894 101.878 12.946 101.914 ;
               RECT 12.894 103.078 12.946 103.114 ;
               RECT 12.894 104.278 12.946 104.314 ;
               RECT 12.974 0.281 13.026 0.317 ;
               RECT 12.974 104.803 13.026 104.839 ;
               RECT 13.054 0.806 13.106 0.842 ;
               RECT 13.054 2.006 13.106 2.042 ;
               RECT 13.054 3.206 13.106 3.242 ;
               RECT 13.054 4.406 13.106 4.442 ;
               RECT 13.054 5.606 13.106 5.642 ;
               RECT 13.054 6.806 13.106 6.842 ;
               RECT 13.054 8.006 13.106 8.042 ;
               RECT 13.054 9.206 13.106 9.242 ;
               RECT 13.054 10.406 13.106 10.442 ;
               RECT 13.054 11.606 13.106 11.642 ;
               RECT 13.054 12.806 13.106 12.842 ;
               RECT 13.054 14.006 13.106 14.042 ;
               RECT 13.054 15.206 13.106 15.242 ;
               RECT 13.054 16.406 13.106 16.442 ;
               RECT 13.054 17.606 13.106 17.642 ;
               RECT 13.054 18.806 13.106 18.842 ;
               RECT 13.054 20.006 13.106 20.042 ;
               RECT 13.054 21.206 13.106 21.242 ;
               RECT 13.054 22.406 13.106 22.442 ;
               RECT 13.054 23.606 13.106 23.642 ;
               RECT 13.054 24.806 13.106 24.842 ;
               RECT 13.054 26.006 13.106 26.042 ;
               RECT 13.054 27.206 13.106 27.242 ;
               RECT 13.054 28.406 13.106 28.442 ;
               RECT 13.054 29.606 13.106 29.642 ;
               RECT 13.054 30.806 13.106 30.842 ;
               RECT 13.054 32.006 13.106 32.042 ;
               RECT 13.054 33.206 13.106 33.242 ;
               RECT 13.054 34.406 13.106 34.442 ;
               RECT 13.054 35.606 13.106 35.642 ;
               RECT 13.054 36.806 13.106 36.842 ;
               RECT 13.054 38.006 13.106 38.042 ;
               RECT 13.054 39.206 13.106 39.242 ;
               RECT 13.054 40.406 13.106 40.442 ;
               RECT 13.054 41.606 13.106 41.642 ;
               RECT 13.054 42.806 13.106 42.842 ;
               RECT 13.054 44.006 13.106 44.042 ;
               RECT 13.054 45.206 13.106 45.242 ;
               RECT 13.054 46.406 13.106 46.442 ;
               RECT 13.054 47.606 13.106 47.642 ;
               RECT 13.054 49.422 13.106 49.458 ;
               RECT 13.054 49.662 13.106 49.698 ;
               RECT 13.054 51.102 13.106 51.138 ;
               RECT 13.054 51.582 13.106 51.618 ;
               RECT 13.054 53.502 13.106 53.538 ;
               RECT 13.054 53.982 13.106 54.018 ;
               RECT 13.054 55.422 13.106 55.458 ;
               RECT 13.054 55.662 13.106 55.698 ;
               RECT 13.054 56.726 13.106 56.762 ;
               RECT 13.054 57.926 13.106 57.962 ;
               RECT 13.054 59.126 13.106 59.162 ;
               RECT 13.054 60.326 13.106 60.362 ;
               RECT 13.054 61.526 13.106 61.562 ;
               RECT 13.054 62.726 13.106 62.762 ;
               RECT 13.054 63.926 13.106 63.962 ;
               RECT 13.054 65.126 13.106 65.162 ;
               RECT 13.054 66.326 13.106 66.362 ;
               RECT 13.054 67.526 13.106 67.562 ;
               RECT 13.054 68.726 13.106 68.762 ;
               RECT 13.054 69.926 13.106 69.962 ;
               RECT 13.054 71.126 13.106 71.162 ;
               RECT 13.054 72.326 13.106 72.362 ;
               RECT 13.054 73.526 13.106 73.562 ;
               RECT 13.054 74.726 13.106 74.762 ;
               RECT 13.054 75.926 13.106 75.962 ;
               RECT 13.054 77.126 13.106 77.162 ;
               RECT 13.054 78.326 13.106 78.362 ;
               RECT 13.054 79.526 13.106 79.562 ;
               RECT 13.054 80.726 13.106 80.762 ;
               RECT 13.054 81.926 13.106 81.962 ;
               RECT 13.054 83.126 13.106 83.162 ;
               RECT 13.054 84.326 13.106 84.362 ;
               RECT 13.054 85.526 13.106 85.562 ;
               RECT 13.054 86.726 13.106 86.762 ;
               RECT 13.054 87.926 13.106 87.962 ;
               RECT 13.054 89.126 13.106 89.162 ;
               RECT 13.054 90.326 13.106 90.362 ;
               RECT 13.054 91.526 13.106 91.562 ;
               RECT 13.054 92.726 13.106 92.762 ;
               RECT 13.054 93.926 13.106 93.962 ;
               RECT 13.054 95.126 13.106 95.162 ;
               RECT 13.054 96.326 13.106 96.362 ;
               RECT 13.054 97.526 13.106 97.562 ;
               RECT 13.054 98.726 13.106 98.762 ;
               RECT 13.054 99.926 13.106 99.962 ;
               RECT 13.054 101.126 13.106 101.162 ;
               RECT 13.054 102.326 13.106 102.362 ;
               RECT 13.054 103.526 13.106 103.562 ;
               RECT 13.134 1.558 13.186 1.594 ;
               RECT 13.134 2.758 13.186 2.794 ;
               RECT 13.134 3.958 13.186 3.994 ;
               RECT 13.134 5.158 13.186 5.194 ;
               RECT 13.134 6.358 13.186 6.394 ;
               RECT 13.134 7.558 13.186 7.594 ;
               RECT 13.134 8.758 13.186 8.794 ;
               RECT 13.134 9.958 13.186 9.994 ;
               RECT 13.134 11.158 13.186 11.194 ;
               RECT 13.134 12.358 13.186 12.394 ;
               RECT 13.134 13.558 13.186 13.594 ;
               RECT 13.134 14.758 13.186 14.794 ;
               RECT 13.134 15.958 13.186 15.994 ;
               RECT 13.134 17.158 13.186 17.194 ;
               RECT 13.134 18.358 13.186 18.394 ;
               RECT 13.134 19.558 13.186 19.594 ;
               RECT 13.134 20.758 13.186 20.794 ;
               RECT 13.134 21.958 13.186 21.994 ;
               RECT 13.134 23.158 13.186 23.194 ;
               RECT 13.134 24.358 13.186 24.394 ;
               RECT 13.134 25.558 13.186 25.594 ;
               RECT 13.134 26.758 13.186 26.794 ;
               RECT 13.134 27.958 13.186 27.994 ;
               RECT 13.134 29.158 13.186 29.194 ;
               RECT 13.134 30.358 13.186 30.394 ;
               RECT 13.134 31.558 13.186 31.594 ;
               RECT 13.134 32.758 13.186 32.794 ;
               RECT 13.134 33.958 13.186 33.994 ;
               RECT 13.134 35.158 13.186 35.194 ;
               RECT 13.134 36.358 13.186 36.394 ;
               RECT 13.134 37.558 13.186 37.594 ;
               RECT 13.134 38.758 13.186 38.794 ;
               RECT 13.134 39.958 13.186 39.994 ;
               RECT 13.134 41.158 13.186 41.194 ;
               RECT 13.134 42.358 13.186 42.394 ;
               RECT 13.134 43.558 13.186 43.594 ;
               RECT 13.134 44.758 13.186 44.794 ;
               RECT 13.134 45.958 13.186 45.994 ;
               RECT 13.134 47.158 13.186 47.194 ;
               RECT 13.134 48.358 13.186 48.394 ;
               RECT 13.134 50.142 13.186 50.178 ;
               RECT 13.134 50.382 13.186 50.418 ;
               RECT 13.134 54.702 13.186 54.738 ;
               RECT 13.134 54.942 13.186 54.978 ;
               RECT 13.134 57.478 13.186 57.514 ;
               RECT 13.134 58.678 13.186 58.714 ;
               RECT 13.134 59.878 13.186 59.914 ;
               RECT 13.134 61.078 13.186 61.114 ;
               RECT 13.134 62.278 13.186 62.314 ;
               RECT 13.134 63.478 13.186 63.514 ;
               RECT 13.134 64.678 13.186 64.714 ;
               RECT 13.134 65.878 13.186 65.914 ;
               RECT 13.134 67.078 13.186 67.114 ;
               RECT 13.134 68.278 13.186 68.314 ;
               RECT 13.134 69.478 13.186 69.514 ;
               RECT 13.134 70.678 13.186 70.714 ;
               RECT 13.134 71.878 13.186 71.914 ;
               RECT 13.134 73.078 13.186 73.114 ;
               RECT 13.134 74.278 13.186 74.314 ;
               RECT 13.134 75.478 13.186 75.514 ;
               RECT 13.134 76.678 13.186 76.714 ;
               RECT 13.134 77.878 13.186 77.914 ;
               RECT 13.134 79.078 13.186 79.114 ;
               RECT 13.134 80.278 13.186 80.314 ;
               RECT 13.134 81.478 13.186 81.514 ;
               RECT 13.134 82.678 13.186 82.714 ;
               RECT 13.134 83.878 13.186 83.914 ;
               RECT 13.134 85.078 13.186 85.114 ;
               RECT 13.134 86.278 13.186 86.314 ;
               RECT 13.134 87.478 13.186 87.514 ;
               RECT 13.134 88.678 13.186 88.714 ;
               RECT 13.134 89.878 13.186 89.914 ;
               RECT 13.134 91.078 13.186 91.114 ;
               RECT 13.134 92.278 13.186 92.314 ;
               RECT 13.134 93.478 13.186 93.514 ;
               RECT 13.134 94.678 13.186 94.714 ;
               RECT 13.134 95.878 13.186 95.914 ;
               RECT 13.134 97.078 13.186 97.114 ;
               RECT 13.134 98.278 13.186 98.314 ;
               RECT 13.134 99.478 13.186 99.514 ;
               RECT 13.134 100.678 13.186 100.714 ;
               RECT 13.134 101.878 13.186 101.914 ;
               RECT 13.134 103.078 13.186 103.114 ;
               RECT 13.134 104.278 13.186 104.314 ;
               RECT 13.214 0.806 13.266 0.842 ;
               RECT 13.214 2.006 13.266 2.042 ;
               RECT 13.214 3.206 13.266 3.242 ;
               RECT 13.214 4.406 13.266 4.442 ;
               RECT 13.214 5.606 13.266 5.642 ;
               RECT 13.214 6.806 13.266 6.842 ;
               RECT 13.214 8.006 13.266 8.042 ;
               RECT 13.214 9.206 13.266 9.242 ;
               RECT 13.214 10.406 13.266 10.442 ;
               RECT 13.214 11.606 13.266 11.642 ;
               RECT 13.214 12.806 13.266 12.842 ;
               RECT 13.214 14.006 13.266 14.042 ;
               RECT 13.214 15.206 13.266 15.242 ;
               RECT 13.214 16.406 13.266 16.442 ;
               RECT 13.214 17.606 13.266 17.642 ;
               RECT 13.214 18.806 13.266 18.842 ;
               RECT 13.214 20.006 13.266 20.042 ;
               RECT 13.214 21.206 13.266 21.242 ;
               RECT 13.214 22.406 13.266 22.442 ;
               RECT 13.214 23.606 13.266 23.642 ;
               RECT 13.214 24.806 13.266 24.842 ;
               RECT 13.214 26.006 13.266 26.042 ;
               RECT 13.214 27.206 13.266 27.242 ;
               RECT 13.214 28.406 13.266 28.442 ;
               RECT 13.214 29.606 13.266 29.642 ;
               RECT 13.214 30.806 13.266 30.842 ;
               RECT 13.214 32.006 13.266 32.042 ;
               RECT 13.214 33.206 13.266 33.242 ;
               RECT 13.214 34.406 13.266 34.442 ;
               RECT 13.214 35.606 13.266 35.642 ;
               RECT 13.214 36.806 13.266 36.842 ;
               RECT 13.214 38.006 13.266 38.042 ;
               RECT 13.214 39.206 13.266 39.242 ;
               RECT 13.214 40.406 13.266 40.442 ;
               RECT 13.214 41.606 13.266 41.642 ;
               RECT 13.214 42.806 13.266 42.842 ;
               RECT 13.214 44.006 13.266 44.042 ;
               RECT 13.214 45.206 13.266 45.242 ;
               RECT 13.214 46.406 13.266 46.442 ;
               RECT 13.214 47.606 13.266 47.642 ;
               RECT 13.214 49.422 13.266 49.458 ;
               RECT 13.214 49.662 13.266 49.698 ;
               RECT 13.214 55.422 13.266 55.458 ;
               RECT 13.214 55.662 13.266 55.698 ;
               RECT 13.214 56.726 13.266 56.762 ;
               RECT 13.214 57.926 13.266 57.962 ;
               RECT 13.214 59.126 13.266 59.162 ;
               RECT 13.214 60.326 13.266 60.362 ;
               RECT 13.214 61.526 13.266 61.562 ;
               RECT 13.214 62.726 13.266 62.762 ;
               RECT 13.214 63.926 13.266 63.962 ;
               RECT 13.214 65.126 13.266 65.162 ;
               RECT 13.214 66.326 13.266 66.362 ;
               RECT 13.214 67.526 13.266 67.562 ;
               RECT 13.214 68.726 13.266 68.762 ;
               RECT 13.214 69.926 13.266 69.962 ;
               RECT 13.214 71.126 13.266 71.162 ;
               RECT 13.214 72.326 13.266 72.362 ;
               RECT 13.214 73.526 13.266 73.562 ;
               RECT 13.214 74.726 13.266 74.762 ;
               RECT 13.214 75.926 13.266 75.962 ;
               RECT 13.214 77.126 13.266 77.162 ;
               RECT 13.214 78.326 13.266 78.362 ;
               RECT 13.214 79.526 13.266 79.562 ;
               RECT 13.214 80.726 13.266 80.762 ;
               RECT 13.214 81.926 13.266 81.962 ;
               RECT 13.214 83.126 13.266 83.162 ;
               RECT 13.214 84.326 13.266 84.362 ;
               RECT 13.214 85.526 13.266 85.562 ;
               RECT 13.214 86.726 13.266 86.762 ;
               RECT 13.214 87.926 13.266 87.962 ;
               RECT 13.214 89.126 13.266 89.162 ;
               RECT 13.214 90.326 13.266 90.362 ;
               RECT 13.214 91.526 13.266 91.562 ;
               RECT 13.214 92.726 13.266 92.762 ;
               RECT 13.214 93.926 13.266 93.962 ;
               RECT 13.214 95.126 13.266 95.162 ;
               RECT 13.214 96.326 13.266 96.362 ;
               RECT 13.214 97.526 13.266 97.562 ;
               RECT 13.214 98.726 13.266 98.762 ;
               RECT 13.214 99.926 13.266 99.962 ;
               RECT 13.214 101.126 13.266 101.162 ;
               RECT 13.214 102.326 13.266 102.362 ;
               RECT 13.214 103.526 13.266 103.562 ;
               RECT 13.294 1.558 13.346 1.594 ;
               RECT 13.294 2.758 13.346 2.794 ;
               RECT 13.294 3.958 13.346 3.994 ;
               RECT 13.294 5.158 13.346 5.194 ;
               RECT 13.294 6.358 13.346 6.394 ;
               RECT 13.294 7.558 13.346 7.594 ;
               RECT 13.294 8.758 13.346 8.794 ;
               RECT 13.294 9.958 13.346 9.994 ;
               RECT 13.294 11.158 13.346 11.194 ;
               RECT 13.294 12.358 13.346 12.394 ;
               RECT 13.294 13.558 13.346 13.594 ;
               RECT 13.294 14.758 13.346 14.794 ;
               RECT 13.294 15.958 13.346 15.994 ;
               RECT 13.294 17.158 13.346 17.194 ;
               RECT 13.294 18.358 13.346 18.394 ;
               RECT 13.294 19.558 13.346 19.594 ;
               RECT 13.294 20.758 13.346 20.794 ;
               RECT 13.294 21.958 13.346 21.994 ;
               RECT 13.294 23.158 13.346 23.194 ;
               RECT 13.294 24.358 13.346 24.394 ;
               RECT 13.294 25.558 13.346 25.594 ;
               RECT 13.294 26.758 13.346 26.794 ;
               RECT 13.294 27.958 13.346 27.994 ;
               RECT 13.294 29.158 13.346 29.194 ;
               RECT 13.294 30.358 13.346 30.394 ;
               RECT 13.294 31.558 13.346 31.594 ;
               RECT 13.294 32.758 13.346 32.794 ;
               RECT 13.294 33.958 13.346 33.994 ;
               RECT 13.294 35.158 13.346 35.194 ;
               RECT 13.294 36.358 13.346 36.394 ;
               RECT 13.294 37.558 13.346 37.594 ;
               RECT 13.294 38.758 13.346 38.794 ;
               RECT 13.294 39.958 13.346 39.994 ;
               RECT 13.294 41.158 13.346 41.194 ;
               RECT 13.294 42.358 13.346 42.394 ;
               RECT 13.294 43.558 13.346 43.594 ;
               RECT 13.294 44.758 13.346 44.794 ;
               RECT 13.294 45.958 13.346 45.994 ;
               RECT 13.294 47.158 13.346 47.194 ;
               RECT 13.294 48.358 13.346 48.394 ;
               RECT 13.294 50.142 13.346 50.178 ;
               RECT 13.294 50.382 13.346 50.418 ;
               RECT 13.294 54.702 13.346 54.738 ;
               RECT 13.294 54.942 13.346 54.978 ;
               RECT 13.294 57.478 13.346 57.514 ;
               RECT 13.294 58.678 13.346 58.714 ;
               RECT 13.294 59.878 13.346 59.914 ;
               RECT 13.294 61.078 13.346 61.114 ;
               RECT 13.294 62.278 13.346 62.314 ;
               RECT 13.294 63.478 13.346 63.514 ;
               RECT 13.294 64.678 13.346 64.714 ;
               RECT 13.294 65.878 13.346 65.914 ;
               RECT 13.294 67.078 13.346 67.114 ;
               RECT 13.294 68.278 13.346 68.314 ;
               RECT 13.294 69.478 13.346 69.514 ;
               RECT 13.294 70.678 13.346 70.714 ;
               RECT 13.294 71.878 13.346 71.914 ;
               RECT 13.294 73.078 13.346 73.114 ;
               RECT 13.294 74.278 13.346 74.314 ;
               RECT 13.294 75.478 13.346 75.514 ;
               RECT 13.294 76.678 13.346 76.714 ;
               RECT 13.294 77.878 13.346 77.914 ;
               RECT 13.294 79.078 13.346 79.114 ;
               RECT 13.294 80.278 13.346 80.314 ;
               RECT 13.294 81.478 13.346 81.514 ;
               RECT 13.294 82.678 13.346 82.714 ;
               RECT 13.294 83.878 13.346 83.914 ;
               RECT 13.294 85.078 13.346 85.114 ;
               RECT 13.294 86.278 13.346 86.314 ;
               RECT 13.294 87.478 13.346 87.514 ;
               RECT 13.294 88.678 13.346 88.714 ;
               RECT 13.294 89.878 13.346 89.914 ;
               RECT 13.294 91.078 13.346 91.114 ;
               RECT 13.294 92.278 13.346 92.314 ;
               RECT 13.294 93.478 13.346 93.514 ;
               RECT 13.294 94.678 13.346 94.714 ;
               RECT 13.294 95.878 13.346 95.914 ;
               RECT 13.294 97.078 13.346 97.114 ;
               RECT 13.294 98.278 13.346 98.314 ;
               RECT 13.294 99.478 13.346 99.514 ;
               RECT 13.294 100.678 13.346 100.714 ;
               RECT 13.294 101.878 13.346 101.914 ;
               RECT 13.294 103.078 13.346 103.114 ;
               RECT 13.294 104.278 13.346 104.314 ;
               RECT 13.374 0.281 13.426 0.317 ;
               RECT 13.374 104.803 13.426 104.839 ;
               RECT 13.778 49.8435 13.814 49.8795 ;
               RECT 13.778 50.982 13.814 51.018 ;
               RECT 13.778 54.102 13.814 54.138 ;
               RECT 13.778 55.2405 13.814 55.2765 ;
               RECT 13.978 0.582 14.022 0.618 ;
               RECT 13.978 1.182 14.022 1.218 ;
               RECT 13.978 1.782 14.022 1.818 ;
               RECT 13.978 2.382 14.022 2.418 ;
               RECT 13.978 2.982 14.022 3.018 ;
               RECT 13.978 3.582 14.022 3.618 ;
               RECT 13.978 4.182 14.022 4.218 ;
               RECT 13.978 4.782 14.022 4.818 ;
               RECT 13.978 5.382 14.022 5.418 ;
               RECT 13.978 5.982 14.022 6.018 ;
               RECT 13.978 6.582 14.022 6.618 ;
               RECT 13.978 7.182 14.022 7.218 ;
               RECT 13.978 7.782 14.022 7.818 ;
               RECT 13.978 8.382 14.022 8.418 ;
               RECT 13.978 8.982 14.022 9.018 ;
               RECT 13.978 9.582 14.022 9.618 ;
               RECT 13.978 10.182 14.022 10.218 ;
               RECT 13.978 10.782 14.022 10.818 ;
               RECT 13.978 11.382 14.022 11.418 ;
               RECT 13.978 11.982 14.022 12.018 ;
               RECT 13.978 12.582 14.022 12.618 ;
               RECT 13.978 13.182 14.022 13.218 ;
               RECT 13.978 13.782 14.022 13.818 ;
               RECT 13.978 14.382 14.022 14.418 ;
               RECT 13.978 14.982 14.022 15.018 ;
               RECT 13.978 15.582 14.022 15.618 ;
               RECT 13.978 16.182 14.022 16.218 ;
               RECT 13.978 16.782 14.022 16.818 ;
               RECT 13.978 17.382 14.022 17.418 ;
               RECT 13.978 17.982 14.022 18.018 ;
               RECT 13.978 18.582 14.022 18.618 ;
               RECT 13.978 19.182 14.022 19.218 ;
               RECT 13.978 19.782 14.022 19.818 ;
               RECT 13.978 20.382 14.022 20.418 ;
               RECT 13.978 20.982 14.022 21.018 ;
               RECT 13.978 21.582 14.022 21.618 ;
               RECT 13.978 22.182 14.022 22.218 ;
               RECT 13.978 22.782 14.022 22.818 ;
               RECT 13.978 23.382 14.022 23.418 ;
               RECT 13.978 23.982 14.022 24.018 ;
               RECT 13.978 24.582 14.022 24.618 ;
               RECT 13.978 25.182 14.022 25.218 ;
               RECT 13.978 25.782 14.022 25.818 ;
               RECT 13.978 26.382 14.022 26.418 ;
               RECT 13.978 26.982 14.022 27.018 ;
               RECT 13.978 27.582 14.022 27.618 ;
               RECT 13.978 28.182 14.022 28.218 ;
               RECT 13.978 28.782 14.022 28.818 ;
               RECT 13.978 29.382 14.022 29.418 ;
               RECT 13.978 29.982 14.022 30.018 ;
               RECT 13.978 30.582 14.022 30.618 ;
               RECT 13.978 31.182 14.022 31.218 ;
               RECT 13.978 31.782 14.022 31.818 ;
               RECT 13.978 32.382 14.022 32.418 ;
               RECT 13.978 32.982 14.022 33.018 ;
               RECT 13.978 33.582 14.022 33.618 ;
               RECT 13.978 34.182 14.022 34.218 ;
               RECT 13.978 34.782 14.022 34.818 ;
               RECT 13.978 35.382 14.022 35.418 ;
               RECT 13.978 35.982 14.022 36.018 ;
               RECT 13.978 36.582 14.022 36.618 ;
               RECT 13.978 37.182 14.022 37.218 ;
               RECT 13.978 37.782 14.022 37.818 ;
               RECT 13.978 38.382 14.022 38.418 ;
               RECT 13.978 38.982 14.022 39.018 ;
               RECT 13.978 39.582 14.022 39.618 ;
               RECT 13.978 40.182 14.022 40.218 ;
               RECT 13.978 40.782 14.022 40.818 ;
               RECT 13.978 41.382 14.022 41.418 ;
               RECT 13.978 41.982 14.022 42.018 ;
               RECT 13.978 42.582 14.022 42.618 ;
               RECT 13.978 43.182 14.022 43.218 ;
               RECT 13.978 43.782 14.022 43.818 ;
               RECT 13.978 44.382 14.022 44.418 ;
               RECT 13.978 44.982 14.022 45.018 ;
               RECT 13.978 45.582 14.022 45.618 ;
               RECT 13.978 46.182 14.022 46.218 ;
               RECT 13.978 46.782 14.022 46.818 ;
               RECT 13.978 47.382 14.022 47.418 ;
               RECT 13.978 47.982 14.022 48.018 ;
               RECT 13.978 48.582 14.022 48.618 ;
               RECT 13.978 48.942 14.022 48.978 ;
               RECT 13.978 49.422 14.022 49.458 ;
               RECT 13.978 49.902 14.022 49.938 ;
               RECT 13.978 50.382 14.022 50.418 ;
               RECT 13.978 50.862 14.022 50.898 ;
               RECT 13.978 51.342 14.022 51.378 ;
               RECT 13.978 51.822 14.022 51.858 ;
               RECT 13.978 52.302 14.022 52.338 ;
               RECT 13.978 52.782 14.022 52.818 ;
               RECT 13.978 53.262 14.022 53.298 ;
               RECT 13.978 53.742 14.022 53.778 ;
               RECT 13.978 54.222 14.022 54.258 ;
               RECT 13.978 54.702 14.022 54.738 ;
               RECT 13.978 55.182 14.022 55.218 ;
               RECT 13.978 55.662 14.022 55.698 ;
               RECT 13.978 56.142 14.022 56.178 ;
               RECT 13.978 56.502 14.022 56.538 ;
               RECT 13.978 57.102 14.022 57.138 ;
               RECT 13.978 57.702 14.022 57.738 ;
               RECT 13.978 58.302 14.022 58.338 ;
               RECT 13.978 58.902 14.022 58.938 ;
               RECT 13.978 59.502 14.022 59.538 ;
               RECT 13.978 60.102 14.022 60.138 ;
               RECT 13.978 60.702 14.022 60.738 ;
               RECT 13.978 61.302 14.022 61.338 ;
               RECT 13.978 61.902 14.022 61.938 ;
               RECT 13.978 62.502 14.022 62.538 ;
               RECT 13.978 63.102 14.022 63.138 ;
               RECT 13.978 63.702 14.022 63.738 ;
               RECT 13.978 64.302 14.022 64.338 ;
               RECT 13.978 64.902 14.022 64.938 ;
               RECT 13.978 65.502 14.022 65.538 ;
               RECT 13.978 66.102 14.022 66.138 ;
               RECT 13.978 66.702 14.022 66.738 ;
               RECT 13.978 67.302 14.022 67.338 ;
               RECT 13.978 67.902 14.022 67.938 ;
               RECT 13.978 68.502 14.022 68.538 ;
               RECT 13.978 69.102 14.022 69.138 ;
               RECT 13.978 69.702 14.022 69.738 ;
               RECT 13.978 70.302 14.022 70.338 ;
               RECT 13.978 70.902 14.022 70.938 ;
               RECT 13.978 71.502 14.022 71.538 ;
               RECT 13.978 72.102 14.022 72.138 ;
               RECT 13.978 72.702 14.022 72.738 ;
               RECT 13.978 73.302 14.022 73.338 ;
               RECT 13.978 73.902 14.022 73.938 ;
               RECT 13.978 74.502 14.022 74.538 ;
               RECT 13.978 75.102 14.022 75.138 ;
               RECT 13.978 75.702 14.022 75.738 ;
               RECT 13.978 76.302 14.022 76.338 ;
               RECT 13.978 76.902 14.022 76.938 ;
               RECT 13.978 77.502 14.022 77.538 ;
               RECT 13.978 78.102 14.022 78.138 ;
               RECT 13.978 78.702 14.022 78.738 ;
               RECT 13.978 79.302 14.022 79.338 ;
               RECT 13.978 79.902 14.022 79.938 ;
               RECT 13.978 80.502 14.022 80.538 ;
               RECT 13.978 81.102 14.022 81.138 ;
               RECT 13.978 81.702 14.022 81.738 ;
               RECT 13.978 82.302 14.022 82.338 ;
               RECT 13.978 82.902 14.022 82.938 ;
               RECT 13.978 83.502 14.022 83.538 ;
               RECT 13.978 84.102 14.022 84.138 ;
               RECT 13.978 84.702 14.022 84.738 ;
               RECT 13.978 85.302 14.022 85.338 ;
               RECT 13.978 85.902 14.022 85.938 ;
               RECT 13.978 86.502 14.022 86.538 ;
               RECT 13.978 87.102 14.022 87.138 ;
               RECT 13.978 87.702 14.022 87.738 ;
               RECT 13.978 88.302 14.022 88.338 ;
               RECT 13.978 88.902 14.022 88.938 ;
               RECT 13.978 89.502 14.022 89.538 ;
               RECT 13.978 90.102 14.022 90.138 ;
               RECT 13.978 90.702 14.022 90.738 ;
               RECT 13.978 91.302 14.022 91.338 ;
               RECT 13.978 91.902 14.022 91.938 ;
               RECT 13.978 92.502 14.022 92.538 ;
               RECT 13.978 93.102 14.022 93.138 ;
               RECT 13.978 93.702 14.022 93.738 ;
               RECT 13.978 94.302 14.022 94.338 ;
               RECT 13.978 94.902 14.022 94.938 ;
               RECT 13.978 95.502 14.022 95.538 ;
               RECT 13.978 96.102 14.022 96.138 ;
               RECT 13.978 96.702 14.022 96.738 ;
               RECT 13.978 97.302 14.022 97.338 ;
               RECT 13.978 97.902 14.022 97.938 ;
               RECT 13.978 98.502 14.022 98.538 ;
               RECT 13.978 99.102 14.022 99.138 ;
               RECT 13.978 99.702 14.022 99.738 ;
               RECT 13.978 100.302 14.022 100.338 ;
               RECT 13.978 100.902 14.022 100.938 ;
               RECT 13.978 101.502 14.022 101.538 ;
               RECT 13.978 102.102 14.022 102.138 ;
               RECT 13.978 102.702 14.022 102.738 ;
               RECT 13.978 103.302 14.022 103.338 ;
               RECT 13.978 103.902 14.022 103.938 ;
               RECT 13.978 104.502 14.022 104.538 ;
               RECT 14.132 1.558 14.186 1.594 ;
               RECT 14.132 2.758 14.186 2.794 ;
               RECT 14.132 3.958 14.186 3.994 ;
               RECT 14.132 5.158 14.186 5.194 ;
               RECT 14.132 6.358 14.186 6.394 ;
               RECT 14.132 7.558 14.186 7.594 ;
               RECT 14.132 8.758 14.186 8.794 ;
               RECT 14.132 9.958 14.186 9.994 ;
               RECT 14.132 11.158 14.186 11.194 ;
               RECT 14.132 12.358 14.186 12.394 ;
               RECT 14.132 13.558 14.186 13.594 ;
               RECT 14.132 14.758 14.186 14.794 ;
               RECT 14.132 15.958 14.186 15.994 ;
               RECT 14.132 17.158 14.186 17.194 ;
               RECT 14.132 18.358 14.186 18.394 ;
               RECT 14.132 19.558 14.186 19.594 ;
               RECT 14.132 20.758 14.186 20.794 ;
               RECT 14.132 21.958 14.186 21.994 ;
               RECT 14.132 23.158 14.186 23.194 ;
               RECT 14.132 24.358 14.186 24.394 ;
               RECT 14.132 25.558 14.186 25.594 ;
               RECT 14.132 26.758 14.186 26.794 ;
               RECT 14.132 27.958 14.186 27.994 ;
               RECT 14.132 29.158 14.186 29.194 ;
               RECT 14.132 30.358 14.186 30.394 ;
               RECT 14.132 31.558 14.186 31.594 ;
               RECT 14.132 32.758 14.186 32.794 ;
               RECT 14.132 33.958 14.186 33.994 ;
               RECT 14.132 35.158 14.186 35.194 ;
               RECT 14.132 36.358 14.186 36.394 ;
               RECT 14.132 37.558 14.186 37.594 ;
               RECT 14.132 38.758 14.186 38.794 ;
               RECT 14.132 39.958 14.186 39.994 ;
               RECT 14.132 41.158 14.186 41.194 ;
               RECT 14.132 42.358 14.186 42.394 ;
               RECT 14.132 43.558 14.186 43.594 ;
               RECT 14.132 44.758 14.186 44.794 ;
               RECT 14.132 45.958 14.186 45.994 ;
               RECT 14.132 47.158 14.186 47.194 ;
               RECT 14.132 48.358 14.186 48.394 ;
               RECT 14.132 50.9205 14.186 50.9565 ;
               RECT 14.132 51.1605 14.186 51.1965 ;
               RECT 14.132 52.7235 14.186 52.7595 ;
               RECT 14.132 54.1635 14.186 54.1995 ;
               RECT 14.132 57.478 14.186 57.514 ;
               RECT 14.132 58.678 14.186 58.714 ;
               RECT 14.132 59.878 14.186 59.914 ;
               RECT 14.132 61.078 14.186 61.114 ;
               RECT 14.132 62.278 14.186 62.314 ;
               RECT 14.132 63.478 14.186 63.514 ;
               RECT 14.132 64.678 14.186 64.714 ;
               RECT 14.132 65.878 14.186 65.914 ;
               RECT 14.132 67.078 14.186 67.114 ;
               RECT 14.132 68.278 14.186 68.314 ;
               RECT 14.132 69.478 14.186 69.514 ;
               RECT 14.132 70.678 14.186 70.714 ;
               RECT 14.132 71.878 14.186 71.914 ;
               RECT 14.132 73.078 14.186 73.114 ;
               RECT 14.132 74.278 14.186 74.314 ;
               RECT 14.132 75.478 14.186 75.514 ;
               RECT 14.132 76.678 14.186 76.714 ;
               RECT 14.132 77.878 14.186 77.914 ;
               RECT 14.132 79.078 14.186 79.114 ;
               RECT 14.132 80.278 14.186 80.314 ;
               RECT 14.132 81.478 14.186 81.514 ;
               RECT 14.132 82.678 14.186 82.714 ;
               RECT 14.132 83.878 14.186 83.914 ;
               RECT 14.132 85.078 14.186 85.114 ;
               RECT 14.132 86.278 14.186 86.314 ;
               RECT 14.132 87.478 14.186 87.514 ;
               RECT 14.132 88.678 14.186 88.714 ;
               RECT 14.132 89.878 14.186 89.914 ;
               RECT 14.132 91.078 14.186 91.114 ;
               RECT 14.132 92.278 14.186 92.314 ;
               RECT 14.132 93.478 14.186 93.514 ;
               RECT 14.132 94.678 14.186 94.714 ;
               RECT 14.132 95.878 14.186 95.914 ;
               RECT 14.132 97.078 14.186 97.114 ;
               RECT 14.132 98.278 14.186 98.314 ;
               RECT 14.132 99.478 14.186 99.514 ;
               RECT 14.132 100.678 14.186 100.714 ;
               RECT 14.132 101.878 14.186 101.914 ;
               RECT 14.132 103.078 14.186 103.114 ;
               RECT 14.132 104.278 14.186 104.314 ;
               RECT 14.214 0.806 14.268 0.842 ;
               RECT 14.214 2.006 14.268 2.042 ;
               RECT 14.214 3.206 14.268 3.242 ;
               RECT 14.214 4.406 14.268 4.442 ;
               RECT 14.214 5.606 14.268 5.642 ;
               RECT 14.214 6.806 14.268 6.842 ;
               RECT 14.214 8.006 14.268 8.042 ;
               RECT 14.214 9.206 14.268 9.242 ;
               RECT 14.214 10.406 14.268 10.442 ;
               RECT 14.214 11.606 14.268 11.642 ;
               RECT 14.214 12.806 14.268 12.842 ;
               RECT 14.214 14.006 14.268 14.042 ;
               RECT 14.214 15.206 14.268 15.242 ;
               RECT 14.214 16.406 14.268 16.442 ;
               RECT 14.214 17.606 14.268 17.642 ;
               RECT 14.214 18.806 14.268 18.842 ;
               RECT 14.214 20.006 14.268 20.042 ;
               RECT 14.214 21.206 14.268 21.242 ;
               RECT 14.214 22.406 14.268 22.442 ;
               RECT 14.214 23.606 14.268 23.642 ;
               RECT 14.214 24.806 14.268 24.842 ;
               RECT 14.214 26.006 14.268 26.042 ;
               RECT 14.214 27.206 14.268 27.242 ;
               RECT 14.214 28.406 14.268 28.442 ;
               RECT 14.214 29.606 14.268 29.642 ;
               RECT 14.214 30.806 14.268 30.842 ;
               RECT 14.214 32.006 14.268 32.042 ;
               RECT 14.214 33.206 14.268 33.242 ;
               RECT 14.214 34.406 14.268 34.442 ;
               RECT 14.214 35.606 14.268 35.642 ;
               RECT 14.214 36.806 14.268 36.842 ;
               RECT 14.214 38.006 14.268 38.042 ;
               RECT 14.214 39.206 14.268 39.242 ;
               RECT 14.214 40.406 14.268 40.442 ;
               RECT 14.214 41.606 14.268 41.642 ;
               RECT 14.214 42.806 14.268 42.842 ;
               RECT 14.214 44.006 14.268 44.042 ;
               RECT 14.214 45.206 14.268 45.242 ;
               RECT 14.214 46.406 14.268 46.442 ;
               RECT 14.214 47.606 14.268 47.642 ;
               RECT 14.214 50.8035 14.268 50.8395 ;
               RECT 14.214 53.8005 14.268 53.8365 ;
               RECT 14.214 56.726 14.268 56.762 ;
               RECT 14.214 57.926 14.268 57.962 ;
               RECT 14.214 59.126 14.268 59.162 ;
               RECT 14.214 60.326 14.268 60.362 ;
               RECT 14.214 61.526 14.268 61.562 ;
               RECT 14.214 62.726 14.268 62.762 ;
               RECT 14.214 63.926 14.268 63.962 ;
               RECT 14.214 65.126 14.268 65.162 ;
               RECT 14.214 66.326 14.268 66.362 ;
               RECT 14.214 67.526 14.268 67.562 ;
               RECT 14.214 68.726 14.268 68.762 ;
               RECT 14.214 69.926 14.268 69.962 ;
               RECT 14.214 71.126 14.268 71.162 ;
               RECT 14.214 72.326 14.268 72.362 ;
               RECT 14.214 73.526 14.268 73.562 ;
               RECT 14.214 74.726 14.268 74.762 ;
               RECT 14.214 75.926 14.268 75.962 ;
               RECT 14.214 77.126 14.268 77.162 ;
               RECT 14.214 78.326 14.268 78.362 ;
               RECT 14.214 79.526 14.268 79.562 ;
               RECT 14.214 80.726 14.268 80.762 ;
               RECT 14.214 81.926 14.268 81.962 ;
               RECT 14.214 83.126 14.268 83.162 ;
               RECT 14.214 84.326 14.268 84.362 ;
               RECT 14.214 85.526 14.268 85.562 ;
               RECT 14.214 86.726 14.268 86.762 ;
               RECT 14.214 87.926 14.268 87.962 ;
               RECT 14.214 89.126 14.268 89.162 ;
               RECT 14.214 90.326 14.268 90.362 ;
               RECT 14.214 91.526 14.268 91.562 ;
               RECT 14.214 92.726 14.268 92.762 ;
               RECT 14.214 93.926 14.268 93.962 ;
               RECT 14.214 95.126 14.268 95.162 ;
               RECT 14.214 96.326 14.268 96.362 ;
               RECT 14.214 97.526 14.268 97.562 ;
               RECT 14.214 98.726 14.268 98.762 ;
               RECT 14.214 99.926 14.268 99.962 ;
               RECT 14.214 101.126 14.268 101.162 ;
               RECT 14.214 102.326 14.268 102.362 ;
               RECT 14.214 103.526 14.268 103.562 ;
               RECT 14.378 50.982 14.422 51.018 ;
               RECT 14.378 51.222 14.422 51.258 ;
               RECT 14.378 53.142 14.422 53.178 ;
               RECT 14.378 54.102 14.422 54.138 ;
               RECT 14.532 1.482 14.586 1.518 ;
               RECT 14.532 2.682 14.586 2.718 ;
               RECT 14.532 3.882 14.586 3.918 ;
               RECT 14.532 5.082 14.586 5.118 ;
               RECT 14.532 6.282 14.586 6.318 ;
               RECT 14.532 7.482 14.586 7.518 ;
               RECT 14.532 8.682 14.586 8.718 ;
               RECT 14.532 9.882 14.586 9.918 ;
               RECT 14.532 11.082 14.586 11.118 ;
               RECT 14.532 12.282 14.586 12.318 ;
               RECT 14.532 13.482 14.586 13.518 ;
               RECT 14.532 14.682 14.586 14.718 ;
               RECT 14.532 15.882 14.586 15.918 ;
               RECT 14.532 17.082 14.586 17.118 ;
               RECT 14.532 18.282 14.586 18.318 ;
               RECT 14.532 19.482 14.586 19.518 ;
               RECT 14.532 20.682 14.586 20.718 ;
               RECT 14.532 21.882 14.586 21.918 ;
               RECT 14.532 23.082 14.586 23.118 ;
               RECT 14.532 24.282 14.586 24.318 ;
               RECT 14.532 25.482 14.586 25.518 ;
               RECT 14.532 26.682 14.586 26.718 ;
               RECT 14.532 27.882 14.586 27.918 ;
               RECT 14.532 29.082 14.586 29.118 ;
               RECT 14.532 30.282 14.586 30.318 ;
               RECT 14.532 31.482 14.586 31.518 ;
               RECT 14.532 32.682 14.586 32.718 ;
               RECT 14.532 33.882 14.586 33.918 ;
               RECT 14.532 35.082 14.586 35.118 ;
               RECT 14.532 36.282 14.586 36.318 ;
               RECT 14.532 37.482 14.586 37.518 ;
               RECT 14.532 38.682 14.586 38.718 ;
               RECT 14.532 39.882 14.586 39.918 ;
               RECT 14.532 41.082 14.586 41.118 ;
               RECT 14.532 42.282 14.586 42.318 ;
               RECT 14.532 43.482 14.586 43.518 ;
               RECT 14.532 44.682 14.586 44.718 ;
               RECT 14.532 45.882 14.586 45.918 ;
               RECT 14.532 47.082 14.586 47.118 ;
               RECT 14.532 48.282 14.586 48.318 ;
               RECT 14.532 49.1235 14.586 49.1595 ;
               RECT 14.532 49.2405 14.586 49.2765 ;
               RECT 14.532 54.4035 14.586 54.4395 ;
               RECT 14.532 55.782 14.586 55.818 ;
               RECT 14.532 56.022 14.586 56.058 ;
               RECT 14.532 57.402 14.586 57.438 ;
               RECT 14.532 58.602 14.586 58.638 ;
               RECT 14.532 59.802 14.586 59.838 ;
               RECT 14.532 61.002 14.586 61.038 ;
               RECT 14.532 62.202 14.586 62.238 ;
               RECT 14.532 63.402 14.586 63.438 ;
               RECT 14.532 64.602 14.586 64.638 ;
               RECT 14.532 65.802 14.586 65.838 ;
               RECT 14.532 67.002 14.586 67.038 ;
               RECT 14.532 68.202 14.586 68.238 ;
               RECT 14.532 69.402 14.586 69.438 ;
               RECT 14.532 70.602 14.586 70.638 ;
               RECT 14.532 71.802 14.586 71.838 ;
               RECT 14.532 73.002 14.586 73.038 ;
               RECT 14.532 74.202 14.586 74.238 ;
               RECT 14.532 75.402 14.586 75.438 ;
               RECT 14.532 76.602 14.586 76.638 ;
               RECT 14.532 77.802 14.586 77.838 ;
               RECT 14.532 79.002 14.586 79.038 ;
               RECT 14.532 80.202 14.586 80.238 ;
               RECT 14.532 81.402 14.586 81.438 ;
               RECT 14.532 82.602 14.586 82.638 ;
               RECT 14.532 83.802 14.586 83.838 ;
               RECT 14.532 85.002 14.586 85.038 ;
               RECT 14.532 86.202 14.586 86.238 ;
               RECT 14.532 87.402 14.586 87.438 ;
               RECT 14.532 88.602 14.586 88.638 ;
               RECT 14.532 89.802 14.586 89.838 ;
               RECT 14.532 91.002 14.586 91.038 ;
               RECT 14.532 92.202 14.586 92.238 ;
               RECT 14.532 93.402 14.586 93.438 ;
               RECT 14.532 94.602 14.586 94.638 ;
               RECT 14.532 95.802 14.586 95.838 ;
               RECT 14.532 97.002 14.586 97.038 ;
               RECT 14.532 98.202 14.586 98.238 ;
               RECT 14.532 99.402 14.586 99.438 ;
               RECT 14.532 100.602 14.586 100.638 ;
               RECT 14.532 101.802 14.586 101.838 ;
               RECT 14.532 103.002 14.586 103.038 ;
               RECT 14.532 104.202 14.586 104.238 ;
               RECT 14.614 0.806 14.668 0.842 ;
               RECT 14.614 2.006 14.668 2.042 ;
               RECT 14.614 3.206 14.668 3.242 ;
               RECT 14.614 4.406 14.668 4.442 ;
               RECT 14.614 5.606 14.668 5.642 ;
               RECT 14.614 6.806 14.668 6.842 ;
               RECT 14.614 8.006 14.668 8.042 ;
               RECT 14.614 9.206 14.668 9.242 ;
               RECT 14.614 10.406 14.668 10.442 ;
               RECT 14.614 11.606 14.668 11.642 ;
               RECT 14.614 12.806 14.668 12.842 ;
               RECT 14.614 14.006 14.668 14.042 ;
               RECT 14.614 15.206 14.668 15.242 ;
               RECT 14.614 16.406 14.668 16.442 ;
               RECT 14.614 17.606 14.668 17.642 ;
               RECT 14.614 18.806 14.668 18.842 ;
               RECT 14.614 20.006 14.668 20.042 ;
               RECT 14.614 21.206 14.668 21.242 ;
               RECT 14.614 22.406 14.668 22.442 ;
               RECT 14.614 23.606 14.668 23.642 ;
               RECT 14.614 24.806 14.668 24.842 ;
               RECT 14.614 26.006 14.668 26.042 ;
               RECT 14.614 27.206 14.668 27.242 ;
               RECT 14.614 28.406 14.668 28.442 ;
               RECT 14.614 29.606 14.668 29.642 ;
               RECT 14.614 30.806 14.668 30.842 ;
               RECT 14.614 32.006 14.668 32.042 ;
               RECT 14.614 33.206 14.668 33.242 ;
               RECT 14.614 34.406 14.668 34.442 ;
               RECT 14.614 35.606 14.668 35.642 ;
               RECT 14.614 36.806 14.668 36.842 ;
               RECT 14.614 38.006 14.668 38.042 ;
               RECT 14.614 39.206 14.668 39.242 ;
               RECT 14.614 40.406 14.668 40.442 ;
               RECT 14.614 41.606 14.668 41.642 ;
               RECT 14.614 42.806 14.668 42.842 ;
               RECT 14.614 44.006 14.668 44.042 ;
               RECT 14.614 45.206 14.668 45.242 ;
               RECT 14.614 46.406 14.668 46.442 ;
               RECT 14.614 47.606 14.668 47.642 ;
               RECT 14.614 49.0005 14.668 49.0365 ;
               RECT 14.614 49.4805 14.668 49.5165 ;
               RECT 14.614 54.6435 14.668 54.6795 ;
               RECT 14.614 55.486 14.668 55.511 ;
               RECT 14.614 55.609 14.668 55.634 ;
               RECT 14.614 56.726 14.668 56.762 ;
               RECT 14.614 57.926 14.668 57.962 ;
               RECT 14.614 59.126 14.668 59.162 ;
               RECT 14.614 60.326 14.668 60.362 ;
               RECT 14.614 61.526 14.668 61.562 ;
               RECT 14.614 62.726 14.668 62.762 ;
               RECT 14.614 63.926 14.668 63.962 ;
               RECT 14.614 65.126 14.668 65.162 ;
               RECT 14.614 66.326 14.668 66.362 ;
               RECT 14.614 67.526 14.668 67.562 ;
               RECT 14.614 68.726 14.668 68.762 ;
               RECT 14.614 69.926 14.668 69.962 ;
               RECT 14.614 71.126 14.668 71.162 ;
               RECT 14.614 72.326 14.668 72.362 ;
               RECT 14.614 73.526 14.668 73.562 ;
               RECT 14.614 74.726 14.668 74.762 ;
               RECT 14.614 75.926 14.668 75.962 ;
               RECT 14.614 77.126 14.668 77.162 ;
               RECT 14.614 78.326 14.668 78.362 ;
               RECT 14.614 79.526 14.668 79.562 ;
               RECT 14.614 80.726 14.668 80.762 ;
               RECT 14.614 81.926 14.668 81.962 ;
               RECT 14.614 83.126 14.668 83.162 ;
               RECT 14.614 84.326 14.668 84.362 ;
               RECT 14.614 85.526 14.668 85.562 ;
               RECT 14.614 86.726 14.668 86.762 ;
               RECT 14.614 87.926 14.668 87.962 ;
               RECT 14.614 89.126 14.668 89.162 ;
               RECT 14.614 90.326 14.668 90.362 ;
               RECT 14.614 91.526 14.668 91.562 ;
               RECT 14.614 92.726 14.668 92.762 ;
               RECT 14.614 93.926 14.668 93.962 ;
               RECT 14.614 95.126 14.668 95.162 ;
               RECT 14.614 96.326 14.668 96.362 ;
               RECT 14.614 97.526 14.668 97.562 ;
               RECT 14.614 98.726 14.668 98.762 ;
               RECT 14.614 99.926 14.668 99.962 ;
               RECT 14.614 101.126 14.668 101.162 ;
               RECT 14.614 102.326 14.668 102.362 ;
               RECT 14.614 103.526 14.668 103.562 ;
               RECT 14.696 1.482 14.75 1.518 ;
               RECT 14.696 2.682 14.75 2.718 ;
               RECT 14.696 3.882 14.75 3.918 ;
               RECT 14.696 5.082 14.75 5.118 ;
               RECT 14.696 6.282 14.75 6.318 ;
               RECT 14.696 7.482 14.75 7.518 ;
               RECT 14.696 8.682 14.75 8.718 ;
               RECT 14.696 9.882 14.75 9.918 ;
               RECT 14.696 11.082 14.75 11.118 ;
               RECT 14.696 12.282 14.75 12.318 ;
               RECT 14.696 13.482 14.75 13.518 ;
               RECT 14.696 14.682 14.75 14.718 ;
               RECT 14.696 15.882 14.75 15.918 ;
               RECT 14.696 17.082 14.75 17.118 ;
               RECT 14.696 18.282 14.75 18.318 ;
               RECT 14.696 19.482 14.75 19.518 ;
               RECT 14.696 20.682 14.75 20.718 ;
               RECT 14.696 21.882 14.75 21.918 ;
               RECT 14.696 23.082 14.75 23.118 ;
               RECT 14.696 24.282 14.75 24.318 ;
               RECT 14.696 25.482 14.75 25.518 ;
               RECT 14.696 26.682 14.75 26.718 ;
               RECT 14.696 27.882 14.75 27.918 ;
               RECT 14.696 29.082 14.75 29.118 ;
               RECT 14.696 30.282 14.75 30.318 ;
               RECT 14.696 31.482 14.75 31.518 ;
               RECT 14.696 32.682 14.75 32.718 ;
               RECT 14.696 33.882 14.75 33.918 ;
               RECT 14.696 35.082 14.75 35.118 ;
               RECT 14.696 36.282 14.75 36.318 ;
               RECT 14.696 37.482 14.75 37.518 ;
               RECT 14.696 38.682 14.75 38.718 ;
               RECT 14.696 39.882 14.75 39.918 ;
               RECT 14.696 41.082 14.75 41.118 ;
               RECT 14.696 42.282 14.75 42.318 ;
               RECT 14.696 43.482 14.75 43.518 ;
               RECT 14.696 44.682 14.75 44.718 ;
               RECT 14.696 45.882 14.75 45.918 ;
               RECT 14.696 47.082 14.75 47.118 ;
               RECT 14.696 48.282 14.75 48.318 ;
               RECT 14.696 49.3635 14.75 49.3995 ;
               RECT 14.696 49.6035 14.75 49.6395 ;
               RECT 14.696 54.4035 14.75 54.4395 ;
               RECT 14.696 55.3635 14.75 55.3995 ;
               RECT 14.696 55.7205 14.75 55.7565 ;
               RECT 14.696 57.402 14.75 57.438 ;
               RECT 14.696 58.602 14.75 58.638 ;
               RECT 14.696 59.802 14.75 59.838 ;
               RECT 14.696 61.002 14.75 61.038 ;
               RECT 14.696 62.202 14.75 62.238 ;
               RECT 14.696 63.402 14.75 63.438 ;
               RECT 14.696 64.602 14.75 64.638 ;
               RECT 14.696 65.802 14.75 65.838 ;
               RECT 14.696 67.002 14.75 67.038 ;
               RECT 14.696 68.202 14.75 68.238 ;
               RECT 14.696 69.402 14.75 69.438 ;
               RECT 14.696 70.602 14.75 70.638 ;
               RECT 14.696 71.802 14.75 71.838 ;
               RECT 14.696 73.002 14.75 73.038 ;
               RECT 14.696 74.202 14.75 74.238 ;
               RECT 14.696 75.402 14.75 75.438 ;
               RECT 14.696 76.602 14.75 76.638 ;
               RECT 14.696 77.802 14.75 77.838 ;
               RECT 14.696 79.002 14.75 79.038 ;
               RECT 14.696 80.202 14.75 80.238 ;
               RECT 14.696 81.402 14.75 81.438 ;
               RECT 14.696 82.602 14.75 82.638 ;
               RECT 14.696 83.802 14.75 83.838 ;
               RECT 14.696 85.002 14.75 85.038 ;
               RECT 14.696 86.202 14.75 86.238 ;
               RECT 14.696 87.402 14.75 87.438 ;
               RECT 14.696 88.602 14.75 88.638 ;
               RECT 14.696 89.802 14.75 89.838 ;
               RECT 14.696 91.002 14.75 91.038 ;
               RECT 14.696 92.202 14.75 92.238 ;
               RECT 14.696 93.402 14.75 93.438 ;
               RECT 14.696 94.602 14.75 94.638 ;
               RECT 14.696 95.802 14.75 95.838 ;
               RECT 14.696 97.002 14.75 97.038 ;
               RECT 14.696 98.202 14.75 98.238 ;
               RECT 14.696 99.402 14.75 99.438 ;
               RECT 14.696 100.602 14.75 100.638 ;
               RECT 14.696 101.802 14.75 101.838 ;
               RECT 14.696 103.002 14.75 103.038 ;
               RECT 14.696 104.202 14.75 104.238 ;
               RECT 14.778 0.806 14.832 0.842 ;
               RECT 14.778 2.006 14.832 2.042 ;
               RECT 14.778 3.206 14.832 3.242 ;
               RECT 14.778 4.406 14.832 4.442 ;
               RECT 14.778 5.606 14.832 5.642 ;
               RECT 14.778 6.806 14.832 6.842 ;
               RECT 14.778 8.006 14.832 8.042 ;
               RECT 14.778 9.206 14.832 9.242 ;
               RECT 14.778 10.406 14.832 10.442 ;
               RECT 14.778 11.606 14.832 11.642 ;
               RECT 14.778 12.806 14.832 12.842 ;
               RECT 14.778 14.006 14.832 14.042 ;
               RECT 14.778 15.206 14.832 15.242 ;
               RECT 14.778 16.406 14.832 16.442 ;
               RECT 14.778 17.606 14.832 17.642 ;
               RECT 14.778 18.806 14.832 18.842 ;
               RECT 14.778 20.006 14.832 20.042 ;
               RECT 14.778 21.206 14.832 21.242 ;
               RECT 14.778 22.406 14.832 22.442 ;
               RECT 14.778 23.606 14.832 23.642 ;
               RECT 14.778 24.806 14.832 24.842 ;
               RECT 14.778 26.006 14.832 26.042 ;
               RECT 14.778 27.206 14.832 27.242 ;
               RECT 14.778 28.406 14.832 28.442 ;
               RECT 14.778 29.606 14.832 29.642 ;
               RECT 14.778 30.806 14.832 30.842 ;
               RECT 14.778 32.006 14.832 32.042 ;
               RECT 14.778 33.206 14.832 33.242 ;
               RECT 14.778 34.406 14.832 34.442 ;
               RECT 14.778 35.606 14.832 35.642 ;
               RECT 14.778 36.806 14.832 36.842 ;
               RECT 14.778 38.006 14.832 38.042 ;
               RECT 14.778 39.206 14.832 39.242 ;
               RECT 14.778 40.406 14.832 40.442 ;
               RECT 14.778 41.606 14.832 41.642 ;
               RECT 14.778 42.806 14.832 42.842 ;
               RECT 14.778 44.006 14.832 44.042 ;
               RECT 14.778 45.206 14.832 45.242 ;
               RECT 14.778 46.406 14.832 46.442 ;
               RECT 14.778 47.606 14.832 47.642 ;
               RECT 14.778 49.7205 14.832 49.7565 ;
               RECT 14.778 50.022 14.832 50.058 ;
               RECT 14.778 54.582 14.832 54.618 ;
               RECT 14.778 55.062 14.832 55.098 ;
               RECT 14.778 55.4805 14.832 55.5165 ;
               RECT 14.778 56.726 14.832 56.762 ;
               RECT 14.778 57.926 14.832 57.962 ;
               RECT 14.778 59.126 14.832 59.162 ;
               RECT 14.778 60.326 14.832 60.362 ;
               RECT 14.778 61.526 14.832 61.562 ;
               RECT 14.778 62.726 14.832 62.762 ;
               RECT 14.778 63.926 14.832 63.962 ;
               RECT 14.778 65.126 14.832 65.162 ;
               RECT 14.778 66.326 14.832 66.362 ;
               RECT 14.778 67.526 14.832 67.562 ;
               RECT 14.778 68.726 14.832 68.762 ;
               RECT 14.778 69.926 14.832 69.962 ;
               RECT 14.778 71.126 14.832 71.162 ;
               RECT 14.778 72.326 14.832 72.362 ;
               RECT 14.778 73.526 14.832 73.562 ;
               RECT 14.778 74.726 14.832 74.762 ;
               RECT 14.778 75.926 14.832 75.962 ;
               RECT 14.778 77.126 14.832 77.162 ;
               RECT 14.778 78.326 14.832 78.362 ;
               RECT 14.778 79.526 14.832 79.562 ;
               RECT 14.778 80.726 14.832 80.762 ;
               RECT 14.778 81.926 14.832 81.962 ;
               RECT 14.778 83.126 14.832 83.162 ;
               RECT 14.778 84.326 14.832 84.362 ;
               RECT 14.778 85.526 14.832 85.562 ;
               RECT 14.778 86.726 14.832 86.762 ;
               RECT 14.778 87.926 14.832 87.962 ;
               RECT 14.778 89.126 14.832 89.162 ;
               RECT 14.778 90.326 14.832 90.362 ;
               RECT 14.778 91.526 14.832 91.562 ;
               RECT 14.778 92.726 14.832 92.762 ;
               RECT 14.778 93.926 14.832 93.962 ;
               RECT 14.778 95.126 14.832 95.162 ;
               RECT 14.778 96.326 14.832 96.362 ;
               RECT 14.778 97.526 14.832 97.562 ;
               RECT 14.778 98.726 14.832 98.762 ;
               RECT 14.778 99.926 14.832 99.962 ;
               RECT 14.778 101.126 14.832 101.162 ;
               RECT 14.778 102.326 14.832 102.362 ;
               RECT 14.778 103.526 14.832 103.562 ;
               RECT 14.86 0.582 14.904 0.618 ;
               RECT 14.86 1.782 14.904 1.818 ;
               RECT 14.86 2.982 14.904 3.018 ;
               RECT 14.86 4.182 14.904 4.218 ;
               RECT 14.86 5.382 14.904 5.418 ;
               RECT 14.86 6.582 14.904 6.618 ;
               RECT 14.86 7.782 14.904 7.818 ;
               RECT 14.86 8.982 14.904 9.018 ;
               RECT 14.86 10.182 14.904 10.218 ;
               RECT 14.86 11.382 14.904 11.418 ;
               RECT 14.86 12.582 14.904 12.618 ;
               RECT 14.86 13.782 14.904 13.818 ;
               RECT 14.86 14.982 14.904 15.018 ;
               RECT 14.86 16.182 14.904 16.218 ;
               RECT 14.86 17.382 14.904 17.418 ;
               RECT 14.86 18.582 14.904 18.618 ;
               RECT 14.86 19.782 14.904 19.818 ;
               RECT 14.86 20.982 14.904 21.018 ;
               RECT 14.86 22.182 14.904 22.218 ;
               RECT 14.86 23.382 14.904 23.418 ;
               RECT 14.86 24.582 14.904 24.618 ;
               RECT 14.86 25.782 14.904 25.818 ;
               RECT 14.86 26.982 14.904 27.018 ;
               RECT 14.86 28.182 14.904 28.218 ;
               RECT 14.86 29.382 14.904 29.418 ;
               RECT 14.86 30.582 14.904 30.618 ;
               RECT 14.86 31.782 14.904 31.818 ;
               RECT 14.86 32.982 14.904 33.018 ;
               RECT 14.86 34.182 14.904 34.218 ;
               RECT 14.86 35.382 14.904 35.418 ;
               RECT 14.86 36.582 14.904 36.618 ;
               RECT 14.86 37.782 14.904 37.818 ;
               RECT 14.86 38.982 14.904 39.018 ;
               RECT 14.86 40.182 14.904 40.218 ;
               RECT 14.86 41.382 14.904 41.418 ;
               RECT 14.86 42.582 14.904 42.618 ;
               RECT 14.86 43.782 14.904 43.818 ;
               RECT 14.86 44.982 14.904 45.018 ;
               RECT 14.86 46.182 14.904 46.218 ;
               RECT 14.86 47.382 14.904 47.418 ;
               RECT 14.86 48.582 14.904 48.618 ;
               RECT 14.86 48.942 14.904 48.978 ;
               RECT 14.86 49.422 14.904 49.458 ;
               RECT 14.86 49.902 14.904 49.938 ;
               RECT 14.86 50.382 14.904 50.418 ;
               RECT 14.86 50.862 14.904 50.898 ;
               RECT 14.86 51.342 14.904 51.378 ;
               RECT 14.86 51.822 14.904 51.858 ;
               RECT 14.86 52.302 14.904 52.338 ;
               RECT 14.86 52.782 14.904 52.818 ;
               RECT 14.86 53.262 14.904 53.298 ;
               RECT 14.86 53.742 14.904 53.778 ;
               RECT 14.86 54.222 14.904 54.258 ;
               RECT 14.86 54.702 14.904 54.738 ;
               RECT 14.86 55.182 14.904 55.218 ;
               RECT 14.86 55.662 14.904 55.698 ;
               RECT 14.86 56.142 14.904 56.178 ;
               RECT 14.86 56.502 14.904 56.538 ;
               RECT 14.86 57.702 14.904 57.738 ;
               RECT 14.86 58.902 14.904 58.938 ;
               RECT 14.86 60.102 14.904 60.138 ;
               RECT 14.86 61.302 14.904 61.338 ;
               RECT 14.86 62.502 14.904 62.538 ;
               RECT 14.86 63.702 14.904 63.738 ;
               RECT 14.86 64.902 14.904 64.938 ;
               RECT 14.86 66.102 14.904 66.138 ;
               RECT 14.86 67.302 14.904 67.338 ;
               RECT 14.86 68.502 14.904 68.538 ;
               RECT 14.86 69.702 14.904 69.738 ;
               RECT 14.86 70.902 14.904 70.938 ;
               RECT 14.86 72.102 14.904 72.138 ;
               RECT 14.86 73.302 14.904 73.338 ;
               RECT 14.86 74.502 14.904 74.538 ;
               RECT 14.86 75.702 14.904 75.738 ;
               RECT 14.86 76.902 14.904 76.938 ;
               RECT 14.86 78.102 14.904 78.138 ;
               RECT 14.86 79.302 14.904 79.338 ;
               RECT 14.86 80.502 14.904 80.538 ;
               RECT 14.86 81.702 14.904 81.738 ;
               RECT 14.86 82.902 14.904 82.938 ;
               RECT 14.86 84.102 14.904 84.138 ;
               RECT 14.86 85.302 14.904 85.338 ;
               RECT 14.86 86.502 14.904 86.538 ;
               RECT 14.86 87.702 14.904 87.738 ;
               RECT 14.86 88.902 14.904 88.938 ;
               RECT 14.86 90.102 14.904 90.138 ;
               RECT 14.86 91.302 14.904 91.338 ;
               RECT 14.86 92.502 14.904 92.538 ;
               RECT 14.86 93.702 14.904 93.738 ;
               RECT 14.86 94.902 14.904 94.938 ;
               RECT 14.86 96.102 14.904 96.138 ;
               RECT 14.86 97.302 14.904 97.338 ;
               RECT 14.86 98.502 14.904 98.538 ;
               RECT 14.86 99.702 14.904 99.738 ;
               RECT 14.86 100.902 14.904 100.938 ;
               RECT 14.86 102.102 14.904 102.138 ;
               RECT 14.86 103.302 14.904 103.338 ;
               RECT 14.86 104.502 14.904 104.538 ;
               RECT 15.014 51.2835 15.068 51.3195 ;
               RECT 15.014 54.1635 15.068 54.1995 ;
               RECT 15.178 0.582 15.222 0.618 ;
               RECT 15.178 1.182 15.222 1.218 ;
               RECT 15.178 1.782 15.222 1.818 ;
               RECT 15.178 2.382 15.222 2.418 ;
               RECT 15.178 2.982 15.222 3.018 ;
               RECT 15.178 3.582 15.222 3.618 ;
               RECT 15.178 4.182 15.222 4.218 ;
               RECT 15.178 4.782 15.222 4.818 ;
               RECT 15.178 5.382 15.222 5.418 ;
               RECT 15.178 5.982 15.222 6.018 ;
               RECT 15.178 6.582 15.222 6.618 ;
               RECT 15.178 7.182 15.222 7.218 ;
               RECT 15.178 7.782 15.222 7.818 ;
               RECT 15.178 8.382 15.222 8.418 ;
               RECT 15.178 8.982 15.222 9.018 ;
               RECT 15.178 9.582 15.222 9.618 ;
               RECT 15.178 10.182 15.222 10.218 ;
               RECT 15.178 10.782 15.222 10.818 ;
               RECT 15.178 11.382 15.222 11.418 ;
               RECT 15.178 11.982 15.222 12.018 ;
               RECT 15.178 12.582 15.222 12.618 ;
               RECT 15.178 13.182 15.222 13.218 ;
               RECT 15.178 13.782 15.222 13.818 ;
               RECT 15.178 14.382 15.222 14.418 ;
               RECT 15.178 14.982 15.222 15.018 ;
               RECT 15.178 15.582 15.222 15.618 ;
               RECT 15.178 16.182 15.222 16.218 ;
               RECT 15.178 16.782 15.222 16.818 ;
               RECT 15.178 17.382 15.222 17.418 ;
               RECT 15.178 17.982 15.222 18.018 ;
               RECT 15.178 18.582 15.222 18.618 ;
               RECT 15.178 19.182 15.222 19.218 ;
               RECT 15.178 19.782 15.222 19.818 ;
               RECT 15.178 20.382 15.222 20.418 ;
               RECT 15.178 20.982 15.222 21.018 ;
               RECT 15.178 21.582 15.222 21.618 ;
               RECT 15.178 22.182 15.222 22.218 ;
               RECT 15.178 22.782 15.222 22.818 ;
               RECT 15.178 23.382 15.222 23.418 ;
               RECT 15.178 23.982 15.222 24.018 ;
               RECT 15.178 24.582 15.222 24.618 ;
               RECT 15.178 25.182 15.222 25.218 ;
               RECT 15.178 25.782 15.222 25.818 ;
               RECT 15.178 26.382 15.222 26.418 ;
               RECT 15.178 26.982 15.222 27.018 ;
               RECT 15.178 27.582 15.222 27.618 ;
               RECT 15.178 28.182 15.222 28.218 ;
               RECT 15.178 28.782 15.222 28.818 ;
               RECT 15.178 29.382 15.222 29.418 ;
               RECT 15.178 29.982 15.222 30.018 ;
               RECT 15.178 30.582 15.222 30.618 ;
               RECT 15.178 31.182 15.222 31.218 ;
               RECT 15.178 31.782 15.222 31.818 ;
               RECT 15.178 32.382 15.222 32.418 ;
               RECT 15.178 32.982 15.222 33.018 ;
               RECT 15.178 33.582 15.222 33.618 ;
               RECT 15.178 34.182 15.222 34.218 ;
               RECT 15.178 34.782 15.222 34.818 ;
               RECT 15.178 35.382 15.222 35.418 ;
               RECT 15.178 35.982 15.222 36.018 ;
               RECT 15.178 36.582 15.222 36.618 ;
               RECT 15.178 37.182 15.222 37.218 ;
               RECT 15.178 37.782 15.222 37.818 ;
               RECT 15.178 38.382 15.222 38.418 ;
               RECT 15.178 38.982 15.222 39.018 ;
               RECT 15.178 39.582 15.222 39.618 ;
               RECT 15.178 40.182 15.222 40.218 ;
               RECT 15.178 40.782 15.222 40.818 ;
               RECT 15.178 41.382 15.222 41.418 ;
               RECT 15.178 41.982 15.222 42.018 ;
               RECT 15.178 42.582 15.222 42.618 ;
               RECT 15.178 43.182 15.222 43.218 ;
               RECT 15.178 43.782 15.222 43.818 ;
               RECT 15.178 44.382 15.222 44.418 ;
               RECT 15.178 44.982 15.222 45.018 ;
               RECT 15.178 45.582 15.222 45.618 ;
               RECT 15.178 46.182 15.222 46.218 ;
               RECT 15.178 46.782 15.222 46.818 ;
               RECT 15.178 47.382 15.222 47.418 ;
               RECT 15.178 47.982 15.222 48.018 ;
               RECT 15.178 48.582 15.222 48.618 ;
               RECT 15.178 48.942 15.222 48.978 ;
               RECT 15.178 49.422 15.222 49.458 ;
               RECT 15.178 49.902 15.222 49.938 ;
               RECT 15.178 50.0835 15.222 50.1195 ;
               RECT 15.178 50.382 15.222 50.418 ;
               RECT 15.178 50.862 15.222 50.898 ;
               RECT 15.178 51.342 15.222 51.378 ;
               RECT 15.178 51.822 15.222 51.858 ;
               RECT 15.178 52.302 15.222 52.338 ;
               RECT 15.178 52.782 15.222 52.818 ;
               RECT 15.178 53.262 15.222 53.298 ;
               RECT 15.178 53.742 15.222 53.778 ;
               RECT 15.178 54.2275 15.222 54.2525 ;
               RECT 15.178 54.7075 15.222 54.7325 ;
               RECT 15.178 55.182 15.222 55.218 ;
               RECT 15.178 55.6675 15.222 55.6925 ;
               RECT 15.178 56.142 15.222 56.178 ;
               RECT 15.178 56.502 15.222 56.538 ;
               RECT 15.178 57.102 15.222 57.138 ;
               RECT 15.178 57.702 15.222 57.738 ;
               RECT 15.178 58.302 15.222 58.338 ;
               RECT 15.178 58.902 15.222 58.938 ;
               RECT 15.178 59.502 15.222 59.538 ;
               RECT 15.178 60.102 15.222 60.138 ;
               RECT 15.178 60.702 15.222 60.738 ;
               RECT 15.178 61.302 15.222 61.338 ;
               RECT 15.178 61.902 15.222 61.938 ;
               RECT 15.178 62.502 15.222 62.538 ;
               RECT 15.178 63.102 15.222 63.138 ;
               RECT 15.178 63.702 15.222 63.738 ;
               RECT 15.178 64.302 15.222 64.338 ;
               RECT 15.178 64.902 15.222 64.938 ;
               RECT 15.178 65.502 15.222 65.538 ;
               RECT 15.178 66.102 15.222 66.138 ;
               RECT 15.178 66.702 15.222 66.738 ;
               RECT 15.178 67.302 15.222 67.338 ;
               RECT 15.178 67.902 15.222 67.938 ;
               RECT 15.178 68.502 15.222 68.538 ;
               RECT 15.178 69.102 15.222 69.138 ;
               RECT 15.178 69.702 15.222 69.738 ;
               RECT 15.178 70.302 15.222 70.338 ;
               RECT 15.178 70.902 15.222 70.938 ;
               RECT 15.178 71.502 15.222 71.538 ;
               RECT 15.178 72.102 15.222 72.138 ;
               RECT 15.178 72.702 15.222 72.738 ;
               RECT 15.178 73.302 15.222 73.338 ;
               RECT 15.178 73.902 15.222 73.938 ;
               RECT 15.178 74.502 15.222 74.538 ;
               RECT 15.178 75.102 15.222 75.138 ;
               RECT 15.178 75.702 15.222 75.738 ;
               RECT 15.178 76.302 15.222 76.338 ;
               RECT 15.178 76.902 15.222 76.938 ;
               RECT 15.178 77.502 15.222 77.538 ;
               RECT 15.178 78.102 15.222 78.138 ;
               RECT 15.178 78.702 15.222 78.738 ;
               RECT 15.178 79.302 15.222 79.338 ;
               RECT 15.178 79.902 15.222 79.938 ;
               RECT 15.178 80.502 15.222 80.538 ;
               RECT 15.178 81.102 15.222 81.138 ;
               RECT 15.178 81.702 15.222 81.738 ;
               RECT 15.178 82.302 15.222 82.338 ;
               RECT 15.178 82.902 15.222 82.938 ;
               RECT 15.178 83.502 15.222 83.538 ;
               RECT 15.178 84.102 15.222 84.138 ;
               RECT 15.178 84.702 15.222 84.738 ;
               RECT 15.178 85.302 15.222 85.338 ;
               RECT 15.178 85.902 15.222 85.938 ;
               RECT 15.178 86.502 15.222 86.538 ;
               RECT 15.178 87.102 15.222 87.138 ;
               RECT 15.178 87.702 15.222 87.738 ;
               RECT 15.178 88.302 15.222 88.338 ;
               RECT 15.178 88.902 15.222 88.938 ;
               RECT 15.178 89.502 15.222 89.538 ;
               RECT 15.178 90.102 15.222 90.138 ;
               RECT 15.178 90.702 15.222 90.738 ;
               RECT 15.178 91.302 15.222 91.338 ;
               RECT 15.178 91.902 15.222 91.938 ;
               RECT 15.178 92.502 15.222 92.538 ;
               RECT 15.178 93.102 15.222 93.138 ;
               RECT 15.178 93.702 15.222 93.738 ;
               RECT 15.178 94.302 15.222 94.338 ;
               RECT 15.178 94.902 15.222 94.938 ;
               RECT 15.178 95.502 15.222 95.538 ;
               RECT 15.178 96.102 15.222 96.138 ;
               RECT 15.178 96.702 15.222 96.738 ;
               RECT 15.178 97.302 15.222 97.338 ;
               RECT 15.178 97.902 15.222 97.938 ;
               RECT 15.178 98.502 15.222 98.538 ;
               RECT 15.178 99.102 15.222 99.138 ;
               RECT 15.178 99.702 15.222 99.738 ;
               RECT 15.178 100.302 15.222 100.338 ;
               RECT 15.178 100.902 15.222 100.938 ;
               RECT 15.178 101.502 15.222 101.538 ;
               RECT 15.178 102.102 15.222 102.138 ;
               RECT 15.178 102.702 15.222 102.738 ;
               RECT 15.178 103.302 15.222 103.338 ;
               RECT 15.178 103.902 15.222 103.938 ;
               RECT 15.178 104.502 15.222 104.538 ;
               RECT 15.398 51.4005 15.45 51.4365 ;
               RECT 15.398 52.902 15.45 52.938 ;
               RECT 15.478 50.502 15.53 50.538 ;
               RECT 15.478 54.8835 15.53 54.9195 ;
               RECT 15.558 1.3345 15.63 1.3595 ;
               RECT 15.558 2.5345 15.63 2.5595 ;
               RECT 15.558 3.7345 15.63 3.7595 ;
               RECT 15.558 4.9345 15.63 4.9595 ;
               RECT 15.558 6.1345 15.63 6.1595 ;
               RECT 15.558 7.3345 15.63 7.3595 ;
               RECT 15.558 8.5345 15.63 8.5595 ;
               RECT 15.558 9.7345 15.63 9.7595 ;
               RECT 15.558 10.9345 15.63 10.9595 ;
               RECT 15.558 12.1345 15.63 12.1595 ;
               RECT 15.558 13.3345 15.63 13.3595 ;
               RECT 15.558 14.5345 15.63 14.5595 ;
               RECT 15.558 15.7345 15.63 15.7595 ;
               RECT 15.558 16.9345 15.63 16.9595 ;
               RECT 15.558 18.1345 15.63 18.1595 ;
               RECT 15.558 19.3345 15.63 19.3595 ;
               RECT 15.558 20.5345 15.63 20.5595 ;
               RECT 15.558 21.7345 15.63 21.7595 ;
               RECT 15.558 22.9345 15.63 22.9595 ;
               RECT 15.558 24.1345 15.63 24.1595 ;
               RECT 15.558 25.3345 15.63 25.3595 ;
               RECT 15.558 26.5345 15.63 26.5595 ;
               RECT 15.558 27.7345 15.63 27.7595 ;
               RECT 15.558 28.9345 15.63 28.9595 ;
               RECT 15.558 30.1345 15.63 30.1595 ;
               RECT 15.558 31.3345 15.63 31.3595 ;
               RECT 15.558 32.5345 15.63 32.5595 ;
               RECT 15.558 33.7345 15.63 33.7595 ;
               RECT 15.558 34.9345 15.63 34.9595 ;
               RECT 15.558 36.1345 15.63 36.1595 ;
               RECT 15.558 37.3345 15.63 37.3595 ;
               RECT 15.558 38.5345 15.63 38.5595 ;
               RECT 15.558 39.7345 15.63 39.7595 ;
               RECT 15.558 40.9345 15.63 40.9595 ;
               RECT 15.558 42.1345 15.63 42.1595 ;
               RECT 15.558 43.3345 15.63 43.3595 ;
               RECT 15.558 44.5345 15.63 44.5595 ;
               RECT 15.558 45.7345 15.63 45.7595 ;
               RECT 15.558 46.9345 15.63 46.9595 ;
               RECT 15.558 48.1345 15.63 48.1595 ;
               RECT 15.558 49.0675 15.63 49.0925 ;
               RECT 15.558 50.2675 15.63 50.2925 ;
               RECT 15.558 54.5875 15.63 54.6125 ;
               RECT 15.558 56.0275 15.63 56.0525 ;
               RECT 15.558 57.2545 15.63 57.2795 ;
               RECT 15.558 58.4545 15.63 58.4795 ;
               RECT 15.558 59.6545 15.63 59.6795 ;
               RECT 15.558 60.8545 15.63 60.8795 ;
               RECT 15.558 62.0545 15.63 62.0795 ;
               RECT 15.558 63.2545 15.63 63.2795 ;
               RECT 15.558 64.4545 15.63 64.4795 ;
               RECT 15.558 65.6545 15.63 65.6795 ;
               RECT 15.558 66.8545 15.63 66.8795 ;
               RECT 15.558 68.0545 15.63 68.0795 ;
               RECT 15.558 69.2545 15.63 69.2795 ;
               RECT 15.558 70.4545 15.63 70.4795 ;
               RECT 15.558 71.6545 15.63 71.6795 ;
               RECT 15.558 72.8545 15.63 72.8795 ;
               RECT 15.558 74.0545 15.63 74.0795 ;
               RECT 15.558 75.2545 15.63 75.2795 ;
               RECT 15.558 76.4545 15.63 76.4795 ;
               RECT 15.558 77.6545 15.63 77.6795 ;
               RECT 15.558 78.8545 15.63 78.8795 ;
               RECT 15.558 80.0545 15.63 80.0795 ;
               RECT 15.558 81.2545 15.63 81.2795 ;
               RECT 15.558 82.4545 15.63 82.4795 ;
               RECT 15.558 83.6545 15.63 83.6795 ;
               RECT 15.558 84.8545 15.63 84.8795 ;
               RECT 15.558 86.0545 15.63 86.0795 ;
               RECT 15.558 87.2545 15.63 87.2795 ;
               RECT 15.558 88.4545 15.63 88.4795 ;
               RECT 15.558 89.6545 15.63 89.6795 ;
               RECT 15.558 90.8545 15.63 90.8795 ;
               RECT 15.558 92.0545 15.63 92.0795 ;
               RECT 15.558 93.2545 15.63 93.2795 ;
               RECT 15.558 94.4545 15.63 94.4795 ;
               RECT 15.558 95.6545 15.63 95.6795 ;
               RECT 15.558 96.8545 15.63 96.8795 ;
               RECT 15.558 98.0545 15.63 98.0795 ;
               RECT 15.558 99.2545 15.63 99.2795 ;
               RECT 15.558 100.4545 15.63 100.4795 ;
               RECT 15.558 101.6545 15.63 101.6795 ;
               RECT 15.558 102.8545 15.63 102.8795 ;
               RECT 15.558 104.0545 15.63 104.0795 ;
               RECT 15.738 50.022 15.778 50.058 ;
               RECT 15.738 52.4835 15.778 52.5195 ;
               RECT 15.738 55.062 15.778 55.098 ;
               RECT 15.806 49.782 15.846 49.818 ;
               RECT 15.806 54.102 15.846 54.138 ;
               RECT 16.114 1.558 16.162 1.594 ;
               RECT 16.114 2.758 16.162 2.794 ;
               RECT 16.114 3.958 16.162 3.994 ;
               RECT 16.114 5.158 16.162 5.194 ;
               RECT 16.114 6.358 16.162 6.394 ;
               RECT 16.114 7.558 16.162 7.594 ;
               RECT 16.114 8.758 16.162 8.794 ;
               RECT 16.114 9.958 16.162 9.994 ;
               RECT 16.114 11.158 16.162 11.194 ;
               RECT 16.114 12.358 16.162 12.394 ;
               RECT 16.114 13.558 16.162 13.594 ;
               RECT 16.114 14.758 16.162 14.794 ;
               RECT 16.114 15.958 16.162 15.994 ;
               RECT 16.114 17.158 16.162 17.194 ;
               RECT 16.114 18.358 16.162 18.394 ;
               RECT 16.114 19.558 16.162 19.594 ;
               RECT 16.114 20.758 16.162 20.794 ;
               RECT 16.114 21.958 16.162 21.994 ;
               RECT 16.114 23.158 16.162 23.194 ;
               RECT 16.114 24.358 16.162 24.394 ;
               RECT 16.114 25.558 16.162 25.594 ;
               RECT 16.114 26.758 16.162 26.794 ;
               RECT 16.114 27.958 16.162 27.994 ;
               RECT 16.114 29.158 16.162 29.194 ;
               RECT 16.114 30.358 16.162 30.394 ;
               RECT 16.114 31.558 16.162 31.594 ;
               RECT 16.114 32.758 16.162 32.794 ;
               RECT 16.114 33.958 16.162 33.994 ;
               RECT 16.114 35.158 16.162 35.194 ;
               RECT 16.114 36.358 16.162 36.394 ;
               RECT 16.114 37.558 16.162 37.594 ;
               RECT 16.114 38.758 16.162 38.794 ;
               RECT 16.114 39.958 16.162 39.994 ;
               RECT 16.114 41.158 16.162 41.194 ;
               RECT 16.114 42.358 16.162 42.394 ;
               RECT 16.114 43.558 16.162 43.594 ;
               RECT 16.114 44.758 16.162 44.794 ;
               RECT 16.114 45.958 16.162 45.994 ;
               RECT 16.114 47.158 16.162 47.194 ;
               RECT 16.114 48.358 16.162 48.394 ;
               RECT 16.114 49.542 16.162 49.578 ;
               RECT 16.114 55.7205 16.162 55.7565 ;
               RECT 16.114 57.478 16.162 57.514 ;
               RECT 16.114 58.678 16.162 58.714 ;
               RECT 16.114 59.878 16.162 59.914 ;
               RECT 16.114 61.078 16.162 61.114 ;
               RECT 16.114 62.278 16.162 62.314 ;
               RECT 16.114 63.478 16.162 63.514 ;
               RECT 16.114 64.678 16.162 64.714 ;
               RECT 16.114 65.878 16.162 65.914 ;
               RECT 16.114 67.078 16.162 67.114 ;
               RECT 16.114 68.278 16.162 68.314 ;
               RECT 16.114 69.478 16.162 69.514 ;
               RECT 16.114 70.678 16.162 70.714 ;
               RECT 16.114 71.878 16.162 71.914 ;
               RECT 16.114 73.078 16.162 73.114 ;
               RECT 16.114 74.278 16.162 74.314 ;
               RECT 16.114 75.478 16.162 75.514 ;
               RECT 16.114 76.678 16.162 76.714 ;
               RECT 16.114 77.878 16.162 77.914 ;
               RECT 16.114 79.078 16.162 79.114 ;
               RECT 16.114 80.278 16.162 80.314 ;
               RECT 16.114 81.478 16.162 81.514 ;
               RECT 16.114 82.678 16.162 82.714 ;
               RECT 16.114 83.878 16.162 83.914 ;
               RECT 16.114 85.078 16.162 85.114 ;
               RECT 16.114 86.278 16.162 86.314 ;
               RECT 16.114 87.478 16.162 87.514 ;
               RECT 16.114 88.678 16.162 88.714 ;
               RECT 16.114 89.878 16.162 89.914 ;
               RECT 16.114 91.078 16.162 91.114 ;
               RECT 16.114 92.278 16.162 92.314 ;
               RECT 16.114 93.478 16.162 93.514 ;
               RECT 16.114 94.678 16.162 94.714 ;
               RECT 16.114 95.878 16.162 95.914 ;
               RECT 16.114 97.078 16.162 97.114 ;
               RECT 16.114 98.278 16.162 98.314 ;
               RECT 16.114 99.478 16.162 99.514 ;
               RECT 16.114 100.678 16.162 100.714 ;
               RECT 16.114 101.878 16.162 101.914 ;
               RECT 16.114 103.078 16.162 103.114 ;
               RECT 16.114 104.278 16.162 104.314 ;
               RECT 16.19 1.035 16.238 1.071 ;
               RECT 16.19 2.235 16.238 2.271 ;
               RECT 16.19 3.435 16.238 3.471 ;
               RECT 16.19 4.635 16.238 4.671 ;
               RECT 16.19 5.835 16.238 5.871 ;
               RECT 16.19 7.035 16.238 7.071 ;
               RECT 16.19 8.235 16.238 8.271 ;
               RECT 16.19 9.435 16.238 9.471 ;
               RECT 16.19 10.635 16.238 10.671 ;
               RECT 16.19 11.835 16.238 11.871 ;
               RECT 16.19 13.035 16.238 13.071 ;
               RECT 16.19 14.235 16.238 14.271 ;
               RECT 16.19 15.435 16.238 15.471 ;
               RECT 16.19 16.635 16.238 16.671 ;
               RECT 16.19 17.835 16.238 17.871 ;
               RECT 16.19 19.035 16.238 19.071 ;
               RECT 16.19 20.235 16.238 20.271 ;
               RECT 16.19 21.435 16.238 21.471 ;
               RECT 16.19 22.635 16.238 22.671 ;
               RECT 16.19 23.835 16.238 23.871 ;
               RECT 16.19 25.035 16.238 25.071 ;
               RECT 16.19 26.235 16.238 26.271 ;
               RECT 16.19 27.435 16.238 27.471 ;
               RECT 16.19 28.635 16.238 28.671 ;
               RECT 16.19 29.835 16.238 29.871 ;
               RECT 16.19 31.035 16.238 31.071 ;
               RECT 16.19 32.235 16.238 32.271 ;
               RECT 16.19 33.435 16.238 33.471 ;
               RECT 16.19 34.635 16.238 34.671 ;
               RECT 16.19 35.835 16.238 35.871 ;
               RECT 16.19 37.035 16.238 37.071 ;
               RECT 16.19 38.235 16.238 38.271 ;
               RECT 16.19 39.435 16.238 39.471 ;
               RECT 16.19 40.635 16.238 40.671 ;
               RECT 16.19 41.835 16.238 41.871 ;
               RECT 16.19 43.035 16.238 43.071 ;
               RECT 16.19 44.235 16.238 44.271 ;
               RECT 16.19 45.435 16.238 45.471 ;
               RECT 16.19 46.635 16.238 46.671 ;
               RECT 16.19 47.835 16.238 47.871 ;
               RECT 16.19 49.302 16.238 49.338 ;
               RECT 16.19 50.022 16.238 50.058 ;
               RECT 16.19 54.0405 16.238 54.0765 ;
               RECT 16.19 55.2405 16.238 55.2765 ;
               RECT 16.19 55.542 16.238 55.578 ;
               RECT 16.19 56.955 16.238 56.991 ;
               RECT 16.19 58.155 16.238 58.191 ;
               RECT 16.19 59.355 16.238 59.391 ;
               RECT 16.19 60.555 16.238 60.591 ;
               RECT 16.19 61.755 16.238 61.791 ;
               RECT 16.19 62.955 16.238 62.991 ;
               RECT 16.19 64.155 16.238 64.191 ;
               RECT 16.19 65.355 16.238 65.391 ;
               RECT 16.19 66.555 16.238 66.591 ;
               RECT 16.19 67.755 16.238 67.791 ;
               RECT 16.19 68.955 16.238 68.991 ;
               RECT 16.19 70.155 16.238 70.191 ;
               RECT 16.19 71.355 16.238 71.391 ;
               RECT 16.19 72.555 16.238 72.591 ;
               RECT 16.19 73.755 16.238 73.791 ;
               RECT 16.19 74.955 16.238 74.991 ;
               RECT 16.19 76.155 16.238 76.191 ;
               RECT 16.19 77.355 16.238 77.391 ;
               RECT 16.19 78.555 16.238 78.591 ;
               RECT 16.19 79.755 16.238 79.791 ;
               RECT 16.19 80.955 16.238 80.991 ;
               RECT 16.19 82.155 16.238 82.191 ;
               RECT 16.19 83.355 16.238 83.391 ;
               RECT 16.19 84.555 16.238 84.591 ;
               RECT 16.19 85.755 16.238 85.791 ;
               RECT 16.19 86.955 16.238 86.991 ;
               RECT 16.19 88.155 16.238 88.191 ;
               RECT 16.19 89.355 16.238 89.391 ;
               RECT 16.19 90.555 16.238 90.591 ;
               RECT 16.19 91.755 16.238 91.791 ;
               RECT 16.19 92.955 16.238 92.991 ;
               RECT 16.19 94.155 16.238 94.191 ;
               RECT 16.19 95.355 16.238 95.391 ;
               RECT 16.19 96.555 16.238 96.591 ;
               RECT 16.19 97.755 16.238 97.791 ;
               RECT 16.19 98.955 16.238 98.991 ;
               RECT 16.19 100.155 16.238 100.191 ;
               RECT 16.19 101.355 16.238 101.391 ;
               RECT 16.19 102.555 16.238 102.591 ;
               RECT 16.19 103.755 16.238 103.791 ;
               RECT 16.346 1.329 16.394 1.365 ;
               RECT 16.346 2.529 16.394 2.565 ;
               RECT 16.346 3.729 16.394 3.765 ;
               RECT 16.346 4.929 16.394 4.965 ;
               RECT 16.346 6.129 16.394 6.165 ;
               RECT 16.346 7.329 16.394 7.365 ;
               RECT 16.346 8.529 16.394 8.565 ;
               RECT 16.346 9.729 16.394 9.765 ;
               RECT 16.346 10.929 16.394 10.965 ;
               RECT 16.346 12.129 16.394 12.165 ;
               RECT 16.346 13.329 16.394 13.365 ;
               RECT 16.346 14.529 16.394 14.565 ;
               RECT 16.346 15.729 16.394 15.765 ;
               RECT 16.346 16.929 16.394 16.965 ;
               RECT 16.346 18.129 16.394 18.165 ;
               RECT 16.346 19.329 16.394 19.365 ;
               RECT 16.346 20.529 16.394 20.565 ;
               RECT 16.346 21.729 16.394 21.765 ;
               RECT 16.346 22.929 16.394 22.965 ;
               RECT 16.346 24.129 16.394 24.165 ;
               RECT 16.346 25.329 16.394 25.365 ;
               RECT 16.346 26.529 16.394 26.565 ;
               RECT 16.346 27.729 16.394 27.765 ;
               RECT 16.346 28.929 16.394 28.965 ;
               RECT 16.346 30.129 16.394 30.165 ;
               RECT 16.346 31.329 16.394 31.365 ;
               RECT 16.346 32.529 16.394 32.565 ;
               RECT 16.346 33.729 16.394 33.765 ;
               RECT 16.346 34.929 16.394 34.965 ;
               RECT 16.346 36.129 16.394 36.165 ;
               RECT 16.346 37.329 16.394 37.365 ;
               RECT 16.346 38.529 16.394 38.565 ;
               RECT 16.346 39.729 16.394 39.765 ;
               RECT 16.346 40.929 16.394 40.965 ;
               RECT 16.346 42.129 16.394 42.165 ;
               RECT 16.346 43.329 16.394 43.365 ;
               RECT 16.346 44.529 16.394 44.565 ;
               RECT 16.346 45.729 16.394 45.765 ;
               RECT 16.346 46.929 16.394 46.965 ;
               RECT 16.346 48.129 16.394 48.165 ;
               RECT 16.346 49.4805 16.394 49.5165 ;
               RECT 16.346 50.022 16.394 50.058 ;
               RECT 16.346 52.422 16.394 52.458 ;
               RECT 16.346 55.062 16.394 55.098 ;
               RECT 16.346 55.782 16.394 55.818 ;
               RECT 16.346 57.249 16.394 57.285 ;
               RECT 16.346 58.449 16.394 58.485 ;
               RECT 16.346 59.649 16.394 59.685 ;
               RECT 16.346 60.849 16.394 60.885 ;
               RECT 16.346 62.049 16.394 62.085 ;
               RECT 16.346 63.249 16.394 63.285 ;
               RECT 16.346 64.449 16.394 64.485 ;
               RECT 16.346 65.649 16.394 65.685 ;
               RECT 16.346 66.849 16.394 66.885 ;
               RECT 16.346 68.049 16.394 68.085 ;
               RECT 16.346 69.249 16.394 69.285 ;
               RECT 16.346 70.449 16.394 70.485 ;
               RECT 16.346 71.649 16.394 71.685 ;
               RECT 16.346 72.849 16.394 72.885 ;
               RECT 16.346 74.049 16.394 74.085 ;
               RECT 16.346 75.249 16.394 75.285 ;
               RECT 16.346 76.449 16.394 76.485 ;
               RECT 16.346 77.649 16.394 77.685 ;
               RECT 16.346 78.849 16.394 78.885 ;
               RECT 16.346 80.049 16.394 80.085 ;
               RECT 16.346 81.249 16.394 81.285 ;
               RECT 16.346 82.449 16.394 82.485 ;
               RECT 16.346 83.649 16.394 83.685 ;
               RECT 16.346 84.849 16.394 84.885 ;
               RECT 16.346 86.049 16.394 86.085 ;
               RECT 16.346 87.249 16.394 87.285 ;
               RECT 16.346 88.449 16.394 88.485 ;
               RECT 16.346 89.649 16.394 89.685 ;
               RECT 16.346 90.849 16.394 90.885 ;
               RECT 16.346 92.049 16.394 92.085 ;
               RECT 16.346 93.249 16.394 93.285 ;
               RECT 16.346 94.449 16.394 94.485 ;
               RECT 16.346 95.649 16.394 95.685 ;
               RECT 16.346 96.849 16.394 96.885 ;
               RECT 16.346 98.049 16.394 98.085 ;
               RECT 16.346 99.249 16.394 99.285 ;
               RECT 16.346 100.449 16.394 100.485 ;
               RECT 16.346 101.649 16.394 101.685 ;
               RECT 16.346 102.849 16.394 102.885 ;
               RECT 16.346 104.049 16.394 104.085 ;
               RECT 16.422 1.558 16.47 1.594 ;
               RECT 16.422 2.758 16.47 2.794 ;
               RECT 16.422 3.958 16.47 3.994 ;
               RECT 16.422 5.158 16.47 5.194 ;
               RECT 16.422 6.358 16.47 6.394 ;
               RECT 16.422 7.558 16.47 7.594 ;
               RECT 16.422 8.758 16.47 8.794 ;
               RECT 16.422 9.958 16.47 9.994 ;
               RECT 16.422 11.158 16.47 11.194 ;
               RECT 16.422 12.358 16.47 12.394 ;
               RECT 16.422 13.558 16.47 13.594 ;
               RECT 16.422 14.758 16.47 14.794 ;
               RECT 16.422 15.958 16.47 15.994 ;
               RECT 16.422 17.158 16.47 17.194 ;
               RECT 16.422 18.358 16.47 18.394 ;
               RECT 16.422 19.558 16.47 19.594 ;
               RECT 16.422 20.758 16.47 20.794 ;
               RECT 16.422 21.958 16.47 21.994 ;
               RECT 16.422 23.158 16.47 23.194 ;
               RECT 16.422 24.358 16.47 24.394 ;
               RECT 16.422 25.558 16.47 25.594 ;
               RECT 16.422 26.758 16.47 26.794 ;
               RECT 16.422 27.958 16.47 27.994 ;
               RECT 16.422 29.158 16.47 29.194 ;
               RECT 16.422 30.358 16.47 30.394 ;
               RECT 16.422 31.558 16.47 31.594 ;
               RECT 16.422 32.758 16.47 32.794 ;
               RECT 16.422 33.958 16.47 33.994 ;
               RECT 16.422 35.158 16.47 35.194 ;
               RECT 16.422 36.358 16.47 36.394 ;
               RECT 16.422 37.558 16.47 37.594 ;
               RECT 16.422 38.758 16.47 38.794 ;
               RECT 16.422 39.958 16.47 39.994 ;
               RECT 16.422 41.158 16.47 41.194 ;
               RECT 16.422 42.358 16.47 42.394 ;
               RECT 16.422 43.558 16.47 43.594 ;
               RECT 16.422 44.758 16.47 44.794 ;
               RECT 16.422 45.958 16.47 45.994 ;
               RECT 16.422 47.158 16.47 47.194 ;
               RECT 16.422 48.358 16.47 48.394 ;
               RECT 16.422 49.2405 16.47 49.2765 ;
               RECT 16.422 51.702 16.47 51.738 ;
               RECT 16.422 53.9235 16.47 53.9595 ;
               RECT 16.422 55.4805 16.47 55.5165 ;
               RECT 16.422 57.478 16.47 57.514 ;
               RECT 16.422 58.678 16.47 58.714 ;
               RECT 16.422 59.878 16.47 59.914 ;
               RECT 16.422 61.078 16.47 61.114 ;
               RECT 16.422 62.278 16.47 62.314 ;
               RECT 16.422 63.478 16.47 63.514 ;
               RECT 16.422 64.678 16.47 64.714 ;
               RECT 16.422 65.878 16.47 65.914 ;
               RECT 16.422 67.078 16.47 67.114 ;
               RECT 16.422 68.278 16.47 68.314 ;
               RECT 16.422 69.478 16.47 69.514 ;
               RECT 16.422 70.678 16.47 70.714 ;
               RECT 16.422 71.878 16.47 71.914 ;
               RECT 16.422 73.078 16.47 73.114 ;
               RECT 16.422 74.278 16.47 74.314 ;
               RECT 16.422 75.478 16.47 75.514 ;
               RECT 16.422 76.678 16.47 76.714 ;
               RECT 16.422 77.878 16.47 77.914 ;
               RECT 16.422 79.078 16.47 79.114 ;
               RECT 16.422 80.278 16.47 80.314 ;
               RECT 16.422 81.478 16.47 81.514 ;
               RECT 16.422 82.678 16.47 82.714 ;
               RECT 16.422 83.878 16.47 83.914 ;
               RECT 16.422 85.078 16.47 85.114 ;
               RECT 16.422 86.278 16.47 86.314 ;
               RECT 16.422 87.478 16.47 87.514 ;
               RECT 16.422 88.678 16.47 88.714 ;
               RECT 16.422 89.878 16.47 89.914 ;
               RECT 16.422 91.078 16.47 91.114 ;
               RECT 16.422 92.278 16.47 92.314 ;
               RECT 16.422 93.478 16.47 93.514 ;
               RECT 16.422 94.678 16.47 94.714 ;
               RECT 16.422 95.878 16.47 95.914 ;
               RECT 16.422 97.078 16.47 97.114 ;
               RECT 16.422 98.278 16.47 98.314 ;
               RECT 16.422 99.478 16.47 99.514 ;
               RECT 16.422 100.678 16.47 100.714 ;
               RECT 16.422 101.878 16.47 101.914 ;
               RECT 16.422 103.078 16.47 103.114 ;
               RECT 16.422 104.278 16.47 104.314 ;
               RECT 16.65 49.7205 16.69 49.7565 ;
               RECT 16.718 1.329 16.772 1.365 ;
               RECT 16.718 2.529 16.772 2.565 ;
               RECT 16.718 3.729 16.772 3.765 ;
               RECT 16.718 4.929 16.772 4.965 ;
               RECT 16.718 6.129 16.772 6.165 ;
               RECT 16.718 7.329 16.772 7.365 ;
               RECT 16.718 8.529 16.772 8.565 ;
               RECT 16.718 9.729 16.772 9.765 ;
               RECT 16.718 10.929 16.772 10.965 ;
               RECT 16.718 12.129 16.772 12.165 ;
               RECT 16.718 13.329 16.772 13.365 ;
               RECT 16.718 14.529 16.772 14.565 ;
               RECT 16.718 15.729 16.772 15.765 ;
               RECT 16.718 16.929 16.772 16.965 ;
               RECT 16.718 18.129 16.772 18.165 ;
               RECT 16.718 19.329 16.772 19.365 ;
               RECT 16.718 20.529 16.772 20.565 ;
               RECT 16.718 21.729 16.772 21.765 ;
               RECT 16.718 22.929 16.772 22.965 ;
               RECT 16.718 24.129 16.772 24.165 ;
               RECT 16.718 25.329 16.772 25.365 ;
               RECT 16.718 26.529 16.772 26.565 ;
               RECT 16.718 27.729 16.772 27.765 ;
               RECT 16.718 28.929 16.772 28.965 ;
               RECT 16.718 30.129 16.772 30.165 ;
               RECT 16.718 31.329 16.772 31.365 ;
               RECT 16.718 32.529 16.772 32.565 ;
               RECT 16.718 33.729 16.772 33.765 ;
               RECT 16.718 34.929 16.772 34.965 ;
               RECT 16.718 36.129 16.772 36.165 ;
               RECT 16.718 37.329 16.772 37.365 ;
               RECT 16.718 38.529 16.772 38.565 ;
               RECT 16.718 39.729 16.772 39.765 ;
               RECT 16.718 40.929 16.772 40.965 ;
               RECT 16.718 42.129 16.772 42.165 ;
               RECT 16.718 43.329 16.772 43.365 ;
               RECT 16.718 44.529 16.772 44.565 ;
               RECT 16.718 45.729 16.772 45.765 ;
               RECT 16.718 46.929 16.772 46.965 ;
               RECT 16.718 48.129 16.772 48.165 ;
               RECT 16.718 49.0005 16.772 49.0365 ;
               RECT 16.718 56.0835 16.772 56.1195 ;
               RECT 16.718 57.249 16.772 57.285 ;
               RECT 16.718 58.449 16.772 58.485 ;
               RECT 16.718 59.649 16.772 59.685 ;
               RECT 16.718 60.849 16.772 60.885 ;
               RECT 16.718 62.049 16.772 62.085 ;
               RECT 16.718 63.249 16.772 63.285 ;
               RECT 16.718 64.449 16.772 64.485 ;
               RECT 16.718 65.649 16.772 65.685 ;
               RECT 16.718 66.849 16.772 66.885 ;
               RECT 16.718 68.049 16.772 68.085 ;
               RECT 16.718 69.249 16.772 69.285 ;
               RECT 16.718 70.449 16.772 70.485 ;
               RECT 16.718 71.649 16.772 71.685 ;
               RECT 16.718 72.849 16.772 72.885 ;
               RECT 16.718 74.049 16.772 74.085 ;
               RECT 16.718 75.249 16.772 75.285 ;
               RECT 16.718 76.449 16.772 76.485 ;
               RECT 16.718 77.649 16.772 77.685 ;
               RECT 16.718 78.849 16.772 78.885 ;
               RECT 16.718 80.049 16.772 80.085 ;
               RECT 16.718 81.249 16.772 81.285 ;
               RECT 16.718 82.449 16.772 82.485 ;
               RECT 16.718 83.649 16.772 83.685 ;
               RECT 16.718 84.849 16.772 84.885 ;
               RECT 16.718 86.049 16.772 86.085 ;
               RECT 16.718 87.249 16.772 87.285 ;
               RECT 16.718 88.449 16.772 88.485 ;
               RECT 16.718 89.649 16.772 89.685 ;
               RECT 16.718 90.849 16.772 90.885 ;
               RECT 16.718 92.049 16.772 92.085 ;
               RECT 16.718 93.249 16.772 93.285 ;
               RECT 16.718 94.449 16.772 94.485 ;
               RECT 16.718 95.649 16.772 95.685 ;
               RECT 16.718 96.849 16.772 96.885 ;
               RECT 16.718 98.049 16.772 98.085 ;
               RECT 16.718 99.249 16.772 99.285 ;
               RECT 16.718 100.449 16.772 100.485 ;
               RECT 16.718 101.649 16.772 101.685 ;
               RECT 16.718 102.849 16.772 102.885 ;
               RECT 16.718 104.049 16.772 104.085 ;
               RECT 16.882 1.558 16.936 1.594 ;
               RECT 16.882 2.758 16.936 2.794 ;
               RECT 16.882 3.958 16.936 3.994 ;
               RECT 16.882 5.158 16.936 5.194 ;
               RECT 16.882 6.358 16.936 6.394 ;
               RECT 16.882 7.558 16.936 7.594 ;
               RECT 16.882 8.758 16.936 8.794 ;
               RECT 16.882 9.958 16.936 9.994 ;
               RECT 16.882 11.158 16.936 11.194 ;
               RECT 16.882 12.358 16.936 12.394 ;
               RECT 16.882 13.558 16.936 13.594 ;
               RECT 16.882 14.758 16.936 14.794 ;
               RECT 16.882 15.958 16.936 15.994 ;
               RECT 16.882 17.158 16.936 17.194 ;
               RECT 16.882 18.358 16.936 18.394 ;
               RECT 16.882 19.558 16.936 19.594 ;
               RECT 16.882 20.758 16.936 20.794 ;
               RECT 16.882 21.958 16.936 21.994 ;
               RECT 16.882 23.158 16.936 23.194 ;
               RECT 16.882 24.358 16.936 24.394 ;
               RECT 16.882 25.558 16.936 25.594 ;
               RECT 16.882 26.758 16.936 26.794 ;
               RECT 16.882 27.958 16.936 27.994 ;
               RECT 16.882 29.158 16.936 29.194 ;
               RECT 16.882 30.358 16.936 30.394 ;
               RECT 16.882 31.558 16.936 31.594 ;
               RECT 16.882 32.758 16.936 32.794 ;
               RECT 16.882 33.958 16.936 33.994 ;
               RECT 16.882 35.158 16.936 35.194 ;
               RECT 16.882 36.358 16.936 36.394 ;
               RECT 16.882 37.558 16.936 37.594 ;
               RECT 16.882 38.758 16.936 38.794 ;
               RECT 16.882 39.958 16.936 39.994 ;
               RECT 16.882 41.158 16.936 41.194 ;
               RECT 16.882 42.358 16.936 42.394 ;
               RECT 16.882 43.558 16.936 43.594 ;
               RECT 16.882 44.758 16.936 44.794 ;
               RECT 16.882 45.958 16.936 45.994 ;
               RECT 16.882 47.158 16.936 47.194 ;
               RECT 16.882 48.358 16.936 48.394 ;
               RECT 16.882 49.0005 16.936 49.0365 ;
               RECT 16.882 56.0835 16.936 56.1195 ;
               RECT 16.882 57.478 16.936 57.514 ;
               RECT 16.882 58.678 16.936 58.714 ;
               RECT 16.882 59.878 16.936 59.914 ;
               RECT 16.882 61.078 16.936 61.114 ;
               RECT 16.882 62.278 16.936 62.314 ;
               RECT 16.882 63.478 16.936 63.514 ;
               RECT 16.882 64.678 16.936 64.714 ;
               RECT 16.882 65.878 16.936 65.914 ;
               RECT 16.882 67.078 16.936 67.114 ;
               RECT 16.882 68.278 16.936 68.314 ;
               RECT 16.882 69.478 16.936 69.514 ;
               RECT 16.882 70.678 16.936 70.714 ;
               RECT 16.882 71.878 16.936 71.914 ;
               RECT 16.882 73.078 16.936 73.114 ;
               RECT 16.882 74.278 16.936 74.314 ;
               RECT 16.882 75.478 16.936 75.514 ;
               RECT 16.882 76.678 16.936 76.714 ;
               RECT 16.882 77.878 16.936 77.914 ;
               RECT 16.882 79.078 16.936 79.114 ;
               RECT 16.882 80.278 16.936 80.314 ;
               RECT 16.882 81.478 16.936 81.514 ;
               RECT 16.882 82.678 16.936 82.714 ;
               RECT 16.882 83.878 16.936 83.914 ;
               RECT 16.882 85.078 16.936 85.114 ;
               RECT 16.882 86.278 16.936 86.314 ;
               RECT 16.882 87.478 16.936 87.514 ;
               RECT 16.882 88.678 16.936 88.714 ;
               RECT 16.882 89.878 16.936 89.914 ;
               RECT 16.882 91.078 16.936 91.114 ;
               RECT 16.882 92.278 16.936 92.314 ;
               RECT 16.882 93.478 16.936 93.514 ;
               RECT 16.882 94.678 16.936 94.714 ;
               RECT 16.882 95.878 16.936 95.914 ;
               RECT 16.882 97.078 16.936 97.114 ;
               RECT 16.882 98.278 16.936 98.314 ;
               RECT 16.882 99.478 16.936 99.514 ;
               RECT 16.882 100.678 16.936 100.714 ;
               RECT 16.882 101.878 16.936 101.914 ;
               RECT 16.882 103.078 16.936 103.114 ;
               RECT 16.882 104.278 16.936 104.314 ;
               RECT 17.136 49.422 17.176 49.458 ;
               RECT 17.136 49.542 17.176 49.578 ;
               RECT 17.548 1.035 17.588 1.071 ;
               RECT 17.548 2.235 17.588 2.271 ;
               RECT 17.548 3.435 17.588 3.471 ;
               RECT 17.548 4.635 17.588 4.671 ;
               RECT 17.548 5.835 17.588 5.871 ;
               RECT 17.548 7.035 17.588 7.071 ;
               RECT 17.548 8.235 17.588 8.271 ;
               RECT 17.548 9.435 17.588 9.471 ;
               RECT 17.548 10.635 17.588 10.671 ;
               RECT 17.548 11.835 17.588 11.871 ;
               RECT 17.548 13.035 17.588 13.071 ;
               RECT 17.548 14.235 17.588 14.271 ;
               RECT 17.548 15.435 17.588 15.471 ;
               RECT 17.548 16.635 17.588 16.671 ;
               RECT 17.548 17.835 17.588 17.871 ;
               RECT 17.548 19.035 17.588 19.071 ;
               RECT 17.548 20.235 17.588 20.271 ;
               RECT 17.548 21.435 17.588 21.471 ;
               RECT 17.548 22.635 17.588 22.671 ;
               RECT 17.548 23.835 17.588 23.871 ;
               RECT 17.548 25.035 17.588 25.071 ;
               RECT 17.548 26.235 17.588 26.271 ;
               RECT 17.548 27.435 17.588 27.471 ;
               RECT 17.548 28.635 17.588 28.671 ;
               RECT 17.548 29.835 17.588 29.871 ;
               RECT 17.548 31.035 17.588 31.071 ;
               RECT 17.548 32.235 17.588 32.271 ;
               RECT 17.548 33.435 17.588 33.471 ;
               RECT 17.548 34.635 17.588 34.671 ;
               RECT 17.548 35.835 17.588 35.871 ;
               RECT 17.548 37.035 17.588 37.071 ;
               RECT 17.548 38.235 17.588 38.271 ;
               RECT 17.548 39.435 17.588 39.471 ;
               RECT 17.548 40.635 17.588 40.671 ;
               RECT 17.548 41.835 17.588 41.871 ;
               RECT 17.548 43.035 17.588 43.071 ;
               RECT 17.548 44.235 17.588 44.271 ;
               RECT 17.548 45.435 17.588 45.471 ;
               RECT 17.548 46.635 17.588 46.671 ;
               RECT 17.548 47.835 17.588 47.871 ;
               RECT 17.548 55.782 17.588 55.818 ;
               RECT 17.548 56.955 17.588 56.991 ;
               RECT 17.548 58.155 17.588 58.191 ;
               RECT 17.548 59.355 17.588 59.391 ;
               RECT 17.548 60.555 17.588 60.591 ;
               RECT 17.548 61.755 17.588 61.791 ;
               RECT 17.548 62.955 17.588 62.991 ;
               RECT 17.548 64.155 17.588 64.191 ;
               RECT 17.548 65.355 17.588 65.391 ;
               RECT 17.548 66.555 17.588 66.591 ;
               RECT 17.548 67.755 17.588 67.791 ;
               RECT 17.548 68.955 17.588 68.991 ;
               RECT 17.548 70.155 17.588 70.191 ;
               RECT 17.548 71.355 17.588 71.391 ;
               RECT 17.548 72.555 17.588 72.591 ;
               RECT 17.548 73.755 17.588 73.791 ;
               RECT 17.548 74.955 17.588 74.991 ;
               RECT 17.548 76.155 17.588 76.191 ;
               RECT 17.548 77.355 17.588 77.391 ;
               RECT 17.548 78.555 17.588 78.591 ;
               RECT 17.548 79.755 17.588 79.791 ;
               RECT 17.548 80.955 17.588 80.991 ;
               RECT 17.548 82.155 17.588 82.191 ;
               RECT 17.548 83.355 17.588 83.391 ;
               RECT 17.548 84.555 17.588 84.591 ;
               RECT 17.548 85.755 17.588 85.791 ;
               RECT 17.548 86.955 17.588 86.991 ;
               RECT 17.548 88.155 17.588 88.191 ;
               RECT 17.548 89.355 17.588 89.391 ;
               RECT 17.548 90.555 17.588 90.591 ;
               RECT 17.548 91.755 17.588 91.791 ;
               RECT 17.548 92.955 17.588 92.991 ;
               RECT 17.548 94.155 17.588 94.191 ;
               RECT 17.548 95.355 17.588 95.391 ;
               RECT 17.548 96.555 17.588 96.591 ;
               RECT 17.548 97.755 17.588 97.791 ;
               RECT 17.548 98.955 17.588 98.991 ;
               RECT 17.548 100.155 17.588 100.191 ;
               RECT 17.548 101.355 17.588 101.391 ;
               RECT 17.548 102.555 17.588 102.591 ;
               RECT 17.548 103.755 17.588 103.791 ;
               RECT 17.616 1.035 17.656 1.071 ;
               RECT 17.616 2.235 17.656 2.271 ;
               RECT 17.616 3.435 17.656 3.471 ;
               RECT 17.616 4.635 17.656 4.671 ;
               RECT 17.616 5.835 17.656 5.871 ;
               RECT 17.616 7.035 17.656 7.071 ;
               RECT 17.616 8.235 17.656 8.271 ;
               RECT 17.616 9.435 17.656 9.471 ;
               RECT 17.616 10.635 17.656 10.671 ;
               RECT 17.616 11.835 17.656 11.871 ;
               RECT 17.616 13.035 17.656 13.071 ;
               RECT 17.616 14.235 17.656 14.271 ;
               RECT 17.616 15.435 17.656 15.471 ;
               RECT 17.616 16.635 17.656 16.671 ;
               RECT 17.616 17.835 17.656 17.871 ;
               RECT 17.616 19.035 17.656 19.071 ;
               RECT 17.616 20.235 17.656 20.271 ;
               RECT 17.616 21.435 17.656 21.471 ;
               RECT 17.616 22.635 17.656 22.671 ;
               RECT 17.616 23.835 17.656 23.871 ;
               RECT 17.616 25.035 17.656 25.071 ;
               RECT 17.616 26.235 17.656 26.271 ;
               RECT 17.616 27.435 17.656 27.471 ;
               RECT 17.616 28.635 17.656 28.671 ;
               RECT 17.616 29.835 17.656 29.871 ;
               RECT 17.616 31.035 17.656 31.071 ;
               RECT 17.616 32.235 17.656 32.271 ;
               RECT 17.616 33.435 17.656 33.471 ;
               RECT 17.616 34.635 17.656 34.671 ;
               RECT 17.616 35.835 17.656 35.871 ;
               RECT 17.616 37.035 17.656 37.071 ;
               RECT 17.616 38.235 17.656 38.271 ;
               RECT 17.616 39.435 17.656 39.471 ;
               RECT 17.616 40.635 17.656 40.671 ;
               RECT 17.616 41.835 17.656 41.871 ;
               RECT 17.616 43.035 17.656 43.071 ;
               RECT 17.616 44.235 17.656 44.271 ;
               RECT 17.616 45.435 17.656 45.471 ;
               RECT 17.616 46.635 17.656 46.671 ;
               RECT 17.616 47.835 17.656 47.871 ;
               RECT 17.616 55.782 17.656 55.818 ;
               RECT 17.616 56.955 17.656 56.991 ;
               RECT 17.616 58.155 17.656 58.191 ;
               RECT 17.616 59.355 17.656 59.391 ;
               RECT 17.616 60.555 17.656 60.591 ;
               RECT 17.616 61.755 17.656 61.791 ;
               RECT 17.616 62.955 17.656 62.991 ;
               RECT 17.616 64.155 17.656 64.191 ;
               RECT 17.616 65.355 17.656 65.391 ;
               RECT 17.616 66.555 17.656 66.591 ;
               RECT 17.616 67.755 17.656 67.791 ;
               RECT 17.616 68.955 17.656 68.991 ;
               RECT 17.616 70.155 17.656 70.191 ;
               RECT 17.616 71.355 17.656 71.391 ;
               RECT 17.616 72.555 17.656 72.591 ;
               RECT 17.616 73.755 17.656 73.791 ;
               RECT 17.616 74.955 17.656 74.991 ;
               RECT 17.616 76.155 17.656 76.191 ;
               RECT 17.616 77.355 17.656 77.391 ;
               RECT 17.616 78.555 17.656 78.591 ;
               RECT 17.616 79.755 17.656 79.791 ;
               RECT 17.616 80.955 17.656 80.991 ;
               RECT 17.616 82.155 17.656 82.191 ;
               RECT 17.616 83.355 17.656 83.391 ;
               RECT 17.616 84.555 17.656 84.591 ;
               RECT 17.616 85.755 17.656 85.791 ;
               RECT 17.616 86.955 17.656 86.991 ;
               RECT 17.616 88.155 17.656 88.191 ;
               RECT 17.616 89.355 17.656 89.391 ;
               RECT 17.616 90.555 17.656 90.591 ;
               RECT 17.616 91.755 17.656 91.791 ;
               RECT 17.616 92.955 17.656 92.991 ;
               RECT 17.616 94.155 17.656 94.191 ;
               RECT 17.616 95.355 17.656 95.391 ;
               RECT 17.616 96.555 17.656 96.591 ;
               RECT 17.616 97.755 17.656 97.791 ;
               RECT 17.616 98.955 17.656 98.991 ;
               RECT 17.616 100.155 17.656 100.191 ;
               RECT 17.616 101.355 17.656 101.391 ;
               RECT 17.616 102.555 17.656 102.591 ;
               RECT 17.616 103.755 17.656 103.791 ;
               RECT 17.944 49.302 17.984 49.338 ;
               RECT 17.944 49.422 17.984 49.458 ;
               RECT 17.944 49.7205 17.984 49.7565 ;
               RECT 17.944 51.222 17.984 51.258 ;
               RECT 17.944 51.342 17.984 51.378 ;
               RECT 17.944 51.822 17.984 51.858 ;
               RECT 18.012 1.329 18.052 1.365 ;
               RECT 18.012 2.529 18.052 2.565 ;
               RECT 18.012 3.729 18.052 3.765 ;
               RECT 18.012 4.929 18.052 4.965 ;
               RECT 18.012 6.129 18.052 6.165 ;
               RECT 18.012 7.329 18.052 7.365 ;
               RECT 18.012 8.529 18.052 8.565 ;
               RECT 18.012 9.729 18.052 9.765 ;
               RECT 18.012 10.929 18.052 10.965 ;
               RECT 18.012 12.129 18.052 12.165 ;
               RECT 18.012 13.329 18.052 13.365 ;
               RECT 18.012 14.529 18.052 14.565 ;
               RECT 18.012 15.729 18.052 15.765 ;
               RECT 18.012 16.929 18.052 16.965 ;
               RECT 18.012 18.129 18.052 18.165 ;
               RECT 18.012 19.329 18.052 19.365 ;
               RECT 18.012 20.529 18.052 20.565 ;
               RECT 18.012 21.729 18.052 21.765 ;
               RECT 18.012 22.929 18.052 22.965 ;
               RECT 18.012 24.129 18.052 24.165 ;
               RECT 18.012 25.329 18.052 25.365 ;
               RECT 18.012 26.529 18.052 26.565 ;
               RECT 18.012 27.729 18.052 27.765 ;
               RECT 18.012 28.929 18.052 28.965 ;
               RECT 18.012 30.129 18.052 30.165 ;
               RECT 18.012 31.329 18.052 31.365 ;
               RECT 18.012 32.529 18.052 32.565 ;
               RECT 18.012 33.729 18.052 33.765 ;
               RECT 18.012 34.929 18.052 34.965 ;
               RECT 18.012 36.129 18.052 36.165 ;
               RECT 18.012 37.329 18.052 37.365 ;
               RECT 18.012 38.529 18.052 38.565 ;
               RECT 18.012 39.729 18.052 39.765 ;
               RECT 18.012 40.929 18.052 40.965 ;
               RECT 18.012 42.129 18.052 42.165 ;
               RECT 18.012 43.329 18.052 43.365 ;
               RECT 18.012 44.529 18.052 44.565 ;
               RECT 18.012 45.729 18.052 45.765 ;
               RECT 18.012 46.929 18.052 46.965 ;
               RECT 18.012 48.129 18.052 48.165 ;
               RECT 18.012 55.782 18.052 55.818 ;
               RECT 18.012 57.249 18.052 57.285 ;
               RECT 18.012 58.449 18.052 58.485 ;
               RECT 18.012 59.649 18.052 59.685 ;
               RECT 18.012 60.849 18.052 60.885 ;
               RECT 18.012 62.049 18.052 62.085 ;
               RECT 18.012 63.249 18.052 63.285 ;
               RECT 18.012 64.449 18.052 64.485 ;
               RECT 18.012 65.649 18.052 65.685 ;
               RECT 18.012 66.849 18.052 66.885 ;
               RECT 18.012 68.049 18.052 68.085 ;
               RECT 18.012 69.249 18.052 69.285 ;
               RECT 18.012 70.449 18.052 70.485 ;
               RECT 18.012 71.649 18.052 71.685 ;
               RECT 18.012 72.849 18.052 72.885 ;
               RECT 18.012 74.049 18.052 74.085 ;
               RECT 18.012 75.249 18.052 75.285 ;
               RECT 18.012 76.449 18.052 76.485 ;
               RECT 18.012 77.649 18.052 77.685 ;
               RECT 18.012 78.849 18.052 78.885 ;
               RECT 18.012 80.049 18.052 80.085 ;
               RECT 18.012 81.249 18.052 81.285 ;
               RECT 18.012 82.449 18.052 82.485 ;
               RECT 18.012 83.649 18.052 83.685 ;
               RECT 18.012 84.849 18.052 84.885 ;
               RECT 18.012 86.049 18.052 86.085 ;
               RECT 18.012 87.249 18.052 87.285 ;
               RECT 18.012 88.449 18.052 88.485 ;
               RECT 18.012 89.649 18.052 89.685 ;
               RECT 18.012 90.849 18.052 90.885 ;
               RECT 18.012 92.049 18.052 92.085 ;
               RECT 18.012 93.249 18.052 93.285 ;
               RECT 18.012 94.449 18.052 94.485 ;
               RECT 18.012 95.649 18.052 95.685 ;
               RECT 18.012 96.849 18.052 96.885 ;
               RECT 18.012 98.049 18.052 98.085 ;
               RECT 18.012 99.249 18.052 99.285 ;
               RECT 18.012 100.449 18.052 100.485 ;
               RECT 18.012 101.649 18.052 101.685 ;
               RECT 18.012 102.849 18.052 102.885 ;
               RECT 18.012 104.049 18.052 104.085 ;
               RECT 18.08 1.329 18.12 1.365 ;
               RECT 18.08 2.529 18.12 2.565 ;
               RECT 18.08 3.729 18.12 3.765 ;
               RECT 18.08 4.929 18.12 4.965 ;
               RECT 18.08 6.129 18.12 6.165 ;
               RECT 18.08 7.329 18.12 7.365 ;
               RECT 18.08 8.529 18.12 8.565 ;
               RECT 18.08 9.729 18.12 9.765 ;
               RECT 18.08 10.929 18.12 10.965 ;
               RECT 18.08 12.129 18.12 12.165 ;
               RECT 18.08 13.329 18.12 13.365 ;
               RECT 18.08 14.529 18.12 14.565 ;
               RECT 18.08 15.729 18.12 15.765 ;
               RECT 18.08 16.929 18.12 16.965 ;
               RECT 18.08 18.129 18.12 18.165 ;
               RECT 18.08 19.329 18.12 19.365 ;
               RECT 18.08 20.529 18.12 20.565 ;
               RECT 18.08 21.729 18.12 21.765 ;
               RECT 18.08 22.929 18.12 22.965 ;
               RECT 18.08 24.129 18.12 24.165 ;
               RECT 18.08 25.329 18.12 25.365 ;
               RECT 18.08 26.529 18.12 26.565 ;
               RECT 18.08 27.729 18.12 27.765 ;
               RECT 18.08 28.929 18.12 28.965 ;
               RECT 18.08 30.129 18.12 30.165 ;
               RECT 18.08 31.329 18.12 31.365 ;
               RECT 18.08 32.529 18.12 32.565 ;
               RECT 18.08 33.729 18.12 33.765 ;
               RECT 18.08 34.929 18.12 34.965 ;
               RECT 18.08 36.129 18.12 36.165 ;
               RECT 18.08 37.329 18.12 37.365 ;
               RECT 18.08 38.529 18.12 38.565 ;
               RECT 18.08 39.729 18.12 39.765 ;
               RECT 18.08 40.929 18.12 40.965 ;
               RECT 18.08 42.129 18.12 42.165 ;
               RECT 18.08 43.329 18.12 43.365 ;
               RECT 18.08 44.529 18.12 44.565 ;
               RECT 18.08 45.729 18.12 45.765 ;
               RECT 18.08 46.929 18.12 46.965 ;
               RECT 18.08 48.129 18.12 48.165 ;
               RECT 18.08 55.782 18.12 55.818 ;
               RECT 18.08 57.249 18.12 57.285 ;
               RECT 18.08 58.449 18.12 58.485 ;
               RECT 18.08 59.649 18.12 59.685 ;
               RECT 18.08 60.849 18.12 60.885 ;
               RECT 18.08 62.049 18.12 62.085 ;
               RECT 18.08 63.249 18.12 63.285 ;
               RECT 18.08 64.449 18.12 64.485 ;
               RECT 18.08 65.649 18.12 65.685 ;
               RECT 18.08 66.849 18.12 66.885 ;
               RECT 18.08 68.049 18.12 68.085 ;
               RECT 18.08 69.249 18.12 69.285 ;
               RECT 18.08 70.449 18.12 70.485 ;
               RECT 18.08 71.649 18.12 71.685 ;
               RECT 18.08 72.849 18.12 72.885 ;
               RECT 18.08 74.049 18.12 74.085 ;
               RECT 18.08 75.249 18.12 75.285 ;
               RECT 18.08 76.449 18.12 76.485 ;
               RECT 18.08 77.649 18.12 77.685 ;
               RECT 18.08 78.849 18.12 78.885 ;
               RECT 18.08 80.049 18.12 80.085 ;
               RECT 18.08 81.249 18.12 81.285 ;
               RECT 18.08 82.449 18.12 82.485 ;
               RECT 18.08 83.649 18.12 83.685 ;
               RECT 18.08 84.849 18.12 84.885 ;
               RECT 18.08 86.049 18.12 86.085 ;
               RECT 18.08 87.249 18.12 87.285 ;
               RECT 18.08 88.449 18.12 88.485 ;
               RECT 18.08 89.649 18.12 89.685 ;
               RECT 18.08 90.849 18.12 90.885 ;
               RECT 18.08 92.049 18.12 92.085 ;
               RECT 18.08 93.249 18.12 93.285 ;
               RECT 18.08 94.449 18.12 94.485 ;
               RECT 18.08 95.649 18.12 95.685 ;
               RECT 18.08 96.849 18.12 96.885 ;
               RECT 18.08 98.049 18.12 98.085 ;
               RECT 18.08 99.249 18.12 99.285 ;
               RECT 18.08 100.449 18.12 100.485 ;
               RECT 18.08 101.649 18.12 101.685 ;
               RECT 18.08 102.849 18.12 102.885 ;
               RECT 18.08 104.049 18.12 104.085 ;
               RECT 18.492 49.302 18.536 49.338 ;
               RECT 18.764 1.1875 18.836 1.2125 ;
               RECT 18.764 1.3345 18.836 1.3595 ;
               RECT 18.764 3.5875 18.836 3.6125 ;
               RECT 18.764 3.7345 18.836 3.7595 ;
               RECT 18.764 5.9875 18.836 6.0125 ;
               RECT 18.764 6.1345 18.836 6.1595 ;
               RECT 18.764 8.3875 18.836 8.4125 ;
               RECT 18.764 8.5345 18.836 8.5595 ;
               RECT 18.764 10.7875 18.836 10.8125 ;
               RECT 18.764 10.9345 18.836 10.9595 ;
               RECT 18.764 13.1875 18.836 13.2125 ;
               RECT 18.764 13.3345 18.836 13.3595 ;
               RECT 18.764 15.5875 18.836 15.6125 ;
               RECT 18.764 15.7345 18.836 15.7595 ;
               RECT 18.764 17.9875 18.836 18.0125 ;
               RECT 18.764 18.1345 18.836 18.1595 ;
               RECT 18.764 20.3875 18.836 20.4125 ;
               RECT 18.764 20.5345 18.836 20.5595 ;
               RECT 18.764 22.7875 18.836 22.8125 ;
               RECT 18.764 22.9345 18.836 22.9595 ;
               RECT 18.764 25.1875 18.836 25.2125 ;
               RECT 18.764 25.3345 18.836 25.3595 ;
               RECT 18.764 27.5875 18.836 27.6125 ;
               RECT 18.764 27.7345 18.836 27.7595 ;
               RECT 18.764 29.9875 18.836 30.0125 ;
               RECT 18.764 30.1345 18.836 30.1595 ;
               RECT 18.764 32.3875 18.836 32.4125 ;
               RECT 18.764 32.5345 18.836 32.5595 ;
               RECT 18.764 34.7875 18.836 34.8125 ;
               RECT 18.764 34.9345 18.836 34.9595 ;
               RECT 18.764 37.1875 18.836 37.2125 ;
               RECT 18.764 37.3345 18.836 37.3595 ;
               RECT 18.764 39.5875 18.836 39.6125 ;
               RECT 18.764 39.7345 18.836 39.7595 ;
               RECT 18.764 41.9875 18.836 42.0125 ;
               RECT 18.764 42.1345 18.836 42.1595 ;
               RECT 18.764 44.3875 18.836 44.4125 ;
               RECT 18.764 44.5345 18.836 44.5595 ;
               RECT 18.764 46.7875 18.836 46.8125 ;
               RECT 18.764 46.9345 18.836 46.9595 ;
               RECT 18.764 57.1075 18.836 57.1325 ;
               RECT 18.764 57.2545 18.836 57.2795 ;
               RECT 18.764 59.5075 18.836 59.5325 ;
               RECT 18.764 59.6545 18.836 59.6795 ;
               RECT 18.764 61.9075 18.836 61.9325 ;
               RECT 18.764 62.0545 18.836 62.0795 ;
               RECT 18.764 64.3075 18.836 64.3325 ;
               RECT 18.764 64.4545 18.836 64.4795 ;
               RECT 18.764 66.7075 18.836 66.7325 ;
               RECT 18.764 66.8545 18.836 66.8795 ;
               RECT 18.764 69.1075 18.836 69.1325 ;
               RECT 18.764 69.2545 18.836 69.2795 ;
               RECT 18.764 71.5075 18.836 71.5325 ;
               RECT 18.764 71.6545 18.836 71.6795 ;
               RECT 18.764 73.9075 18.836 73.9325 ;
               RECT 18.764 74.0545 18.836 74.0795 ;
               RECT 18.764 76.3075 18.836 76.3325 ;
               RECT 18.764 76.4545 18.836 76.4795 ;
               RECT 18.764 78.7075 18.836 78.7325 ;
               RECT 18.764 78.8545 18.836 78.8795 ;
               RECT 18.764 81.1075 18.836 81.1325 ;
               RECT 18.764 81.2545 18.836 81.2795 ;
               RECT 18.764 83.5075 18.836 83.5325 ;
               RECT 18.764 83.6545 18.836 83.6795 ;
               RECT 18.764 85.9075 18.836 85.9325 ;
               RECT 18.764 86.0545 18.836 86.0795 ;
               RECT 18.764 88.3075 18.836 88.3325 ;
               RECT 18.764 88.4545 18.836 88.4795 ;
               RECT 18.764 90.7075 18.836 90.7325 ;
               RECT 18.764 90.8545 18.836 90.8795 ;
               RECT 18.764 93.1075 18.836 93.1325 ;
               RECT 18.764 93.2545 18.836 93.2795 ;
               RECT 18.764 95.5075 18.836 95.5325 ;
               RECT 18.764 95.6545 18.836 95.6795 ;
               RECT 18.764 97.9075 18.836 97.9325 ;
               RECT 18.764 98.0545 18.836 98.0795 ;
               RECT 18.764 100.3075 18.836 100.3325 ;
               RECT 18.764 100.4545 18.836 100.4795 ;
               RECT 18.764 102.7075 18.836 102.7325 ;
               RECT 18.764 102.8545 18.836 102.8795 ;
               RECT 19.53 1.558 19.578 1.594 ;
               RECT 19.53 2.758 19.578 2.794 ;
               RECT 19.53 3.958 19.578 3.994 ;
               RECT 19.53 5.158 19.578 5.194 ;
               RECT 19.53 6.358 19.578 6.394 ;
               RECT 19.53 7.558 19.578 7.594 ;
               RECT 19.53 8.758 19.578 8.794 ;
               RECT 19.53 9.958 19.578 9.994 ;
               RECT 19.53 11.158 19.578 11.194 ;
               RECT 19.53 12.358 19.578 12.394 ;
               RECT 19.53 13.558 19.578 13.594 ;
               RECT 19.53 14.758 19.578 14.794 ;
               RECT 19.53 15.958 19.578 15.994 ;
               RECT 19.53 17.158 19.578 17.194 ;
               RECT 19.53 18.358 19.578 18.394 ;
               RECT 19.53 19.558 19.578 19.594 ;
               RECT 19.53 20.758 19.578 20.794 ;
               RECT 19.53 21.958 19.578 21.994 ;
               RECT 19.53 23.158 19.578 23.194 ;
               RECT 19.53 24.358 19.578 24.394 ;
               RECT 19.53 25.558 19.578 25.594 ;
               RECT 19.53 26.758 19.578 26.794 ;
               RECT 19.53 27.958 19.578 27.994 ;
               RECT 19.53 29.158 19.578 29.194 ;
               RECT 19.53 30.358 19.578 30.394 ;
               RECT 19.53 31.558 19.578 31.594 ;
               RECT 19.53 32.758 19.578 32.794 ;
               RECT 19.53 33.958 19.578 33.994 ;
               RECT 19.53 35.158 19.578 35.194 ;
               RECT 19.53 36.358 19.578 36.394 ;
               RECT 19.53 37.558 19.578 37.594 ;
               RECT 19.53 38.758 19.578 38.794 ;
               RECT 19.53 39.958 19.578 39.994 ;
               RECT 19.53 41.158 19.578 41.194 ;
               RECT 19.53 42.358 19.578 42.394 ;
               RECT 19.53 43.558 19.578 43.594 ;
               RECT 19.53 44.758 19.578 44.794 ;
               RECT 19.53 45.958 19.578 45.994 ;
               RECT 19.53 47.158 19.578 47.194 ;
               RECT 19.53 48.358 19.578 48.394 ;
               RECT 19.53 49.1235 19.578 49.1595 ;
               RECT 19.53 55.4805 19.578 55.5165 ;
               RECT 19.53 57.478 19.578 57.514 ;
               RECT 19.53 58.678 19.578 58.714 ;
               RECT 19.53 59.878 19.578 59.914 ;
               RECT 19.53 61.078 19.578 61.114 ;
               RECT 19.53 62.278 19.578 62.314 ;
               RECT 19.53 63.478 19.578 63.514 ;
               RECT 19.53 64.678 19.578 64.714 ;
               RECT 19.53 65.878 19.578 65.914 ;
               RECT 19.53 67.078 19.578 67.114 ;
               RECT 19.53 68.278 19.578 68.314 ;
               RECT 19.53 69.478 19.578 69.514 ;
               RECT 19.53 70.678 19.578 70.714 ;
               RECT 19.53 71.878 19.578 71.914 ;
               RECT 19.53 73.078 19.578 73.114 ;
               RECT 19.53 74.278 19.578 74.314 ;
               RECT 19.53 75.478 19.578 75.514 ;
               RECT 19.53 76.678 19.578 76.714 ;
               RECT 19.53 77.878 19.578 77.914 ;
               RECT 19.53 79.078 19.578 79.114 ;
               RECT 19.53 80.278 19.578 80.314 ;
               RECT 19.53 81.478 19.578 81.514 ;
               RECT 19.53 82.678 19.578 82.714 ;
               RECT 19.53 83.878 19.578 83.914 ;
               RECT 19.53 85.078 19.578 85.114 ;
               RECT 19.53 86.278 19.578 86.314 ;
               RECT 19.53 87.478 19.578 87.514 ;
               RECT 19.53 88.678 19.578 88.714 ;
               RECT 19.53 89.878 19.578 89.914 ;
               RECT 19.53 91.078 19.578 91.114 ;
               RECT 19.53 92.278 19.578 92.314 ;
               RECT 19.53 93.478 19.578 93.514 ;
               RECT 19.53 94.678 19.578 94.714 ;
               RECT 19.53 95.878 19.578 95.914 ;
               RECT 19.53 97.078 19.578 97.114 ;
               RECT 19.53 98.278 19.578 98.314 ;
               RECT 19.53 99.478 19.578 99.514 ;
               RECT 19.53 100.678 19.578 100.714 ;
               RECT 19.53 101.878 19.578 101.914 ;
               RECT 19.53 103.078 19.578 103.114 ;
               RECT 19.53 104.278 19.578 104.314 ;
               RECT 19.606 1.329 19.654 1.365 ;
               RECT 19.606 2.529 19.654 2.565 ;
               RECT 19.606 3.729 19.654 3.765 ;
               RECT 19.606 4.929 19.654 4.965 ;
               RECT 19.606 6.129 19.654 6.165 ;
               RECT 19.606 7.329 19.654 7.365 ;
               RECT 19.606 8.529 19.654 8.565 ;
               RECT 19.606 9.729 19.654 9.765 ;
               RECT 19.606 10.929 19.654 10.965 ;
               RECT 19.606 12.129 19.654 12.165 ;
               RECT 19.606 13.329 19.654 13.365 ;
               RECT 19.606 14.529 19.654 14.565 ;
               RECT 19.606 15.729 19.654 15.765 ;
               RECT 19.606 16.929 19.654 16.965 ;
               RECT 19.606 18.129 19.654 18.165 ;
               RECT 19.606 19.329 19.654 19.365 ;
               RECT 19.606 20.529 19.654 20.565 ;
               RECT 19.606 21.729 19.654 21.765 ;
               RECT 19.606 22.929 19.654 22.965 ;
               RECT 19.606 24.129 19.654 24.165 ;
               RECT 19.606 25.329 19.654 25.365 ;
               RECT 19.606 26.529 19.654 26.565 ;
               RECT 19.606 27.729 19.654 27.765 ;
               RECT 19.606 28.929 19.654 28.965 ;
               RECT 19.606 30.129 19.654 30.165 ;
               RECT 19.606 31.329 19.654 31.365 ;
               RECT 19.606 32.529 19.654 32.565 ;
               RECT 19.606 33.729 19.654 33.765 ;
               RECT 19.606 34.929 19.654 34.965 ;
               RECT 19.606 36.129 19.654 36.165 ;
               RECT 19.606 37.329 19.654 37.365 ;
               RECT 19.606 38.529 19.654 38.565 ;
               RECT 19.606 39.729 19.654 39.765 ;
               RECT 19.606 40.929 19.654 40.965 ;
               RECT 19.606 42.129 19.654 42.165 ;
               RECT 19.606 43.329 19.654 43.365 ;
               RECT 19.606 44.529 19.654 44.565 ;
               RECT 19.606 45.729 19.654 45.765 ;
               RECT 19.606 46.929 19.654 46.965 ;
               RECT 19.606 48.129 19.654 48.165 ;
               RECT 19.606 49.542 19.654 49.578 ;
               RECT 19.606 50.022 19.654 50.058 ;
               RECT 19.606 52.6005 19.654 52.6365 ;
               RECT 19.606 55.062 19.654 55.098 ;
               RECT 19.606 55.782 19.654 55.818 ;
               RECT 19.606 57.249 19.654 57.285 ;
               RECT 19.606 58.449 19.654 58.485 ;
               RECT 19.606 59.649 19.654 59.685 ;
               RECT 19.606 60.849 19.654 60.885 ;
               RECT 19.606 62.049 19.654 62.085 ;
               RECT 19.606 63.249 19.654 63.285 ;
               RECT 19.606 64.449 19.654 64.485 ;
               RECT 19.606 65.649 19.654 65.685 ;
               RECT 19.606 66.849 19.654 66.885 ;
               RECT 19.606 68.049 19.654 68.085 ;
               RECT 19.606 69.249 19.654 69.285 ;
               RECT 19.606 70.449 19.654 70.485 ;
               RECT 19.606 71.649 19.654 71.685 ;
               RECT 19.606 72.849 19.654 72.885 ;
               RECT 19.606 74.049 19.654 74.085 ;
               RECT 19.606 75.249 19.654 75.285 ;
               RECT 19.606 76.449 19.654 76.485 ;
               RECT 19.606 77.649 19.654 77.685 ;
               RECT 19.606 78.849 19.654 78.885 ;
               RECT 19.606 80.049 19.654 80.085 ;
               RECT 19.606 81.249 19.654 81.285 ;
               RECT 19.606 82.449 19.654 82.485 ;
               RECT 19.606 83.649 19.654 83.685 ;
               RECT 19.606 84.849 19.654 84.885 ;
               RECT 19.606 86.049 19.654 86.085 ;
               RECT 19.606 87.249 19.654 87.285 ;
               RECT 19.606 88.449 19.654 88.485 ;
               RECT 19.606 89.649 19.654 89.685 ;
               RECT 19.606 90.849 19.654 90.885 ;
               RECT 19.606 92.049 19.654 92.085 ;
               RECT 19.606 93.249 19.654 93.285 ;
               RECT 19.606 94.449 19.654 94.485 ;
               RECT 19.606 95.649 19.654 95.685 ;
               RECT 19.606 96.849 19.654 96.885 ;
               RECT 19.606 98.049 19.654 98.085 ;
               RECT 19.606 99.249 19.654 99.285 ;
               RECT 19.606 100.449 19.654 100.485 ;
               RECT 19.606 101.649 19.654 101.685 ;
               RECT 19.606 102.849 19.654 102.885 ;
               RECT 19.606 104.049 19.654 104.085 ;
               RECT 19.762 1.035 19.81 1.071 ;
               RECT 19.762 2.235 19.81 2.271 ;
               RECT 19.762 3.435 19.81 3.471 ;
               RECT 19.762 4.635 19.81 4.671 ;
               RECT 19.762 5.835 19.81 5.871 ;
               RECT 19.762 7.035 19.81 7.071 ;
               RECT 19.762 8.235 19.81 8.271 ;
               RECT 19.762 9.435 19.81 9.471 ;
               RECT 19.762 10.635 19.81 10.671 ;
               RECT 19.762 11.835 19.81 11.871 ;
               RECT 19.762 13.035 19.81 13.071 ;
               RECT 19.762 14.235 19.81 14.271 ;
               RECT 19.762 15.435 19.81 15.471 ;
               RECT 19.762 16.635 19.81 16.671 ;
               RECT 19.762 17.835 19.81 17.871 ;
               RECT 19.762 19.035 19.81 19.071 ;
               RECT 19.762 20.235 19.81 20.271 ;
               RECT 19.762 21.435 19.81 21.471 ;
               RECT 19.762 22.635 19.81 22.671 ;
               RECT 19.762 23.835 19.81 23.871 ;
               RECT 19.762 25.035 19.81 25.071 ;
               RECT 19.762 26.235 19.81 26.271 ;
               RECT 19.762 27.435 19.81 27.471 ;
               RECT 19.762 28.635 19.81 28.671 ;
               RECT 19.762 29.835 19.81 29.871 ;
               RECT 19.762 31.035 19.81 31.071 ;
               RECT 19.762 32.235 19.81 32.271 ;
               RECT 19.762 33.435 19.81 33.471 ;
               RECT 19.762 34.635 19.81 34.671 ;
               RECT 19.762 35.835 19.81 35.871 ;
               RECT 19.762 37.035 19.81 37.071 ;
               RECT 19.762 38.235 19.81 38.271 ;
               RECT 19.762 39.435 19.81 39.471 ;
               RECT 19.762 40.635 19.81 40.671 ;
               RECT 19.762 41.835 19.81 41.871 ;
               RECT 19.762 43.035 19.81 43.071 ;
               RECT 19.762 44.235 19.81 44.271 ;
               RECT 19.762 45.435 19.81 45.471 ;
               RECT 19.762 46.635 19.81 46.671 ;
               RECT 19.762 47.835 19.81 47.871 ;
               RECT 19.762 49.062 19.81 49.098 ;
               RECT 19.762 50.022 19.81 50.058 ;
               RECT 19.762 53.9235 19.81 53.9595 ;
               RECT 19.762 55.2405 19.81 55.2765 ;
               RECT 19.762 55.542 19.81 55.578 ;
               RECT 19.762 56.955 19.81 56.991 ;
               RECT 19.762 58.155 19.81 58.191 ;
               RECT 19.762 59.355 19.81 59.391 ;
               RECT 19.762 60.555 19.81 60.591 ;
               RECT 19.762 61.755 19.81 61.791 ;
               RECT 19.762 62.955 19.81 62.991 ;
               RECT 19.762 64.155 19.81 64.191 ;
               RECT 19.762 65.355 19.81 65.391 ;
               RECT 19.762 66.555 19.81 66.591 ;
               RECT 19.762 67.755 19.81 67.791 ;
               RECT 19.762 68.955 19.81 68.991 ;
               RECT 19.762 70.155 19.81 70.191 ;
               RECT 19.762 71.355 19.81 71.391 ;
               RECT 19.762 72.555 19.81 72.591 ;
               RECT 19.762 73.755 19.81 73.791 ;
               RECT 19.762 74.955 19.81 74.991 ;
               RECT 19.762 76.155 19.81 76.191 ;
               RECT 19.762 77.355 19.81 77.391 ;
               RECT 19.762 78.555 19.81 78.591 ;
               RECT 19.762 79.755 19.81 79.791 ;
               RECT 19.762 80.955 19.81 80.991 ;
               RECT 19.762 82.155 19.81 82.191 ;
               RECT 19.762 83.355 19.81 83.391 ;
               RECT 19.762 84.555 19.81 84.591 ;
               RECT 19.762 85.755 19.81 85.791 ;
               RECT 19.762 86.955 19.81 86.991 ;
               RECT 19.762 88.155 19.81 88.191 ;
               RECT 19.762 89.355 19.81 89.391 ;
               RECT 19.762 90.555 19.81 90.591 ;
               RECT 19.762 91.755 19.81 91.791 ;
               RECT 19.762 92.955 19.81 92.991 ;
               RECT 19.762 94.155 19.81 94.191 ;
               RECT 19.762 95.355 19.81 95.391 ;
               RECT 19.762 96.555 19.81 96.591 ;
               RECT 19.762 97.755 19.81 97.791 ;
               RECT 19.762 98.955 19.81 98.991 ;
               RECT 19.762 100.155 19.81 100.191 ;
               RECT 19.762 101.355 19.81 101.391 ;
               RECT 19.762 102.555 19.81 102.591 ;
               RECT 19.762 103.755 19.81 103.791 ;
               RECT 19.838 1.558 19.886 1.594 ;
               RECT 19.838 2.758 19.886 2.794 ;
               RECT 19.838 3.958 19.886 3.994 ;
               RECT 19.838 5.158 19.886 5.194 ;
               RECT 19.838 6.358 19.886 6.394 ;
               RECT 19.838 7.558 19.886 7.594 ;
               RECT 19.838 8.758 19.886 8.794 ;
               RECT 19.838 9.958 19.886 9.994 ;
               RECT 19.838 11.158 19.886 11.194 ;
               RECT 19.838 12.358 19.886 12.394 ;
               RECT 19.838 13.558 19.886 13.594 ;
               RECT 19.838 14.758 19.886 14.794 ;
               RECT 19.838 15.958 19.886 15.994 ;
               RECT 19.838 17.158 19.886 17.194 ;
               RECT 19.838 18.358 19.886 18.394 ;
               RECT 19.838 19.558 19.886 19.594 ;
               RECT 19.838 20.758 19.886 20.794 ;
               RECT 19.838 21.958 19.886 21.994 ;
               RECT 19.838 23.158 19.886 23.194 ;
               RECT 19.838 24.358 19.886 24.394 ;
               RECT 19.838 25.558 19.886 25.594 ;
               RECT 19.838 26.758 19.886 26.794 ;
               RECT 19.838 27.958 19.886 27.994 ;
               RECT 19.838 29.158 19.886 29.194 ;
               RECT 19.838 30.358 19.886 30.394 ;
               RECT 19.838 31.558 19.886 31.594 ;
               RECT 19.838 32.758 19.886 32.794 ;
               RECT 19.838 33.958 19.886 33.994 ;
               RECT 19.838 35.158 19.886 35.194 ;
               RECT 19.838 36.358 19.886 36.394 ;
               RECT 19.838 37.558 19.886 37.594 ;
               RECT 19.838 38.758 19.886 38.794 ;
               RECT 19.838 39.958 19.886 39.994 ;
               RECT 19.838 41.158 19.886 41.194 ;
               RECT 19.838 42.358 19.886 42.394 ;
               RECT 19.838 43.558 19.886 43.594 ;
               RECT 19.838 44.758 19.886 44.794 ;
               RECT 19.838 45.958 19.886 45.994 ;
               RECT 19.838 47.158 19.886 47.194 ;
               RECT 19.838 48.358 19.886 48.394 ;
               RECT 19.838 49.302 19.886 49.338 ;
               RECT 19.838 51.702 19.886 51.738 ;
               RECT 19.838 52.182 19.886 52.218 ;
               RECT 19.838 53.8005 19.886 53.8365 ;
               RECT 19.838 55.7205 19.886 55.7565 ;
               RECT 19.838 57.478 19.886 57.514 ;
               RECT 19.838 58.678 19.886 58.714 ;
               RECT 19.838 59.878 19.886 59.914 ;
               RECT 19.838 61.078 19.886 61.114 ;
               RECT 19.838 62.278 19.886 62.314 ;
               RECT 19.838 63.478 19.886 63.514 ;
               RECT 19.838 64.678 19.886 64.714 ;
               RECT 19.838 65.878 19.886 65.914 ;
               RECT 19.838 67.078 19.886 67.114 ;
               RECT 19.838 68.278 19.886 68.314 ;
               RECT 19.838 69.478 19.886 69.514 ;
               RECT 19.838 70.678 19.886 70.714 ;
               RECT 19.838 71.878 19.886 71.914 ;
               RECT 19.838 73.078 19.886 73.114 ;
               RECT 19.838 74.278 19.886 74.314 ;
               RECT 19.838 75.478 19.886 75.514 ;
               RECT 19.838 76.678 19.886 76.714 ;
               RECT 19.838 77.878 19.886 77.914 ;
               RECT 19.838 79.078 19.886 79.114 ;
               RECT 19.838 80.278 19.886 80.314 ;
               RECT 19.838 81.478 19.886 81.514 ;
               RECT 19.838 82.678 19.886 82.714 ;
               RECT 19.838 83.878 19.886 83.914 ;
               RECT 19.838 85.078 19.886 85.114 ;
               RECT 19.838 86.278 19.886 86.314 ;
               RECT 19.838 87.478 19.886 87.514 ;
               RECT 19.838 88.678 19.886 88.714 ;
               RECT 19.838 89.878 19.886 89.914 ;
               RECT 19.838 91.078 19.886 91.114 ;
               RECT 19.838 92.278 19.886 92.314 ;
               RECT 19.838 93.478 19.886 93.514 ;
               RECT 19.838 94.678 19.886 94.714 ;
               RECT 19.838 95.878 19.886 95.914 ;
               RECT 19.838 97.078 19.886 97.114 ;
               RECT 19.838 98.278 19.886 98.314 ;
               RECT 19.838 99.478 19.886 99.514 ;
               RECT 19.838 100.678 19.886 100.714 ;
               RECT 19.838 101.878 19.886 101.914 ;
               RECT 19.838 103.078 19.886 103.114 ;
               RECT 19.838 104.278 19.886 104.314 ;
               RECT 20.154 49.782 20.194 49.818 ;
               RECT 20.154 54.102 20.194 54.138 ;
               RECT 20.222 50.022 20.262 50.058 ;
               RECT 20.222 52.4835 20.262 52.5195 ;
               RECT 20.222 55.062 20.262 55.098 ;
               RECT 20.37 1.3345 20.442 1.3595 ;
               RECT 20.37 2.5345 20.442 2.5595 ;
               RECT 20.37 3.7345 20.442 3.7595 ;
               RECT 20.37 4.9345 20.442 4.9595 ;
               RECT 20.37 6.1345 20.442 6.1595 ;
               RECT 20.37 7.3345 20.442 7.3595 ;
               RECT 20.37 8.5345 20.442 8.5595 ;
               RECT 20.37 9.7345 20.442 9.7595 ;
               RECT 20.37 10.9345 20.442 10.9595 ;
               RECT 20.37 12.1345 20.442 12.1595 ;
               RECT 20.37 13.3345 20.442 13.3595 ;
               RECT 20.37 14.5345 20.442 14.5595 ;
               RECT 20.37 15.7345 20.442 15.7595 ;
               RECT 20.37 16.9345 20.442 16.9595 ;
               RECT 20.37 18.1345 20.442 18.1595 ;
               RECT 20.37 19.3345 20.442 19.3595 ;
               RECT 20.37 20.5345 20.442 20.5595 ;
               RECT 20.37 21.7345 20.442 21.7595 ;
               RECT 20.37 22.9345 20.442 22.9595 ;
               RECT 20.37 24.1345 20.442 24.1595 ;
               RECT 20.37 25.3345 20.442 25.3595 ;
               RECT 20.37 26.5345 20.442 26.5595 ;
               RECT 20.37 27.7345 20.442 27.7595 ;
               RECT 20.37 28.9345 20.442 28.9595 ;
               RECT 20.37 30.1345 20.442 30.1595 ;
               RECT 20.37 31.3345 20.442 31.3595 ;
               RECT 20.37 32.5345 20.442 32.5595 ;
               RECT 20.37 33.7345 20.442 33.7595 ;
               RECT 20.37 34.9345 20.442 34.9595 ;
               RECT 20.37 36.1345 20.442 36.1595 ;
               RECT 20.37 37.3345 20.442 37.3595 ;
               RECT 20.37 38.5345 20.442 38.5595 ;
               RECT 20.37 39.7345 20.442 39.7595 ;
               RECT 20.37 40.9345 20.442 40.9595 ;
               RECT 20.37 42.1345 20.442 42.1595 ;
               RECT 20.37 43.3345 20.442 43.3595 ;
               RECT 20.37 44.5345 20.442 44.5595 ;
               RECT 20.37 45.7345 20.442 45.7595 ;
               RECT 20.37 46.9345 20.442 46.9595 ;
               RECT 20.37 48.1345 20.442 48.1595 ;
               RECT 20.37 49.0675 20.442 49.0925 ;
               RECT 20.37 50.206 20.442 50.231 ;
               RECT 20.37 54.5875 20.442 54.6125 ;
               RECT 20.37 56.0275 20.442 56.0525 ;
               RECT 20.37 57.2545 20.442 57.2795 ;
               RECT 20.37 58.4545 20.442 58.4795 ;
               RECT 20.37 59.6545 20.442 59.6795 ;
               RECT 20.37 60.8545 20.442 60.8795 ;
               RECT 20.37 62.0545 20.442 62.0795 ;
               RECT 20.37 63.2545 20.442 63.2795 ;
               RECT 20.37 64.4545 20.442 64.4795 ;
               RECT 20.37 65.6545 20.442 65.6795 ;
               RECT 20.37 66.8545 20.442 66.8795 ;
               RECT 20.37 68.0545 20.442 68.0795 ;
               RECT 20.37 69.2545 20.442 69.2795 ;
               RECT 20.37 70.4545 20.442 70.4795 ;
               RECT 20.37 71.6545 20.442 71.6795 ;
               RECT 20.37 72.8545 20.442 72.8795 ;
               RECT 20.37 74.0545 20.442 74.0795 ;
               RECT 20.37 75.2545 20.442 75.2795 ;
               RECT 20.37 76.4545 20.442 76.4795 ;
               RECT 20.37 77.6545 20.442 77.6795 ;
               RECT 20.37 78.8545 20.442 78.8795 ;
               RECT 20.37 80.0545 20.442 80.0795 ;
               RECT 20.37 81.2545 20.442 81.2795 ;
               RECT 20.37 82.4545 20.442 82.4795 ;
               RECT 20.37 83.6545 20.442 83.6795 ;
               RECT 20.37 84.8545 20.442 84.8795 ;
               RECT 20.37 86.0545 20.442 86.0795 ;
               RECT 20.37 87.2545 20.442 87.2795 ;
               RECT 20.37 88.4545 20.442 88.4795 ;
               RECT 20.37 89.6545 20.442 89.6795 ;
               RECT 20.37 90.8545 20.442 90.8795 ;
               RECT 20.37 92.0545 20.442 92.0795 ;
               RECT 20.37 93.2545 20.442 93.2795 ;
               RECT 20.37 94.4545 20.442 94.4795 ;
               RECT 20.37 95.6545 20.442 95.6795 ;
               RECT 20.37 96.8545 20.442 96.8795 ;
               RECT 20.37 98.0545 20.442 98.0795 ;
               RECT 20.37 99.2545 20.442 99.2795 ;
               RECT 20.37 100.4545 20.442 100.4795 ;
               RECT 20.37 101.6545 20.442 101.6795 ;
               RECT 20.37 102.8545 20.442 102.8795 ;
               RECT 20.37 104.0545 20.442 104.0795 ;
               RECT 20.47 50.502 20.522 50.538 ;
               RECT 20.47 54.8835 20.522 54.9195 ;
               RECT 20.55 51.4005 20.602 51.4365 ;
               RECT 20.55 52.902 20.602 52.938 ;
               RECT 20.778 0.582 20.822 0.618 ;
               RECT 20.778 1.182 20.822 1.218 ;
               RECT 20.778 1.782 20.822 1.818 ;
               RECT 20.778 2.382 20.822 2.418 ;
               RECT 20.778 2.982 20.822 3.018 ;
               RECT 20.778 3.582 20.822 3.618 ;
               RECT 20.778 4.182 20.822 4.218 ;
               RECT 20.778 4.782 20.822 4.818 ;
               RECT 20.778 5.382 20.822 5.418 ;
               RECT 20.778 5.982 20.822 6.018 ;
               RECT 20.778 6.582 20.822 6.618 ;
               RECT 20.778 7.182 20.822 7.218 ;
               RECT 20.778 7.782 20.822 7.818 ;
               RECT 20.778 8.382 20.822 8.418 ;
               RECT 20.778 8.982 20.822 9.018 ;
               RECT 20.778 9.582 20.822 9.618 ;
               RECT 20.778 10.182 20.822 10.218 ;
               RECT 20.778 10.782 20.822 10.818 ;
               RECT 20.778 11.382 20.822 11.418 ;
               RECT 20.778 11.982 20.822 12.018 ;
               RECT 20.778 12.582 20.822 12.618 ;
               RECT 20.778 13.182 20.822 13.218 ;
               RECT 20.778 13.782 20.822 13.818 ;
               RECT 20.778 14.382 20.822 14.418 ;
               RECT 20.778 14.982 20.822 15.018 ;
               RECT 20.778 15.582 20.822 15.618 ;
               RECT 20.778 16.182 20.822 16.218 ;
               RECT 20.778 16.782 20.822 16.818 ;
               RECT 20.778 17.382 20.822 17.418 ;
               RECT 20.778 17.982 20.822 18.018 ;
               RECT 20.778 18.582 20.822 18.618 ;
               RECT 20.778 19.182 20.822 19.218 ;
               RECT 20.778 19.782 20.822 19.818 ;
               RECT 20.778 20.382 20.822 20.418 ;
               RECT 20.778 20.982 20.822 21.018 ;
               RECT 20.778 21.582 20.822 21.618 ;
               RECT 20.778 22.182 20.822 22.218 ;
               RECT 20.778 22.782 20.822 22.818 ;
               RECT 20.778 23.382 20.822 23.418 ;
               RECT 20.778 23.982 20.822 24.018 ;
               RECT 20.778 24.582 20.822 24.618 ;
               RECT 20.778 25.182 20.822 25.218 ;
               RECT 20.778 25.782 20.822 25.818 ;
               RECT 20.778 26.382 20.822 26.418 ;
               RECT 20.778 26.982 20.822 27.018 ;
               RECT 20.778 27.582 20.822 27.618 ;
               RECT 20.778 28.182 20.822 28.218 ;
               RECT 20.778 28.782 20.822 28.818 ;
               RECT 20.778 29.382 20.822 29.418 ;
               RECT 20.778 29.982 20.822 30.018 ;
               RECT 20.778 30.582 20.822 30.618 ;
               RECT 20.778 31.182 20.822 31.218 ;
               RECT 20.778 31.782 20.822 31.818 ;
               RECT 20.778 32.382 20.822 32.418 ;
               RECT 20.778 32.982 20.822 33.018 ;
               RECT 20.778 33.582 20.822 33.618 ;
               RECT 20.778 34.182 20.822 34.218 ;
               RECT 20.778 34.782 20.822 34.818 ;
               RECT 20.778 35.382 20.822 35.418 ;
               RECT 20.778 35.982 20.822 36.018 ;
               RECT 20.778 36.582 20.822 36.618 ;
               RECT 20.778 37.182 20.822 37.218 ;
               RECT 20.778 37.782 20.822 37.818 ;
               RECT 20.778 38.382 20.822 38.418 ;
               RECT 20.778 38.982 20.822 39.018 ;
               RECT 20.778 39.582 20.822 39.618 ;
               RECT 20.778 40.182 20.822 40.218 ;
               RECT 20.778 40.782 20.822 40.818 ;
               RECT 20.778 41.382 20.822 41.418 ;
               RECT 20.778 41.982 20.822 42.018 ;
               RECT 20.778 42.582 20.822 42.618 ;
               RECT 20.778 43.182 20.822 43.218 ;
               RECT 20.778 43.782 20.822 43.818 ;
               RECT 20.778 44.382 20.822 44.418 ;
               RECT 20.778 44.982 20.822 45.018 ;
               RECT 20.778 45.582 20.822 45.618 ;
               RECT 20.778 46.182 20.822 46.218 ;
               RECT 20.778 46.782 20.822 46.818 ;
               RECT 20.778 47.382 20.822 47.418 ;
               RECT 20.778 47.982 20.822 48.018 ;
               RECT 20.778 48.582 20.822 48.618 ;
               RECT 20.778 48.942 20.822 48.978 ;
               RECT 20.778 49.422 20.822 49.458 ;
               RECT 20.778 49.902 20.822 49.938 ;
               RECT 20.778 50.382 20.822 50.418 ;
               RECT 20.778 50.862 20.822 50.898 ;
               RECT 20.778 51.342 20.822 51.378 ;
               RECT 20.778 51.822 20.822 51.858 ;
               RECT 20.778 52.302 20.822 52.338 ;
               RECT 20.778 52.782 20.822 52.818 ;
               RECT 20.778 53.262 20.822 53.298 ;
               RECT 20.778 53.742 20.822 53.778 ;
               RECT 20.778 54.2275 20.822 54.2525 ;
               RECT 20.778 54.7075 20.822 54.7325 ;
               RECT 20.778 55.182 20.822 55.218 ;
               RECT 20.778 55.6675 20.822 55.6925 ;
               RECT 20.778 56.142 20.822 56.178 ;
               RECT 20.778 56.502 20.822 56.538 ;
               RECT 20.778 57.102 20.822 57.138 ;
               RECT 20.778 57.702 20.822 57.738 ;
               RECT 20.778 58.302 20.822 58.338 ;
               RECT 20.778 58.902 20.822 58.938 ;
               RECT 20.778 59.502 20.822 59.538 ;
               RECT 20.778 60.102 20.822 60.138 ;
               RECT 20.778 60.702 20.822 60.738 ;
               RECT 20.778 61.302 20.822 61.338 ;
               RECT 20.778 61.902 20.822 61.938 ;
               RECT 20.778 62.502 20.822 62.538 ;
               RECT 20.778 63.102 20.822 63.138 ;
               RECT 20.778 63.702 20.822 63.738 ;
               RECT 20.778 64.302 20.822 64.338 ;
               RECT 20.778 64.902 20.822 64.938 ;
               RECT 20.778 65.502 20.822 65.538 ;
               RECT 20.778 66.102 20.822 66.138 ;
               RECT 20.778 66.702 20.822 66.738 ;
               RECT 20.778 67.302 20.822 67.338 ;
               RECT 20.778 67.902 20.822 67.938 ;
               RECT 20.778 68.502 20.822 68.538 ;
               RECT 20.778 69.102 20.822 69.138 ;
               RECT 20.778 69.702 20.822 69.738 ;
               RECT 20.778 70.302 20.822 70.338 ;
               RECT 20.778 70.902 20.822 70.938 ;
               RECT 20.778 71.502 20.822 71.538 ;
               RECT 20.778 72.102 20.822 72.138 ;
               RECT 20.778 72.702 20.822 72.738 ;
               RECT 20.778 73.302 20.822 73.338 ;
               RECT 20.778 73.902 20.822 73.938 ;
               RECT 20.778 74.502 20.822 74.538 ;
               RECT 20.778 75.102 20.822 75.138 ;
               RECT 20.778 75.702 20.822 75.738 ;
               RECT 20.778 76.302 20.822 76.338 ;
               RECT 20.778 76.902 20.822 76.938 ;
               RECT 20.778 77.502 20.822 77.538 ;
               RECT 20.778 78.102 20.822 78.138 ;
               RECT 20.778 78.702 20.822 78.738 ;
               RECT 20.778 79.302 20.822 79.338 ;
               RECT 20.778 79.902 20.822 79.938 ;
               RECT 20.778 80.502 20.822 80.538 ;
               RECT 20.778 81.102 20.822 81.138 ;
               RECT 20.778 81.702 20.822 81.738 ;
               RECT 20.778 82.302 20.822 82.338 ;
               RECT 20.778 82.902 20.822 82.938 ;
               RECT 20.778 83.502 20.822 83.538 ;
               RECT 20.778 84.102 20.822 84.138 ;
               RECT 20.778 84.702 20.822 84.738 ;
               RECT 20.778 85.302 20.822 85.338 ;
               RECT 20.778 85.902 20.822 85.938 ;
               RECT 20.778 86.502 20.822 86.538 ;
               RECT 20.778 87.102 20.822 87.138 ;
               RECT 20.778 87.702 20.822 87.738 ;
               RECT 20.778 88.302 20.822 88.338 ;
               RECT 20.778 88.902 20.822 88.938 ;
               RECT 20.778 89.502 20.822 89.538 ;
               RECT 20.778 90.102 20.822 90.138 ;
               RECT 20.778 90.702 20.822 90.738 ;
               RECT 20.778 91.302 20.822 91.338 ;
               RECT 20.778 91.902 20.822 91.938 ;
               RECT 20.778 92.502 20.822 92.538 ;
               RECT 20.778 93.102 20.822 93.138 ;
               RECT 20.778 93.702 20.822 93.738 ;
               RECT 20.778 94.302 20.822 94.338 ;
               RECT 20.778 94.902 20.822 94.938 ;
               RECT 20.778 95.502 20.822 95.538 ;
               RECT 20.778 96.102 20.822 96.138 ;
               RECT 20.778 96.702 20.822 96.738 ;
               RECT 20.778 97.302 20.822 97.338 ;
               RECT 20.778 97.902 20.822 97.938 ;
               RECT 20.778 98.502 20.822 98.538 ;
               RECT 20.778 99.102 20.822 99.138 ;
               RECT 20.778 99.702 20.822 99.738 ;
               RECT 20.778 100.302 20.822 100.338 ;
               RECT 20.778 100.902 20.822 100.938 ;
               RECT 20.778 101.502 20.822 101.538 ;
               RECT 20.778 102.102 20.822 102.138 ;
               RECT 20.778 102.702 20.822 102.738 ;
               RECT 20.778 103.302 20.822 103.338 ;
               RECT 20.778 103.902 20.822 103.938 ;
               RECT 20.778 104.502 20.822 104.538 ;
               RECT 20.932 51.2835 20.986 51.3195 ;
               RECT 20.932 54.1635 20.986 54.1995 ;
               RECT 21.096 0.582 21.14 0.618 ;
               RECT 21.096 1.782 21.14 1.818 ;
               RECT 21.096 2.982 21.14 3.018 ;
               RECT 21.096 4.182 21.14 4.218 ;
               RECT 21.096 5.382 21.14 5.418 ;
               RECT 21.096 6.582 21.14 6.618 ;
               RECT 21.096 7.782 21.14 7.818 ;
               RECT 21.096 8.982 21.14 9.018 ;
               RECT 21.096 10.182 21.14 10.218 ;
               RECT 21.096 11.382 21.14 11.418 ;
               RECT 21.096 12.582 21.14 12.618 ;
               RECT 21.096 13.782 21.14 13.818 ;
               RECT 21.096 14.982 21.14 15.018 ;
               RECT 21.096 16.182 21.14 16.218 ;
               RECT 21.096 17.382 21.14 17.418 ;
               RECT 21.096 18.582 21.14 18.618 ;
               RECT 21.096 19.782 21.14 19.818 ;
               RECT 21.096 20.982 21.14 21.018 ;
               RECT 21.096 22.182 21.14 22.218 ;
               RECT 21.096 23.382 21.14 23.418 ;
               RECT 21.096 24.582 21.14 24.618 ;
               RECT 21.096 25.782 21.14 25.818 ;
               RECT 21.096 26.982 21.14 27.018 ;
               RECT 21.096 28.182 21.14 28.218 ;
               RECT 21.096 29.382 21.14 29.418 ;
               RECT 21.096 30.582 21.14 30.618 ;
               RECT 21.096 31.782 21.14 31.818 ;
               RECT 21.096 32.982 21.14 33.018 ;
               RECT 21.096 34.182 21.14 34.218 ;
               RECT 21.096 35.382 21.14 35.418 ;
               RECT 21.096 36.582 21.14 36.618 ;
               RECT 21.096 37.782 21.14 37.818 ;
               RECT 21.096 38.982 21.14 39.018 ;
               RECT 21.096 40.182 21.14 40.218 ;
               RECT 21.096 41.382 21.14 41.418 ;
               RECT 21.096 42.582 21.14 42.618 ;
               RECT 21.096 43.782 21.14 43.818 ;
               RECT 21.096 44.982 21.14 45.018 ;
               RECT 21.096 46.182 21.14 46.218 ;
               RECT 21.096 47.382 21.14 47.418 ;
               RECT 21.096 48.582 21.14 48.618 ;
               RECT 21.096 48.942 21.14 48.978 ;
               RECT 21.096 49.422 21.14 49.458 ;
               RECT 21.096 49.902 21.14 49.938 ;
               RECT 21.096 50.382 21.14 50.418 ;
               RECT 21.096 50.862 21.14 50.898 ;
               RECT 21.096 51.342 21.14 51.378 ;
               RECT 21.096 51.822 21.14 51.858 ;
               RECT 21.096 52.302 21.14 52.338 ;
               RECT 21.096 52.782 21.14 52.818 ;
               RECT 21.096 53.262 21.14 53.298 ;
               RECT 21.096 53.742 21.14 53.778 ;
               RECT 21.096 54.222 21.14 54.258 ;
               RECT 21.096 54.702 21.14 54.738 ;
               RECT 21.096 55.182 21.14 55.218 ;
               RECT 21.096 55.662 21.14 55.698 ;
               RECT 21.096 56.142 21.14 56.178 ;
               RECT 21.096 56.502 21.14 56.538 ;
               RECT 21.096 57.702 21.14 57.738 ;
               RECT 21.096 58.902 21.14 58.938 ;
               RECT 21.096 60.102 21.14 60.138 ;
               RECT 21.096 61.302 21.14 61.338 ;
               RECT 21.096 62.502 21.14 62.538 ;
               RECT 21.096 63.702 21.14 63.738 ;
               RECT 21.096 64.902 21.14 64.938 ;
               RECT 21.096 66.102 21.14 66.138 ;
               RECT 21.096 67.302 21.14 67.338 ;
               RECT 21.096 68.502 21.14 68.538 ;
               RECT 21.096 69.702 21.14 69.738 ;
               RECT 21.096 70.902 21.14 70.938 ;
               RECT 21.096 72.102 21.14 72.138 ;
               RECT 21.096 73.302 21.14 73.338 ;
               RECT 21.096 74.502 21.14 74.538 ;
               RECT 21.096 75.702 21.14 75.738 ;
               RECT 21.096 76.902 21.14 76.938 ;
               RECT 21.096 78.102 21.14 78.138 ;
               RECT 21.096 79.302 21.14 79.338 ;
               RECT 21.096 80.502 21.14 80.538 ;
               RECT 21.096 81.702 21.14 81.738 ;
               RECT 21.096 82.902 21.14 82.938 ;
               RECT 21.096 84.102 21.14 84.138 ;
               RECT 21.096 85.302 21.14 85.338 ;
               RECT 21.096 86.502 21.14 86.538 ;
               RECT 21.096 87.702 21.14 87.738 ;
               RECT 21.096 88.902 21.14 88.938 ;
               RECT 21.096 90.102 21.14 90.138 ;
               RECT 21.096 91.302 21.14 91.338 ;
               RECT 21.096 92.502 21.14 92.538 ;
               RECT 21.096 93.702 21.14 93.738 ;
               RECT 21.096 94.902 21.14 94.938 ;
               RECT 21.096 96.102 21.14 96.138 ;
               RECT 21.096 97.302 21.14 97.338 ;
               RECT 21.096 98.502 21.14 98.538 ;
               RECT 21.096 99.702 21.14 99.738 ;
               RECT 21.096 100.902 21.14 100.938 ;
               RECT 21.096 102.102 21.14 102.138 ;
               RECT 21.096 103.302 21.14 103.338 ;
               RECT 21.096 104.502 21.14 104.538 ;
               RECT 21.168 0.806 21.222 0.842 ;
               RECT 21.168 2.006 21.222 2.042 ;
               RECT 21.168 3.206 21.222 3.242 ;
               RECT 21.168 4.406 21.222 4.442 ;
               RECT 21.168 5.606 21.222 5.642 ;
               RECT 21.168 6.806 21.222 6.842 ;
               RECT 21.168 8.006 21.222 8.042 ;
               RECT 21.168 9.206 21.222 9.242 ;
               RECT 21.168 10.406 21.222 10.442 ;
               RECT 21.168 11.606 21.222 11.642 ;
               RECT 21.168 12.806 21.222 12.842 ;
               RECT 21.168 14.006 21.222 14.042 ;
               RECT 21.168 15.206 21.222 15.242 ;
               RECT 21.168 16.406 21.222 16.442 ;
               RECT 21.168 17.606 21.222 17.642 ;
               RECT 21.168 18.806 21.222 18.842 ;
               RECT 21.168 20.006 21.222 20.042 ;
               RECT 21.168 21.206 21.222 21.242 ;
               RECT 21.168 22.406 21.222 22.442 ;
               RECT 21.168 23.606 21.222 23.642 ;
               RECT 21.168 24.806 21.222 24.842 ;
               RECT 21.168 26.006 21.222 26.042 ;
               RECT 21.168 27.206 21.222 27.242 ;
               RECT 21.168 28.406 21.222 28.442 ;
               RECT 21.168 29.606 21.222 29.642 ;
               RECT 21.168 30.806 21.222 30.842 ;
               RECT 21.168 32.006 21.222 32.042 ;
               RECT 21.168 33.206 21.222 33.242 ;
               RECT 21.168 34.406 21.222 34.442 ;
               RECT 21.168 35.606 21.222 35.642 ;
               RECT 21.168 36.806 21.222 36.842 ;
               RECT 21.168 38.006 21.222 38.042 ;
               RECT 21.168 39.206 21.222 39.242 ;
               RECT 21.168 40.406 21.222 40.442 ;
               RECT 21.168 41.606 21.222 41.642 ;
               RECT 21.168 42.806 21.222 42.842 ;
               RECT 21.168 44.006 21.222 44.042 ;
               RECT 21.168 45.206 21.222 45.242 ;
               RECT 21.168 46.406 21.222 46.442 ;
               RECT 21.168 47.606 21.222 47.642 ;
               RECT 21.168 49.7205 21.222 49.7565 ;
               RECT 21.168 50.022 21.222 50.058 ;
               RECT 21.168 54.582 21.222 54.618 ;
               RECT 21.168 55.062 21.222 55.098 ;
               RECT 21.168 55.4805 21.222 55.5165 ;
               RECT 21.168 56.726 21.222 56.762 ;
               RECT 21.168 57.926 21.222 57.962 ;
               RECT 21.168 59.126 21.222 59.162 ;
               RECT 21.168 60.326 21.222 60.362 ;
               RECT 21.168 61.526 21.222 61.562 ;
               RECT 21.168 62.726 21.222 62.762 ;
               RECT 21.168 63.926 21.222 63.962 ;
               RECT 21.168 65.126 21.222 65.162 ;
               RECT 21.168 66.326 21.222 66.362 ;
               RECT 21.168 67.526 21.222 67.562 ;
               RECT 21.168 68.726 21.222 68.762 ;
               RECT 21.168 69.926 21.222 69.962 ;
               RECT 21.168 71.126 21.222 71.162 ;
               RECT 21.168 72.326 21.222 72.362 ;
               RECT 21.168 73.526 21.222 73.562 ;
               RECT 21.168 74.726 21.222 74.762 ;
               RECT 21.168 75.926 21.222 75.962 ;
               RECT 21.168 77.126 21.222 77.162 ;
               RECT 21.168 78.326 21.222 78.362 ;
               RECT 21.168 79.526 21.222 79.562 ;
               RECT 21.168 80.726 21.222 80.762 ;
               RECT 21.168 81.926 21.222 81.962 ;
               RECT 21.168 83.126 21.222 83.162 ;
               RECT 21.168 84.326 21.222 84.362 ;
               RECT 21.168 85.526 21.222 85.562 ;
               RECT 21.168 86.726 21.222 86.762 ;
               RECT 21.168 87.926 21.222 87.962 ;
               RECT 21.168 89.126 21.222 89.162 ;
               RECT 21.168 90.326 21.222 90.362 ;
               RECT 21.168 91.526 21.222 91.562 ;
               RECT 21.168 92.726 21.222 92.762 ;
               RECT 21.168 93.926 21.222 93.962 ;
               RECT 21.168 95.126 21.222 95.162 ;
               RECT 21.168 96.326 21.222 96.362 ;
               RECT 21.168 97.526 21.222 97.562 ;
               RECT 21.168 98.726 21.222 98.762 ;
               RECT 21.168 99.926 21.222 99.962 ;
               RECT 21.168 101.126 21.222 101.162 ;
               RECT 21.168 102.326 21.222 102.362 ;
               RECT 21.168 103.526 21.222 103.562 ;
               RECT 21.25 1.482 21.304 1.518 ;
               RECT 21.25 2.682 21.304 2.718 ;
               RECT 21.25 3.882 21.304 3.918 ;
               RECT 21.25 5.082 21.304 5.118 ;
               RECT 21.25 6.282 21.304 6.318 ;
               RECT 21.25 7.482 21.304 7.518 ;
               RECT 21.25 8.682 21.304 8.718 ;
               RECT 21.25 9.882 21.304 9.918 ;
               RECT 21.25 11.082 21.304 11.118 ;
               RECT 21.25 12.282 21.304 12.318 ;
               RECT 21.25 13.482 21.304 13.518 ;
               RECT 21.25 14.682 21.304 14.718 ;
               RECT 21.25 15.882 21.304 15.918 ;
               RECT 21.25 17.082 21.304 17.118 ;
               RECT 21.25 18.282 21.304 18.318 ;
               RECT 21.25 19.482 21.304 19.518 ;
               RECT 21.25 20.682 21.304 20.718 ;
               RECT 21.25 21.882 21.304 21.918 ;
               RECT 21.25 23.082 21.304 23.118 ;
               RECT 21.25 24.282 21.304 24.318 ;
               RECT 21.25 25.482 21.304 25.518 ;
               RECT 21.25 26.682 21.304 26.718 ;
               RECT 21.25 27.882 21.304 27.918 ;
               RECT 21.25 29.082 21.304 29.118 ;
               RECT 21.25 30.282 21.304 30.318 ;
               RECT 21.25 31.482 21.304 31.518 ;
               RECT 21.25 32.682 21.304 32.718 ;
               RECT 21.25 33.882 21.304 33.918 ;
               RECT 21.25 35.082 21.304 35.118 ;
               RECT 21.25 36.282 21.304 36.318 ;
               RECT 21.25 37.482 21.304 37.518 ;
               RECT 21.25 38.682 21.304 38.718 ;
               RECT 21.25 39.882 21.304 39.918 ;
               RECT 21.25 41.082 21.304 41.118 ;
               RECT 21.25 42.282 21.304 42.318 ;
               RECT 21.25 43.482 21.304 43.518 ;
               RECT 21.25 44.682 21.304 44.718 ;
               RECT 21.25 45.882 21.304 45.918 ;
               RECT 21.25 47.082 21.304 47.118 ;
               RECT 21.25 48.282 21.304 48.318 ;
               RECT 21.25 49.3635 21.304 49.3995 ;
               RECT 21.25 49.6035 21.304 49.6395 ;
               RECT 21.25 54.4035 21.304 54.4395 ;
               RECT 21.25 55.3635 21.304 55.3995 ;
               RECT 21.25 55.7205 21.304 55.7565 ;
               RECT 21.25 57.402 21.304 57.438 ;
               RECT 21.25 58.602 21.304 58.638 ;
               RECT 21.25 59.802 21.304 59.838 ;
               RECT 21.25 61.002 21.304 61.038 ;
               RECT 21.25 62.202 21.304 62.238 ;
               RECT 21.25 63.402 21.304 63.438 ;
               RECT 21.25 64.602 21.304 64.638 ;
               RECT 21.25 65.802 21.304 65.838 ;
               RECT 21.25 67.002 21.304 67.038 ;
               RECT 21.25 68.202 21.304 68.238 ;
               RECT 21.25 69.402 21.304 69.438 ;
               RECT 21.25 70.602 21.304 70.638 ;
               RECT 21.25 71.802 21.304 71.838 ;
               RECT 21.25 73.002 21.304 73.038 ;
               RECT 21.25 74.202 21.304 74.238 ;
               RECT 21.25 75.402 21.304 75.438 ;
               RECT 21.25 76.602 21.304 76.638 ;
               RECT 21.25 77.802 21.304 77.838 ;
               RECT 21.25 79.002 21.304 79.038 ;
               RECT 21.25 80.202 21.304 80.238 ;
               RECT 21.25 81.402 21.304 81.438 ;
               RECT 21.25 82.602 21.304 82.638 ;
               RECT 21.25 83.802 21.304 83.838 ;
               RECT 21.25 85.002 21.304 85.038 ;
               RECT 21.25 86.202 21.304 86.238 ;
               RECT 21.25 87.402 21.304 87.438 ;
               RECT 21.25 88.602 21.304 88.638 ;
               RECT 21.25 89.802 21.304 89.838 ;
               RECT 21.25 91.002 21.304 91.038 ;
               RECT 21.25 92.202 21.304 92.238 ;
               RECT 21.25 93.402 21.304 93.438 ;
               RECT 21.25 94.602 21.304 94.638 ;
               RECT 21.25 95.802 21.304 95.838 ;
               RECT 21.25 97.002 21.304 97.038 ;
               RECT 21.25 98.202 21.304 98.238 ;
               RECT 21.25 99.402 21.304 99.438 ;
               RECT 21.25 100.602 21.304 100.638 ;
               RECT 21.25 101.802 21.304 101.838 ;
               RECT 21.25 103.002 21.304 103.038 ;
               RECT 21.25 104.202 21.304 104.238 ;
               RECT 21.332 0.806 21.386 0.842 ;
               RECT 21.332 2.006 21.386 2.042 ;
               RECT 21.332 3.206 21.386 3.242 ;
               RECT 21.332 4.406 21.386 4.442 ;
               RECT 21.332 5.606 21.386 5.642 ;
               RECT 21.332 6.806 21.386 6.842 ;
               RECT 21.332 8.006 21.386 8.042 ;
               RECT 21.332 9.206 21.386 9.242 ;
               RECT 21.332 10.406 21.386 10.442 ;
               RECT 21.332 11.606 21.386 11.642 ;
               RECT 21.332 12.806 21.386 12.842 ;
               RECT 21.332 14.006 21.386 14.042 ;
               RECT 21.332 15.206 21.386 15.242 ;
               RECT 21.332 16.406 21.386 16.442 ;
               RECT 21.332 17.606 21.386 17.642 ;
               RECT 21.332 18.806 21.386 18.842 ;
               RECT 21.332 20.006 21.386 20.042 ;
               RECT 21.332 21.206 21.386 21.242 ;
               RECT 21.332 22.406 21.386 22.442 ;
               RECT 21.332 23.606 21.386 23.642 ;
               RECT 21.332 24.806 21.386 24.842 ;
               RECT 21.332 26.006 21.386 26.042 ;
               RECT 21.332 27.206 21.386 27.242 ;
               RECT 21.332 28.406 21.386 28.442 ;
               RECT 21.332 29.606 21.386 29.642 ;
               RECT 21.332 30.806 21.386 30.842 ;
               RECT 21.332 32.006 21.386 32.042 ;
               RECT 21.332 33.206 21.386 33.242 ;
               RECT 21.332 34.406 21.386 34.442 ;
               RECT 21.332 35.606 21.386 35.642 ;
               RECT 21.332 36.806 21.386 36.842 ;
               RECT 21.332 38.006 21.386 38.042 ;
               RECT 21.332 39.206 21.386 39.242 ;
               RECT 21.332 40.406 21.386 40.442 ;
               RECT 21.332 41.606 21.386 41.642 ;
               RECT 21.332 42.806 21.386 42.842 ;
               RECT 21.332 44.006 21.386 44.042 ;
               RECT 21.332 45.206 21.386 45.242 ;
               RECT 21.332 46.406 21.386 46.442 ;
               RECT 21.332 47.606 21.386 47.642 ;
               RECT 21.332 49.0005 21.386 49.0365 ;
               RECT 21.332 49.4805 21.386 49.5165 ;
               RECT 21.332 54.6435 21.386 54.6795 ;
               RECT 21.332 55.486 21.386 55.511 ;
               RECT 21.332 55.609 21.386 55.634 ;
               RECT 21.332 56.726 21.386 56.762 ;
               RECT 21.332 57.926 21.386 57.962 ;
               RECT 21.332 59.126 21.386 59.162 ;
               RECT 21.332 60.326 21.386 60.362 ;
               RECT 21.332 61.526 21.386 61.562 ;
               RECT 21.332 62.726 21.386 62.762 ;
               RECT 21.332 63.926 21.386 63.962 ;
               RECT 21.332 65.126 21.386 65.162 ;
               RECT 21.332 66.326 21.386 66.362 ;
               RECT 21.332 67.526 21.386 67.562 ;
               RECT 21.332 68.726 21.386 68.762 ;
               RECT 21.332 69.926 21.386 69.962 ;
               RECT 21.332 71.126 21.386 71.162 ;
               RECT 21.332 72.326 21.386 72.362 ;
               RECT 21.332 73.526 21.386 73.562 ;
               RECT 21.332 74.726 21.386 74.762 ;
               RECT 21.332 75.926 21.386 75.962 ;
               RECT 21.332 77.126 21.386 77.162 ;
               RECT 21.332 78.326 21.386 78.362 ;
               RECT 21.332 79.526 21.386 79.562 ;
               RECT 21.332 80.726 21.386 80.762 ;
               RECT 21.332 81.926 21.386 81.962 ;
               RECT 21.332 83.126 21.386 83.162 ;
               RECT 21.332 84.326 21.386 84.362 ;
               RECT 21.332 85.526 21.386 85.562 ;
               RECT 21.332 86.726 21.386 86.762 ;
               RECT 21.332 87.926 21.386 87.962 ;
               RECT 21.332 89.126 21.386 89.162 ;
               RECT 21.332 90.326 21.386 90.362 ;
               RECT 21.332 91.526 21.386 91.562 ;
               RECT 21.332 92.726 21.386 92.762 ;
               RECT 21.332 93.926 21.386 93.962 ;
               RECT 21.332 95.126 21.386 95.162 ;
               RECT 21.332 96.326 21.386 96.362 ;
               RECT 21.332 97.526 21.386 97.562 ;
               RECT 21.332 98.726 21.386 98.762 ;
               RECT 21.332 99.926 21.386 99.962 ;
               RECT 21.332 101.126 21.386 101.162 ;
               RECT 21.332 102.326 21.386 102.362 ;
               RECT 21.332 103.526 21.386 103.562 ;
               RECT 21.414 1.482 21.468 1.518 ;
               RECT 21.414 2.682 21.468 2.718 ;
               RECT 21.414 3.882 21.468 3.918 ;
               RECT 21.414 5.082 21.468 5.118 ;
               RECT 21.414 6.282 21.468 6.318 ;
               RECT 21.414 7.482 21.468 7.518 ;
               RECT 21.414 8.682 21.468 8.718 ;
               RECT 21.414 9.882 21.468 9.918 ;
               RECT 21.414 11.082 21.468 11.118 ;
               RECT 21.414 12.282 21.468 12.318 ;
               RECT 21.414 13.482 21.468 13.518 ;
               RECT 21.414 14.682 21.468 14.718 ;
               RECT 21.414 15.882 21.468 15.918 ;
               RECT 21.414 17.082 21.468 17.118 ;
               RECT 21.414 18.282 21.468 18.318 ;
               RECT 21.414 19.482 21.468 19.518 ;
               RECT 21.414 20.682 21.468 20.718 ;
               RECT 21.414 21.882 21.468 21.918 ;
               RECT 21.414 23.082 21.468 23.118 ;
               RECT 21.414 24.282 21.468 24.318 ;
               RECT 21.414 25.482 21.468 25.518 ;
               RECT 21.414 26.682 21.468 26.718 ;
               RECT 21.414 27.882 21.468 27.918 ;
               RECT 21.414 29.082 21.468 29.118 ;
               RECT 21.414 30.282 21.468 30.318 ;
               RECT 21.414 31.482 21.468 31.518 ;
               RECT 21.414 32.682 21.468 32.718 ;
               RECT 21.414 33.882 21.468 33.918 ;
               RECT 21.414 35.082 21.468 35.118 ;
               RECT 21.414 36.282 21.468 36.318 ;
               RECT 21.414 37.482 21.468 37.518 ;
               RECT 21.414 38.682 21.468 38.718 ;
               RECT 21.414 39.882 21.468 39.918 ;
               RECT 21.414 41.082 21.468 41.118 ;
               RECT 21.414 42.282 21.468 42.318 ;
               RECT 21.414 43.482 21.468 43.518 ;
               RECT 21.414 44.682 21.468 44.718 ;
               RECT 21.414 45.882 21.468 45.918 ;
               RECT 21.414 47.082 21.468 47.118 ;
               RECT 21.414 48.282 21.468 48.318 ;
               RECT 21.414 49.1235 21.468 49.1595 ;
               RECT 21.414 49.2405 21.468 49.2765 ;
               RECT 21.414 54.4035 21.468 54.4395 ;
               RECT 21.414 55.782 21.468 55.818 ;
               RECT 21.414 56.022 21.468 56.058 ;
               RECT 21.414 57.402 21.468 57.438 ;
               RECT 21.414 58.602 21.468 58.638 ;
               RECT 21.414 59.802 21.468 59.838 ;
               RECT 21.414 61.002 21.468 61.038 ;
               RECT 21.414 62.202 21.468 62.238 ;
               RECT 21.414 63.402 21.468 63.438 ;
               RECT 21.414 64.602 21.468 64.638 ;
               RECT 21.414 65.802 21.468 65.838 ;
               RECT 21.414 67.002 21.468 67.038 ;
               RECT 21.414 68.202 21.468 68.238 ;
               RECT 21.414 69.402 21.468 69.438 ;
               RECT 21.414 70.602 21.468 70.638 ;
               RECT 21.414 71.802 21.468 71.838 ;
               RECT 21.414 73.002 21.468 73.038 ;
               RECT 21.414 74.202 21.468 74.238 ;
               RECT 21.414 75.402 21.468 75.438 ;
               RECT 21.414 76.602 21.468 76.638 ;
               RECT 21.414 77.802 21.468 77.838 ;
               RECT 21.414 79.002 21.468 79.038 ;
               RECT 21.414 80.202 21.468 80.238 ;
               RECT 21.414 81.402 21.468 81.438 ;
               RECT 21.414 82.602 21.468 82.638 ;
               RECT 21.414 83.802 21.468 83.838 ;
               RECT 21.414 85.002 21.468 85.038 ;
               RECT 21.414 86.202 21.468 86.238 ;
               RECT 21.414 87.402 21.468 87.438 ;
               RECT 21.414 88.602 21.468 88.638 ;
               RECT 21.414 89.802 21.468 89.838 ;
               RECT 21.414 91.002 21.468 91.038 ;
               RECT 21.414 92.202 21.468 92.238 ;
               RECT 21.414 93.402 21.468 93.438 ;
               RECT 21.414 94.602 21.468 94.638 ;
               RECT 21.414 95.802 21.468 95.838 ;
               RECT 21.414 97.002 21.468 97.038 ;
               RECT 21.414 98.202 21.468 98.238 ;
               RECT 21.414 99.402 21.468 99.438 ;
               RECT 21.414 100.602 21.468 100.638 ;
               RECT 21.414 101.802 21.468 101.838 ;
               RECT 21.414 103.002 21.468 103.038 ;
               RECT 21.414 104.202 21.468 104.238 ;
               RECT 21.578 50.982 21.622 51.018 ;
               RECT 21.578 51.222 21.622 51.258 ;
               RECT 21.578 53.142 21.622 53.178 ;
               RECT 21.578 54.102 21.622 54.138 ;
               RECT 21.732 0.806 21.786 0.842 ;
               RECT 21.732 2.006 21.786 2.042 ;
               RECT 21.732 3.206 21.786 3.242 ;
               RECT 21.732 4.406 21.786 4.442 ;
               RECT 21.732 5.606 21.786 5.642 ;
               RECT 21.732 6.806 21.786 6.842 ;
               RECT 21.732 8.006 21.786 8.042 ;
               RECT 21.732 9.206 21.786 9.242 ;
               RECT 21.732 10.406 21.786 10.442 ;
               RECT 21.732 11.606 21.786 11.642 ;
               RECT 21.732 12.806 21.786 12.842 ;
               RECT 21.732 14.006 21.786 14.042 ;
               RECT 21.732 15.206 21.786 15.242 ;
               RECT 21.732 16.406 21.786 16.442 ;
               RECT 21.732 17.606 21.786 17.642 ;
               RECT 21.732 18.806 21.786 18.842 ;
               RECT 21.732 20.006 21.786 20.042 ;
               RECT 21.732 21.206 21.786 21.242 ;
               RECT 21.732 22.406 21.786 22.442 ;
               RECT 21.732 23.606 21.786 23.642 ;
               RECT 21.732 24.806 21.786 24.842 ;
               RECT 21.732 26.006 21.786 26.042 ;
               RECT 21.732 27.206 21.786 27.242 ;
               RECT 21.732 28.406 21.786 28.442 ;
               RECT 21.732 29.606 21.786 29.642 ;
               RECT 21.732 30.806 21.786 30.842 ;
               RECT 21.732 32.006 21.786 32.042 ;
               RECT 21.732 33.206 21.786 33.242 ;
               RECT 21.732 34.406 21.786 34.442 ;
               RECT 21.732 35.606 21.786 35.642 ;
               RECT 21.732 36.806 21.786 36.842 ;
               RECT 21.732 38.006 21.786 38.042 ;
               RECT 21.732 39.206 21.786 39.242 ;
               RECT 21.732 40.406 21.786 40.442 ;
               RECT 21.732 41.606 21.786 41.642 ;
               RECT 21.732 42.806 21.786 42.842 ;
               RECT 21.732 44.006 21.786 44.042 ;
               RECT 21.732 45.206 21.786 45.242 ;
               RECT 21.732 46.406 21.786 46.442 ;
               RECT 21.732 47.606 21.786 47.642 ;
               RECT 21.732 50.8035 21.786 50.8395 ;
               RECT 21.732 53.8005 21.786 53.8365 ;
               RECT 21.732 56.726 21.786 56.762 ;
               RECT 21.732 57.926 21.786 57.962 ;
               RECT 21.732 59.126 21.786 59.162 ;
               RECT 21.732 60.326 21.786 60.362 ;
               RECT 21.732 61.526 21.786 61.562 ;
               RECT 21.732 62.726 21.786 62.762 ;
               RECT 21.732 63.926 21.786 63.962 ;
               RECT 21.732 65.126 21.786 65.162 ;
               RECT 21.732 66.326 21.786 66.362 ;
               RECT 21.732 67.526 21.786 67.562 ;
               RECT 21.732 68.726 21.786 68.762 ;
               RECT 21.732 69.926 21.786 69.962 ;
               RECT 21.732 71.126 21.786 71.162 ;
               RECT 21.732 72.326 21.786 72.362 ;
               RECT 21.732 73.526 21.786 73.562 ;
               RECT 21.732 74.726 21.786 74.762 ;
               RECT 21.732 75.926 21.786 75.962 ;
               RECT 21.732 77.126 21.786 77.162 ;
               RECT 21.732 78.326 21.786 78.362 ;
               RECT 21.732 79.526 21.786 79.562 ;
               RECT 21.732 80.726 21.786 80.762 ;
               RECT 21.732 81.926 21.786 81.962 ;
               RECT 21.732 83.126 21.786 83.162 ;
               RECT 21.732 84.326 21.786 84.362 ;
               RECT 21.732 85.526 21.786 85.562 ;
               RECT 21.732 86.726 21.786 86.762 ;
               RECT 21.732 87.926 21.786 87.962 ;
               RECT 21.732 89.126 21.786 89.162 ;
               RECT 21.732 90.326 21.786 90.362 ;
               RECT 21.732 91.526 21.786 91.562 ;
               RECT 21.732 92.726 21.786 92.762 ;
               RECT 21.732 93.926 21.786 93.962 ;
               RECT 21.732 95.126 21.786 95.162 ;
               RECT 21.732 96.326 21.786 96.362 ;
               RECT 21.732 97.526 21.786 97.562 ;
               RECT 21.732 98.726 21.786 98.762 ;
               RECT 21.732 99.926 21.786 99.962 ;
               RECT 21.732 101.126 21.786 101.162 ;
               RECT 21.732 102.326 21.786 102.362 ;
               RECT 21.732 103.526 21.786 103.562 ;
               RECT 21.814 1.558 21.868 1.594 ;
               RECT 21.814 2.758 21.868 2.794 ;
               RECT 21.814 3.958 21.868 3.994 ;
               RECT 21.814 5.158 21.868 5.194 ;
               RECT 21.814 6.358 21.868 6.394 ;
               RECT 21.814 7.558 21.868 7.594 ;
               RECT 21.814 8.758 21.868 8.794 ;
               RECT 21.814 9.958 21.868 9.994 ;
               RECT 21.814 11.158 21.868 11.194 ;
               RECT 21.814 12.358 21.868 12.394 ;
               RECT 21.814 13.558 21.868 13.594 ;
               RECT 21.814 14.758 21.868 14.794 ;
               RECT 21.814 15.958 21.868 15.994 ;
               RECT 21.814 17.158 21.868 17.194 ;
               RECT 21.814 18.358 21.868 18.394 ;
               RECT 21.814 19.558 21.868 19.594 ;
               RECT 21.814 20.758 21.868 20.794 ;
               RECT 21.814 21.958 21.868 21.994 ;
               RECT 21.814 23.158 21.868 23.194 ;
               RECT 21.814 24.358 21.868 24.394 ;
               RECT 21.814 25.558 21.868 25.594 ;
               RECT 21.814 26.758 21.868 26.794 ;
               RECT 21.814 27.958 21.868 27.994 ;
               RECT 21.814 29.158 21.868 29.194 ;
               RECT 21.814 30.358 21.868 30.394 ;
               RECT 21.814 31.558 21.868 31.594 ;
               RECT 21.814 32.758 21.868 32.794 ;
               RECT 21.814 33.958 21.868 33.994 ;
               RECT 21.814 35.158 21.868 35.194 ;
               RECT 21.814 36.358 21.868 36.394 ;
               RECT 21.814 37.558 21.868 37.594 ;
               RECT 21.814 38.758 21.868 38.794 ;
               RECT 21.814 39.958 21.868 39.994 ;
               RECT 21.814 41.158 21.868 41.194 ;
               RECT 21.814 42.358 21.868 42.394 ;
               RECT 21.814 43.558 21.868 43.594 ;
               RECT 21.814 44.758 21.868 44.794 ;
               RECT 21.814 45.958 21.868 45.994 ;
               RECT 21.814 47.158 21.868 47.194 ;
               RECT 21.814 48.358 21.868 48.394 ;
               RECT 21.814 50.9205 21.868 50.9565 ;
               RECT 21.814 51.1605 21.868 51.1965 ;
               RECT 21.814 52.7235 21.868 52.7595 ;
               RECT 21.814 54.1635 21.868 54.1995 ;
               RECT 21.814 57.478 21.868 57.514 ;
               RECT 21.814 58.678 21.868 58.714 ;
               RECT 21.814 59.878 21.868 59.914 ;
               RECT 21.814 61.078 21.868 61.114 ;
               RECT 21.814 62.278 21.868 62.314 ;
               RECT 21.814 63.478 21.868 63.514 ;
               RECT 21.814 64.678 21.868 64.714 ;
               RECT 21.814 65.878 21.868 65.914 ;
               RECT 21.814 67.078 21.868 67.114 ;
               RECT 21.814 68.278 21.868 68.314 ;
               RECT 21.814 69.478 21.868 69.514 ;
               RECT 21.814 70.678 21.868 70.714 ;
               RECT 21.814 71.878 21.868 71.914 ;
               RECT 21.814 73.078 21.868 73.114 ;
               RECT 21.814 74.278 21.868 74.314 ;
               RECT 21.814 75.478 21.868 75.514 ;
               RECT 21.814 76.678 21.868 76.714 ;
               RECT 21.814 77.878 21.868 77.914 ;
               RECT 21.814 79.078 21.868 79.114 ;
               RECT 21.814 80.278 21.868 80.314 ;
               RECT 21.814 81.478 21.868 81.514 ;
               RECT 21.814 82.678 21.868 82.714 ;
               RECT 21.814 83.878 21.868 83.914 ;
               RECT 21.814 85.078 21.868 85.114 ;
               RECT 21.814 86.278 21.868 86.314 ;
               RECT 21.814 87.478 21.868 87.514 ;
               RECT 21.814 88.678 21.868 88.714 ;
               RECT 21.814 89.878 21.868 89.914 ;
               RECT 21.814 91.078 21.868 91.114 ;
               RECT 21.814 92.278 21.868 92.314 ;
               RECT 21.814 93.478 21.868 93.514 ;
               RECT 21.814 94.678 21.868 94.714 ;
               RECT 21.814 95.878 21.868 95.914 ;
               RECT 21.814 97.078 21.868 97.114 ;
               RECT 21.814 98.278 21.868 98.314 ;
               RECT 21.814 99.478 21.868 99.514 ;
               RECT 21.814 100.678 21.868 100.714 ;
               RECT 21.814 101.878 21.868 101.914 ;
               RECT 21.814 103.078 21.868 103.114 ;
               RECT 21.814 104.278 21.868 104.314 ;
               RECT 21.978 0.582 22.022 0.618 ;
               RECT 21.978 1.182 22.022 1.218 ;
               RECT 21.978 1.782 22.022 1.818 ;
               RECT 21.978 2.382 22.022 2.418 ;
               RECT 21.978 2.982 22.022 3.018 ;
               RECT 21.978 3.582 22.022 3.618 ;
               RECT 21.978 4.182 22.022 4.218 ;
               RECT 21.978 4.782 22.022 4.818 ;
               RECT 21.978 5.382 22.022 5.418 ;
               RECT 21.978 5.982 22.022 6.018 ;
               RECT 21.978 6.582 22.022 6.618 ;
               RECT 21.978 7.182 22.022 7.218 ;
               RECT 21.978 7.782 22.022 7.818 ;
               RECT 21.978 8.382 22.022 8.418 ;
               RECT 21.978 8.982 22.022 9.018 ;
               RECT 21.978 9.582 22.022 9.618 ;
               RECT 21.978 10.182 22.022 10.218 ;
               RECT 21.978 10.782 22.022 10.818 ;
               RECT 21.978 11.382 22.022 11.418 ;
               RECT 21.978 11.982 22.022 12.018 ;
               RECT 21.978 12.582 22.022 12.618 ;
               RECT 21.978 13.182 22.022 13.218 ;
               RECT 21.978 13.782 22.022 13.818 ;
               RECT 21.978 14.382 22.022 14.418 ;
               RECT 21.978 14.982 22.022 15.018 ;
               RECT 21.978 15.582 22.022 15.618 ;
               RECT 21.978 16.182 22.022 16.218 ;
               RECT 21.978 16.782 22.022 16.818 ;
               RECT 21.978 17.382 22.022 17.418 ;
               RECT 21.978 17.982 22.022 18.018 ;
               RECT 21.978 18.582 22.022 18.618 ;
               RECT 21.978 19.182 22.022 19.218 ;
               RECT 21.978 19.782 22.022 19.818 ;
               RECT 21.978 20.382 22.022 20.418 ;
               RECT 21.978 20.982 22.022 21.018 ;
               RECT 21.978 21.582 22.022 21.618 ;
               RECT 21.978 22.182 22.022 22.218 ;
               RECT 21.978 22.782 22.022 22.818 ;
               RECT 21.978 23.382 22.022 23.418 ;
               RECT 21.978 23.982 22.022 24.018 ;
               RECT 21.978 24.582 22.022 24.618 ;
               RECT 21.978 25.182 22.022 25.218 ;
               RECT 21.978 25.782 22.022 25.818 ;
               RECT 21.978 26.382 22.022 26.418 ;
               RECT 21.978 26.982 22.022 27.018 ;
               RECT 21.978 27.582 22.022 27.618 ;
               RECT 21.978 28.182 22.022 28.218 ;
               RECT 21.978 28.782 22.022 28.818 ;
               RECT 21.978 29.382 22.022 29.418 ;
               RECT 21.978 29.982 22.022 30.018 ;
               RECT 21.978 30.582 22.022 30.618 ;
               RECT 21.978 31.182 22.022 31.218 ;
               RECT 21.978 31.782 22.022 31.818 ;
               RECT 21.978 32.382 22.022 32.418 ;
               RECT 21.978 32.982 22.022 33.018 ;
               RECT 21.978 33.582 22.022 33.618 ;
               RECT 21.978 34.182 22.022 34.218 ;
               RECT 21.978 34.782 22.022 34.818 ;
               RECT 21.978 35.382 22.022 35.418 ;
               RECT 21.978 35.982 22.022 36.018 ;
               RECT 21.978 36.582 22.022 36.618 ;
               RECT 21.978 37.182 22.022 37.218 ;
               RECT 21.978 37.782 22.022 37.818 ;
               RECT 21.978 38.382 22.022 38.418 ;
               RECT 21.978 38.982 22.022 39.018 ;
               RECT 21.978 39.582 22.022 39.618 ;
               RECT 21.978 40.182 22.022 40.218 ;
               RECT 21.978 40.782 22.022 40.818 ;
               RECT 21.978 41.382 22.022 41.418 ;
               RECT 21.978 41.982 22.022 42.018 ;
               RECT 21.978 42.582 22.022 42.618 ;
               RECT 21.978 43.182 22.022 43.218 ;
               RECT 21.978 43.782 22.022 43.818 ;
               RECT 21.978 44.382 22.022 44.418 ;
               RECT 21.978 44.982 22.022 45.018 ;
               RECT 21.978 45.582 22.022 45.618 ;
               RECT 21.978 46.182 22.022 46.218 ;
               RECT 21.978 46.782 22.022 46.818 ;
               RECT 21.978 47.382 22.022 47.418 ;
               RECT 21.978 47.982 22.022 48.018 ;
               RECT 21.978 48.582 22.022 48.618 ;
               RECT 21.978 48.942 22.022 48.978 ;
               RECT 21.978 49.422 22.022 49.458 ;
               RECT 21.978 49.902 22.022 49.938 ;
               RECT 21.978 50.382 22.022 50.418 ;
               RECT 21.978 50.862 22.022 50.898 ;
               RECT 21.978 51.342 22.022 51.378 ;
               RECT 21.978 51.822 22.022 51.858 ;
               RECT 21.978 52.302 22.022 52.338 ;
               RECT 21.978 52.782 22.022 52.818 ;
               RECT 21.978 53.262 22.022 53.298 ;
               RECT 21.978 53.742 22.022 53.778 ;
               RECT 21.978 54.222 22.022 54.258 ;
               RECT 21.978 54.702 22.022 54.738 ;
               RECT 21.978 55.182 22.022 55.218 ;
               RECT 21.978 55.662 22.022 55.698 ;
               RECT 21.978 56.142 22.022 56.178 ;
               RECT 21.978 56.502 22.022 56.538 ;
               RECT 21.978 57.102 22.022 57.138 ;
               RECT 21.978 57.702 22.022 57.738 ;
               RECT 21.978 58.302 22.022 58.338 ;
               RECT 21.978 58.902 22.022 58.938 ;
               RECT 21.978 59.502 22.022 59.538 ;
               RECT 21.978 60.102 22.022 60.138 ;
               RECT 21.978 60.702 22.022 60.738 ;
               RECT 21.978 61.302 22.022 61.338 ;
               RECT 21.978 61.902 22.022 61.938 ;
               RECT 21.978 62.502 22.022 62.538 ;
               RECT 21.978 63.102 22.022 63.138 ;
               RECT 21.978 63.702 22.022 63.738 ;
               RECT 21.978 64.302 22.022 64.338 ;
               RECT 21.978 64.902 22.022 64.938 ;
               RECT 21.978 65.502 22.022 65.538 ;
               RECT 21.978 66.102 22.022 66.138 ;
               RECT 21.978 66.702 22.022 66.738 ;
               RECT 21.978 67.302 22.022 67.338 ;
               RECT 21.978 67.902 22.022 67.938 ;
               RECT 21.978 68.502 22.022 68.538 ;
               RECT 21.978 69.102 22.022 69.138 ;
               RECT 21.978 69.702 22.022 69.738 ;
               RECT 21.978 70.302 22.022 70.338 ;
               RECT 21.978 70.902 22.022 70.938 ;
               RECT 21.978 71.502 22.022 71.538 ;
               RECT 21.978 72.102 22.022 72.138 ;
               RECT 21.978 72.702 22.022 72.738 ;
               RECT 21.978 73.302 22.022 73.338 ;
               RECT 21.978 73.902 22.022 73.938 ;
               RECT 21.978 74.502 22.022 74.538 ;
               RECT 21.978 75.102 22.022 75.138 ;
               RECT 21.978 75.702 22.022 75.738 ;
               RECT 21.978 76.302 22.022 76.338 ;
               RECT 21.978 76.902 22.022 76.938 ;
               RECT 21.978 77.502 22.022 77.538 ;
               RECT 21.978 78.102 22.022 78.138 ;
               RECT 21.978 78.702 22.022 78.738 ;
               RECT 21.978 79.302 22.022 79.338 ;
               RECT 21.978 79.902 22.022 79.938 ;
               RECT 21.978 80.502 22.022 80.538 ;
               RECT 21.978 81.102 22.022 81.138 ;
               RECT 21.978 81.702 22.022 81.738 ;
               RECT 21.978 82.302 22.022 82.338 ;
               RECT 21.978 82.902 22.022 82.938 ;
               RECT 21.978 83.502 22.022 83.538 ;
               RECT 21.978 84.102 22.022 84.138 ;
               RECT 21.978 84.702 22.022 84.738 ;
               RECT 21.978 85.302 22.022 85.338 ;
               RECT 21.978 85.902 22.022 85.938 ;
               RECT 21.978 86.502 22.022 86.538 ;
               RECT 21.978 87.102 22.022 87.138 ;
               RECT 21.978 87.702 22.022 87.738 ;
               RECT 21.978 88.302 22.022 88.338 ;
               RECT 21.978 88.902 22.022 88.938 ;
               RECT 21.978 89.502 22.022 89.538 ;
               RECT 21.978 90.102 22.022 90.138 ;
               RECT 21.978 90.702 22.022 90.738 ;
               RECT 21.978 91.302 22.022 91.338 ;
               RECT 21.978 91.902 22.022 91.938 ;
               RECT 21.978 92.502 22.022 92.538 ;
               RECT 21.978 93.102 22.022 93.138 ;
               RECT 21.978 93.702 22.022 93.738 ;
               RECT 21.978 94.302 22.022 94.338 ;
               RECT 21.978 94.902 22.022 94.938 ;
               RECT 21.978 95.502 22.022 95.538 ;
               RECT 21.978 96.102 22.022 96.138 ;
               RECT 21.978 96.702 22.022 96.738 ;
               RECT 21.978 97.302 22.022 97.338 ;
               RECT 21.978 97.902 22.022 97.938 ;
               RECT 21.978 98.502 22.022 98.538 ;
               RECT 21.978 99.102 22.022 99.138 ;
               RECT 21.978 99.702 22.022 99.738 ;
               RECT 21.978 100.302 22.022 100.338 ;
               RECT 21.978 100.902 22.022 100.938 ;
               RECT 21.978 101.502 22.022 101.538 ;
               RECT 21.978 102.102 22.022 102.138 ;
               RECT 21.978 102.702 22.022 102.738 ;
               RECT 21.978 103.302 22.022 103.338 ;
               RECT 21.978 103.902 22.022 103.938 ;
               RECT 21.978 104.502 22.022 104.538 ;
               RECT 22.186 49.8435 22.222 49.8795 ;
               RECT 22.186 50.982 22.222 51.018 ;
               RECT 22.186 54.102 22.222 54.138 ;
               RECT 22.186 55.2405 22.222 55.2765 ;
               RECT 22.614 1.558 22.666 1.594 ;
               RECT 22.614 2.758 22.666 2.794 ;
               RECT 22.614 3.958 22.666 3.994 ;
               RECT 22.614 5.158 22.666 5.194 ;
               RECT 22.614 6.358 22.666 6.394 ;
               RECT 22.614 7.558 22.666 7.594 ;
               RECT 22.614 8.758 22.666 8.794 ;
               RECT 22.614 9.958 22.666 9.994 ;
               RECT 22.614 11.158 22.666 11.194 ;
               RECT 22.614 12.358 22.666 12.394 ;
               RECT 22.614 13.558 22.666 13.594 ;
               RECT 22.614 14.758 22.666 14.794 ;
               RECT 22.614 15.958 22.666 15.994 ;
               RECT 22.614 17.158 22.666 17.194 ;
               RECT 22.614 18.358 22.666 18.394 ;
               RECT 22.614 19.558 22.666 19.594 ;
               RECT 22.614 20.758 22.666 20.794 ;
               RECT 22.614 21.958 22.666 21.994 ;
               RECT 22.614 23.158 22.666 23.194 ;
               RECT 22.614 24.358 22.666 24.394 ;
               RECT 22.614 25.558 22.666 25.594 ;
               RECT 22.614 26.758 22.666 26.794 ;
               RECT 22.614 27.958 22.666 27.994 ;
               RECT 22.614 29.158 22.666 29.194 ;
               RECT 22.614 30.358 22.666 30.394 ;
               RECT 22.614 31.558 22.666 31.594 ;
               RECT 22.614 32.758 22.666 32.794 ;
               RECT 22.614 33.958 22.666 33.994 ;
               RECT 22.614 35.158 22.666 35.194 ;
               RECT 22.614 36.358 22.666 36.394 ;
               RECT 22.614 37.558 22.666 37.594 ;
               RECT 22.614 38.758 22.666 38.794 ;
               RECT 22.614 39.958 22.666 39.994 ;
               RECT 22.614 41.158 22.666 41.194 ;
               RECT 22.614 42.358 22.666 42.394 ;
               RECT 22.614 43.558 22.666 43.594 ;
               RECT 22.614 44.758 22.666 44.794 ;
               RECT 22.614 45.958 22.666 45.994 ;
               RECT 22.614 47.158 22.666 47.194 ;
               RECT 22.614 48.358 22.666 48.394 ;
               RECT 22.614 49.422 22.666 49.458 ;
               RECT 22.614 49.662 22.666 49.698 ;
               RECT 22.614 55.422 22.666 55.458 ;
               RECT 22.614 55.662 22.666 55.698 ;
               RECT 22.614 57.478 22.666 57.514 ;
               RECT 22.614 58.678 22.666 58.714 ;
               RECT 22.614 59.878 22.666 59.914 ;
               RECT 22.614 61.078 22.666 61.114 ;
               RECT 22.614 62.278 22.666 62.314 ;
               RECT 22.614 63.478 22.666 63.514 ;
               RECT 22.614 64.678 22.666 64.714 ;
               RECT 22.614 65.878 22.666 65.914 ;
               RECT 22.614 67.078 22.666 67.114 ;
               RECT 22.614 68.278 22.666 68.314 ;
               RECT 22.614 69.478 22.666 69.514 ;
               RECT 22.614 70.678 22.666 70.714 ;
               RECT 22.614 71.878 22.666 71.914 ;
               RECT 22.614 73.078 22.666 73.114 ;
               RECT 22.614 74.278 22.666 74.314 ;
               RECT 22.614 75.478 22.666 75.514 ;
               RECT 22.614 76.678 22.666 76.714 ;
               RECT 22.614 77.878 22.666 77.914 ;
               RECT 22.614 79.078 22.666 79.114 ;
               RECT 22.614 80.278 22.666 80.314 ;
               RECT 22.614 81.478 22.666 81.514 ;
               RECT 22.614 82.678 22.666 82.714 ;
               RECT 22.614 83.878 22.666 83.914 ;
               RECT 22.614 85.078 22.666 85.114 ;
               RECT 22.614 86.278 22.666 86.314 ;
               RECT 22.614 87.478 22.666 87.514 ;
               RECT 22.614 88.678 22.666 88.714 ;
               RECT 22.614 89.878 22.666 89.914 ;
               RECT 22.614 91.078 22.666 91.114 ;
               RECT 22.614 92.278 22.666 92.314 ;
               RECT 22.614 93.478 22.666 93.514 ;
               RECT 22.614 94.678 22.666 94.714 ;
               RECT 22.614 95.878 22.666 95.914 ;
               RECT 22.614 97.078 22.666 97.114 ;
               RECT 22.614 98.278 22.666 98.314 ;
               RECT 22.614 99.478 22.666 99.514 ;
               RECT 22.614 100.678 22.666 100.714 ;
               RECT 22.614 101.878 22.666 101.914 ;
               RECT 22.614 103.078 22.666 103.114 ;
               RECT 22.614 104.278 22.666 104.314 ;
               RECT 22.694 0.806 22.746 0.842 ;
               RECT 22.694 2.006 22.746 2.042 ;
               RECT 22.694 3.206 22.746 3.242 ;
               RECT 22.694 4.406 22.746 4.442 ;
               RECT 22.694 5.606 22.746 5.642 ;
               RECT 22.694 6.806 22.746 6.842 ;
               RECT 22.694 8.006 22.746 8.042 ;
               RECT 22.694 9.206 22.746 9.242 ;
               RECT 22.694 10.406 22.746 10.442 ;
               RECT 22.694 11.606 22.746 11.642 ;
               RECT 22.694 12.806 22.746 12.842 ;
               RECT 22.694 14.006 22.746 14.042 ;
               RECT 22.694 15.206 22.746 15.242 ;
               RECT 22.694 16.406 22.746 16.442 ;
               RECT 22.694 17.606 22.746 17.642 ;
               RECT 22.694 18.806 22.746 18.842 ;
               RECT 22.694 20.006 22.746 20.042 ;
               RECT 22.694 21.206 22.746 21.242 ;
               RECT 22.694 22.406 22.746 22.442 ;
               RECT 22.694 23.606 22.746 23.642 ;
               RECT 22.694 24.806 22.746 24.842 ;
               RECT 22.694 26.006 22.746 26.042 ;
               RECT 22.694 27.206 22.746 27.242 ;
               RECT 22.694 28.406 22.746 28.442 ;
               RECT 22.694 29.606 22.746 29.642 ;
               RECT 22.694 30.806 22.746 30.842 ;
               RECT 22.694 32.006 22.746 32.042 ;
               RECT 22.694 33.206 22.746 33.242 ;
               RECT 22.694 34.406 22.746 34.442 ;
               RECT 22.694 35.606 22.746 35.642 ;
               RECT 22.694 36.806 22.746 36.842 ;
               RECT 22.694 38.006 22.746 38.042 ;
               RECT 22.694 39.206 22.746 39.242 ;
               RECT 22.694 40.406 22.746 40.442 ;
               RECT 22.694 41.606 22.746 41.642 ;
               RECT 22.694 42.806 22.746 42.842 ;
               RECT 22.694 44.006 22.746 44.042 ;
               RECT 22.694 45.206 22.746 45.242 ;
               RECT 22.694 46.406 22.746 46.442 ;
               RECT 22.694 47.606 22.746 47.642 ;
               RECT 22.694 50.142 22.746 50.178 ;
               RECT 22.694 50.382 22.746 50.418 ;
               RECT 22.694 54.702 22.746 54.738 ;
               RECT 22.694 54.942 22.746 54.978 ;
               RECT 22.694 56.726 22.746 56.762 ;
               RECT 22.694 57.926 22.746 57.962 ;
               RECT 22.694 59.126 22.746 59.162 ;
               RECT 22.694 60.326 22.746 60.362 ;
               RECT 22.694 61.526 22.746 61.562 ;
               RECT 22.694 62.726 22.746 62.762 ;
               RECT 22.694 63.926 22.746 63.962 ;
               RECT 22.694 65.126 22.746 65.162 ;
               RECT 22.694 66.326 22.746 66.362 ;
               RECT 22.694 67.526 22.746 67.562 ;
               RECT 22.694 68.726 22.746 68.762 ;
               RECT 22.694 69.926 22.746 69.962 ;
               RECT 22.694 71.126 22.746 71.162 ;
               RECT 22.694 72.326 22.746 72.362 ;
               RECT 22.694 73.526 22.746 73.562 ;
               RECT 22.694 74.726 22.746 74.762 ;
               RECT 22.694 75.926 22.746 75.962 ;
               RECT 22.694 77.126 22.746 77.162 ;
               RECT 22.694 78.326 22.746 78.362 ;
               RECT 22.694 79.526 22.746 79.562 ;
               RECT 22.694 80.726 22.746 80.762 ;
               RECT 22.694 81.926 22.746 81.962 ;
               RECT 22.694 83.126 22.746 83.162 ;
               RECT 22.694 84.326 22.746 84.362 ;
               RECT 22.694 85.526 22.746 85.562 ;
               RECT 22.694 86.726 22.746 86.762 ;
               RECT 22.694 87.926 22.746 87.962 ;
               RECT 22.694 89.126 22.746 89.162 ;
               RECT 22.694 90.326 22.746 90.362 ;
               RECT 22.694 91.526 22.746 91.562 ;
               RECT 22.694 92.726 22.746 92.762 ;
               RECT 22.694 93.926 22.746 93.962 ;
               RECT 22.694 95.126 22.746 95.162 ;
               RECT 22.694 96.326 22.746 96.362 ;
               RECT 22.694 97.526 22.746 97.562 ;
               RECT 22.694 98.726 22.746 98.762 ;
               RECT 22.694 99.926 22.746 99.962 ;
               RECT 22.694 101.126 22.746 101.162 ;
               RECT 22.694 102.326 22.746 102.362 ;
               RECT 22.694 103.526 22.746 103.562 ;
               RECT 22.774 0.281 22.826 0.317 ;
               RECT 22.774 104.803 22.826 104.839 ;
               RECT 22.854 0.806 22.906 0.842 ;
               RECT 22.854 2.006 22.906 2.042 ;
               RECT 22.854 3.206 22.906 3.242 ;
               RECT 22.854 4.406 22.906 4.442 ;
               RECT 22.854 5.606 22.906 5.642 ;
               RECT 22.854 6.806 22.906 6.842 ;
               RECT 22.854 8.006 22.906 8.042 ;
               RECT 22.854 9.206 22.906 9.242 ;
               RECT 22.854 10.406 22.906 10.442 ;
               RECT 22.854 11.606 22.906 11.642 ;
               RECT 22.854 12.806 22.906 12.842 ;
               RECT 22.854 14.006 22.906 14.042 ;
               RECT 22.854 15.206 22.906 15.242 ;
               RECT 22.854 16.406 22.906 16.442 ;
               RECT 22.854 17.606 22.906 17.642 ;
               RECT 22.854 18.806 22.906 18.842 ;
               RECT 22.854 20.006 22.906 20.042 ;
               RECT 22.854 21.206 22.906 21.242 ;
               RECT 22.854 22.406 22.906 22.442 ;
               RECT 22.854 23.606 22.906 23.642 ;
               RECT 22.854 24.806 22.906 24.842 ;
               RECT 22.854 26.006 22.906 26.042 ;
               RECT 22.854 27.206 22.906 27.242 ;
               RECT 22.854 28.406 22.906 28.442 ;
               RECT 22.854 29.606 22.906 29.642 ;
               RECT 22.854 30.806 22.906 30.842 ;
               RECT 22.854 32.006 22.906 32.042 ;
               RECT 22.854 33.206 22.906 33.242 ;
               RECT 22.854 34.406 22.906 34.442 ;
               RECT 22.854 35.606 22.906 35.642 ;
               RECT 22.854 36.806 22.906 36.842 ;
               RECT 22.854 38.006 22.906 38.042 ;
               RECT 22.854 39.206 22.906 39.242 ;
               RECT 22.854 40.406 22.906 40.442 ;
               RECT 22.854 41.606 22.906 41.642 ;
               RECT 22.854 42.806 22.906 42.842 ;
               RECT 22.854 44.006 22.906 44.042 ;
               RECT 22.854 45.206 22.906 45.242 ;
               RECT 22.854 46.406 22.906 46.442 ;
               RECT 22.854 47.606 22.906 47.642 ;
               RECT 22.854 49.422 22.906 49.458 ;
               RECT 22.854 49.662 22.906 49.698 ;
               RECT 22.854 55.422 22.906 55.458 ;
               RECT 22.854 55.662 22.906 55.698 ;
               RECT 22.854 56.726 22.906 56.762 ;
               RECT 22.854 57.926 22.906 57.962 ;
               RECT 22.854 59.126 22.906 59.162 ;
               RECT 22.854 60.326 22.906 60.362 ;
               RECT 22.854 61.526 22.906 61.562 ;
               RECT 22.854 62.726 22.906 62.762 ;
               RECT 22.854 63.926 22.906 63.962 ;
               RECT 22.854 65.126 22.906 65.162 ;
               RECT 22.854 66.326 22.906 66.362 ;
               RECT 22.854 67.526 22.906 67.562 ;
               RECT 22.854 68.726 22.906 68.762 ;
               RECT 22.854 69.926 22.906 69.962 ;
               RECT 22.854 71.126 22.906 71.162 ;
               RECT 22.854 72.326 22.906 72.362 ;
               RECT 22.854 73.526 22.906 73.562 ;
               RECT 22.854 74.726 22.906 74.762 ;
               RECT 22.854 75.926 22.906 75.962 ;
               RECT 22.854 77.126 22.906 77.162 ;
               RECT 22.854 78.326 22.906 78.362 ;
               RECT 22.854 79.526 22.906 79.562 ;
               RECT 22.854 80.726 22.906 80.762 ;
               RECT 22.854 81.926 22.906 81.962 ;
               RECT 22.854 83.126 22.906 83.162 ;
               RECT 22.854 84.326 22.906 84.362 ;
               RECT 22.854 85.526 22.906 85.562 ;
               RECT 22.854 86.726 22.906 86.762 ;
               RECT 22.854 87.926 22.906 87.962 ;
               RECT 22.854 89.126 22.906 89.162 ;
               RECT 22.854 90.326 22.906 90.362 ;
               RECT 22.854 91.526 22.906 91.562 ;
               RECT 22.854 92.726 22.906 92.762 ;
               RECT 22.854 93.926 22.906 93.962 ;
               RECT 22.854 95.126 22.906 95.162 ;
               RECT 22.854 96.326 22.906 96.362 ;
               RECT 22.854 97.526 22.906 97.562 ;
               RECT 22.854 98.726 22.906 98.762 ;
               RECT 22.854 99.926 22.906 99.962 ;
               RECT 22.854 101.126 22.906 101.162 ;
               RECT 22.854 102.326 22.906 102.362 ;
               RECT 22.854 103.526 22.906 103.562 ;
               RECT 22.934 1.558 22.986 1.594 ;
               RECT 22.934 2.758 22.986 2.794 ;
               RECT 22.934 3.958 22.986 3.994 ;
               RECT 22.934 5.158 22.986 5.194 ;
               RECT 22.934 6.358 22.986 6.394 ;
               RECT 22.934 7.558 22.986 7.594 ;
               RECT 22.934 8.758 22.986 8.794 ;
               RECT 22.934 9.958 22.986 9.994 ;
               RECT 22.934 11.158 22.986 11.194 ;
               RECT 22.934 12.358 22.986 12.394 ;
               RECT 22.934 13.558 22.986 13.594 ;
               RECT 22.934 14.758 22.986 14.794 ;
               RECT 22.934 15.958 22.986 15.994 ;
               RECT 22.934 17.158 22.986 17.194 ;
               RECT 22.934 18.358 22.986 18.394 ;
               RECT 22.934 19.558 22.986 19.594 ;
               RECT 22.934 20.758 22.986 20.794 ;
               RECT 22.934 21.958 22.986 21.994 ;
               RECT 22.934 23.158 22.986 23.194 ;
               RECT 22.934 24.358 22.986 24.394 ;
               RECT 22.934 25.558 22.986 25.594 ;
               RECT 22.934 26.758 22.986 26.794 ;
               RECT 22.934 27.958 22.986 27.994 ;
               RECT 22.934 29.158 22.986 29.194 ;
               RECT 22.934 30.358 22.986 30.394 ;
               RECT 22.934 31.558 22.986 31.594 ;
               RECT 22.934 32.758 22.986 32.794 ;
               RECT 22.934 33.958 22.986 33.994 ;
               RECT 22.934 35.158 22.986 35.194 ;
               RECT 22.934 36.358 22.986 36.394 ;
               RECT 22.934 37.558 22.986 37.594 ;
               RECT 22.934 38.758 22.986 38.794 ;
               RECT 22.934 39.958 22.986 39.994 ;
               RECT 22.934 41.158 22.986 41.194 ;
               RECT 22.934 42.358 22.986 42.394 ;
               RECT 22.934 43.558 22.986 43.594 ;
               RECT 22.934 44.758 22.986 44.794 ;
               RECT 22.934 45.958 22.986 45.994 ;
               RECT 22.934 47.158 22.986 47.194 ;
               RECT 22.934 48.358 22.986 48.394 ;
               RECT 22.934 50.142 22.986 50.178 ;
               RECT 22.934 50.382 22.986 50.418 ;
               RECT 22.934 54.702 22.986 54.738 ;
               RECT 22.934 54.942 22.986 54.978 ;
               RECT 22.934 57.478 22.986 57.514 ;
               RECT 22.934 58.678 22.986 58.714 ;
               RECT 22.934 59.878 22.986 59.914 ;
               RECT 22.934 61.078 22.986 61.114 ;
               RECT 22.934 62.278 22.986 62.314 ;
               RECT 22.934 63.478 22.986 63.514 ;
               RECT 22.934 64.678 22.986 64.714 ;
               RECT 22.934 65.878 22.986 65.914 ;
               RECT 22.934 67.078 22.986 67.114 ;
               RECT 22.934 68.278 22.986 68.314 ;
               RECT 22.934 69.478 22.986 69.514 ;
               RECT 22.934 70.678 22.986 70.714 ;
               RECT 22.934 71.878 22.986 71.914 ;
               RECT 22.934 73.078 22.986 73.114 ;
               RECT 22.934 74.278 22.986 74.314 ;
               RECT 22.934 75.478 22.986 75.514 ;
               RECT 22.934 76.678 22.986 76.714 ;
               RECT 22.934 77.878 22.986 77.914 ;
               RECT 22.934 79.078 22.986 79.114 ;
               RECT 22.934 80.278 22.986 80.314 ;
               RECT 22.934 81.478 22.986 81.514 ;
               RECT 22.934 82.678 22.986 82.714 ;
               RECT 22.934 83.878 22.986 83.914 ;
               RECT 22.934 85.078 22.986 85.114 ;
               RECT 22.934 86.278 22.986 86.314 ;
               RECT 22.934 87.478 22.986 87.514 ;
               RECT 22.934 88.678 22.986 88.714 ;
               RECT 22.934 89.878 22.986 89.914 ;
               RECT 22.934 91.078 22.986 91.114 ;
               RECT 22.934 92.278 22.986 92.314 ;
               RECT 22.934 93.478 22.986 93.514 ;
               RECT 22.934 94.678 22.986 94.714 ;
               RECT 22.934 95.878 22.986 95.914 ;
               RECT 22.934 97.078 22.986 97.114 ;
               RECT 22.934 98.278 22.986 98.314 ;
               RECT 22.934 99.478 22.986 99.514 ;
               RECT 22.934 100.678 22.986 100.714 ;
               RECT 22.934 101.878 22.986 101.914 ;
               RECT 22.934 103.078 22.986 103.114 ;
               RECT 22.934 104.278 22.986 104.314 ;
               RECT 23.014 0.806 23.066 0.842 ;
               RECT 23.014 2.006 23.066 2.042 ;
               RECT 23.014 3.206 23.066 3.242 ;
               RECT 23.014 4.406 23.066 4.442 ;
               RECT 23.014 5.606 23.066 5.642 ;
               RECT 23.014 6.806 23.066 6.842 ;
               RECT 23.014 8.006 23.066 8.042 ;
               RECT 23.014 9.206 23.066 9.242 ;
               RECT 23.014 10.406 23.066 10.442 ;
               RECT 23.014 11.606 23.066 11.642 ;
               RECT 23.014 12.806 23.066 12.842 ;
               RECT 23.014 14.006 23.066 14.042 ;
               RECT 23.014 15.206 23.066 15.242 ;
               RECT 23.014 16.406 23.066 16.442 ;
               RECT 23.014 17.606 23.066 17.642 ;
               RECT 23.014 18.806 23.066 18.842 ;
               RECT 23.014 20.006 23.066 20.042 ;
               RECT 23.014 21.206 23.066 21.242 ;
               RECT 23.014 22.406 23.066 22.442 ;
               RECT 23.014 23.606 23.066 23.642 ;
               RECT 23.014 24.806 23.066 24.842 ;
               RECT 23.014 26.006 23.066 26.042 ;
               RECT 23.014 27.206 23.066 27.242 ;
               RECT 23.014 28.406 23.066 28.442 ;
               RECT 23.014 29.606 23.066 29.642 ;
               RECT 23.014 30.806 23.066 30.842 ;
               RECT 23.014 32.006 23.066 32.042 ;
               RECT 23.014 33.206 23.066 33.242 ;
               RECT 23.014 34.406 23.066 34.442 ;
               RECT 23.014 35.606 23.066 35.642 ;
               RECT 23.014 36.806 23.066 36.842 ;
               RECT 23.014 38.006 23.066 38.042 ;
               RECT 23.014 39.206 23.066 39.242 ;
               RECT 23.014 40.406 23.066 40.442 ;
               RECT 23.014 41.606 23.066 41.642 ;
               RECT 23.014 42.806 23.066 42.842 ;
               RECT 23.014 44.006 23.066 44.042 ;
               RECT 23.014 45.206 23.066 45.242 ;
               RECT 23.014 46.406 23.066 46.442 ;
               RECT 23.014 47.606 23.066 47.642 ;
               RECT 23.014 49.422 23.066 49.458 ;
               RECT 23.014 49.662 23.066 49.698 ;
               RECT 23.014 55.422 23.066 55.458 ;
               RECT 23.014 55.662 23.066 55.698 ;
               RECT 23.014 56.726 23.066 56.762 ;
               RECT 23.014 57.926 23.066 57.962 ;
               RECT 23.014 59.126 23.066 59.162 ;
               RECT 23.014 60.326 23.066 60.362 ;
               RECT 23.014 61.526 23.066 61.562 ;
               RECT 23.014 62.726 23.066 62.762 ;
               RECT 23.014 63.926 23.066 63.962 ;
               RECT 23.014 65.126 23.066 65.162 ;
               RECT 23.014 66.326 23.066 66.362 ;
               RECT 23.014 67.526 23.066 67.562 ;
               RECT 23.014 68.726 23.066 68.762 ;
               RECT 23.014 69.926 23.066 69.962 ;
               RECT 23.014 71.126 23.066 71.162 ;
               RECT 23.014 72.326 23.066 72.362 ;
               RECT 23.014 73.526 23.066 73.562 ;
               RECT 23.014 74.726 23.066 74.762 ;
               RECT 23.014 75.926 23.066 75.962 ;
               RECT 23.014 77.126 23.066 77.162 ;
               RECT 23.014 78.326 23.066 78.362 ;
               RECT 23.014 79.526 23.066 79.562 ;
               RECT 23.014 80.726 23.066 80.762 ;
               RECT 23.014 81.926 23.066 81.962 ;
               RECT 23.014 83.126 23.066 83.162 ;
               RECT 23.014 84.326 23.066 84.362 ;
               RECT 23.014 85.526 23.066 85.562 ;
               RECT 23.014 86.726 23.066 86.762 ;
               RECT 23.014 87.926 23.066 87.962 ;
               RECT 23.014 89.126 23.066 89.162 ;
               RECT 23.014 90.326 23.066 90.362 ;
               RECT 23.014 91.526 23.066 91.562 ;
               RECT 23.014 92.726 23.066 92.762 ;
               RECT 23.014 93.926 23.066 93.962 ;
               RECT 23.014 95.126 23.066 95.162 ;
               RECT 23.014 96.326 23.066 96.362 ;
               RECT 23.014 97.526 23.066 97.562 ;
               RECT 23.014 98.726 23.066 98.762 ;
               RECT 23.014 99.926 23.066 99.962 ;
               RECT 23.014 101.126 23.066 101.162 ;
               RECT 23.014 102.326 23.066 102.362 ;
               RECT 23.014 103.526 23.066 103.562 ;
               RECT 23.094 1.558 23.146 1.594 ;
               RECT 23.094 2.758 23.146 2.794 ;
               RECT 23.094 3.958 23.146 3.994 ;
               RECT 23.094 5.158 23.146 5.194 ;
               RECT 23.094 6.358 23.146 6.394 ;
               RECT 23.094 7.558 23.146 7.594 ;
               RECT 23.094 8.758 23.146 8.794 ;
               RECT 23.094 9.958 23.146 9.994 ;
               RECT 23.094 11.158 23.146 11.194 ;
               RECT 23.094 12.358 23.146 12.394 ;
               RECT 23.094 13.558 23.146 13.594 ;
               RECT 23.094 14.758 23.146 14.794 ;
               RECT 23.094 15.958 23.146 15.994 ;
               RECT 23.094 17.158 23.146 17.194 ;
               RECT 23.094 18.358 23.146 18.394 ;
               RECT 23.094 19.558 23.146 19.594 ;
               RECT 23.094 20.758 23.146 20.794 ;
               RECT 23.094 21.958 23.146 21.994 ;
               RECT 23.094 23.158 23.146 23.194 ;
               RECT 23.094 24.358 23.146 24.394 ;
               RECT 23.094 25.558 23.146 25.594 ;
               RECT 23.094 26.758 23.146 26.794 ;
               RECT 23.094 27.958 23.146 27.994 ;
               RECT 23.094 29.158 23.146 29.194 ;
               RECT 23.094 30.358 23.146 30.394 ;
               RECT 23.094 31.558 23.146 31.594 ;
               RECT 23.094 32.758 23.146 32.794 ;
               RECT 23.094 33.958 23.146 33.994 ;
               RECT 23.094 35.158 23.146 35.194 ;
               RECT 23.094 36.358 23.146 36.394 ;
               RECT 23.094 37.558 23.146 37.594 ;
               RECT 23.094 38.758 23.146 38.794 ;
               RECT 23.094 39.958 23.146 39.994 ;
               RECT 23.094 41.158 23.146 41.194 ;
               RECT 23.094 42.358 23.146 42.394 ;
               RECT 23.094 43.558 23.146 43.594 ;
               RECT 23.094 44.758 23.146 44.794 ;
               RECT 23.094 45.958 23.146 45.994 ;
               RECT 23.094 47.158 23.146 47.194 ;
               RECT 23.094 48.358 23.146 48.394 ;
               RECT 23.094 50.142 23.146 50.178 ;
               RECT 23.094 50.382 23.146 50.418 ;
               RECT 23.094 54.702 23.146 54.738 ;
               RECT 23.094 54.942 23.146 54.978 ;
               RECT 23.094 57.478 23.146 57.514 ;
               RECT 23.094 58.678 23.146 58.714 ;
               RECT 23.094 59.878 23.146 59.914 ;
               RECT 23.094 61.078 23.146 61.114 ;
               RECT 23.094 62.278 23.146 62.314 ;
               RECT 23.094 63.478 23.146 63.514 ;
               RECT 23.094 64.678 23.146 64.714 ;
               RECT 23.094 65.878 23.146 65.914 ;
               RECT 23.094 67.078 23.146 67.114 ;
               RECT 23.094 68.278 23.146 68.314 ;
               RECT 23.094 69.478 23.146 69.514 ;
               RECT 23.094 70.678 23.146 70.714 ;
               RECT 23.094 71.878 23.146 71.914 ;
               RECT 23.094 73.078 23.146 73.114 ;
               RECT 23.094 74.278 23.146 74.314 ;
               RECT 23.094 75.478 23.146 75.514 ;
               RECT 23.094 76.678 23.146 76.714 ;
               RECT 23.094 77.878 23.146 77.914 ;
               RECT 23.094 79.078 23.146 79.114 ;
               RECT 23.094 80.278 23.146 80.314 ;
               RECT 23.094 81.478 23.146 81.514 ;
               RECT 23.094 82.678 23.146 82.714 ;
               RECT 23.094 83.878 23.146 83.914 ;
               RECT 23.094 85.078 23.146 85.114 ;
               RECT 23.094 86.278 23.146 86.314 ;
               RECT 23.094 87.478 23.146 87.514 ;
               RECT 23.094 88.678 23.146 88.714 ;
               RECT 23.094 89.878 23.146 89.914 ;
               RECT 23.094 91.078 23.146 91.114 ;
               RECT 23.094 92.278 23.146 92.314 ;
               RECT 23.094 93.478 23.146 93.514 ;
               RECT 23.094 94.678 23.146 94.714 ;
               RECT 23.094 95.878 23.146 95.914 ;
               RECT 23.094 97.078 23.146 97.114 ;
               RECT 23.094 98.278 23.146 98.314 ;
               RECT 23.094 99.478 23.146 99.514 ;
               RECT 23.094 100.678 23.146 100.714 ;
               RECT 23.094 101.878 23.146 101.914 ;
               RECT 23.094 103.078 23.146 103.114 ;
               RECT 23.094 104.278 23.146 104.314 ;
               RECT 23.174 0.281 23.226 0.317 ;
               RECT 23.174 104.803 23.226 104.839 ;
               RECT 23.254 0.806 23.306 0.842 ;
               RECT 23.254 2.006 23.306 2.042 ;
               RECT 23.254 3.206 23.306 3.242 ;
               RECT 23.254 4.406 23.306 4.442 ;
               RECT 23.254 5.606 23.306 5.642 ;
               RECT 23.254 6.806 23.306 6.842 ;
               RECT 23.254 8.006 23.306 8.042 ;
               RECT 23.254 9.206 23.306 9.242 ;
               RECT 23.254 10.406 23.306 10.442 ;
               RECT 23.254 11.606 23.306 11.642 ;
               RECT 23.254 12.806 23.306 12.842 ;
               RECT 23.254 14.006 23.306 14.042 ;
               RECT 23.254 15.206 23.306 15.242 ;
               RECT 23.254 16.406 23.306 16.442 ;
               RECT 23.254 17.606 23.306 17.642 ;
               RECT 23.254 18.806 23.306 18.842 ;
               RECT 23.254 20.006 23.306 20.042 ;
               RECT 23.254 21.206 23.306 21.242 ;
               RECT 23.254 22.406 23.306 22.442 ;
               RECT 23.254 23.606 23.306 23.642 ;
               RECT 23.254 24.806 23.306 24.842 ;
               RECT 23.254 26.006 23.306 26.042 ;
               RECT 23.254 27.206 23.306 27.242 ;
               RECT 23.254 28.406 23.306 28.442 ;
               RECT 23.254 29.606 23.306 29.642 ;
               RECT 23.254 30.806 23.306 30.842 ;
               RECT 23.254 32.006 23.306 32.042 ;
               RECT 23.254 33.206 23.306 33.242 ;
               RECT 23.254 34.406 23.306 34.442 ;
               RECT 23.254 35.606 23.306 35.642 ;
               RECT 23.254 36.806 23.306 36.842 ;
               RECT 23.254 38.006 23.306 38.042 ;
               RECT 23.254 39.206 23.306 39.242 ;
               RECT 23.254 40.406 23.306 40.442 ;
               RECT 23.254 41.606 23.306 41.642 ;
               RECT 23.254 42.806 23.306 42.842 ;
               RECT 23.254 44.006 23.306 44.042 ;
               RECT 23.254 45.206 23.306 45.242 ;
               RECT 23.254 46.406 23.306 46.442 ;
               RECT 23.254 47.606 23.306 47.642 ;
               RECT 23.254 49.422 23.306 49.458 ;
               RECT 23.254 49.662 23.306 49.698 ;
               RECT 23.254 51.102 23.306 51.138 ;
               RECT 23.254 51.582 23.306 51.618 ;
               RECT 23.254 53.502 23.306 53.538 ;
               RECT 23.254 53.982 23.306 54.018 ;
               RECT 23.254 55.422 23.306 55.458 ;
               RECT 23.254 55.662 23.306 55.698 ;
               RECT 23.254 56.726 23.306 56.762 ;
               RECT 23.254 57.926 23.306 57.962 ;
               RECT 23.254 59.126 23.306 59.162 ;
               RECT 23.254 60.326 23.306 60.362 ;
               RECT 23.254 61.526 23.306 61.562 ;
               RECT 23.254 62.726 23.306 62.762 ;
               RECT 23.254 63.926 23.306 63.962 ;
               RECT 23.254 65.126 23.306 65.162 ;
               RECT 23.254 66.326 23.306 66.362 ;
               RECT 23.254 67.526 23.306 67.562 ;
               RECT 23.254 68.726 23.306 68.762 ;
               RECT 23.254 69.926 23.306 69.962 ;
               RECT 23.254 71.126 23.306 71.162 ;
               RECT 23.254 72.326 23.306 72.362 ;
               RECT 23.254 73.526 23.306 73.562 ;
               RECT 23.254 74.726 23.306 74.762 ;
               RECT 23.254 75.926 23.306 75.962 ;
               RECT 23.254 77.126 23.306 77.162 ;
               RECT 23.254 78.326 23.306 78.362 ;
               RECT 23.254 79.526 23.306 79.562 ;
               RECT 23.254 80.726 23.306 80.762 ;
               RECT 23.254 81.926 23.306 81.962 ;
               RECT 23.254 83.126 23.306 83.162 ;
               RECT 23.254 84.326 23.306 84.362 ;
               RECT 23.254 85.526 23.306 85.562 ;
               RECT 23.254 86.726 23.306 86.762 ;
               RECT 23.254 87.926 23.306 87.962 ;
               RECT 23.254 89.126 23.306 89.162 ;
               RECT 23.254 90.326 23.306 90.362 ;
               RECT 23.254 91.526 23.306 91.562 ;
               RECT 23.254 92.726 23.306 92.762 ;
               RECT 23.254 93.926 23.306 93.962 ;
               RECT 23.254 95.126 23.306 95.162 ;
               RECT 23.254 96.326 23.306 96.362 ;
               RECT 23.254 97.526 23.306 97.562 ;
               RECT 23.254 98.726 23.306 98.762 ;
               RECT 23.254 99.926 23.306 99.962 ;
               RECT 23.254 101.126 23.306 101.162 ;
               RECT 23.254 102.326 23.306 102.362 ;
               RECT 23.254 103.526 23.306 103.562 ;
               RECT 23.334 1.558 23.386 1.594 ;
               RECT 23.334 2.758 23.386 2.794 ;
               RECT 23.334 3.958 23.386 3.994 ;
               RECT 23.334 5.158 23.386 5.194 ;
               RECT 23.334 6.358 23.386 6.394 ;
               RECT 23.334 7.558 23.386 7.594 ;
               RECT 23.334 8.758 23.386 8.794 ;
               RECT 23.334 9.958 23.386 9.994 ;
               RECT 23.334 11.158 23.386 11.194 ;
               RECT 23.334 12.358 23.386 12.394 ;
               RECT 23.334 13.558 23.386 13.594 ;
               RECT 23.334 14.758 23.386 14.794 ;
               RECT 23.334 15.958 23.386 15.994 ;
               RECT 23.334 17.158 23.386 17.194 ;
               RECT 23.334 18.358 23.386 18.394 ;
               RECT 23.334 19.558 23.386 19.594 ;
               RECT 23.334 20.758 23.386 20.794 ;
               RECT 23.334 21.958 23.386 21.994 ;
               RECT 23.334 23.158 23.386 23.194 ;
               RECT 23.334 24.358 23.386 24.394 ;
               RECT 23.334 25.558 23.386 25.594 ;
               RECT 23.334 26.758 23.386 26.794 ;
               RECT 23.334 27.958 23.386 27.994 ;
               RECT 23.334 29.158 23.386 29.194 ;
               RECT 23.334 30.358 23.386 30.394 ;
               RECT 23.334 31.558 23.386 31.594 ;
               RECT 23.334 32.758 23.386 32.794 ;
               RECT 23.334 33.958 23.386 33.994 ;
               RECT 23.334 35.158 23.386 35.194 ;
               RECT 23.334 36.358 23.386 36.394 ;
               RECT 23.334 37.558 23.386 37.594 ;
               RECT 23.334 38.758 23.386 38.794 ;
               RECT 23.334 39.958 23.386 39.994 ;
               RECT 23.334 41.158 23.386 41.194 ;
               RECT 23.334 42.358 23.386 42.394 ;
               RECT 23.334 43.558 23.386 43.594 ;
               RECT 23.334 44.758 23.386 44.794 ;
               RECT 23.334 45.958 23.386 45.994 ;
               RECT 23.334 47.158 23.386 47.194 ;
               RECT 23.334 48.358 23.386 48.394 ;
               RECT 23.334 50.142 23.386 50.178 ;
               RECT 23.334 50.382 23.386 50.418 ;
               RECT 23.334 54.702 23.386 54.738 ;
               RECT 23.334 54.942 23.386 54.978 ;
               RECT 23.334 57.478 23.386 57.514 ;
               RECT 23.334 58.678 23.386 58.714 ;
               RECT 23.334 59.878 23.386 59.914 ;
               RECT 23.334 61.078 23.386 61.114 ;
               RECT 23.334 62.278 23.386 62.314 ;
               RECT 23.334 63.478 23.386 63.514 ;
               RECT 23.334 64.678 23.386 64.714 ;
               RECT 23.334 65.878 23.386 65.914 ;
               RECT 23.334 67.078 23.386 67.114 ;
               RECT 23.334 68.278 23.386 68.314 ;
               RECT 23.334 69.478 23.386 69.514 ;
               RECT 23.334 70.678 23.386 70.714 ;
               RECT 23.334 71.878 23.386 71.914 ;
               RECT 23.334 73.078 23.386 73.114 ;
               RECT 23.334 74.278 23.386 74.314 ;
               RECT 23.334 75.478 23.386 75.514 ;
               RECT 23.334 76.678 23.386 76.714 ;
               RECT 23.334 77.878 23.386 77.914 ;
               RECT 23.334 79.078 23.386 79.114 ;
               RECT 23.334 80.278 23.386 80.314 ;
               RECT 23.334 81.478 23.386 81.514 ;
               RECT 23.334 82.678 23.386 82.714 ;
               RECT 23.334 83.878 23.386 83.914 ;
               RECT 23.334 85.078 23.386 85.114 ;
               RECT 23.334 86.278 23.386 86.314 ;
               RECT 23.334 87.478 23.386 87.514 ;
               RECT 23.334 88.678 23.386 88.714 ;
               RECT 23.334 89.878 23.386 89.914 ;
               RECT 23.334 91.078 23.386 91.114 ;
               RECT 23.334 92.278 23.386 92.314 ;
               RECT 23.334 93.478 23.386 93.514 ;
               RECT 23.334 94.678 23.386 94.714 ;
               RECT 23.334 95.878 23.386 95.914 ;
               RECT 23.334 97.078 23.386 97.114 ;
               RECT 23.334 98.278 23.386 98.314 ;
               RECT 23.334 99.478 23.386 99.514 ;
               RECT 23.334 100.678 23.386 100.714 ;
               RECT 23.334 101.878 23.386 101.914 ;
               RECT 23.334 103.078 23.386 103.114 ;
               RECT 23.334 104.278 23.386 104.314 ;
               RECT 23.414 0.806 23.466 0.842 ;
               RECT 23.414 2.006 23.466 2.042 ;
               RECT 23.414 3.206 23.466 3.242 ;
               RECT 23.414 4.406 23.466 4.442 ;
               RECT 23.414 5.606 23.466 5.642 ;
               RECT 23.414 6.806 23.466 6.842 ;
               RECT 23.414 8.006 23.466 8.042 ;
               RECT 23.414 9.206 23.466 9.242 ;
               RECT 23.414 10.406 23.466 10.442 ;
               RECT 23.414 11.606 23.466 11.642 ;
               RECT 23.414 12.806 23.466 12.842 ;
               RECT 23.414 14.006 23.466 14.042 ;
               RECT 23.414 15.206 23.466 15.242 ;
               RECT 23.414 16.406 23.466 16.442 ;
               RECT 23.414 17.606 23.466 17.642 ;
               RECT 23.414 18.806 23.466 18.842 ;
               RECT 23.414 20.006 23.466 20.042 ;
               RECT 23.414 21.206 23.466 21.242 ;
               RECT 23.414 22.406 23.466 22.442 ;
               RECT 23.414 23.606 23.466 23.642 ;
               RECT 23.414 24.806 23.466 24.842 ;
               RECT 23.414 26.006 23.466 26.042 ;
               RECT 23.414 27.206 23.466 27.242 ;
               RECT 23.414 28.406 23.466 28.442 ;
               RECT 23.414 29.606 23.466 29.642 ;
               RECT 23.414 30.806 23.466 30.842 ;
               RECT 23.414 32.006 23.466 32.042 ;
               RECT 23.414 33.206 23.466 33.242 ;
               RECT 23.414 34.406 23.466 34.442 ;
               RECT 23.414 35.606 23.466 35.642 ;
               RECT 23.414 36.806 23.466 36.842 ;
               RECT 23.414 38.006 23.466 38.042 ;
               RECT 23.414 39.206 23.466 39.242 ;
               RECT 23.414 40.406 23.466 40.442 ;
               RECT 23.414 41.606 23.466 41.642 ;
               RECT 23.414 42.806 23.466 42.842 ;
               RECT 23.414 44.006 23.466 44.042 ;
               RECT 23.414 45.206 23.466 45.242 ;
               RECT 23.414 46.406 23.466 46.442 ;
               RECT 23.414 47.606 23.466 47.642 ;
               RECT 23.414 49.422 23.466 49.458 ;
               RECT 23.414 49.662 23.466 49.698 ;
               RECT 23.414 55.422 23.466 55.458 ;
               RECT 23.414 55.662 23.466 55.698 ;
               RECT 23.414 56.726 23.466 56.762 ;
               RECT 23.414 57.926 23.466 57.962 ;
               RECT 23.414 59.126 23.466 59.162 ;
               RECT 23.414 60.326 23.466 60.362 ;
               RECT 23.414 61.526 23.466 61.562 ;
               RECT 23.414 62.726 23.466 62.762 ;
               RECT 23.414 63.926 23.466 63.962 ;
               RECT 23.414 65.126 23.466 65.162 ;
               RECT 23.414 66.326 23.466 66.362 ;
               RECT 23.414 67.526 23.466 67.562 ;
               RECT 23.414 68.726 23.466 68.762 ;
               RECT 23.414 69.926 23.466 69.962 ;
               RECT 23.414 71.126 23.466 71.162 ;
               RECT 23.414 72.326 23.466 72.362 ;
               RECT 23.414 73.526 23.466 73.562 ;
               RECT 23.414 74.726 23.466 74.762 ;
               RECT 23.414 75.926 23.466 75.962 ;
               RECT 23.414 77.126 23.466 77.162 ;
               RECT 23.414 78.326 23.466 78.362 ;
               RECT 23.414 79.526 23.466 79.562 ;
               RECT 23.414 80.726 23.466 80.762 ;
               RECT 23.414 81.926 23.466 81.962 ;
               RECT 23.414 83.126 23.466 83.162 ;
               RECT 23.414 84.326 23.466 84.362 ;
               RECT 23.414 85.526 23.466 85.562 ;
               RECT 23.414 86.726 23.466 86.762 ;
               RECT 23.414 87.926 23.466 87.962 ;
               RECT 23.414 89.126 23.466 89.162 ;
               RECT 23.414 90.326 23.466 90.362 ;
               RECT 23.414 91.526 23.466 91.562 ;
               RECT 23.414 92.726 23.466 92.762 ;
               RECT 23.414 93.926 23.466 93.962 ;
               RECT 23.414 95.126 23.466 95.162 ;
               RECT 23.414 96.326 23.466 96.362 ;
               RECT 23.414 97.526 23.466 97.562 ;
               RECT 23.414 98.726 23.466 98.762 ;
               RECT 23.414 99.926 23.466 99.962 ;
               RECT 23.414 101.126 23.466 101.162 ;
               RECT 23.414 102.326 23.466 102.362 ;
               RECT 23.414 103.526 23.466 103.562 ;
               RECT 23.494 1.558 23.546 1.594 ;
               RECT 23.494 2.758 23.546 2.794 ;
               RECT 23.494 3.958 23.546 3.994 ;
               RECT 23.494 5.158 23.546 5.194 ;
               RECT 23.494 6.358 23.546 6.394 ;
               RECT 23.494 7.558 23.546 7.594 ;
               RECT 23.494 8.758 23.546 8.794 ;
               RECT 23.494 9.958 23.546 9.994 ;
               RECT 23.494 11.158 23.546 11.194 ;
               RECT 23.494 12.358 23.546 12.394 ;
               RECT 23.494 13.558 23.546 13.594 ;
               RECT 23.494 14.758 23.546 14.794 ;
               RECT 23.494 15.958 23.546 15.994 ;
               RECT 23.494 17.158 23.546 17.194 ;
               RECT 23.494 18.358 23.546 18.394 ;
               RECT 23.494 19.558 23.546 19.594 ;
               RECT 23.494 20.758 23.546 20.794 ;
               RECT 23.494 21.958 23.546 21.994 ;
               RECT 23.494 23.158 23.546 23.194 ;
               RECT 23.494 24.358 23.546 24.394 ;
               RECT 23.494 25.558 23.546 25.594 ;
               RECT 23.494 26.758 23.546 26.794 ;
               RECT 23.494 27.958 23.546 27.994 ;
               RECT 23.494 29.158 23.546 29.194 ;
               RECT 23.494 30.358 23.546 30.394 ;
               RECT 23.494 31.558 23.546 31.594 ;
               RECT 23.494 32.758 23.546 32.794 ;
               RECT 23.494 33.958 23.546 33.994 ;
               RECT 23.494 35.158 23.546 35.194 ;
               RECT 23.494 36.358 23.546 36.394 ;
               RECT 23.494 37.558 23.546 37.594 ;
               RECT 23.494 38.758 23.546 38.794 ;
               RECT 23.494 39.958 23.546 39.994 ;
               RECT 23.494 41.158 23.546 41.194 ;
               RECT 23.494 42.358 23.546 42.394 ;
               RECT 23.494 43.558 23.546 43.594 ;
               RECT 23.494 44.758 23.546 44.794 ;
               RECT 23.494 45.958 23.546 45.994 ;
               RECT 23.494 47.158 23.546 47.194 ;
               RECT 23.494 48.358 23.546 48.394 ;
               RECT 23.494 50.142 23.546 50.178 ;
               RECT 23.494 50.382 23.546 50.418 ;
               RECT 23.494 54.702 23.546 54.738 ;
               RECT 23.494 54.942 23.546 54.978 ;
               RECT 23.494 57.478 23.546 57.514 ;
               RECT 23.494 58.678 23.546 58.714 ;
               RECT 23.494 59.878 23.546 59.914 ;
               RECT 23.494 61.078 23.546 61.114 ;
               RECT 23.494 62.278 23.546 62.314 ;
               RECT 23.494 63.478 23.546 63.514 ;
               RECT 23.494 64.678 23.546 64.714 ;
               RECT 23.494 65.878 23.546 65.914 ;
               RECT 23.494 67.078 23.546 67.114 ;
               RECT 23.494 68.278 23.546 68.314 ;
               RECT 23.494 69.478 23.546 69.514 ;
               RECT 23.494 70.678 23.546 70.714 ;
               RECT 23.494 71.878 23.546 71.914 ;
               RECT 23.494 73.078 23.546 73.114 ;
               RECT 23.494 74.278 23.546 74.314 ;
               RECT 23.494 75.478 23.546 75.514 ;
               RECT 23.494 76.678 23.546 76.714 ;
               RECT 23.494 77.878 23.546 77.914 ;
               RECT 23.494 79.078 23.546 79.114 ;
               RECT 23.494 80.278 23.546 80.314 ;
               RECT 23.494 81.478 23.546 81.514 ;
               RECT 23.494 82.678 23.546 82.714 ;
               RECT 23.494 83.878 23.546 83.914 ;
               RECT 23.494 85.078 23.546 85.114 ;
               RECT 23.494 86.278 23.546 86.314 ;
               RECT 23.494 87.478 23.546 87.514 ;
               RECT 23.494 88.678 23.546 88.714 ;
               RECT 23.494 89.878 23.546 89.914 ;
               RECT 23.494 91.078 23.546 91.114 ;
               RECT 23.494 92.278 23.546 92.314 ;
               RECT 23.494 93.478 23.546 93.514 ;
               RECT 23.494 94.678 23.546 94.714 ;
               RECT 23.494 95.878 23.546 95.914 ;
               RECT 23.494 97.078 23.546 97.114 ;
               RECT 23.494 98.278 23.546 98.314 ;
               RECT 23.494 99.478 23.546 99.514 ;
               RECT 23.494 100.678 23.546 100.714 ;
               RECT 23.494 101.878 23.546 101.914 ;
               RECT 23.494 103.078 23.546 103.114 ;
               RECT 23.494 104.278 23.546 104.314 ;
               RECT 23.574 0.281 23.626 0.317 ;
               RECT 23.574 104.803 23.626 104.839 ;
               RECT 23.654 0.806 23.706 0.842 ;
               RECT 23.654 2.006 23.706 2.042 ;
               RECT 23.654 3.206 23.706 3.242 ;
               RECT 23.654 4.406 23.706 4.442 ;
               RECT 23.654 5.606 23.706 5.642 ;
               RECT 23.654 6.806 23.706 6.842 ;
               RECT 23.654 8.006 23.706 8.042 ;
               RECT 23.654 9.206 23.706 9.242 ;
               RECT 23.654 10.406 23.706 10.442 ;
               RECT 23.654 11.606 23.706 11.642 ;
               RECT 23.654 12.806 23.706 12.842 ;
               RECT 23.654 14.006 23.706 14.042 ;
               RECT 23.654 15.206 23.706 15.242 ;
               RECT 23.654 16.406 23.706 16.442 ;
               RECT 23.654 17.606 23.706 17.642 ;
               RECT 23.654 18.806 23.706 18.842 ;
               RECT 23.654 20.006 23.706 20.042 ;
               RECT 23.654 21.206 23.706 21.242 ;
               RECT 23.654 22.406 23.706 22.442 ;
               RECT 23.654 23.606 23.706 23.642 ;
               RECT 23.654 24.806 23.706 24.842 ;
               RECT 23.654 26.006 23.706 26.042 ;
               RECT 23.654 27.206 23.706 27.242 ;
               RECT 23.654 28.406 23.706 28.442 ;
               RECT 23.654 29.606 23.706 29.642 ;
               RECT 23.654 30.806 23.706 30.842 ;
               RECT 23.654 32.006 23.706 32.042 ;
               RECT 23.654 33.206 23.706 33.242 ;
               RECT 23.654 34.406 23.706 34.442 ;
               RECT 23.654 35.606 23.706 35.642 ;
               RECT 23.654 36.806 23.706 36.842 ;
               RECT 23.654 38.006 23.706 38.042 ;
               RECT 23.654 39.206 23.706 39.242 ;
               RECT 23.654 40.406 23.706 40.442 ;
               RECT 23.654 41.606 23.706 41.642 ;
               RECT 23.654 42.806 23.706 42.842 ;
               RECT 23.654 44.006 23.706 44.042 ;
               RECT 23.654 45.206 23.706 45.242 ;
               RECT 23.654 46.406 23.706 46.442 ;
               RECT 23.654 47.606 23.706 47.642 ;
               RECT 23.654 49.422 23.706 49.458 ;
               RECT 23.654 49.662 23.706 49.698 ;
               RECT 23.654 55.422 23.706 55.458 ;
               RECT 23.654 55.662 23.706 55.698 ;
               RECT 23.654 56.726 23.706 56.762 ;
               RECT 23.654 57.926 23.706 57.962 ;
               RECT 23.654 59.126 23.706 59.162 ;
               RECT 23.654 60.326 23.706 60.362 ;
               RECT 23.654 61.526 23.706 61.562 ;
               RECT 23.654 62.726 23.706 62.762 ;
               RECT 23.654 63.926 23.706 63.962 ;
               RECT 23.654 65.126 23.706 65.162 ;
               RECT 23.654 66.326 23.706 66.362 ;
               RECT 23.654 67.526 23.706 67.562 ;
               RECT 23.654 68.726 23.706 68.762 ;
               RECT 23.654 69.926 23.706 69.962 ;
               RECT 23.654 71.126 23.706 71.162 ;
               RECT 23.654 72.326 23.706 72.362 ;
               RECT 23.654 73.526 23.706 73.562 ;
               RECT 23.654 74.726 23.706 74.762 ;
               RECT 23.654 75.926 23.706 75.962 ;
               RECT 23.654 77.126 23.706 77.162 ;
               RECT 23.654 78.326 23.706 78.362 ;
               RECT 23.654 79.526 23.706 79.562 ;
               RECT 23.654 80.726 23.706 80.762 ;
               RECT 23.654 81.926 23.706 81.962 ;
               RECT 23.654 83.126 23.706 83.162 ;
               RECT 23.654 84.326 23.706 84.362 ;
               RECT 23.654 85.526 23.706 85.562 ;
               RECT 23.654 86.726 23.706 86.762 ;
               RECT 23.654 87.926 23.706 87.962 ;
               RECT 23.654 89.126 23.706 89.162 ;
               RECT 23.654 90.326 23.706 90.362 ;
               RECT 23.654 91.526 23.706 91.562 ;
               RECT 23.654 92.726 23.706 92.762 ;
               RECT 23.654 93.926 23.706 93.962 ;
               RECT 23.654 95.126 23.706 95.162 ;
               RECT 23.654 96.326 23.706 96.362 ;
               RECT 23.654 97.526 23.706 97.562 ;
               RECT 23.654 98.726 23.706 98.762 ;
               RECT 23.654 99.926 23.706 99.962 ;
               RECT 23.654 101.126 23.706 101.162 ;
               RECT 23.654 102.326 23.706 102.362 ;
               RECT 23.654 103.526 23.706 103.562 ;
               RECT 23.734 1.558 23.786 1.594 ;
               RECT 23.734 2.758 23.786 2.794 ;
               RECT 23.734 3.958 23.786 3.994 ;
               RECT 23.734 5.158 23.786 5.194 ;
               RECT 23.734 6.358 23.786 6.394 ;
               RECT 23.734 7.558 23.786 7.594 ;
               RECT 23.734 8.758 23.786 8.794 ;
               RECT 23.734 9.958 23.786 9.994 ;
               RECT 23.734 11.158 23.786 11.194 ;
               RECT 23.734 12.358 23.786 12.394 ;
               RECT 23.734 13.558 23.786 13.594 ;
               RECT 23.734 14.758 23.786 14.794 ;
               RECT 23.734 15.958 23.786 15.994 ;
               RECT 23.734 17.158 23.786 17.194 ;
               RECT 23.734 18.358 23.786 18.394 ;
               RECT 23.734 19.558 23.786 19.594 ;
               RECT 23.734 20.758 23.786 20.794 ;
               RECT 23.734 21.958 23.786 21.994 ;
               RECT 23.734 23.158 23.786 23.194 ;
               RECT 23.734 24.358 23.786 24.394 ;
               RECT 23.734 25.558 23.786 25.594 ;
               RECT 23.734 26.758 23.786 26.794 ;
               RECT 23.734 27.958 23.786 27.994 ;
               RECT 23.734 29.158 23.786 29.194 ;
               RECT 23.734 30.358 23.786 30.394 ;
               RECT 23.734 31.558 23.786 31.594 ;
               RECT 23.734 32.758 23.786 32.794 ;
               RECT 23.734 33.958 23.786 33.994 ;
               RECT 23.734 35.158 23.786 35.194 ;
               RECT 23.734 36.358 23.786 36.394 ;
               RECT 23.734 37.558 23.786 37.594 ;
               RECT 23.734 38.758 23.786 38.794 ;
               RECT 23.734 39.958 23.786 39.994 ;
               RECT 23.734 41.158 23.786 41.194 ;
               RECT 23.734 42.358 23.786 42.394 ;
               RECT 23.734 43.558 23.786 43.594 ;
               RECT 23.734 44.758 23.786 44.794 ;
               RECT 23.734 45.958 23.786 45.994 ;
               RECT 23.734 47.158 23.786 47.194 ;
               RECT 23.734 48.358 23.786 48.394 ;
               RECT 23.734 50.142 23.786 50.178 ;
               RECT 23.734 50.382 23.786 50.418 ;
               RECT 23.734 54.702 23.786 54.738 ;
               RECT 23.734 54.942 23.786 54.978 ;
               RECT 23.734 57.478 23.786 57.514 ;
               RECT 23.734 58.678 23.786 58.714 ;
               RECT 23.734 59.878 23.786 59.914 ;
               RECT 23.734 61.078 23.786 61.114 ;
               RECT 23.734 62.278 23.786 62.314 ;
               RECT 23.734 63.478 23.786 63.514 ;
               RECT 23.734 64.678 23.786 64.714 ;
               RECT 23.734 65.878 23.786 65.914 ;
               RECT 23.734 67.078 23.786 67.114 ;
               RECT 23.734 68.278 23.786 68.314 ;
               RECT 23.734 69.478 23.786 69.514 ;
               RECT 23.734 70.678 23.786 70.714 ;
               RECT 23.734 71.878 23.786 71.914 ;
               RECT 23.734 73.078 23.786 73.114 ;
               RECT 23.734 74.278 23.786 74.314 ;
               RECT 23.734 75.478 23.786 75.514 ;
               RECT 23.734 76.678 23.786 76.714 ;
               RECT 23.734 77.878 23.786 77.914 ;
               RECT 23.734 79.078 23.786 79.114 ;
               RECT 23.734 80.278 23.786 80.314 ;
               RECT 23.734 81.478 23.786 81.514 ;
               RECT 23.734 82.678 23.786 82.714 ;
               RECT 23.734 83.878 23.786 83.914 ;
               RECT 23.734 85.078 23.786 85.114 ;
               RECT 23.734 86.278 23.786 86.314 ;
               RECT 23.734 87.478 23.786 87.514 ;
               RECT 23.734 88.678 23.786 88.714 ;
               RECT 23.734 89.878 23.786 89.914 ;
               RECT 23.734 91.078 23.786 91.114 ;
               RECT 23.734 92.278 23.786 92.314 ;
               RECT 23.734 93.478 23.786 93.514 ;
               RECT 23.734 94.678 23.786 94.714 ;
               RECT 23.734 95.878 23.786 95.914 ;
               RECT 23.734 97.078 23.786 97.114 ;
               RECT 23.734 98.278 23.786 98.314 ;
               RECT 23.734 99.478 23.786 99.514 ;
               RECT 23.734 100.678 23.786 100.714 ;
               RECT 23.734 101.878 23.786 101.914 ;
               RECT 23.734 103.078 23.786 103.114 ;
               RECT 23.734 104.278 23.786 104.314 ;
               RECT 23.814 0.806 23.866 0.842 ;
               RECT 23.814 2.006 23.866 2.042 ;
               RECT 23.814 3.206 23.866 3.242 ;
               RECT 23.814 4.406 23.866 4.442 ;
               RECT 23.814 5.606 23.866 5.642 ;
               RECT 23.814 6.806 23.866 6.842 ;
               RECT 23.814 8.006 23.866 8.042 ;
               RECT 23.814 9.206 23.866 9.242 ;
               RECT 23.814 10.406 23.866 10.442 ;
               RECT 23.814 11.606 23.866 11.642 ;
               RECT 23.814 12.806 23.866 12.842 ;
               RECT 23.814 14.006 23.866 14.042 ;
               RECT 23.814 15.206 23.866 15.242 ;
               RECT 23.814 16.406 23.866 16.442 ;
               RECT 23.814 17.606 23.866 17.642 ;
               RECT 23.814 18.806 23.866 18.842 ;
               RECT 23.814 20.006 23.866 20.042 ;
               RECT 23.814 21.206 23.866 21.242 ;
               RECT 23.814 22.406 23.866 22.442 ;
               RECT 23.814 23.606 23.866 23.642 ;
               RECT 23.814 24.806 23.866 24.842 ;
               RECT 23.814 26.006 23.866 26.042 ;
               RECT 23.814 27.206 23.866 27.242 ;
               RECT 23.814 28.406 23.866 28.442 ;
               RECT 23.814 29.606 23.866 29.642 ;
               RECT 23.814 30.806 23.866 30.842 ;
               RECT 23.814 32.006 23.866 32.042 ;
               RECT 23.814 33.206 23.866 33.242 ;
               RECT 23.814 34.406 23.866 34.442 ;
               RECT 23.814 35.606 23.866 35.642 ;
               RECT 23.814 36.806 23.866 36.842 ;
               RECT 23.814 38.006 23.866 38.042 ;
               RECT 23.814 39.206 23.866 39.242 ;
               RECT 23.814 40.406 23.866 40.442 ;
               RECT 23.814 41.606 23.866 41.642 ;
               RECT 23.814 42.806 23.866 42.842 ;
               RECT 23.814 44.006 23.866 44.042 ;
               RECT 23.814 45.206 23.866 45.242 ;
               RECT 23.814 46.406 23.866 46.442 ;
               RECT 23.814 47.606 23.866 47.642 ;
               RECT 23.814 49.422 23.866 49.458 ;
               RECT 23.814 49.662 23.866 49.698 ;
               RECT 23.814 55.422 23.866 55.458 ;
               RECT 23.814 55.662 23.866 55.698 ;
               RECT 23.814 56.726 23.866 56.762 ;
               RECT 23.814 57.926 23.866 57.962 ;
               RECT 23.814 59.126 23.866 59.162 ;
               RECT 23.814 60.326 23.866 60.362 ;
               RECT 23.814 61.526 23.866 61.562 ;
               RECT 23.814 62.726 23.866 62.762 ;
               RECT 23.814 63.926 23.866 63.962 ;
               RECT 23.814 65.126 23.866 65.162 ;
               RECT 23.814 66.326 23.866 66.362 ;
               RECT 23.814 67.526 23.866 67.562 ;
               RECT 23.814 68.726 23.866 68.762 ;
               RECT 23.814 69.926 23.866 69.962 ;
               RECT 23.814 71.126 23.866 71.162 ;
               RECT 23.814 72.326 23.866 72.362 ;
               RECT 23.814 73.526 23.866 73.562 ;
               RECT 23.814 74.726 23.866 74.762 ;
               RECT 23.814 75.926 23.866 75.962 ;
               RECT 23.814 77.126 23.866 77.162 ;
               RECT 23.814 78.326 23.866 78.362 ;
               RECT 23.814 79.526 23.866 79.562 ;
               RECT 23.814 80.726 23.866 80.762 ;
               RECT 23.814 81.926 23.866 81.962 ;
               RECT 23.814 83.126 23.866 83.162 ;
               RECT 23.814 84.326 23.866 84.362 ;
               RECT 23.814 85.526 23.866 85.562 ;
               RECT 23.814 86.726 23.866 86.762 ;
               RECT 23.814 87.926 23.866 87.962 ;
               RECT 23.814 89.126 23.866 89.162 ;
               RECT 23.814 90.326 23.866 90.362 ;
               RECT 23.814 91.526 23.866 91.562 ;
               RECT 23.814 92.726 23.866 92.762 ;
               RECT 23.814 93.926 23.866 93.962 ;
               RECT 23.814 95.126 23.866 95.162 ;
               RECT 23.814 96.326 23.866 96.362 ;
               RECT 23.814 97.526 23.866 97.562 ;
               RECT 23.814 98.726 23.866 98.762 ;
               RECT 23.814 99.926 23.866 99.962 ;
               RECT 23.814 101.126 23.866 101.162 ;
               RECT 23.814 102.326 23.866 102.362 ;
               RECT 23.814 103.526 23.866 103.562 ;
               RECT 23.894 1.558 23.946 1.594 ;
               RECT 23.894 2.758 23.946 2.794 ;
               RECT 23.894 3.958 23.946 3.994 ;
               RECT 23.894 5.158 23.946 5.194 ;
               RECT 23.894 6.358 23.946 6.394 ;
               RECT 23.894 7.558 23.946 7.594 ;
               RECT 23.894 8.758 23.946 8.794 ;
               RECT 23.894 9.958 23.946 9.994 ;
               RECT 23.894 11.158 23.946 11.194 ;
               RECT 23.894 12.358 23.946 12.394 ;
               RECT 23.894 13.558 23.946 13.594 ;
               RECT 23.894 14.758 23.946 14.794 ;
               RECT 23.894 15.958 23.946 15.994 ;
               RECT 23.894 17.158 23.946 17.194 ;
               RECT 23.894 18.358 23.946 18.394 ;
               RECT 23.894 19.558 23.946 19.594 ;
               RECT 23.894 20.758 23.946 20.794 ;
               RECT 23.894 21.958 23.946 21.994 ;
               RECT 23.894 23.158 23.946 23.194 ;
               RECT 23.894 24.358 23.946 24.394 ;
               RECT 23.894 25.558 23.946 25.594 ;
               RECT 23.894 26.758 23.946 26.794 ;
               RECT 23.894 27.958 23.946 27.994 ;
               RECT 23.894 29.158 23.946 29.194 ;
               RECT 23.894 30.358 23.946 30.394 ;
               RECT 23.894 31.558 23.946 31.594 ;
               RECT 23.894 32.758 23.946 32.794 ;
               RECT 23.894 33.958 23.946 33.994 ;
               RECT 23.894 35.158 23.946 35.194 ;
               RECT 23.894 36.358 23.946 36.394 ;
               RECT 23.894 37.558 23.946 37.594 ;
               RECT 23.894 38.758 23.946 38.794 ;
               RECT 23.894 39.958 23.946 39.994 ;
               RECT 23.894 41.158 23.946 41.194 ;
               RECT 23.894 42.358 23.946 42.394 ;
               RECT 23.894 43.558 23.946 43.594 ;
               RECT 23.894 44.758 23.946 44.794 ;
               RECT 23.894 45.958 23.946 45.994 ;
               RECT 23.894 47.158 23.946 47.194 ;
               RECT 23.894 48.358 23.946 48.394 ;
               RECT 23.894 50.142 23.946 50.178 ;
               RECT 23.894 50.382 23.946 50.418 ;
               RECT 23.894 54.702 23.946 54.738 ;
               RECT 23.894 54.942 23.946 54.978 ;
               RECT 23.894 57.478 23.946 57.514 ;
               RECT 23.894 58.678 23.946 58.714 ;
               RECT 23.894 59.878 23.946 59.914 ;
               RECT 23.894 61.078 23.946 61.114 ;
               RECT 23.894 62.278 23.946 62.314 ;
               RECT 23.894 63.478 23.946 63.514 ;
               RECT 23.894 64.678 23.946 64.714 ;
               RECT 23.894 65.878 23.946 65.914 ;
               RECT 23.894 67.078 23.946 67.114 ;
               RECT 23.894 68.278 23.946 68.314 ;
               RECT 23.894 69.478 23.946 69.514 ;
               RECT 23.894 70.678 23.946 70.714 ;
               RECT 23.894 71.878 23.946 71.914 ;
               RECT 23.894 73.078 23.946 73.114 ;
               RECT 23.894 74.278 23.946 74.314 ;
               RECT 23.894 75.478 23.946 75.514 ;
               RECT 23.894 76.678 23.946 76.714 ;
               RECT 23.894 77.878 23.946 77.914 ;
               RECT 23.894 79.078 23.946 79.114 ;
               RECT 23.894 80.278 23.946 80.314 ;
               RECT 23.894 81.478 23.946 81.514 ;
               RECT 23.894 82.678 23.946 82.714 ;
               RECT 23.894 83.878 23.946 83.914 ;
               RECT 23.894 85.078 23.946 85.114 ;
               RECT 23.894 86.278 23.946 86.314 ;
               RECT 23.894 87.478 23.946 87.514 ;
               RECT 23.894 88.678 23.946 88.714 ;
               RECT 23.894 89.878 23.946 89.914 ;
               RECT 23.894 91.078 23.946 91.114 ;
               RECT 23.894 92.278 23.946 92.314 ;
               RECT 23.894 93.478 23.946 93.514 ;
               RECT 23.894 94.678 23.946 94.714 ;
               RECT 23.894 95.878 23.946 95.914 ;
               RECT 23.894 97.078 23.946 97.114 ;
               RECT 23.894 98.278 23.946 98.314 ;
               RECT 23.894 99.478 23.946 99.514 ;
               RECT 23.894 100.678 23.946 100.714 ;
               RECT 23.894 101.878 23.946 101.914 ;
               RECT 23.894 103.078 23.946 103.114 ;
               RECT 23.894 104.278 23.946 104.314 ;
               RECT 23.974 0.281 24.026 0.317 ;
               RECT 23.974 104.803 24.026 104.839 ;
               RECT 24.054 0.806 24.106 0.842 ;
               RECT 24.054 2.006 24.106 2.042 ;
               RECT 24.054 3.206 24.106 3.242 ;
               RECT 24.054 4.406 24.106 4.442 ;
               RECT 24.054 5.606 24.106 5.642 ;
               RECT 24.054 6.806 24.106 6.842 ;
               RECT 24.054 8.006 24.106 8.042 ;
               RECT 24.054 9.206 24.106 9.242 ;
               RECT 24.054 10.406 24.106 10.442 ;
               RECT 24.054 11.606 24.106 11.642 ;
               RECT 24.054 12.806 24.106 12.842 ;
               RECT 24.054 14.006 24.106 14.042 ;
               RECT 24.054 15.206 24.106 15.242 ;
               RECT 24.054 16.406 24.106 16.442 ;
               RECT 24.054 17.606 24.106 17.642 ;
               RECT 24.054 18.806 24.106 18.842 ;
               RECT 24.054 20.006 24.106 20.042 ;
               RECT 24.054 21.206 24.106 21.242 ;
               RECT 24.054 22.406 24.106 22.442 ;
               RECT 24.054 23.606 24.106 23.642 ;
               RECT 24.054 24.806 24.106 24.842 ;
               RECT 24.054 26.006 24.106 26.042 ;
               RECT 24.054 27.206 24.106 27.242 ;
               RECT 24.054 28.406 24.106 28.442 ;
               RECT 24.054 29.606 24.106 29.642 ;
               RECT 24.054 30.806 24.106 30.842 ;
               RECT 24.054 32.006 24.106 32.042 ;
               RECT 24.054 33.206 24.106 33.242 ;
               RECT 24.054 34.406 24.106 34.442 ;
               RECT 24.054 35.606 24.106 35.642 ;
               RECT 24.054 36.806 24.106 36.842 ;
               RECT 24.054 38.006 24.106 38.042 ;
               RECT 24.054 39.206 24.106 39.242 ;
               RECT 24.054 40.406 24.106 40.442 ;
               RECT 24.054 41.606 24.106 41.642 ;
               RECT 24.054 42.806 24.106 42.842 ;
               RECT 24.054 44.006 24.106 44.042 ;
               RECT 24.054 45.206 24.106 45.242 ;
               RECT 24.054 46.406 24.106 46.442 ;
               RECT 24.054 47.606 24.106 47.642 ;
               RECT 24.054 49.422 24.106 49.458 ;
               RECT 24.054 49.662 24.106 49.698 ;
               RECT 24.054 51.102 24.106 51.138 ;
               RECT 24.054 51.582 24.106 51.618 ;
               RECT 24.054 53.502 24.106 53.538 ;
               RECT 24.054 53.982 24.106 54.018 ;
               RECT 24.054 55.422 24.106 55.458 ;
               RECT 24.054 55.662 24.106 55.698 ;
               RECT 24.054 56.726 24.106 56.762 ;
               RECT 24.054 57.926 24.106 57.962 ;
               RECT 24.054 59.126 24.106 59.162 ;
               RECT 24.054 60.326 24.106 60.362 ;
               RECT 24.054 61.526 24.106 61.562 ;
               RECT 24.054 62.726 24.106 62.762 ;
               RECT 24.054 63.926 24.106 63.962 ;
               RECT 24.054 65.126 24.106 65.162 ;
               RECT 24.054 66.326 24.106 66.362 ;
               RECT 24.054 67.526 24.106 67.562 ;
               RECT 24.054 68.726 24.106 68.762 ;
               RECT 24.054 69.926 24.106 69.962 ;
               RECT 24.054 71.126 24.106 71.162 ;
               RECT 24.054 72.326 24.106 72.362 ;
               RECT 24.054 73.526 24.106 73.562 ;
               RECT 24.054 74.726 24.106 74.762 ;
               RECT 24.054 75.926 24.106 75.962 ;
               RECT 24.054 77.126 24.106 77.162 ;
               RECT 24.054 78.326 24.106 78.362 ;
               RECT 24.054 79.526 24.106 79.562 ;
               RECT 24.054 80.726 24.106 80.762 ;
               RECT 24.054 81.926 24.106 81.962 ;
               RECT 24.054 83.126 24.106 83.162 ;
               RECT 24.054 84.326 24.106 84.362 ;
               RECT 24.054 85.526 24.106 85.562 ;
               RECT 24.054 86.726 24.106 86.762 ;
               RECT 24.054 87.926 24.106 87.962 ;
               RECT 24.054 89.126 24.106 89.162 ;
               RECT 24.054 90.326 24.106 90.362 ;
               RECT 24.054 91.526 24.106 91.562 ;
               RECT 24.054 92.726 24.106 92.762 ;
               RECT 24.054 93.926 24.106 93.962 ;
               RECT 24.054 95.126 24.106 95.162 ;
               RECT 24.054 96.326 24.106 96.362 ;
               RECT 24.054 97.526 24.106 97.562 ;
               RECT 24.054 98.726 24.106 98.762 ;
               RECT 24.054 99.926 24.106 99.962 ;
               RECT 24.054 101.126 24.106 101.162 ;
               RECT 24.054 102.326 24.106 102.362 ;
               RECT 24.054 103.526 24.106 103.562 ;
               RECT 24.134 1.558 24.186 1.594 ;
               RECT 24.134 2.758 24.186 2.794 ;
               RECT 24.134 3.958 24.186 3.994 ;
               RECT 24.134 5.158 24.186 5.194 ;
               RECT 24.134 6.358 24.186 6.394 ;
               RECT 24.134 7.558 24.186 7.594 ;
               RECT 24.134 8.758 24.186 8.794 ;
               RECT 24.134 9.958 24.186 9.994 ;
               RECT 24.134 11.158 24.186 11.194 ;
               RECT 24.134 12.358 24.186 12.394 ;
               RECT 24.134 13.558 24.186 13.594 ;
               RECT 24.134 14.758 24.186 14.794 ;
               RECT 24.134 15.958 24.186 15.994 ;
               RECT 24.134 17.158 24.186 17.194 ;
               RECT 24.134 18.358 24.186 18.394 ;
               RECT 24.134 19.558 24.186 19.594 ;
               RECT 24.134 20.758 24.186 20.794 ;
               RECT 24.134 21.958 24.186 21.994 ;
               RECT 24.134 23.158 24.186 23.194 ;
               RECT 24.134 24.358 24.186 24.394 ;
               RECT 24.134 25.558 24.186 25.594 ;
               RECT 24.134 26.758 24.186 26.794 ;
               RECT 24.134 27.958 24.186 27.994 ;
               RECT 24.134 29.158 24.186 29.194 ;
               RECT 24.134 30.358 24.186 30.394 ;
               RECT 24.134 31.558 24.186 31.594 ;
               RECT 24.134 32.758 24.186 32.794 ;
               RECT 24.134 33.958 24.186 33.994 ;
               RECT 24.134 35.158 24.186 35.194 ;
               RECT 24.134 36.358 24.186 36.394 ;
               RECT 24.134 37.558 24.186 37.594 ;
               RECT 24.134 38.758 24.186 38.794 ;
               RECT 24.134 39.958 24.186 39.994 ;
               RECT 24.134 41.158 24.186 41.194 ;
               RECT 24.134 42.358 24.186 42.394 ;
               RECT 24.134 43.558 24.186 43.594 ;
               RECT 24.134 44.758 24.186 44.794 ;
               RECT 24.134 45.958 24.186 45.994 ;
               RECT 24.134 47.158 24.186 47.194 ;
               RECT 24.134 48.358 24.186 48.394 ;
               RECT 24.134 50.142 24.186 50.178 ;
               RECT 24.134 50.382 24.186 50.418 ;
               RECT 24.134 54.702 24.186 54.738 ;
               RECT 24.134 54.942 24.186 54.978 ;
               RECT 24.134 57.478 24.186 57.514 ;
               RECT 24.134 58.678 24.186 58.714 ;
               RECT 24.134 59.878 24.186 59.914 ;
               RECT 24.134 61.078 24.186 61.114 ;
               RECT 24.134 62.278 24.186 62.314 ;
               RECT 24.134 63.478 24.186 63.514 ;
               RECT 24.134 64.678 24.186 64.714 ;
               RECT 24.134 65.878 24.186 65.914 ;
               RECT 24.134 67.078 24.186 67.114 ;
               RECT 24.134 68.278 24.186 68.314 ;
               RECT 24.134 69.478 24.186 69.514 ;
               RECT 24.134 70.678 24.186 70.714 ;
               RECT 24.134 71.878 24.186 71.914 ;
               RECT 24.134 73.078 24.186 73.114 ;
               RECT 24.134 74.278 24.186 74.314 ;
               RECT 24.134 75.478 24.186 75.514 ;
               RECT 24.134 76.678 24.186 76.714 ;
               RECT 24.134 77.878 24.186 77.914 ;
               RECT 24.134 79.078 24.186 79.114 ;
               RECT 24.134 80.278 24.186 80.314 ;
               RECT 24.134 81.478 24.186 81.514 ;
               RECT 24.134 82.678 24.186 82.714 ;
               RECT 24.134 83.878 24.186 83.914 ;
               RECT 24.134 85.078 24.186 85.114 ;
               RECT 24.134 86.278 24.186 86.314 ;
               RECT 24.134 87.478 24.186 87.514 ;
               RECT 24.134 88.678 24.186 88.714 ;
               RECT 24.134 89.878 24.186 89.914 ;
               RECT 24.134 91.078 24.186 91.114 ;
               RECT 24.134 92.278 24.186 92.314 ;
               RECT 24.134 93.478 24.186 93.514 ;
               RECT 24.134 94.678 24.186 94.714 ;
               RECT 24.134 95.878 24.186 95.914 ;
               RECT 24.134 97.078 24.186 97.114 ;
               RECT 24.134 98.278 24.186 98.314 ;
               RECT 24.134 99.478 24.186 99.514 ;
               RECT 24.134 100.678 24.186 100.714 ;
               RECT 24.134 101.878 24.186 101.914 ;
               RECT 24.134 103.078 24.186 103.114 ;
               RECT 24.134 104.278 24.186 104.314 ;
               RECT 24.214 0.806 24.266 0.842 ;
               RECT 24.214 2.006 24.266 2.042 ;
               RECT 24.214 3.206 24.266 3.242 ;
               RECT 24.214 4.406 24.266 4.442 ;
               RECT 24.214 5.606 24.266 5.642 ;
               RECT 24.214 6.806 24.266 6.842 ;
               RECT 24.214 8.006 24.266 8.042 ;
               RECT 24.214 9.206 24.266 9.242 ;
               RECT 24.214 10.406 24.266 10.442 ;
               RECT 24.214 11.606 24.266 11.642 ;
               RECT 24.214 12.806 24.266 12.842 ;
               RECT 24.214 14.006 24.266 14.042 ;
               RECT 24.214 15.206 24.266 15.242 ;
               RECT 24.214 16.406 24.266 16.442 ;
               RECT 24.214 17.606 24.266 17.642 ;
               RECT 24.214 18.806 24.266 18.842 ;
               RECT 24.214 20.006 24.266 20.042 ;
               RECT 24.214 21.206 24.266 21.242 ;
               RECT 24.214 22.406 24.266 22.442 ;
               RECT 24.214 23.606 24.266 23.642 ;
               RECT 24.214 24.806 24.266 24.842 ;
               RECT 24.214 26.006 24.266 26.042 ;
               RECT 24.214 27.206 24.266 27.242 ;
               RECT 24.214 28.406 24.266 28.442 ;
               RECT 24.214 29.606 24.266 29.642 ;
               RECT 24.214 30.806 24.266 30.842 ;
               RECT 24.214 32.006 24.266 32.042 ;
               RECT 24.214 33.206 24.266 33.242 ;
               RECT 24.214 34.406 24.266 34.442 ;
               RECT 24.214 35.606 24.266 35.642 ;
               RECT 24.214 36.806 24.266 36.842 ;
               RECT 24.214 38.006 24.266 38.042 ;
               RECT 24.214 39.206 24.266 39.242 ;
               RECT 24.214 40.406 24.266 40.442 ;
               RECT 24.214 41.606 24.266 41.642 ;
               RECT 24.214 42.806 24.266 42.842 ;
               RECT 24.214 44.006 24.266 44.042 ;
               RECT 24.214 45.206 24.266 45.242 ;
               RECT 24.214 46.406 24.266 46.442 ;
               RECT 24.214 47.606 24.266 47.642 ;
               RECT 24.214 49.422 24.266 49.458 ;
               RECT 24.214 49.662 24.266 49.698 ;
               RECT 24.214 55.422 24.266 55.458 ;
               RECT 24.214 55.662 24.266 55.698 ;
               RECT 24.214 56.726 24.266 56.762 ;
               RECT 24.214 57.926 24.266 57.962 ;
               RECT 24.214 59.126 24.266 59.162 ;
               RECT 24.214 60.326 24.266 60.362 ;
               RECT 24.214 61.526 24.266 61.562 ;
               RECT 24.214 62.726 24.266 62.762 ;
               RECT 24.214 63.926 24.266 63.962 ;
               RECT 24.214 65.126 24.266 65.162 ;
               RECT 24.214 66.326 24.266 66.362 ;
               RECT 24.214 67.526 24.266 67.562 ;
               RECT 24.214 68.726 24.266 68.762 ;
               RECT 24.214 69.926 24.266 69.962 ;
               RECT 24.214 71.126 24.266 71.162 ;
               RECT 24.214 72.326 24.266 72.362 ;
               RECT 24.214 73.526 24.266 73.562 ;
               RECT 24.214 74.726 24.266 74.762 ;
               RECT 24.214 75.926 24.266 75.962 ;
               RECT 24.214 77.126 24.266 77.162 ;
               RECT 24.214 78.326 24.266 78.362 ;
               RECT 24.214 79.526 24.266 79.562 ;
               RECT 24.214 80.726 24.266 80.762 ;
               RECT 24.214 81.926 24.266 81.962 ;
               RECT 24.214 83.126 24.266 83.162 ;
               RECT 24.214 84.326 24.266 84.362 ;
               RECT 24.214 85.526 24.266 85.562 ;
               RECT 24.214 86.726 24.266 86.762 ;
               RECT 24.214 87.926 24.266 87.962 ;
               RECT 24.214 89.126 24.266 89.162 ;
               RECT 24.214 90.326 24.266 90.362 ;
               RECT 24.214 91.526 24.266 91.562 ;
               RECT 24.214 92.726 24.266 92.762 ;
               RECT 24.214 93.926 24.266 93.962 ;
               RECT 24.214 95.126 24.266 95.162 ;
               RECT 24.214 96.326 24.266 96.362 ;
               RECT 24.214 97.526 24.266 97.562 ;
               RECT 24.214 98.726 24.266 98.762 ;
               RECT 24.214 99.926 24.266 99.962 ;
               RECT 24.214 101.126 24.266 101.162 ;
               RECT 24.214 102.326 24.266 102.362 ;
               RECT 24.214 103.526 24.266 103.562 ;
               RECT 24.294 1.558 24.346 1.594 ;
               RECT 24.294 2.758 24.346 2.794 ;
               RECT 24.294 3.958 24.346 3.994 ;
               RECT 24.294 5.158 24.346 5.194 ;
               RECT 24.294 6.358 24.346 6.394 ;
               RECT 24.294 7.558 24.346 7.594 ;
               RECT 24.294 8.758 24.346 8.794 ;
               RECT 24.294 9.958 24.346 9.994 ;
               RECT 24.294 11.158 24.346 11.194 ;
               RECT 24.294 12.358 24.346 12.394 ;
               RECT 24.294 13.558 24.346 13.594 ;
               RECT 24.294 14.758 24.346 14.794 ;
               RECT 24.294 15.958 24.346 15.994 ;
               RECT 24.294 17.158 24.346 17.194 ;
               RECT 24.294 18.358 24.346 18.394 ;
               RECT 24.294 19.558 24.346 19.594 ;
               RECT 24.294 20.758 24.346 20.794 ;
               RECT 24.294 21.958 24.346 21.994 ;
               RECT 24.294 23.158 24.346 23.194 ;
               RECT 24.294 24.358 24.346 24.394 ;
               RECT 24.294 25.558 24.346 25.594 ;
               RECT 24.294 26.758 24.346 26.794 ;
               RECT 24.294 27.958 24.346 27.994 ;
               RECT 24.294 29.158 24.346 29.194 ;
               RECT 24.294 30.358 24.346 30.394 ;
               RECT 24.294 31.558 24.346 31.594 ;
               RECT 24.294 32.758 24.346 32.794 ;
               RECT 24.294 33.958 24.346 33.994 ;
               RECT 24.294 35.158 24.346 35.194 ;
               RECT 24.294 36.358 24.346 36.394 ;
               RECT 24.294 37.558 24.346 37.594 ;
               RECT 24.294 38.758 24.346 38.794 ;
               RECT 24.294 39.958 24.346 39.994 ;
               RECT 24.294 41.158 24.346 41.194 ;
               RECT 24.294 42.358 24.346 42.394 ;
               RECT 24.294 43.558 24.346 43.594 ;
               RECT 24.294 44.758 24.346 44.794 ;
               RECT 24.294 45.958 24.346 45.994 ;
               RECT 24.294 47.158 24.346 47.194 ;
               RECT 24.294 48.358 24.346 48.394 ;
               RECT 24.294 50.142 24.346 50.178 ;
               RECT 24.294 50.382 24.346 50.418 ;
               RECT 24.294 54.702 24.346 54.738 ;
               RECT 24.294 54.942 24.346 54.978 ;
               RECT 24.294 57.478 24.346 57.514 ;
               RECT 24.294 58.678 24.346 58.714 ;
               RECT 24.294 59.878 24.346 59.914 ;
               RECT 24.294 61.078 24.346 61.114 ;
               RECT 24.294 62.278 24.346 62.314 ;
               RECT 24.294 63.478 24.346 63.514 ;
               RECT 24.294 64.678 24.346 64.714 ;
               RECT 24.294 65.878 24.346 65.914 ;
               RECT 24.294 67.078 24.346 67.114 ;
               RECT 24.294 68.278 24.346 68.314 ;
               RECT 24.294 69.478 24.346 69.514 ;
               RECT 24.294 70.678 24.346 70.714 ;
               RECT 24.294 71.878 24.346 71.914 ;
               RECT 24.294 73.078 24.346 73.114 ;
               RECT 24.294 74.278 24.346 74.314 ;
               RECT 24.294 75.478 24.346 75.514 ;
               RECT 24.294 76.678 24.346 76.714 ;
               RECT 24.294 77.878 24.346 77.914 ;
               RECT 24.294 79.078 24.346 79.114 ;
               RECT 24.294 80.278 24.346 80.314 ;
               RECT 24.294 81.478 24.346 81.514 ;
               RECT 24.294 82.678 24.346 82.714 ;
               RECT 24.294 83.878 24.346 83.914 ;
               RECT 24.294 85.078 24.346 85.114 ;
               RECT 24.294 86.278 24.346 86.314 ;
               RECT 24.294 87.478 24.346 87.514 ;
               RECT 24.294 88.678 24.346 88.714 ;
               RECT 24.294 89.878 24.346 89.914 ;
               RECT 24.294 91.078 24.346 91.114 ;
               RECT 24.294 92.278 24.346 92.314 ;
               RECT 24.294 93.478 24.346 93.514 ;
               RECT 24.294 94.678 24.346 94.714 ;
               RECT 24.294 95.878 24.346 95.914 ;
               RECT 24.294 97.078 24.346 97.114 ;
               RECT 24.294 98.278 24.346 98.314 ;
               RECT 24.294 99.478 24.346 99.514 ;
               RECT 24.294 100.678 24.346 100.714 ;
               RECT 24.294 101.878 24.346 101.914 ;
               RECT 24.294 103.078 24.346 103.114 ;
               RECT 24.294 104.278 24.346 104.314 ;
               RECT 24.374 0.281 24.426 0.317 ;
               RECT 24.374 104.803 24.426 104.839 ;
               RECT 24.454 0.806 24.506 0.842 ;
               RECT 24.454 2.006 24.506 2.042 ;
               RECT 24.454 3.206 24.506 3.242 ;
               RECT 24.454 4.406 24.506 4.442 ;
               RECT 24.454 5.606 24.506 5.642 ;
               RECT 24.454 6.806 24.506 6.842 ;
               RECT 24.454 8.006 24.506 8.042 ;
               RECT 24.454 9.206 24.506 9.242 ;
               RECT 24.454 10.406 24.506 10.442 ;
               RECT 24.454 11.606 24.506 11.642 ;
               RECT 24.454 12.806 24.506 12.842 ;
               RECT 24.454 14.006 24.506 14.042 ;
               RECT 24.454 15.206 24.506 15.242 ;
               RECT 24.454 16.406 24.506 16.442 ;
               RECT 24.454 17.606 24.506 17.642 ;
               RECT 24.454 18.806 24.506 18.842 ;
               RECT 24.454 20.006 24.506 20.042 ;
               RECT 24.454 21.206 24.506 21.242 ;
               RECT 24.454 22.406 24.506 22.442 ;
               RECT 24.454 23.606 24.506 23.642 ;
               RECT 24.454 24.806 24.506 24.842 ;
               RECT 24.454 26.006 24.506 26.042 ;
               RECT 24.454 27.206 24.506 27.242 ;
               RECT 24.454 28.406 24.506 28.442 ;
               RECT 24.454 29.606 24.506 29.642 ;
               RECT 24.454 30.806 24.506 30.842 ;
               RECT 24.454 32.006 24.506 32.042 ;
               RECT 24.454 33.206 24.506 33.242 ;
               RECT 24.454 34.406 24.506 34.442 ;
               RECT 24.454 35.606 24.506 35.642 ;
               RECT 24.454 36.806 24.506 36.842 ;
               RECT 24.454 38.006 24.506 38.042 ;
               RECT 24.454 39.206 24.506 39.242 ;
               RECT 24.454 40.406 24.506 40.442 ;
               RECT 24.454 41.606 24.506 41.642 ;
               RECT 24.454 42.806 24.506 42.842 ;
               RECT 24.454 44.006 24.506 44.042 ;
               RECT 24.454 45.206 24.506 45.242 ;
               RECT 24.454 46.406 24.506 46.442 ;
               RECT 24.454 47.606 24.506 47.642 ;
               RECT 24.454 49.422 24.506 49.458 ;
               RECT 24.454 49.662 24.506 49.698 ;
               RECT 24.454 55.422 24.506 55.458 ;
               RECT 24.454 55.662 24.506 55.698 ;
               RECT 24.454 56.726 24.506 56.762 ;
               RECT 24.454 57.926 24.506 57.962 ;
               RECT 24.454 59.126 24.506 59.162 ;
               RECT 24.454 60.326 24.506 60.362 ;
               RECT 24.454 61.526 24.506 61.562 ;
               RECT 24.454 62.726 24.506 62.762 ;
               RECT 24.454 63.926 24.506 63.962 ;
               RECT 24.454 65.126 24.506 65.162 ;
               RECT 24.454 66.326 24.506 66.362 ;
               RECT 24.454 67.526 24.506 67.562 ;
               RECT 24.454 68.726 24.506 68.762 ;
               RECT 24.454 69.926 24.506 69.962 ;
               RECT 24.454 71.126 24.506 71.162 ;
               RECT 24.454 72.326 24.506 72.362 ;
               RECT 24.454 73.526 24.506 73.562 ;
               RECT 24.454 74.726 24.506 74.762 ;
               RECT 24.454 75.926 24.506 75.962 ;
               RECT 24.454 77.126 24.506 77.162 ;
               RECT 24.454 78.326 24.506 78.362 ;
               RECT 24.454 79.526 24.506 79.562 ;
               RECT 24.454 80.726 24.506 80.762 ;
               RECT 24.454 81.926 24.506 81.962 ;
               RECT 24.454 83.126 24.506 83.162 ;
               RECT 24.454 84.326 24.506 84.362 ;
               RECT 24.454 85.526 24.506 85.562 ;
               RECT 24.454 86.726 24.506 86.762 ;
               RECT 24.454 87.926 24.506 87.962 ;
               RECT 24.454 89.126 24.506 89.162 ;
               RECT 24.454 90.326 24.506 90.362 ;
               RECT 24.454 91.526 24.506 91.562 ;
               RECT 24.454 92.726 24.506 92.762 ;
               RECT 24.454 93.926 24.506 93.962 ;
               RECT 24.454 95.126 24.506 95.162 ;
               RECT 24.454 96.326 24.506 96.362 ;
               RECT 24.454 97.526 24.506 97.562 ;
               RECT 24.454 98.726 24.506 98.762 ;
               RECT 24.454 99.926 24.506 99.962 ;
               RECT 24.454 101.126 24.506 101.162 ;
               RECT 24.454 102.326 24.506 102.362 ;
               RECT 24.454 103.526 24.506 103.562 ;
               RECT 24.534 1.558 24.586 1.594 ;
               RECT 24.534 2.758 24.586 2.794 ;
               RECT 24.534 3.958 24.586 3.994 ;
               RECT 24.534 5.158 24.586 5.194 ;
               RECT 24.534 6.358 24.586 6.394 ;
               RECT 24.534 7.558 24.586 7.594 ;
               RECT 24.534 8.758 24.586 8.794 ;
               RECT 24.534 9.958 24.586 9.994 ;
               RECT 24.534 11.158 24.586 11.194 ;
               RECT 24.534 12.358 24.586 12.394 ;
               RECT 24.534 13.558 24.586 13.594 ;
               RECT 24.534 14.758 24.586 14.794 ;
               RECT 24.534 15.958 24.586 15.994 ;
               RECT 24.534 17.158 24.586 17.194 ;
               RECT 24.534 18.358 24.586 18.394 ;
               RECT 24.534 19.558 24.586 19.594 ;
               RECT 24.534 20.758 24.586 20.794 ;
               RECT 24.534 21.958 24.586 21.994 ;
               RECT 24.534 23.158 24.586 23.194 ;
               RECT 24.534 24.358 24.586 24.394 ;
               RECT 24.534 25.558 24.586 25.594 ;
               RECT 24.534 26.758 24.586 26.794 ;
               RECT 24.534 27.958 24.586 27.994 ;
               RECT 24.534 29.158 24.586 29.194 ;
               RECT 24.534 30.358 24.586 30.394 ;
               RECT 24.534 31.558 24.586 31.594 ;
               RECT 24.534 32.758 24.586 32.794 ;
               RECT 24.534 33.958 24.586 33.994 ;
               RECT 24.534 35.158 24.586 35.194 ;
               RECT 24.534 36.358 24.586 36.394 ;
               RECT 24.534 37.558 24.586 37.594 ;
               RECT 24.534 38.758 24.586 38.794 ;
               RECT 24.534 39.958 24.586 39.994 ;
               RECT 24.534 41.158 24.586 41.194 ;
               RECT 24.534 42.358 24.586 42.394 ;
               RECT 24.534 43.558 24.586 43.594 ;
               RECT 24.534 44.758 24.586 44.794 ;
               RECT 24.534 45.958 24.586 45.994 ;
               RECT 24.534 47.158 24.586 47.194 ;
               RECT 24.534 48.358 24.586 48.394 ;
               RECT 24.534 50.142 24.586 50.178 ;
               RECT 24.534 50.382 24.586 50.418 ;
               RECT 24.534 54.702 24.586 54.738 ;
               RECT 24.534 54.942 24.586 54.978 ;
               RECT 24.534 57.478 24.586 57.514 ;
               RECT 24.534 58.678 24.586 58.714 ;
               RECT 24.534 59.878 24.586 59.914 ;
               RECT 24.534 61.078 24.586 61.114 ;
               RECT 24.534 62.278 24.586 62.314 ;
               RECT 24.534 63.478 24.586 63.514 ;
               RECT 24.534 64.678 24.586 64.714 ;
               RECT 24.534 65.878 24.586 65.914 ;
               RECT 24.534 67.078 24.586 67.114 ;
               RECT 24.534 68.278 24.586 68.314 ;
               RECT 24.534 69.478 24.586 69.514 ;
               RECT 24.534 70.678 24.586 70.714 ;
               RECT 24.534 71.878 24.586 71.914 ;
               RECT 24.534 73.078 24.586 73.114 ;
               RECT 24.534 74.278 24.586 74.314 ;
               RECT 24.534 75.478 24.586 75.514 ;
               RECT 24.534 76.678 24.586 76.714 ;
               RECT 24.534 77.878 24.586 77.914 ;
               RECT 24.534 79.078 24.586 79.114 ;
               RECT 24.534 80.278 24.586 80.314 ;
               RECT 24.534 81.478 24.586 81.514 ;
               RECT 24.534 82.678 24.586 82.714 ;
               RECT 24.534 83.878 24.586 83.914 ;
               RECT 24.534 85.078 24.586 85.114 ;
               RECT 24.534 86.278 24.586 86.314 ;
               RECT 24.534 87.478 24.586 87.514 ;
               RECT 24.534 88.678 24.586 88.714 ;
               RECT 24.534 89.878 24.586 89.914 ;
               RECT 24.534 91.078 24.586 91.114 ;
               RECT 24.534 92.278 24.586 92.314 ;
               RECT 24.534 93.478 24.586 93.514 ;
               RECT 24.534 94.678 24.586 94.714 ;
               RECT 24.534 95.878 24.586 95.914 ;
               RECT 24.534 97.078 24.586 97.114 ;
               RECT 24.534 98.278 24.586 98.314 ;
               RECT 24.534 99.478 24.586 99.514 ;
               RECT 24.534 100.678 24.586 100.714 ;
               RECT 24.534 101.878 24.586 101.914 ;
               RECT 24.534 103.078 24.586 103.114 ;
               RECT 24.534 104.278 24.586 104.314 ;
               RECT 24.614 0.806 24.666 0.842 ;
               RECT 24.614 2.006 24.666 2.042 ;
               RECT 24.614 3.206 24.666 3.242 ;
               RECT 24.614 4.406 24.666 4.442 ;
               RECT 24.614 5.606 24.666 5.642 ;
               RECT 24.614 6.806 24.666 6.842 ;
               RECT 24.614 8.006 24.666 8.042 ;
               RECT 24.614 9.206 24.666 9.242 ;
               RECT 24.614 10.406 24.666 10.442 ;
               RECT 24.614 11.606 24.666 11.642 ;
               RECT 24.614 12.806 24.666 12.842 ;
               RECT 24.614 14.006 24.666 14.042 ;
               RECT 24.614 15.206 24.666 15.242 ;
               RECT 24.614 16.406 24.666 16.442 ;
               RECT 24.614 17.606 24.666 17.642 ;
               RECT 24.614 18.806 24.666 18.842 ;
               RECT 24.614 20.006 24.666 20.042 ;
               RECT 24.614 21.206 24.666 21.242 ;
               RECT 24.614 22.406 24.666 22.442 ;
               RECT 24.614 23.606 24.666 23.642 ;
               RECT 24.614 24.806 24.666 24.842 ;
               RECT 24.614 26.006 24.666 26.042 ;
               RECT 24.614 27.206 24.666 27.242 ;
               RECT 24.614 28.406 24.666 28.442 ;
               RECT 24.614 29.606 24.666 29.642 ;
               RECT 24.614 30.806 24.666 30.842 ;
               RECT 24.614 32.006 24.666 32.042 ;
               RECT 24.614 33.206 24.666 33.242 ;
               RECT 24.614 34.406 24.666 34.442 ;
               RECT 24.614 35.606 24.666 35.642 ;
               RECT 24.614 36.806 24.666 36.842 ;
               RECT 24.614 38.006 24.666 38.042 ;
               RECT 24.614 39.206 24.666 39.242 ;
               RECT 24.614 40.406 24.666 40.442 ;
               RECT 24.614 41.606 24.666 41.642 ;
               RECT 24.614 42.806 24.666 42.842 ;
               RECT 24.614 44.006 24.666 44.042 ;
               RECT 24.614 45.206 24.666 45.242 ;
               RECT 24.614 46.406 24.666 46.442 ;
               RECT 24.614 47.606 24.666 47.642 ;
               RECT 24.614 49.422 24.666 49.458 ;
               RECT 24.614 49.662 24.666 49.698 ;
               RECT 24.614 55.422 24.666 55.458 ;
               RECT 24.614 55.662 24.666 55.698 ;
               RECT 24.614 56.726 24.666 56.762 ;
               RECT 24.614 57.926 24.666 57.962 ;
               RECT 24.614 59.126 24.666 59.162 ;
               RECT 24.614 60.326 24.666 60.362 ;
               RECT 24.614 61.526 24.666 61.562 ;
               RECT 24.614 62.726 24.666 62.762 ;
               RECT 24.614 63.926 24.666 63.962 ;
               RECT 24.614 65.126 24.666 65.162 ;
               RECT 24.614 66.326 24.666 66.362 ;
               RECT 24.614 67.526 24.666 67.562 ;
               RECT 24.614 68.726 24.666 68.762 ;
               RECT 24.614 69.926 24.666 69.962 ;
               RECT 24.614 71.126 24.666 71.162 ;
               RECT 24.614 72.326 24.666 72.362 ;
               RECT 24.614 73.526 24.666 73.562 ;
               RECT 24.614 74.726 24.666 74.762 ;
               RECT 24.614 75.926 24.666 75.962 ;
               RECT 24.614 77.126 24.666 77.162 ;
               RECT 24.614 78.326 24.666 78.362 ;
               RECT 24.614 79.526 24.666 79.562 ;
               RECT 24.614 80.726 24.666 80.762 ;
               RECT 24.614 81.926 24.666 81.962 ;
               RECT 24.614 83.126 24.666 83.162 ;
               RECT 24.614 84.326 24.666 84.362 ;
               RECT 24.614 85.526 24.666 85.562 ;
               RECT 24.614 86.726 24.666 86.762 ;
               RECT 24.614 87.926 24.666 87.962 ;
               RECT 24.614 89.126 24.666 89.162 ;
               RECT 24.614 90.326 24.666 90.362 ;
               RECT 24.614 91.526 24.666 91.562 ;
               RECT 24.614 92.726 24.666 92.762 ;
               RECT 24.614 93.926 24.666 93.962 ;
               RECT 24.614 95.126 24.666 95.162 ;
               RECT 24.614 96.326 24.666 96.362 ;
               RECT 24.614 97.526 24.666 97.562 ;
               RECT 24.614 98.726 24.666 98.762 ;
               RECT 24.614 99.926 24.666 99.962 ;
               RECT 24.614 101.126 24.666 101.162 ;
               RECT 24.614 102.326 24.666 102.362 ;
               RECT 24.614 103.526 24.666 103.562 ;
               RECT 24.694 1.558 24.746 1.594 ;
               RECT 24.694 2.758 24.746 2.794 ;
               RECT 24.694 3.958 24.746 3.994 ;
               RECT 24.694 5.158 24.746 5.194 ;
               RECT 24.694 6.358 24.746 6.394 ;
               RECT 24.694 7.558 24.746 7.594 ;
               RECT 24.694 8.758 24.746 8.794 ;
               RECT 24.694 9.958 24.746 9.994 ;
               RECT 24.694 11.158 24.746 11.194 ;
               RECT 24.694 12.358 24.746 12.394 ;
               RECT 24.694 13.558 24.746 13.594 ;
               RECT 24.694 14.758 24.746 14.794 ;
               RECT 24.694 15.958 24.746 15.994 ;
               RECT 24.694 17.158 24.746 17.194 ;
               RECT 24.694 18.358 24.746 18.394 ;
               RECT 24.694 19.558 24.746 19.594 ;
               RECT 24.694 20.758 24.746 20.794 ;
               RECT 24.694 21.958 24.746 21.994 ;
               RECT 24.694 23.158 24.746 23.194 ;
               RECT 24.694 24.358 24.746 24.394 ;
               RECT 24.694 25.558 24.746 25.594 ;
               RECT 24.694 26.758 24.746 26.794 ;
               RECT 24.694 27.958 24.746 27.994 ;
               RECT 24.694 29.158 24.746 29.194 ;
               RECT 24.694 30.358 24.746 30.394 ;
               RECT 24.694 31.558 24.746 31.594 ;
               RECT 24.694 32.758 24.746 32.794 ;
               RECT 24.694 33.958 24.746 33.994 ;
               RECT 24.694 35.158 24.746 35.194 ;
               RECT 24.694 36.358 24.746 36.394 ;
               RECT 24.694 37.558 24.746 37.594 ;
               RECT 24.694 38.758 24.746 38.794 ;
               RECT 24.694 39.958 24.746 39.994 ;
               RECT 24.694 41.158 24.746 41.194 ;
               RECT 24.694 42.358 24.746 42.394 ;
               RECT 24.694 43.558 24.746 43.594 ;
               RECT 24.694 44.758 24.746 44.794 ;
               RECT 24.694 45.958 24.746 45.994 ;
               RECT 24.694 47.158 24.746 47.194 ;
               RECT 24.694 48.358 24.746 48.394 ;
               RECT 24.694 50.142 24.746 50.178 ;
               RECT 24.694 50.382 24.746 50.418 ;
               RECT 24.694 54.702 24.746 54.738 ;
               RECT 24.694 54.942 24.746 54.978 ;
               RECT 24.694 57.478 24.746 57.514 ;
               RECT 24.694 58.678 24.746 58.714 ;
               RECT 24.694 59.878 24.746 59.914 ;
               RECT 24.694 61.078 24.746 61.114 ;
               RECT 24.694 62.278 24.746 62.314 ;
               RECT 24.694 63.478 24.746 63.514 ;
               RECT 24.694 64.678 24.746 64.714 ;
               RECT 24.694 65.878 24.746 65.914 ;
               RECT 24.694 67.078 24.746 67.114 ;
               RECT 24.694 68.278 24.746 68.314 ;
               RECT 24.694 69.478 24.746 69.514 ;
               RECT 24.694 70.678 24.746 70.714 ;
               RECT 24.694 71.878 24.746 71.914 ;
               RECT 24.694 73.078 24.746 73.114 ;
               RECT 24.694 74.278 24.746 74.314 ;
               RECT 24.694 75.478 24.746 75.514 ;
               RECT 24.694 76.678 24.746 76.714 ;
               RECT 24.694 77.878 24.746 77.914 ;
               RECT 24.694 79.078 24.746 79.114 ;
               RECT 24.694 80.278 24.746 80.314 ;
               RECT 24.694 81.478 24.746 81.514 ;
               RECT 24.694 82.678 24.746 82.714 ;
               RECT 24.694 83.878 24.746 83.914 ;
               RECT 24.694 85.078 24.746 85.114 ;
               RECT 24.694 86.278 24.746 86.314 ;
               RECT 24.694 87.478 24.746 87.514 ;
               RECT 24.694 88.678 24.746 88.714 ;
               RECT 24.694 89.878 24.746 89.914 ;
               RECT 24.694 91.078 24.746 91.114 ;
               RECT 24.694 92.278 24.746 92.314 ;
               RECT 24.694 93.478 24.746 93.514 ;
               RECT 24.694 94.678 24.746 94.714 ;
               RECT 24.694 95.878 24.746 95.914 ;
               RECT 24.694 97.078 24.746 97.114 ;
               RECT 24.694 98.278 24.746 98.314 ;
               RECT 24.694 99.478 24.746 99.514 ;
               RECT 24.694 100.678 24.746 100.714 ;
               RECT 24.694 101.878 24.746 101.914 ;
               RECT 24.694 103.078 24.746 103.114 ;
               RECT 24.694 104.278 24.746 104.314 ;
               RECT 24.774 0.281 24.826 0.317 ;
               RECT 24.774 104.803 24.826 104.839 ;
               RECT 24.854 0.806 24.906 0.842 ;
               RECT 24.854 2.006 24.906 2.042 ;
               RECT 24.854 3.206 24.906 3.242 ;
               RECT 24.854 4.406 24.906 4.442 ;
               RECT 24.854 5.606 24.906 5.642 ;
               RECT 24.854 6.806 24.906 6.842 ;
               RECT 24.854 8.006 24.906 8.042 ;
               RECT 24.854 9.206 24.906 9.242 ;
               RECT 24.854 10.406 24.906 10.442 ;
               RECT 24.854 11.606 24.906 11.642 ;
               RECT 24.854 12.806 24.906 12.842 ;
               RECT 24.854 14.006 24.906 14.042 ;
               RECT 24.854 15.206 24.906 15.242 ;
               RECT 24.854 16.406 24.906 16.442 ;
               RECT 24.854 17.606 24.906 17.642 ;
               RECT 24.854 18.806 24.906 18.842 ;
               RECT 24.854 20.006 24.906 20.042 ;
               RECT 24.854 21.206 24.906 21.242 ;
               RECT 24.854 22.406 24.906 22.442 ;
               RECT 24.854 23.606 24.906 23.642 ;
               RECT 24.854 24.806 24.906 24.842 ;
               RECT 24.854 26.006 24.906 26.042 ;
               RECT 24.854 27.206 24.906 27.242 ;
               RECT 24.854 28.406 24.906 28.442 ;
               RECT 24.854 29.606 24.906 29.642 ;
               RECT 24.854 30.806 24.906 30.842 ;
               RECT 24.854 32.006 24.906 32.042 ;
               RECT 24.854 33.206 24.906 33.242 ;
               RECT 24.854 34.406 24.906 34.442 ;
               RECT 24.854 35.606 24.906 35.642 ;
               RECT 24.854 36.806 24.906 36.842 ;
               RECT 24.854 38.006 24.906 38.042 ;
               RECT 24.854 39.206 24.906 39.242 ;
               RECT 24.854 40.406 24.906 40.442 ;
               RECT 24.854 41.606 24.906 41.642 ;
               RECT 24.854 42.806 24.906 42.842 ;
               RECT 24.854 44.006 24.906 44.042 ;
               RECT 24.854 45.206 24.906 45.242 ;
               RECT 24.854 46.406 24.906 46.442 ;
               RECT 24.854 47.606 24.906 47.642 ;
               RECT 24.854 49.422 24.906 49.458 ;
               RECT 24.854 49.662 24.906 49.698 ;
               RECT 24.854 51.102 24.906 51.138 ;
               RECT 24.854 51.582 24.906 51.618 ;
               RECT 24.854 53.502 24.906 53.538 ;
               RECT 24.854 53.982 24.906 54.018 ;
               RECT 24.854 55.422 24.906 55.458 ;
               RECT 24.854 55.662 24.906 55.698 ;
               RECT 24.854 56.726 24.906 56.762 ;
               RECT 24.854 57.926 24.906 57.962 ;
               RECT 24.854 59.126 24.906 59.162 ;
               RECT 24.854 60.326 24.906 60.362 ;
               RECT 24.854 61.526 24.906 61.562 ;
               RECT 24.854 62.726 24.906 62.762 ;
               RECT 24.854 63.926 24.906 63.962 ;
               RECT 24.854 65.126 24.906 65.162 ;
               RECT 24.854 66.326 24.906 66.362 ;
               RECT 24.854 67.526 24.906 67.562 ;
               RECT 24.854 68.726 24.906 68.762 ;
               RECT 24.854 69.926 24.906 69.962 ;
               RECT 24.854 71.126 24.906 71.162 ;
               RECT 24.854 72.326 24.906 72.362 ;
               RECT 24.854 73.526 24.906 73.562 ;
               RECT 24.854 74.726 24.906 74.762 ;
               RECT 24.854 75.926 24.906 75.962 ;
               RECT 24.854 77.126 24.906 77.162 ;
               RECT 24.854 78.326 24.906 78.362 ;
               RECT 24.854 79.526 24.906 79.562 ;
               RECT 24.854 80.726 24.906 80.762 ;
               RECT 24.854 81.926 24.906 81.962 ;
               RECT 24.854 83.126 24.906 83.162 ;
               RECT 24.854 84.326 24.906 84.362 ;
               RECT 24.854 85.526 24.906 85.562 ;
               RECT 24.854 86.726 24.906 86.762 ;
               RECT 24.854 87.926 24.906 87.962 ;
               RECT 24.854 89.126 24.906 89.162 ;
               RECT 24.854 90.326 24.906 90.362 ;
               RECT 24.854 91.526 24.906 91.562 ;
               RECT 24.854 92.726 24.906 92.762 ;
               RECT 24.854 93.926 24.906 93.962 ;
               RECT 24.854 95.126 24.906 95.162 ;
               RECT 24.854 96.326 24.906 96.362 ;
               RECT 24.854 97.526 24.906 97.562 ;
               RECT 24.854 98.726 24.906 98.762 ;
               RECT 24.854 99.926 24.906 99.962 ;
               RECT 24.854 101.126 24.906 101.162 ;
               RECT 24.854 102.326 24.906 102.362 ;
               RECT 24.854 103.526 24.906 103.562 ;
               RECT 24.934 1.558 24.986 1.594 ;
               RECT 24.934 2.758 24.986 2.794 ;
               RECT 24.934 3.958 24.986 3.994 ;
               RECT 24.934 5.158 24.986 5.194 ;
               RECT 24.934 6.358 24.986 6.394 ;
               RECT 24.934 7.558 24.986 7.594 ;
               RECT 24.934 8.758 24.986 8.794 ;
               RECT 24.934 9.958 24.986 9.994 ;
               RECT 24.934 11.158 24.986 11.194 ;
               RECT 24.934 12.358 24.986 12.394 ;
               RECT 24.934 13.558 24.986 13.594 ;
               RECT 24.934 14.758 24.986 14.794 ;
               RECT 24.934 15.958 24.986 15.994 ;
               RECT 24.934 17.158 24.986 17.194 ;
               RECT 24.934 18.358 24.986 18.394 ;
               RECT 24.934 19.558 24.986 19.594 ;
               RECT 24.934 20.758 24.986 20.794 ;
               RECT 24.934 21.958 24.986 21.994 ;
               RECT 24.934 23.158 24.986 23.194 ;
               RECT 24.934 24.358 24.986 24.394 ;
               RECT 24.934 25.558 24.986 25.594 ;
               RECT 24.934 26.758 24.986 26.794 ;
               RECT 24.934 27.958 24.986 27.994 ;
               RECT 24.934 29.158 24.986 29.194 ;
               RECT 24.934 30.358 24.986 30.394 ;
               RECT 24.934 31.558 24.986 31.594 ;
               RECT 24.934 32.758 24.986 32.794 ;
               RECT 24.934 33.958 24.986 33.994 ;
               RECT 24.934 35.158 24.986 35.194 ;
               RECT 24.934 36.358 24.986 36.394 ;
               RECT 24.934 37.558 24.986 37.594 ;
               RECT 24.934 38.758 24.986 38.794 ;
               RECT 24.934 39.958 24.986 39.994 ;
               RECT 24.934 41.158 24.986 41.194 ;
               RECT 24.934 42.358 24.986 42.394 ;
               RECT 24.934 43.558 24.986 43.594 ;
               RECT 24.934 44.758 24.986 44.794 ;
               RECT 24.934 45.958 24.986 45.994 ;
               RECT 24.934 47.158 24.986 47.194 ;
               RECT 24.934 48.358 24.986 48.394 ;
               RECT 24.934 50.142 24.986 50.178 ;
               RECT 24.934 50.382 24.986 50.418 ;
               RECT 24.934 54.702 24.986 54.738 ;
               RECT 24.934 54.942 24.986 54.978 ;
               RECT 24.934 57.478 24.986 57.514 ;
               RECT 24.934 58.678 24.986 58.714 ;
               RECT 24.934 59.878 24.986 59.914 ;
               RECT 24.934 61.078 24.986 61.114 ;
               RECT 24.934 62.278 24.986 62.314 ;
               RECT 24.934 63.478 24.986 63.514 ;
               RECT 24.934 64.678 24.986 64.714 ;
               RECT 24.934 65.878 24.986 65.914 ;
               RECT 24.934 67.078 24.986 67.114 ;
               RECT 24.934 68.278 24.986 68.314 ;
               RECT 24.934 69.478 24.986 69.514 ;
               RECT 24.934 70.678 24.986 70.714 ;
               RECT 24.934 71.878 24.986 71.914 ;
               RECT 24.934 73.078 24.986 73.114 ;
               RECT 24.934 74.278 24.986 74.314 ;
               RECT 24.934 75.478 24.986 75.514 ;
               RECT 24.934 76.678 24.986 76.714 ;
               RECT 24.934 77.878 24.986 77.914 ;
               RECT 24.934 79.078 24.986 79.114 ;
               RECT 24.934 80.278 24.986 80.314 ;
               RECT 24.934 81.478 24.986 81.514 ;
               RECT 24.934 82.678 24.986 82.714 ;
               RECT 24.934 83.878 24.986 83.914 ;
               RECT 24.934 85.078 24.986 85.114 ;
               RECT 24.934 86.278 24.986 86.314 ;
               RECT 24.934 87.478 24.986 87.514 ;
               RECT 24.934 88.678 24.986 88.714 ;
               RECT 24.934 89.878 24.986 89.914 ;
               RECT 24.934 91.078 24.986 91.114 ;
               RECT 24.934 92.278 24.986 92.314 ;
               RECT 24.934 93.478 24.986 93.514 ;
               RECT 24.934 94.678 24.986 94.714 ;
               RECT 24.934 95.878 24.986 95.914 ;
               RECT 24.934 97.078 24.986 97.114 ;
               RECT 24.934 98.278 24.986 98.314 ;
               RECT 24.934 99.478 24.986 99.514 ;
               RECT 24.934 100.678 24.986 100.714 ;
               RECT 24.934 101.878 24.986 101.914 ;
               RECT 24.934 103.078 24.986 103.114 ;
               RECT 24.934 104.278 24.986 104.314 ;
               RECT 25.014 0.806 25.066 0.842 ;
               RECT 25.014 2.006 25.066 2.042 ;
               RECT 25.014 3.206 25.066 3.242 ;
               RECT 25.014 4.406 25.066 4.442 ;
               RECT 25.014 5.606 25.066 5.642 ;
               RECT 25.014 6.806 25.066 6.842 ;
               RECT 25.014 8.006 25.066 8.042 ;
               RECT 25.014 9.206 25.066 9.242 ;
               RECT 25.014 10.406 25.066 10.442 ;
               RECT 25.014 11.606 25.066 11.642 ;
               RECT 25.014 12.806 25.066 12.842 ;
               RECT 25.014 14.006 25.066 14.042 ;
               RECT 25.014 15.206 25.066 15.242 ;
               RECT 25.014 16.406 25.066 16.442 ;
               RECT 25.014 17.606 25.066 17.642 ;
               RECT 25.014 18.806 25.066 18.842 ;
               RECT 25.014 20.006 25.066 20.042 ;
               RECT 25.014 21.206 25.066 21.242 ;
               RECT 25.014 22.406 25.066 22.442 ;
               RECT 25.014 23.606 25.066 23.642 ;
               RECT 25.014 24.806 25.066 24.842 ;
               RECT 25.014 26.006 25.066 26.042 ;
               RECT 25.014 27.206 25.066 27.242 ;
               RECT 25.014 28.406 25.066 28.442 ;
               RECT 25.014 29.606 25.066 29.642 ;
               RECT 25.014 30.806 25.066 30.842 ;
               RECT 25.014 32.006 25.066 32.042 ;
               RECT 25.014 33.206 25.066 33.242 ;
               RECT 25.014 34.406 25.066 34.442 ;
               RECT 25.014 35.606 25.066 35.642 ;
               RECT 25.014 36.806 25.066 36.842 ;
               RECT 25.014 38.006 25.066 38.042 ;
               RECT 25.014 39.206 25.066 39.242 ;
               RECT 25.014 40.406 25.066 40.442 ;
               RECT 25.014 41.606 25.066 41.642 ;
               RECT 25.014 42.806 25.066 42.842 ;
               RECT 25.014 44.006 25.066 44.042 ;
               RECT 25.014 45.206 25.066 45.242 ;
               RECT 25.014 46.406 25.066 46.442 ;
               RECT 25.014 47.606 25.066 47.642 ;
               RECT 25.014 49.422 25.066 49.458 ;
               RECT 25.014 49.662 25.066 49.698 ;
               RECT 25.014 55.422 25.066 55.458 ;
               RECT 25.014 55.662 25.066 55.698 ;
               RECT 25.014 56.726 25.066 56.762 ;
               RECT 25.014 57.926 25.066 57.962 ;
               RECT 25.014 59.126 25.066 59.162 ;
               RECT 25.014 60.326 25.066 60.362 ;
               RECT 25.014 61.526 25.066 61.562 ;
               RECT 25.014 62.726 25.066 62.762 ;
               RECT 25.014 63.926 25.066 63.962 ;
               RECT 25.014 65.126 25.066 65.162 ;
               RECT 25.014 66.326 25.066 66.362 ;
               RECT 25.014 67.526 25.066 67.562 ;
               RECT 25.014 68.726 25.066 68.762 ;
               RECT 25.014 69.926 25.066 69.962 ;
               RECT 25.014 71.126 25.066 71.162 ;
               RECT 25.014 72.326 25.066 72.362 ;
               RECT 25.014 73.526 25.066 73.562 ;
               RECT 25.014 74.726 25.066 74.762 ;
               RECT 25.014 75.926 25.066 75.962 ;
               RECT 25.014 77.126 25.066 77.162 ;
               RECT 25.014 78.326 25.066 78.362 ;
               RECT 25.014 79.526 25.066 79.562 ;
               RECT 25.014 80.726 25.066 80.762 ;
               RECT 25.014 81.926 25.066 81.962 ;
               RECT 25.014 83.126 25.066 83.162 ;
               RECT 25.014 84.326 25.066 84.362 ;
               RECT 25.014 85.526 25.066 85.562 ;
               RECT 25.014 86.726 25.066 86.762 ;
               RECT 25.014 87.926 25.066 87.962 ;
               RECT 25.014 89.126 25.066 89.162 ;
               RECT 25.014 90.326 25.066 90.362 ;
               RECT 25.014 91.526 25.066 91.562 ;
               RECT 25.014 92.726 25.066 92.762 ;
               RECT 25.014 93.926 25.066 93.962 ;
               RECT 25.014 95.126 25.066 95.162 ;
               RECT 25.014 96.326 25.066 96.362 ;
               RECT 25.014 97.526 25.066 97.562 ;
               RECT 25.014 98.726 25.066 98.762 ;
               RECT 25.014 99.926 25.066 99.962 ;
               RECT 25.014 101.126 25.066 101.162 ;
               RECT 25.014 102.326 25.066 102.362 ;
               RECT 25.014 103.526 25.066 103.562 ;
               RECT 25.094 1.558 25.146 1.594 ;
               RECT 25.094 2.758 25.146 2.794 ;
               RECT 25.094 3.958 25.146 3.994 ;
               RECT 25.094 5.158 25.146 5.194 ;
               RECT 25.094 6.358 25.146 6.394 ;
               RECT 25.094 7.558 25.146 7.594 ;
               RECT 25.094 8.758 25.146 8.794 ;
               RECT 25.094 9.958 25.146 9.994 ;
               RECT 25.094 11.158 25.146 11.194 ;
               RECT 25.094 12.358 25.146 12.394 ;
               RECT 25.094 13.558 25.146 13.594 ;
               RECT 25.094 14.758 25.146 14.794 ;
               RECT 25.094 15.958 25.146 15.994 ;
               RECT 25.094 17.158 25.146 17.194 ;
               RECT 25.094 18.358 25.146 18.394 ;
               RECT 25.094 19.558 25.146 19.594 ;
               RECT 25.094 20.758 25.146 20.794 ;
               RECT 25.094 21.958 25.146 21.994 ;
               RECT 25.094 23.158 25.146 23.194 ;
               RECT 25.094 24.358 25.146 24.394 ;
               RECT 25.094 25.558 25.146 25.594 ;
               RECT 25.094 26.758 25.146 26.794 ;
               RECT 25.094 27.958 25.146 27.994 ;
               RECT 25.094 29.158 25.146 29.194 ;
               RECT 25.094 30.358 25.146 30.394 ;
               RECT 25.094 31.558 25.146 31.594 ;
               RECT 25.094 32.758 25.146 32.794 ;
               RECT 25.094 33.958 25.146 33.994 ;
               RECT 25.094 35.158 25.146 35.194 ;
               RECT 25.094 36.358 25.146 36.394 ;
               RECT 25.094 37.558 25.146 37.594 ;
               RECT 25.094 38.758 25.146 38.794 ;
               RECT 25.094 39.958 25.146 39.994 ;
               RECT 25.094 41.158 25.146 41.194 ;
               RECT 25.094 42.358 25.146 42.394 ;
               RECT 25.094 43.558 25.146 43.594 ;
               RECT 25.094 44.758 25.146 44.794 ;
               RECT 25.094 45.958 25.146 45.994 ;
               RECT 25.094 47.158 25.146 47.194 ;
               RECT 25.094 48.358 25.146 48.394 ;
               RECT 25.094 50.142 25.146 50.178 ;
               RECT 25.094 50.382 25.146 50.418 ;
               RECT 25.094 54.702 25.146 54.738 ;
               RECT 25.094 54.942 25.146 54.978 ;
               RECT 25.094 57.478 25.146 57.514 ;
               RECT 25.094 58.678 25.146 58.714 ;
               RECT 25.094 59.878 25.146 59.914 ;
               RECT 25.094 61.078 25.146 61.114 ;
               RECT 25.094 62.278 25.146 62.314 ;
               RECT 25.094 63.478 25.146 63.514 ;
               RECT 25.094 64.678 25.146 64.714 ;
               RECT 25.094 65.878 25.146 65.914 ;
               RECT 25.094 67.078 25.146 67.114 ;
               RECT 25.094 68.278 25.146 68.314 ;
               RECT 25.094 69.478 25.146 69.514 ;
               RECT 25.094 70.678 25.146 70.714 ;
               RECT 25.094 71.878 25.146 71.914 ;
               RECT 25.094 73.078 25.146 73.114 ;
               RECT 25.094 74.278 25.146 74.314 ;
               RECT 25.094 75.478 25.146 75.514 ;
               RECT 25.094 76.678 25.146 76.714 ;
               RECT 25.094 77.878 25.146 77.914 ;
               RECT 25.094 79.078 25.146 79.114 ;
               RECT 25.094 80.278 25.146 80.314 ;
               RECT 25.094 81.478 25.146 81.514 ;
               RECT 25.094 82.678 25.146 82.714 ;
               RECT 25.094 83.878 25.146 83.914 ;
               RECT 25.094 85.078 25.146 85.114 ;
               RECT 25.094 86.278 25.146 86.314 ;
               RECT 25.094 87.478 25.146 87.514 ;
               RECT 25.094 88.678 25.146 88.714 ;
               RECT 25.094 89.878 25.146 89.914 ;
               RECT 25.094 91.078 25.146 91.114 ;
               RECT 25.094 92.278 25.146 92.314 ;
               RECT 25.094 93.478 25.146 93.514 ;
               RECT 25.094 94.678 25.146 94.714 ;
               RECT 25.094 95.878 25.146 95.914 ;
               RECT 25.094 97.078 25.146 97.114 ;
               RECT 25.094 98.278 25.146 98.314 ;
               RECT 25.094 99.478 25.146 99.514 ;
               RECT 25.094 100.678 25.146 100.714 ;
               RECT 25.094 101.878 25.146 101.914 ;
               RECT 25.094 103.078 25.146 103.114 ;
               RECT 25.094 104.278 25.146 104.314 ;
               RECT 25.174 0.281 25.226 0.317 ;
               RECT 25.174 104.803 25.226 104.839 ;
               RECT 25.254 0.806 25.306 0.842 ;
               RECT 25.254 2.006 25.306 2.042 ;
               RECT 25.254 3.206 25.306 3.242 ;
               RECT 25.254 4.406 25.306 4.442 ;
               RECT 25.254 5.606 25.306 5.642 ;
               RECT 25.254 6.806 25.306 6.842 ;
               RECT 25.254 8.006 25.306 8.042 ;
               RECT 25.254 9.206 25.306 9.242 ;
               RECT 25.254 10.406 25.306 10.442 ;
               RECT 25.254 11.606 25.306 11.642 ;
               RECT 25.254 12.806 25.306 12.842 ;
               RECT 25.254 14.006 25.306 14.042 ;
               RECT 25.254 15.206 25.306 15.242 ;
               RECT 25.254 16.406 25.306 16.442 ;
               RECT 25.254 17.606 25.306 17.642 ;
               RECT 25.254 18.806 25.306 18.842 ;
               RECT 25.254 20.006 25.306 20.042 ;
               RECT 25.254 21.206 25.306 21.242 ;
               RECT 25.254 22.406 25.306 22.442 ;
               RECT 25.254 23.606 25.306 23.642 ;
               RECT 25.254 24.806 25.306 24.842 ;
               RECT 25.254 26.006 25.306 26.042 ;
               RECT 25.254 27.206 25.306 27.242 ;
               RECT 25.254 28.406 25.306 28.442 ;
               RECT 25.254 29.606 25.306 29.642 ;
               RECT 25.254 30.806 25.306 30.842 ;
               RECT 25.254 32.006 25.306 32.042 ;
               RECT 25.254 33.206 25.306 33.242 ;
               RECT 25.254 34.406 25.306 34.442 ;
               RECT 25.254 35.606 25.306 35.642 ;
               RECT 25.254 36.806 25.306 36.842 ;
               RECT 25.254 38.006 25.306 38.042 ;
               RECT 25.254 39.206 25.306 39.242 ;
               RECT 25.254 40.406 25.306 40.442 ;
               RECT 25.254 41.606 25.306 41.642 ;
               RECT 25.254 42.806 25.306 42.842 ;
               RECT 25.254 44.006 25.306 44.042 ;
               RECT 25.254 45.206 25.306 45.242 ;
               RECT 25.254 46.406 25.306 46.442 ;
               RECT 25.254 47.606 25.306 47.642 ;
               RECT 25.254 49.422 25.306 49.458 ;
               RECT 25.254 49.662 25.306 49.698 ;
               RECT 25.254 55.422 25.306 55.458 ;
               RECT 25.254 55.662 25.306 55.698 ;
               RECT 25.254 56.726 25.306 56.762 ;
               RECT 25.254 57.926 25.306 57.962 ;
               RECT 25.254 59.126 25.306 59.162 ;
               RECT 25.254 60.326 25.306 60.362 ;
               RECT 25.254 61.526 25.306 61.562 ;
               RECT 25.254 62.726 25.306 62.762 ;
               RECT 25.254 63.926 25.306 63.962 ;
               RECT 25.254 65.126 25.306 65.162 ;
               RECT 25.254 66.326 25.306 66.362 ;
               RECT 25.254 67.526 25.306 67.562 ;
               RECT 25.254 68.726 25.306 68.762 ;
               RECT 25.254 69.926 25.306 69.962 ;
               RECT 25.254 71.126 25.306 71.162 ;
               RECT 25.254 72.326 25.306 72.362 ;
               RECT 25.254 73.526 25.306 73.562 ;
               RECT 25.254 74.726 25.306 74.762 ;
               RECT 25.254 75.926 25.306 75.962 ;
               RECT 25.254 77.126 25.306 77.162 ;
               RECT 25.254 78.326 25.306 78.362 ;
               RECT 25.254 79.526 25.306 79.562 ;
               RECT 25.254 80.726 25.306 80.762 ;
               RECT 25.254 81.926 25.306 81.962 ;
               RECT 25.254 83.126 25.306 83.162 ;
               RECT 25.254 84.326 25.306 84.362 ;
               RECT 25.254 85.526 25.306 85.562 ;
               RECT 25.254 86.726 25.306 86.762 ;
               RECT 25.254 87.926 25.306 87.962 ;
               RECT 25.254 89.126 25.306 89.162 ;
               RECT 25.254 90.326 25.306 90.362 ;
               RECT 25.254 91.526 25.306 91.562 ;
               RECT 25.254 92.726 25.306 92.762 ;
               RECT 25.254 93.926 25.306 93.962 ;
               RECT 25.254 95.126 25.306 95.162 ;
               RECT 25.254 96.326 25.306 96.362 ;
               RECT 25.254 97.526 25.306 97.562 ;
               RECT 25.254 98.726 25.306 98.762 ;
               RECT 25.254 99.926 25.306 99.962 ;
               RECT 25.254 101.126 25.306 101.162 ;
               RECT 25.254 102.326 25.306 102.362 ;
               RECT 25.254 103.526 25.306 103.562 ;
               RECT 25.334 1.558 25.386 1.594 ;
               RECT 25.334 2.758 25.386 2.794 ;
               RECT 25.334 3.958 25.386 3.994 ;
               RECT 25.334 5.158 25.386 5.194 ;
               RECT 25.334 6.358 25.386 6.394 ;
               RECT 25.334 7.558 25.386 7.594 ;
               RECT 25.334 8.758 25.386 8.794 ;
               RECT 25.334 9.958 25.386 9.994 ;
               RECT 25.334 11.158 25.386 11.194 ;
               RECT 25.334 12.358 25.386 12.394 ;
               RECT 25.334 13.558 25.386 13.594 ;
               RECT 25.334 14.758 25.386 14.794 ;
               RECT 25.334 15.958 25.386 15.994 ;
               RECT 25.334 17.158 25.386 17.194 ;
               RECT 25.334 18.358 25.386 18.394 ;
               RECT 25.334 19.558 25.386 19.594 ;
               RECT 25.334 20.758 25.386 20.794 ;
               RECT 25.334 21.958 25.386 21.994 ;
               RECT 25.334 23.158 25.386 23.194 ;
               RECT 25.334 24.358 25.386 24.394 ;
               RECT 25.334 25.558 25.386 25.594 ;
               RECT 25.334 26.758 25.386 26.794 ;
               RECT 25.334 27.958 25.386 27.994 ;
               RECT 25.334 29.158 25.386 29.194 ;
               RECT 25.334 30.358 25.386 30.394 ;
               RECT 25.334 31.558 25.386 31.594 ;
               RECT 25.334 32.758 25.386 32.794 ;
               RECT 25.334 33.958 25.386 33.994 ;
               RECT 25.334 35.158 25.386 35.194 ;
               RECT 25.334 36.358 25.386 36.394 ;
               RECT 25.334 37.558 25.386 37.594 ;
               RECT 25.334 38.758 25.386 38.794 ;
               RECT 25.334 39.958 25.386 39.994 ;
               RECT 25.334 41.158 25.386 41.194 ;
               RECT 25.334 42.358 25.386 42.394 ;
               RECT 25.334 43.558 25.386 43.594 ;
               RECT 25.334 44.758 25.386 44.794 ;
               RECT 25.334 45.958 25.386 45.994 ;
               RECT 25.334 47.158 25.386 47.194 ;
               RECT 25.334 48.358 25.386 48.394 ;
               RECT 25.334 50.142 25.386 50.178 ;
               RECT 25.334 50.382 25.386 50.418 ;
               RECT 25.334 54.702 25.386 54.738 ;
               RECT 25.334 54.942 25.386 54.978 ;
               RECT 25.334 57.478 25.386 57.514 ;
               RECT 25.334 58.678 25.386 58.714 ;
               RECT 25.334 59.878 25.386 59.914 ;
               RECT 25.334 61.078 25.386 61.114 ;
               RECT 25.334 62.278 25.386 62.314 ;
               RECT 25.334 63.478 25.386 63.514 ;
               RECT 25.334 64.678 25.386 64.714 ;
               RECT 25.334 65.878 25.386 65.914 ;
               RECT 25.334 67.078 25.386 67.114 ;
               RECT 25.334 68.278 25.386 68.314 ;
               RECT 25.334 69.478 25.386 69.514 ;
               RECT 25.334 70.678 25.386 70.714 ;
               RECT 25.334 71.878 25.386 71.914 ;
               RECT 25.334 73.078 25.386 73.114 ;
               RECT 25.334 74.278 25.386 74.314 ;
               RECT 25.334 75.478 25.386 75.514 ;
               RECT 25.334 76.678 25.386 76.714 ;
               RECT 25.334 77.878 25.386 77.914 ;
               RECT 25.334 79.078 25.386 79.114 ;
               RECT 25.334 80.278 25.386 80.314 ;
               RECT 25.334 81.478 25.386 81.514 ;
               RECT 25.334 82.678 25.386 82.714 ;
               RECT 25.334 83.878 25.386 83.914 ;
               RECT 25.334 85.078 25.386 85.114 ;
               RECT 25.334 86.278 25.386 86.314 ;
               RECT 25.334 87.478 25.386 87.514 ;
               RECT 25.334 88.678 25.386 88.714 ;
               RECT 25.334 89.878 25.386 89.914 ;
               RECT 25.334 91.078 25.386 91.114 ;
               RECT 25.334 92.278 25.386 92.314 ;
               RECT 25.334 93.478 25.386 93.514 ;
               RECT 25.334 94.678 25.386 94.714 ;
               RECT 25.334 95.878 25.386 95.914 ;
               RECT 25.334 97.078 25.386 97.114 ;
               RECT 25.334 98.278 25.386 98.314 ;
               RECT 25.334 99.478 25.386 99.514 ;
               RECT 25.334 100.678 25.386 100.714 ;
               RECT 25.334 101.878 25.386 101.914 ;
               RECT 25.334 103.078 25.386 103.114 ;
               RECT 25.334 104.278 25.386 104.314 ;
               RECT 25.414 0.806 25.466 0.842 ;
               RECT 25.414 2.006 25.466 2.042 ;
               RECT 25.414 3.206 25.466 3.242 ;
               RECT 25.414 4.406 25.466 4.442 ;
               RECT 25.414 5.606 25.466 5.642 ;
               RECT 25.414 6.806 25.466 6.842 ;
               RECT 25.414 8.006 25.466 8.042 ;
               RECT 25.414 9.206 25.466 9.242 ;
               RECT 25.414 10.406 25.466 10.442 ;
               RECT 25.414 11.606 25.466 11.642 ;
               RECT 25.414 12.806 25.466 12.842 ;
               RECT 25.414 14.006 25.466 14.042 ;
               RECT 25.414 15.206 25.466 15.242 ;
               RECT 25.414 16.406 25.466 16.442 ;
               RECT 25.414 17.606 25.466 17.642 ;
               RECT 25.414 18.806 25.466 18.842 ;
               RECT 25.414 20.006 25.466 20.042 ;
               RECT 25.414 21.206 25.466 21.242 ;
               RECT 25.414 22.406 25.466 22.442 ;
               RECT 25.414 23.606 25.466 23.642 ;
               RECT 25.414 24.806 25.466 24.842 ;
               RECT 25.414 26.006 25.466 26.042 ;
               RECT 25.414 27.206 25.466 27.242 ;
               RECT 25.414 28.406 25.466 28.442 ;
               RECT 25.414 29.606 25.466 29.642 ;
               RECT 25.414 30.806 25.466 30.842 ;
               RECT 25.414 32.006 25.466 32.042 ;
               RECT 25.414 33.206 25.466 33.242 ;
               RECT 25.414 34.406 25.466 34.442 ;
               RECT 25.414 35.606 25.466 35.642 ;
               RECT 25.414 36.806 25.466 36.842 ;
               RECT 25.414 38.006 25.466 38.042 ;
               RECT 25.414 39.206 25.466 39.242 ;
               RECT 25.414 40.406 25.466 40.442 ;
               RECT 25.414 41.606 25.466 41.642 ;
               RECT 25.414 42.806 25.466 42.842 ;
               RECT 25.414 44.006 25.466 44.042 ;
               RECT 25.414 45.206 25.466 45.242 ;
               RECT 25.414 46.406 25.466 46.442 ;
               RECT 25.414 47.606 25.466 47.642 ;
               RECT 25.414 49.422 25.466 49.458 ;
               RECT 25.414 49.662 25.466 49.698 ;
               RECT 25.414 55.422 25.466 55.458 ;
               RECT 25.414 55.662 25.466 55.698 ;
               RECT 25.414 56.726 25.466 56.762 ;
               RECT 25.414 57.926 25.466 57.962 ;
               RECT 25.414 59.126 25.466 59.162 ;
               RECT 25.414 60.326 25.466 60.362 ;
               RECT 25.414 61.526 25.466 61.562 ;
               RECT 25.414 62.726 25.466 62.762 ;
               RECT 25.414 63.926 25.466 63.962 ;
               RECT 25.414 65.126 25.466 65.162 ;
               RECT 25.414 66.326 25.466 66.362 ;
               RECT 25.414 67.526 25.466 67.562 ;
               RECT 25.414 68.726 25.466 68.762 ;
               RECT 25.414 69.926 25.466 69.962 ;
               RECT 25.414 71.126 25.466 71.162 ;
               RECT 25.414 72.326 25.466 72.362 ;
               RECT 25.414 73.526 25.466 73.562 ;
               RECT 25.414 74.726 25.466 74.762 ;
               RECT 25.414 75.926 25.466 75.962 ;
               RECT 25.414 77.126 25.466 77.162 ;
               RECT 25.414 78.326 25.466 78.362 ;
               RECT 25.414 79.526 25.466 79.562 ;
               RECT 25.414 80.726 25.466 80.762 ;
               RECT 25.414 81.926 25.466 81.962 ;
               RECT 25.414 83.126 25.466 83.162 ;
               RECT 25.414 84.326 25.466 84.362 ;
               RECT 25.414 85.526 25.466 85.562 ;
               RECT 25.414 86.726 25.466 86.762 ;
               RECT 25.414 87.926 25.466 87.962 ;
               RECT 25.414 89.126 25.466 89.162 ;
               RECT 25.414 90.326 25.466 90.362 ;
               RECT 25.414 91.526 25.466 91.562 ;
               RECT 25.414 92.726 25.466 92.762 ;
               RECT 25.414 93.926 25.466 93.962 ;
               RECT 25.414 95.126 25.466 95.162 ;
               RECT 25.414 96.326 25.466 96.362 ;
               RECT 25.414 97.526 25.466 97.562 ;
               RECT 25.414 98.726 25.466 98.762 ;
               RECT 25.414 99.926 25.466 99.962 ;
               RECT 25.414 101.126 25.466 101.162 ;
               RECT 25.414 102.326 25.466 102.362 ;
               RECT 25.414 103.526 25.466 103.562 ;
               RECT 25.494 1.558 25.546 1.594 ;
               RECT 25.494 2.758 25.546 2.794 ;
               RECT 25.494 3.958 25.546 3.994 ;
               RECT 25.494 5.158 25.546 5.194 ;
               RECT 25.494 6.358 25.546 6.394 ;
               RECT 25.494 7.558 25.546 7.594 ;
               RECT 25.494 8.758 25.546 8.794 ;
               RECT 25.494 9.958 25.546 9.994 ;
               RECT 25.494 11.158 25.546 11.194 ;
               RECT 25.494 12.358 25.546 12.394 ;
               RECT 25.494 13.558 25.546 13.594 ;
               RECT 25.494 14.758 25.546 14.794 ;
               RECT 25.494 15.958 25.546 15.994 ;
               RECT 25.494 17.158 25.546 17.194 ;
               RECT 25.494 18.358 25.546 18.394 ;
               RECT 25.494 19.558 25.546 19.594 ;
               RECT 25.494 20.758 25.546 20.794 ;
               RECT 25.494 21.958 25.546 21.994 ;
               RECT 25.494 23.158 25.546 23.194 ;
               RECT 25.494 24.358 25.546 24.394 ;
               RECT 25.494 25.558 25.546 25.594 ;
               RECT 25.494 26.758 25.546 26.794 ;
               RECT 25.494 27.958 25.546 27.994 ;
               RECT 25.494 29.158 25.546 29.194 ;
               RECT 25.494 30.358 25.546 30.394 ;
               RECT 25.494 31.558 25.546 31.594 ;
               RECT 25.494 32.758 25.546 32.794 ;
               RECT 25.494 33.958 25.546 33.994 ;
               RECT 25.494 35.158 25.546 35.194 ;
               RECT 25.494 36.358 25.546 36.394 ;
               RECT 25.494 37.558 25.546 37.594 ;
               RECT 25.494 38.758 25.546 38.794 ;
               RECT 25.494 39.958 25.546 39.994 ;
               RECT 25.494 41.158 25.546 41.194 ;
               RECT 25.494 42.358 25.546 42.394 ;
               RECT 25.494 43.558 25.546 43.594 ;
               RECT 25.494 44.758 25.546 44.794 ;
               RECT 25.494 45.958 25.546 45.994 ;
               RECT 25.494 47.158 25.546 47.194 ;
               RECT 25.494 48.358 25.546 48.394 ;
               RECT 25.494 50.142 25.546 50.178 ;
               RECT 25.494 50.382 25.546 50.418 ;
               RECT 25.494 54.702 25.546 54.738 ;
               RECT 25.494 54.942 25.546 54.978 ;
               RECT 25.494 57.478 25.546 57.514 ;
               RECT 25.494 58.678 25.546 58.714 ;
               RECT 25.494 59.878 25.546 59.914 ;
               RECT 25.494 61.078 25.546 61.114 ;
               RECT 25.494 62.278 25.546 62.314 ;
               RECT 25.494 63.478 25.546 63.514 ;
               RECT 25.494 64.678 25.546 64.714 ;
               RECT 25.494 65.878 25.546 65.914 ;
               RECT 25.494 67.078 25.546 67.114 ;
               RECT 25.494 68.278 25.546 68.314 ;
               RECT 25.494 69.478 25.546 69.514 ;
               RECT 25.494 70.678 25.546 70.714 ;
               RECT 25.494 71.878 25.546 71.914 ;
               RECT 25.494 73.078 25.546 73.114 ;
               RECT 25.494 74.278 25.546 74.314 ;
               RECT 25.494 75.478 25.546 75.514 ;
               RECT 25.494 76.678 25.546 76.714 ;
               RECT 25.494 77.878 25.546 77.914 ;
               RECT 25.494 79.078 25.546 79.114 ;
               RECT 25.494 80.278 25.546 80.314 ;
               RECT 25.494 81.478 25.546 81.514 ;
               RECT 25.494 82.678 25.546 82.714 ;
               RECT 25.494 83.878 25.546 83.914 ;
               RECT 25.494 85.078 25.546 85.114 ;
               RECT 25.494 86.278 25.546 86.314 ;
               RECT 25.494 87.478 25.546 87.514 ;
               RECT 25.494 88.678 25.546 88.714 ;
               RECT 25.494 89.878 25.546 89.914 ;
               RECT 25.494 91.078 25.546 91.114 ;
               RECT 25.494 92.278 25.546 92.314 ;
               RECT 25.494 93.478 25.546 93.514 ;
               RECT 25.494 94.678 25.546 94.714 ;
               RECT 25.494 95.878 25.546 95.914 ;
               RECT 25.494 97.078 25.546 97.114 ;
               RECT 25.494 98.278 25.546 98.314 ;
               RECT 25.494 99.478 25.546 99.514 ;
               RECT 25.494 100.678 25.546 100.714 ;
               RECT 25.494 101.878 25.546 101.914 ;
               RECT 25.494 103.078 25.546 103.114 ;
               RECT 25.494 104.278 25.546 104.314 ;
               RECT 25.574 0.281 25.626 0.317 ;
               RECT 25.574 104.803 25.626 104.839 ;
               RECT 25.654 0.806 25.706 0.842 ;
               RECT 25.654 2.006 25.706 2.042 ;
               RECT 25.654 3.206 25.706 3.242 ;
               RECT 25.654 4.406 25.706 4.442 ;
               RECT 25.654 5.606 25.706 5.642 ;
               RECT 25.654 6.806 25.706 6.842 ;
               RECT 25.654 8.006 25.706 8.042 ;
               RECT 25.654 9.206 25.706 9.242 ;
               RECT 25.654 10.406 25.706 10.442 ;
               RECT 25.654 11.606 25.706 11.642 ;
               RECT 25.654 12.806 25.706 12.842 ;
               RECT 25.654 14.006 25.706 14.042 ;
               RECT 25.654 15.206 25.706 15.242 ;
               RECT 25.654 16.406 25.706 16.442 ;
               RECT 25.654 17.606 25.706 17.642 ;
               RECT 25.654 18.806 25.706 18.842 ;
               RECT 25.654 20.006 25.706 20.042 ;
               RECT 25.654 21.206 25.706 21.242 ;
               RECT 25.654 22.406 25.706 22.442 ;
               RECT 25.654 23.606 25.706 23.642 ;
               RECT 25.654 24.806 25.706 24.842 ;
               RECT 25.654 26.006 25.706 26.042 ;
               RECT 25.654 27.206 25.706 27.242 ;
               RECT 25.654 28.406 25.706 28.442 ;
               RECT 25.654 29.606 25.706 29.642 ;
               RECT 25.654 30.806 25.706 30.842 ;
               RECT 25.654 32.006 25.706 32.042 ;
               RECT 25.654 33.206 25.706 33.242 ;
               RECT 25.654 34.406 25.706 34.442 ;
               RECT 25.654 35.606 25.706 35.642 ;
               RECT 25.654 36.806 25.706 36.842 ;
               RECT 25.654 38.006 25.706 38.042 ;
               RECT 25.654 39.206 25.706 39.242 ;
               RECT 25.654 40.406 25.706 40.442 ;
               RECT 25.654 41.606 25.706 41.642 ;
               RECT 25.654 42.806 25.706 42.842 ;
               RECT 25.654 44.006 25.706 44.042 ;
               RECT 25.654 45.206 25.706 45.242 ;
               RECT 25.654 46.406 25.706 46.442 ;
               RECT 25.654 47.606 25.706 47.642 ;
               RECT 25.654 49.422 25.706 49.458 ;
               RECT 25.654 49.662 25.706 49.698 ;
               RECT 25.654 51.102 25.706 51.138 ;
               RECT 25.654 51.582 25.706 51.618 ;
               RECT 25.654 53.502 25.706 53.538 ;
               RECT 25.654 53.982 25.706 54.018 ;
               RECT 25.654 55.422 25.706 55.458 ;
               RECT 25.654 55.662 25.706 55.698 ;
               RECT 25.654 56.726 25.706 56.762 ;
               RECT 25.654 57.926 25.706 57.962 ;
               RECT 25.654 59.126 25.706 59.162 ;
               RECT 25.654 60.326 25.706 60.362 ;
               RECT 25.654 61.526 25.706 61.562 ;
               RECT 25.654 62.726 25.706 62.762 ;
               RECT 25.654 63.926 25.706 63.962 ;
               RECT 25.654 65.126 25.706 65.162 ;
               RECT 25.654 66.326 25.706 66.362 ;
               RECT 25.654 67.526 25.706 67.562 ;
               RECT 25.654 68.726 25.706 68.762 ;
               RECT 25.654 69.926 25.706 69.962 ;
               RECT 25.654 71.126 25.706 71.162 ;
               RECT 25.654 72.326 25.706 72.362 ;
               RECT 25.654 73.526 25.706 73.562 ;
               RECT 25.654 74.726 25.706 74.762 ;
               RECT 25.654 75.926 25.706 75.962 ;
               RECT 25.654 77.126 25.706 77.162 ;
               RECT 25.654 78.326 25.706 78.362 ;
               RECT 25.654 79.526 25.706 79.562 ;
               RECT 25.654 80.726 25.706 80.762 ;
               RECT 25.654 81.926 25.706 81.962 ;
               RECT 25.654 83.126 25.706 83.162 ;
               RECT 25.654 84.326 25.706 84.362 ;
               RECT 25.654 85.526 25.706 85.562 ;
               RECT 25.654 86.726 25.706 86.762 ;
               RECT 25.654 87.926 25.706 87.962 ;
               RECT 25.654 89.126 25.706 89.162 ;
               RECT 25.654 90.326 25.706 90.362 ;
               RECT 25.654 91.526 25.706 91.562 ;
               RECT 25.654 92.726 25.706 92.762 ;
               RECT 25.654 93.926 25.706 93.962 ;
               RECT 25.654 95.126 25.706 95.162 ;
               RECT 25.654 96.326 25.706 96.362 ;
               RECT 25.654 97.526 25.706 97.562 ;
               RECT 25.654 98.726 25.706 98.762 ;
               RECT 25.654 99.926 25.706 99.962 ;
               RECT 25.654 101.126 25.706 101.162 ;
               RECT 25.654 102.326 25.706 102.362 ;
               RECT 25.654 103.526 25.706 103.562 ;
               RECT 25.734 1.558 25.786 1.594 ;
               RECT 25.734 2.758 25.786 2.794 ;
               RECT 25.734 3.958 25.786 3.994 ;
               RECT 25.734 5.158 25.786 5.194 ;
               RECT 25.734 6.358 25.786 6.394 ;
               RECT 25.734 7.558 25.786 7.594 ;
               RECT 25.734 8.758 25.786 8.794 ;
               RECT 25.734 9.958 25.786 9.994 ;
               RECT 25.734 11.158 25.786 11.194 ;
               RECT 25.734 12.358 25.786 12.394 ;
               RECT 25.734 13.558 25.786 13.594 ;
               RECT 25.734 14.758 25.786 14.794 ;
               RECT 25.734 15.958 25.786 15.994 ;
               RECT 25.734 17.158 25.786 17.194 ;
               RECT 25.734 18.358 25.786 18.394 ;
               RECT 25.734 19.558 25.786 19.594 ;
               RECT 25.734 20.758 25.786 20.794 ;
               RECT 25.734 21.958 25.786 21.994 ;
               RECT 25.734 23.158 25.786 23.194 ;
               RECT 25.734 24.358 25.786 24.394 ;
               RECT 25.734 25.558 25.786 25.594 ;
               RECT 25.734 26.758 25.786 26.794 ;
               RECT 25.734 27.958 25.786 27.994 ;
               RECT 25.734 29.158 25.786 29.194 ;
               RECT 25.734 30.358 25.786 30.394 ;
               RECT 25.734 31.558 25.786 31.594 ;
               RECT 25.734 32.758 25.786 32.794 ;
               RECT 25.734 33.958 25.786 33.994 ;
               RECT 25.734 35.158 25.786 35.194 ;
               RECT 25.734 36.358 25.786 36.394 ;
               RECT 25.734 37.558 25.786 37.594 ;
               RECT 25.734 38.758 25.786 38.794 ;
               RECT 25.734 39.958 25.786 39.994 ;
               RECT 25.734 41.158 25.786 41.194 ;
               RECT 25.734 42.358 25.786 42.394 ;
               RECT 25.734 43.558 25.786 43.594 ;
               RECT 25.734 44.758 25.786 44.794 ;
               RECT 25.734 45.958 25.786 45.994 ;
               RECT 25.734 47.158 25.786 47.194 ;
               RECT 25.734 48.358 25.786 48.394 ;
               RECT 25.734 50.142 25.786 50.178 ;
               RECT 25.734 50.382 25.786 50.418 ;
               RECT 25.734 54.702 25.786 54.738 ;
               RECT 25.734 54.942 25.786 54.978 ;
               RECT 25.734 57.478 25.786 57.514 ;
               RECT 25.734 58.678 25.786 58.714 ;
               RECT 25.734 59.878 25.786 59.914 ;
               RECT 25.734 61.078 25.786 61.114 ;
               RECT 25.734 62.278 25.786 62.314 ;
               RECT 25.734 63.478 25.786 63.514 ;
               RECT 25.734 64.678 25.786 64.714 ;
               RECT 25.734 65.878 25.786 65.914 ;
               RECT 25.734 67.078 25.786 67.114 ;
               RECT 25.734 68.278 25.786 68.314 ;
               RECT 25.734 69.478 25.786 69.514 ;
               RECT 25.734 70.678 25.786 70.714 ;
               RECT 25.734 71.878 25.786 71.914 ;
               RECT 25.734 73.078 25.786 73.114 ;
               RECT 25.734 74.278 25.786 74.314 ;
               RECT 25.734 75.478 25.786 75.514 ;
               RECT 25.734 76.678 25.786 76.714 ;
               RECT 25.734 77.878 25.786 77.914 ;
               RECT 25.734 79.078 25.786 79.114 ;
               RECT 25.734 80.278 25.786 80.314 ;
               RECT 25.734 81.478 25.786 81.514 ;
               RECT 25.734 82.678 25.786 82.714 ;
               RECT 25.734 83.878 25.786 83.914 ;
               RECT 25.734 85.078 25.786 85.114 ;
               RECT 25.734 86.278 25.786 86.314 ;
               RECT 25.734 87.478 25.786 87.514 ;
               RECT 25.734 88.678 25.786 88.714 ;
               RECT 25.734 89.878 25.786 89.914 ;
               RECT 25.734 91.078 25.786 91.114 ;
               RECT 25.734 92.278 25.786 92.314 ;
               RECT 25.734 93.478 25.786 93.514 ;
               RECT 25.734 94.678 25.786 94.714 ;
               RECT 25.734 95.878 25.786 95.914 ;
               RECT 25.734 97.078 25.786 97.114 ;
               RECT 25.734 98.278 25.786 98.314 ;
               RECT 25.734 99.478 25.786 99.514 ;
               RECT 25.734 100.678 25.786 100.714 ;
               RECT 25.734 101.878 25.786 101.914 ;
               RECT 25.734 103.078 25.786 103.114 ;
               RECT 25.734 104.278 25.786 104.314 ;
               RECT 25.814 0.806 25.866 0.842 ;
               RECT 25.814 2.006 25.866 2.042 ;
               RECT 25.814 3.206 25.866 3.242 ;
               RECT 25.814 4.406 25.866 4.442 ;
               RECT 25.814 5.606 25.866 5.642 ;
               RECT 25.814 6.806 25.866 6.842 ;
               RECT 25.814 8.006 25.866 8.042 ;
               RECT 25.814 9.206 25.866 9.242 ;
               RECT 25.814 10.406 25.866 10.442 ;
               RECT 25.814 11.606 25.866 11.642 ;
               RECT 25.814 12.806 25.866 12.842 ;
               RECT 25.814 14.006 25.866 14.042 ;
               RECT 25.814 15.206 25.866 15.242 ;
               RECT 25.814 16.406 25.866 16.442 ;
               RECT 25.814 17.606 25.866 17.642 ;
               RECT 25.814 18.806 25.866 18.842 ;
               RECT 25.814 20.006 25.866 20.042 ;
               RECT 25.814 21.206 25.866 21.242 ;
               RECT 25.814 22.406 25.866 22.442 ;
               RECT 25.814 23.606 25.866 23.642 ;
               RECT 25.814 24.806 25.866 24.842 ;
               RECT 25.814 26.006 25.866 26.042 ;
               RECT 25.814 27.206 25.866 27.242 ;
               RECT 25.814 28.406 25.866 28.442 ;
               RECT 25.814 29.606 25.866 29.642 ;
               RECT 25.814 30.806 25.866 30.842 ;
               RECT 25.814 32.006 25.866 32.042 ;
               RECT 25.814 33.206 25.866 33.242 ;
               RECT 25.814 34.406 25.866 34.442 ;
               RECT 25.814 35.606 25.866 35.642 ;
               RECT 25.814 36.806 25.866 36.842 ;
               RECT 25.814 38.006 25.866 38.042 ;
               RECT 25.814 39.206 25.866 39.242 ;
               RECT 25.814 40.406 25.866 40.442 ;
               RECT 25.814 41.606 25.866 41.642 ;
               RECT 25.814 42.806 25.866 42.842 ;
               RECT 25.814 44.006 25.866 44.042 ;
               RECT 25.814 45.206 25.866 45.242 ;
               RECT 25.814 46.406 25.866 46.442 ;
               RECT 25.814 47.606 25.866 47.642 ;
               RECT 25.814 49.422 25.866 49.458 ;
               RECT 25.814 49.662 25.866 49.698 ;
               RECT 25.814 55.422 25.866 55.458 ;
               RECT 25.814 55.662 25.866 55.698 ;
               RECT 25.814 56.726 25.866 56.762 ;
               RECT 25.814 57.926 25.866 57.962 ;
               RECT 25.814 59.126 25.866 59.162 ;
               RECT 25.814 60.326 25.866 60.362 ;
               RECT 25.814 61.526 25.866 61.562 ;
               RECT 25.814 62.726 25.866 62.762 ;
               RECT 25.814 63.926 25.866 63.962 ;
               RECT 25.814 65.126 25.866 65.162 ;
               RECT 25.814 66.326 25.866 66.362 ;
               RECT 25.814 67.526 25.866 67.562 ;
               RECT 25.814 68.726 25.866 68.762 ;
               RECT 25.814 69.926 25.866 69.962 ;
               RECT 25.814 71.126 25.866 71.162 ;
               RECT 25.814 72.326 25.866 72.362 ;
               RECT 25.814 73.526 25.866 73.562 ;
               RECT 25.814 74.726 25.866 74.762 ;
               RECT 25.814 75.926 25.866 75.962 ;
               RECT 25.814 77.126 25.866 77.162 ;
               RECT 25.814 78.326 25.866 78.362 ;
               RECT 25.814 79.526 25.866 79.562 ;
               RECT 25.814 80.726 25.866 80.762 ;
               RECT 25.814 81.926 25.866 81.962 ;
               RECT 25.814 83.126 25.866 83.162 ;
               RECT 25.814 84.326 25.866 84.362 ;
               RECT 25.814 85.526 25.866 85.562 ;
               RECT 25.814 86.726 25.866 86.762 ;
               RECT 25.814 87.926 25.866 87.962 ;
               RECT 25.814 89.126 25.866 89.162 ;
               RECT 25.814 90.326 25.866 90.362 ;
               RECT 25.814 91.526 25.866 91.562 ;
               RECT 25.814 92.726 25.866 92.762 ;
               RECT 25.814 93.926 25.866 93.962 ;
               RECT 25.814 95.126 25.866 95.162 ;
               RECT 25.814 96.326 25.866 96.362 ;
               RECT 25.814 97.526 25.866 97.562 ;
               RECT 25.814 98.726 25.866 98.762 ;
               RECT 25.814 99.926 25.866 99.962 ;
               RECT 25.814 101.126 25.866 101.162 ;
               RECT 25.814 102.326 25.866 102.362 ;
               RECT 25.814 103.526 25.866 103.562 ;
               RECT 25.894 1.558 25.946 1.594 ;
               RECT 25.894 2.758 25.946 2.794 ;
               RECT 25.894 3.958 25.946 3.994 ;
               RECT 25.894 5.158 25.946 5.194 ;
               RECT 25.894 6.358 25.946 6.394 ;
               RECT 25.894 7.558 25.946 7.594 ;
               RECT 25.894 8.758 25.946 8.794 ;
               RECT 25.894 9.958 25.946 9.994 ;
               RECT 25.894 11.158 25.946 11.194 ;
               RECT 25.894 12.358 25.946 12.394 ;
               RECT 25.894 13.558 25.946 13.594 ;
               RECT 25.894 14.758 25.946 14.794 ;
               RECT 25.894 15.958 25.946 15.994 ;
               RECT 25.894 17.158 25.946 17.194 ;
               RECT 25.894 18.358 25.946 18.394 ;
               RECT 25.894 19.558 25.946 19.594 ;
               RECT 25.894 20.758 25.946 20.794 ;
               RECT 25.894 21.958 25.946 21.994 ;
               RECT 25.894 23.158 25.946 23.194 ;
               RECT 25.894 24.358 25.946 24.394 ;
               RECT 25.894 25.558 25.946 25.594 ;
               RECT 25.894 26.758 25.946 26.794 ;
               RECT 25.894 27.958 25.946 27.994 ;
               RECT 25.894 29.158 25.946 29.194 ;
               RECT 25.894 30.358 25.946 30.394 ;
               RECT 25.894 31.558 25.946 31.594 ;
               RECT 25.894 32.758 25.946 32.794 ;
               RECT 25.894 33.958 25.946 33.994 ;
               RECT 25.894 35.158 25.946 35.194 ;
               RECT 25.894 36.358 25.946 36.394 ;
               RECT 25.894 37.558 25.946 37.594 ;
               RECT 25.894 38.758 25.946 38.794 ;
               RECT 25.894 39.958 25.946 39.994 ;
               RECT 25.894 41.158 25.946 41.194 ;
               RECT 25.894 42.358 25.946 42.394 ;
               RECT 25.894 43.558 25.946 43.594 ;
               RECT 25.894 44.758 25.946 44.794 ;
               RECT 25.894 45.958 25.946 45.994 ;
               RECT 25.894 47.158 25.946 47.194 ;
               RECT 25.894 48.358 25.946 48.394 ;
               RECT 25.894 50.142 25.946 50.178 ;
               RECT 25.894 50.382 25.946 50.418 ;
               RECT 25.894 54.702 25.946 54.738 ;
               RECT 25.894 54.942 25.946 54.978 ;
               RECT 25.894 57.478 25.946 57.514 ;
               RECT 25.894 58.678 25.946 58.714 ;
               RECT 25.894 59.878 25.946 59.914 ;
               RECT 25.894 61.078 25.946 61.114 ;
               RECT 25.894 62.278 25.946 62.314 ;
               RECT 25.894 63.478 25.946 63.514 ;
               RECT 25.894 64.678 25.946 64.714 ;
               RECT 25.894 65.878 25.946 65.914 ;
               RECT 25.894 67.078 25.946 67.114 ;
               RECT 25.894 68.278 25.946 68.314 ;
               RECT 25.894 69.478 25.946 69.514 ;
               RECT 25.894 70.678 25.946 70.714 ;
               RECT 25.894 71.878 25.946 71.914 ;
               RECT 25.894 73.078 25.946 73.114 ;
               RECT 25.894 74.278 25.946 74.314 ;
               RECT 25.894 75.478 25.946 75.514 ;
               RECT 25.894 76.678 25.946 76.714 ;
               RECT 25.894 77.878 25.946 77.914 ;
               RECT 25.894 79.078 25.946 79.114 ;
               RECT 25.894 80.278 25.946 80.314 ;
               RECT 25.894 81.478 25.946 81.514 ;
               RECT 25.894 82.678 25.946 82.714 ;
               RECT 25.894 83.878 25.946 83.914 ;
               RECT 25.894 85.078 25.946 85.114 ;
               RECT 25.894 86.278 25.946 86.314 ;
               RECT 25.894 87.478 25.946 87.514 ;
               RECT 25.894 88.678 25.946 88.714 ;
               RECT 25.894 89.878 25.946 89.914 ;
               RECT 25.894 91.078 25.946 91.114 ;
               RECT 25.894 92.278 25.946 92.314 ;
               RECT 25.894 93.478 25.946 93.514 ;
               RECT 25.894 94.678 25.946 94.714 ;
               RECT 25.894 95.878 25.946 95.914 ;
               RECT 25.894 97.078 25.946 97.114 ;
               RECT 25.894 98.278 25.946 98.314 ;
               RECT 25.894 99.478 25.946 99.514 ;
               RECT 25.894 100.678 25.946 100.714 ;
               RECT 25.894 101.878 25.946 101.914 ;
               RECT 25.894 103.078 25.946 103.114 ;
               RECT 25.894 104.278 25.946 104.314 ;
               RECT 25.974 0.281 26.026 0.317 ;
               RECT 25.974 104.803 26.026 104.839 ;
               RECT 26.054 0.806 26.106 0.842 ;
               RECT 26.054 2.006 26.106 2.042 ;
               RECT 26.054 3.206 26.106 3.242 ;
               RECT 26.054 4.406 26.106 4.442 ;
               RECT 26.054 5.606 26.106 5.642 ;
               RECT 26.054 6.806 26.106 6.842 ;
               RECT 26.054 8.006 26.106 8.042 ;
               RECT 26.054 9.206 26.106 9.242 ;
               RECT 26.054 10.406 26.106 10.442 ;
               RECT 26.054 11.606 26.106 11.642 ;
               RECT 26.054 12.806 26.106 12.842 ;
               RECT 26.054 14.006 26.106 14.042 ;
               RECT 26.054 15.206 26.106 15.242 ;
               RECT 26.054 16.406 26.106 16.442 ;
               RECT 26.054 17.606 26.106 17.642 ;
               RECT 26.054 18.806 26.106 18.842 ;
               RECT 26.054 20.006 26.106 20.042 ;
               RECT 26.054 21.206 26.106 21.242 ;
               RECT 26.054 22.406 26.106 22.442 ;
               RECT 26.054 23.606 26.106 23.642 ;
               RECT 26.054 24.806 26.106 24.842 ;
               RECT 26.054 26.006 26.106 26.042 ;
               RECT 26.054 27.206 26.106 27.242 ;
               RECT 26.054 28.406 26.106 28.442 ;
               RECT 26.054 29.606 26.106 29.642 ;
               RECT 26.054 30.806 26.106 30.842 ;
               RECT 26.054 32.006 26.106 32.042 ;
               RECT 26.054 33.206 26.106 33.242 ;
               RECT 26.054 34.406 26.106 34.442 ;
               RECT 26.054 35.606 26.106 35.642 ;
               RECT 26.054 36.806 26.106 36.842 ;
               RECT 26.054 38.006 26.106 38.042 ;
               RECT 26.054 39.206 26.106 39.242 ;
               RECT 26.054 40.406 26.106 40.442 ;
               RECT 26.054 41.606 26.106 41.642 ;
               RECT 26.054 42.806 26.106 42.842 ;
               RECT 26.054 44.006 26.106 44.042 ;
               RECT 26.054 45.206 26.106 45.242 ;
               RECT 26.054 46.406 26.106 46.442 ;
               RECT 26.054 47.606 26.106 47.642 ;
               RECT 26.054 49.422 26.106 49.458 ;
               RECT 26.054 49.662 26.106 49.698 ;
               RECT 26.054 55.422 26.106 55.458 ;
               RECT 26.054 55.662 26.106 55.698 ;
               RECT 26.054 56.726 26.106 56.762 ;
               RECT 26.054 57.926 26.106 57.962 ;
               RECT 26.054 59.126 26.106 59.162 ;
               RECT 26.054 60.326 26.106 60.362 ;
               RECT 26.054 61.526 26.106 61.562 ;
               RECT 26.054 62.726 26.106 62.762 ;
               RECT 26.054 63.926 26.106 63.962 ;
               RECT 26.054 65.126 26.106 65.162 ;
               RECT 26.054 66.326 26.106 66.362 ;
               RECT 26.054 67.526 26.106 67.562 ;
               RECT 26.054 68.726 26.106 68.762 ;
               RECT 26.054 69.926 26.106 69.962 ;
               RECT 26.054 71.126 26.106 71.162 ;
               RECT 26.054 72.326 26.106 72.362 ;
               RECT 26.054 73.526 26.106 73.562 ;
               RECT 26.054 74.726 26.106 74.762 ;
               RECT 26.054 75.926 26.106 75.962 ;
               RECT 26.054 77.126 26.106 77.162 ;
               RECT 26.054 78.326 26.106 78.362 ;
               RECT 26.054 79.526 26.106 79.562 ;
               RECT 26.054 80.726 26.106 80.762 ;
               RECT 26.054 81.926 26.106 81.962 ;
               RECT 26.054 83.126 26.106 83.162 ;
               RECT 26.054 84.326 26.106 84.362 ;
               RECT 26.054 85.526 26.106 85.562 ;
               RECT 26.054 86.726 26.106 86.762 ;
               RECT 26.054 87.926 26.106 87.962 ;
               RECT 26.054 89.126 26.106 89.162 ;
               RECT 26.054 90.326 26.106 90.362 ;
               RECT 26.054 91.526 26.106 91.562 ;
               RECT 26.054 92.726 26.106 92.762 ;
               RECT 26.054 93.926 26.106 93.962 ;
               RECT 26.054 95.126 26.106 95.162 ;
               RECT 26.054 96.326 26.106 96.362 ;
               RECT 26.054 97.526 26.106 97.562 ;
               RECT 26.054 98.726 26.106 98.762 ;
               RECT 26.054 99.926 26.106 99.962 ;
               RECT 26.054 101.126 26.106 101.162 ;
               RECT 26.054 102.326 26.106 102.362 ;
               RECT 26.054 103.526 26.106 103.562 ;
               RECT 26.134 1.558 26.186 1.594 ;
               RECT 26.134 2.758 26.186 2.794 ;
               RECT 26.134 3.958 26.186 3.994 ;
               RECT 26.134 5.158 26.186 5.194 ;
               RECT 26.134 6.358 26.186 6.394 ;
               RECT 26.134 7.558 26.186 7.594 ;
               RECT 26.134 8.758 26.186 8.794 ;
               RECT 26.134 9.958 26.186 9.994 ;
               RECT 26.134 11.158 26.186 11.194 ;
               RECT 26.134 12.358 26.186 12.394 ;
               RECT 26.134 13.558 26.186 13.594 ;
               RECT 26.134 14.758 26.186 14.794 ;
               RECT 26.134 15.958 26.186 15.994 ;
               RECT 26.134 17.158 26.186 17.194 ;
               RECT 26.134 18.358 26.186 18.394 ;
               RECT 26.134 19.558 26.186 19.594 ;
               RECT 26.134 20.758 26.186 20.794 ;
               RECT 26.134 21.958 26.186 21.994 ;
               RECT 26.134 23.158 26.186 23.194 ;
               RECT 26.134 24.358 26.186 24.394 ;
               RECT 26.134 25.558 26.186 25.594 ;
               RECT 26.134 26.758 26.186 26.794 ;
               RECT 26.134 27.958 26.186 27.994 ;
               RECT 26.134 29.158 26.186 29.194 ;
               RECT 26.134 30.358 26.186 30.394 ;
               RECT 26.134 31.558 26.186 31.594 ;
               RECT 26.134 32.758 26.186 32.794 ;
               RECT 26.134 33.958 26.186 33.994 ;
               RECT 26.134 35.158 26.186 35.194 ;
               RECT 26.134 36.358 26.186 36.394 ;
               RECT 26.134 37.558 26.186 37.594 ;
               RECT 26.134 38.758 26.186 38.794 ;
               RECT 26.134 39.958 26.186 39.994 ;
               RECT 26.134 41.158 26.186 41.194 ;
               RECT 26.134 42.358 26.186 42.394 ;
               RECT 26.134 43.558 26.186 43.594 ;
               RECT 26.134 44.758 26.186 44.794 ;
               RECT 26.134 45.958 26.186 45.994 ;
               RECT 26.134 47.158 26.186 47.194 ;
               RECT 26.134 48.358 26.186 48.394 ;
               RECT 26.134 50.142 26.186 50.178 ;
               RECT 26.134 50.382 26.186 50.418 ;
               RECT 26.134 54.702 26.186 54.738 ;
               RECT 26.134 54.942 26.186 54.978 ;
               RECT 26.134 57.478 26.186 57.514 ;
               RECT 26.134 58.678 26.186 58.714 ;
               RECT 26.134 59.878 26.186 59.914 ;
               RECT 26.134 61.078 26.186 61.114 ;
               RECT 26.134 62.278 26.186 62.314 ;
               RECT 26.134 63.478 26.186 63.514 ;
               RECT 26.134 64.678 26.186 64.714 ;
               RECT 26.134 65.878 26.186 65.914 ;
               RECT 26.134 67.078 26.186 67.114 ;
               RECT 26.134 68.278 26.186 68.314 ;
               RECT 26.134 69.478 26.186 69.514 ;
               RECT 26.134 70.678 26.186 70.714 ;
               RECT 26.134 71.878 26.186 71.914 ;
               RECT 26.134 73.078 26.186 73.114 ;
               RECT 26.134 74.278 26.186 74.314 ;
               RECT 26.134 75.478 26.186 75.514 ;
               RECT 26.134 76.678 26.186 76.714 ;
               RECT 26.134 77.878 26.186 77.914 ;
               RECT 26.134 79.078 26.186 79.114 ;
               RECT 26.134 80.278 26.186 80.314 ;
               RECT 26.134 81.478 26.186 81.514 ;
               RECT 26.134 82.678 26.186 82.714 ;
               RECT 26.134 83.878 26.186 83.914 ;
               RECT 26.134 85.078 26.186 85.114 ;
               RECT 26.134 86.278 26.186 86.314 ;
               RECT 26.134 87.478 26.186 87.514 ;
               RECT 26.134 88.678 26.186 88.714 ;
               RECT 26.134 89.878 26.186 89.914 ;
               RECT 26.134 91.078 26.186 91.114 ;
               RECT 26.134 92.278 26.186 92.314 ;
               RECT 26.134 93.478 26.186 93.514 ;
               RECT 26.134 94.678 26.186 94.714 ;
               RECT 26.134 95.878 26.186 95.914 ;
               RECT 26.134 97.078 26.186 97.114 ;
               RECT 26.134 98.278 26.186 98.314 ;
               RECT 26.134 99.478 26.186 99.514 ;
               RECT 26.134 100.678 26.186 100.714 ;
               RECT 26.134 101.878 26.186 101.914 ;
               RECT 26.134 103.078 26.186 103.114 ;
               RECT 26.134 104.278 26.186 104.314 ;
               RECT 26.214 0.806 26.266 0.842 ;
               RECT 26.214 2.006 26.266 2.042 ;
               RECT 26.214 3.206 26.266 3.242 ;
               RECT 26.214 4.406 26.266 4.442 ;
               RECT 26.214 5.606 26.266 5.642 ;
               RECT 26.214 6.806 26.266 6.842 ;
               RECT 26.214 8.006 26.266 8.042 ;
               RECT 26.214 9.206 26.266 9.242 ;
               RECT 26.214 10.406 26.266 10.442 ;
               RECT 26.214 11.606 26.266 11.642 ;
               RECT 26.214 12.806 26.266 12.842 ;
               RECT 26.214 14.006 26.266 14.042 ;
               RECT 26.214 15.206 26.266 15.242 ;
               RECT 26.214 16.406 26.266 16.442 ;
               RECT 26.214 17.606 26.266 17.642 ;
               RECT 26.214 18.806 26.266 18.842 ;
               RECT 26.214 20.006 26.266 20.042 ;
               RECT 26.214 21.206 26.266 21.242 ;
               RECT 26.214 22.406 26.266 22.442 ;
               RECT 26.214 23.606 26.266 23.642 ;
               RECT 26.214 24.806 26.266 24.842 ;
               RECT 26.214 26.006 26.266 26.042 ;
               RECT 26.214 27.206 26.266 27.242 ;
               RECT 26.214 28.406 26.266 28.442 ;
               RECT 26.214 29.606 26.266 29.642 ;
               RECT 26.214 30.806 26.266 30.842 ;
               RECT 26.214 32.006 26.266 32.042 ;
               RECT 26.214 33.206 26.266 33.242 ;
               RECT 26.214 34.406 26.266 34.442 ;
               RECT 26.214 35.606 26.266 35.642 ;
               RECT 26.214 36.806 26.266 36.842 ;
               RECT 26.214 38.006 26.266 38.042 ;
               RECT 26.214 39.206 26.266 39.242 ;
               RECT 26.214 40.406 26.266 40.442 ;
               RECT 26.214 41.606 26.266 41.642 ;
               RECT 26.214 42.806 26.266 42.842 ;
               RECT 26.214 44.006 26.266 44.042 ;
               RECT 26.214 45.206 26.266 45.242 ;
               RECT 26.214 46.406 26.266 46.442 ;
               RECT 26.214 47.606 26.266 47.642 ;
               RECT 26.214 49.422 26.266 49.458 ;
               RECT 26.214 49.662 26.266 49.698 ;
               RECT 26.214 55.422 26.266 55.458 ;
               RECT 26.214 55.662 26.266 55.698 ;
               RECT 26.214 56.726 26.266 56.762 ;
               RECT 26.214 57.926 26.266 57.962 ;
               RECT 26.214 59.126 26.266 59.162 ;
               RECT 26.214 60.326 26.266 60.362 ;
               RECT 26.214 61.526 26.266 61.562 ;
               RECT 26.214 62.726 26.266 62.762 ;
               RECT 26.214 63.926 26.266 63.962 ;
               RECT 26.214 65.126 26.266 65.162 ;
               RECT 26.214 66.326 26.266 66.362 ;
               RECT 26.214 67.526 26.266 67.562 ;
               RECT 26.214 68.726 26.266 68.762 ;
               RECT 26.214 69.926 26.266 69.962 ;
               RECT 26.214 71.126 26.266 71.162 ;
               RECT 26.214 72.326 26.266 72.362 ;
               RECT 26.214 73.526 26.266 73.562 ;
               RECT 26.214 74.726 26.266 74.762 ;
               RECT 26.214 75.926 26.266 75.962 ;
               RECT 26.214 77.126 26.266 77.162 ;
               RECT 26.214 78.326 26.266 78.362 ;
               RECT 26.214 79.526 26.266 79.562 ;
               RECT 26.214 80.726 26.266 80.762 ;
               RECT 26.214 81.926 26.266 81.962 ;
               RECT 26.214 83.126 26.266 83.162 ;
               RECT 26.214 84.326 26.266 84.362 ;
               RECT 26.214 85.526 26.266 85.562 ;
               RECT 26.214 86.726 26.266 86.762 ;
               RECT 26.214 87.926 26.266 87.962 ;
               RECT 26.214 89.126 26.266 89.162 ;
               RECT 26.214 90.326 26.266 90.362 ;
               RECT 26.214 91.526 26.266 91.562 ;
               RECT 26.214 92.726 26.266 92.762 ;
               RECT 26.214 93.926 26.266 93.962 ;
               RECT 26.214 95.126 26.266 95.162 ;
               RECT 26.214 96.326 26.266 96.362 ;
               RECT 26.214 97.526 26.266 97.562 ;
               RECT 26.214 98.726 26.266 98.762 ;
               RECT 26.214 99.926 26.266 99.962 ;
               RECT 26.214 101.126 26.266 101.162 ;
               RECT 26.214 102.326 26.266 102.362 ;
               RECT 26.214 103.526 26.266 103.562 ;
               RECT 26.294 1.558 26.346 1.594 ;
               RECT 26.294 2.758 26.346 2.794 ;
               RECT 26.294 3.958 26.346 3.994 ;
               RECT 26.294 5.158 26.346 5.194 ;
               RECT 26.294 6.358 26.346 6.394 ;
               RECT 26.294 7.558 26.346 7.594 ;
               RECT 26.294 8.758 26.346 8.794 ;
               RECT 26.294 9.958 26.346 9.994 ;
               RECT 26.294 11.158 26.346 11.194 ;
               RECT 26.294 12.358 26.346 12.394 ;
               RECT 26.294 13.558 26.346 13.594 ;
               RECT 26.294 14.758 26.346 14.794 ;
               RECT 26.294 15.958 26.346 15.994 ;
               RECT 26.294 17.158 26.346 17.194 ;
               RECT 26.294 18.358 26.346 18.394 ;
               RECT 26.294 19.558 26.346 19.594 ;
               RECT 26.294 20.758 26.346 20.794 ;
               RECT 26.294 21.958 26.346 21.994 ;
               RECT 26.294 23.158 26.346 23.194 ;
               RECT 26.294 24.358 26.346 24.394 ;
               RECT 26.294 25.558 26.346 25.594 ;
               RECT 26.294 26.758 26.346 26.794 ;
               RECT 26.294 27.958 26.346 27.994 ;
               RECT 26.294 29.158 26.346 29.194 ;
               RECT 26.294 30.358 26.346 30.394 ;
               RECT 26.294 31.558 26.346 31.594 ;
               RECT 26.294 32.758 26.346 32.794 ;
               RECT 26.294 33.958 26.346 33.994 ;
               RECT 26.294 35.158 26.346 35.194 ;
               RECT 26.294 36.358 26.346 36.394 ;
               RECT 26.294 37.558 26.346 37.594 ;
               RECT 26.294 38.758 26.346 38.794 ;
               RECT 26.294 39.958 26.346 39.994 ;
               RECT 26.294 41.158 26.346 41.194 ;
               RECT 26.294 42.358 26.346 42.394 ;
               RECT 26.294 43.558 26.346 43.594 ;
               RECT 26.294 44.758 26.346 44.794 ;
               RECT 26.294 45.958 26.346 45.994 ;
               RECT 26.294 47.158 26.346 47.194 ;
               RECT 26.294 48.358 26.346 48.394 ;
               RECT 26.294 50.142 26.346 50.178 ;
               RECT 26.294 50.382 26.346 50.418 ;
               RECT 26.294 54.702 26.346 54.738 ;
               RECT 26.294 54.942 26.346 54.978 ;
               RECT 26.294 57.478 26.346 57.514 ;
               RECT 26.294 58.678 26.346 58.714 ;
               RECT 26.294 59.878 26.346 59.914 ;
               RECT 26.294 61.078 26.346 61.114 ;
               RECT 26.294 62.278 26.346 62.314 ;
               RECT 26.294 63.478 26.346 63.514 ;
               RECT 26.294 64.678 26.346 64.714 ;
               RECT 26.294 65.878 26.346 65.914 ;
               RECT 26.294 67.078 26.346 67.114 ;
               RECT 26.294 68.278 26.346 68.314 ;
               RECT 26.294 69.478 26.346 69.514 ;
               RECT 26.294 70.678 26.346 70.714 ;
               RECT 26.294 71.878 26.346 71.914 ;
               RECT 26.294 73.078 26.346 73.114 ;
               RECT 26.294 74.278 26.346 74.314 ;
               RECT 26.294 75.478 26.346 75.514 ;
               RECT 26.294 76.678 26.346 76.714 ;
               RECT 26.294 77.878 26.346 77.914 ;
               RECT 26.294 79.078 26.346 79.114 ;
               RECT 26.294 80.278 26.346 80.314 ;
               RECT 26.294 81.478 26.346 81.514 ;
               RECT 26.294 82.678 26.346 82.714 ;
               RECT 26.294 83.878 26.346 83.914 ;
               RECT 26.294 85.078 26.346 85.114 ;
               RECT 26.294 86.278 26.346 86.314 ;
               RECT 26.294 87.478 26.346 87.514 ;
               RECT 26.294 88.678 26.346 88.714 ;
               RECT 26.294 89.878 26.346 89.914 ;
               RECT 26.294 91.078 26.346 91.114 ;
               RECT 26.294 92.278 26.346 92.314 ;
               RECT 26.294 93.478 26.346 93.514 ;
               RECT 26.294 94.678 26.346 94.714 ;
               RECT 26.294 95.878 26.346 95.914 ;
               RECT 26.294 97.078 26.346 97.114 ;
               RECT 26.294 98.278 26.346 98.314 ;
               RECT 26.294 99.478 26.346 99.514 ;
               RECT 26.294 100.678 26.346 100.714 ;
               RECT 26.294 101.878 26.346 101.914 ;
               RECT 26.294 103.078 26.346 103.114 ;
               RECT 26.294 104.278 26.346 104.314 ;
               RECT 26.374 0.281 26.426 0.317 ;
               RECT 26.374 104.803 26.426 104.839 ;
               RECT 26.454 0.806 26.506 0.842 ;
               RECT 26.454 2.006 26.506 2.042 ;
               RECT 26.454 3.206 26.506 3.242 ;
               RECT 26.454 4.406 26.506 4.442 ;
               RECT 26.454 5.606 26.506 5.642 ;
               RECT 26.454 6.806 26.506 6.842 ;
               RECT 26.454 8.006 26.506 8.042 ;
               RECT 26.454 9.206 26.506 9.242 ;
               RECT 26.454 10.406 26.506 10.442 ;
               RECT 26.454 11.606 26.506 11.642 ;
               RECT 26.454 12.806 26.506 12.842 ;
               RECT 26.454 14.006 26.506 14.042 ;
               RECT 26.454 15.206 26.506 15.242 ;
               RECT 26.454 16.406 26.506 16.442 ;
               RECT 26.454 17.606 26.506 17.642 ;
               RECT 26.454 18.806 26.506 18.842 ;
               RECT 26.454 20.006 26.506 20.042 ;
               RECT 26.454 21.206 26.506 21.242 ;
               RECT 26.454 22.406 26.506 22.442 ;
               RECT 26.454 23.606 26.506 23.642 ;
               RECT 26.454 24.806 26.506 24.842 ;
               RECT 26.454 26.006 26.506 26.042 ;
               RECT 26.454 27.206 26.506 27.242 ;
               RECT 26.454 28.406 26.506 28.442 ;
               RECT 26.454 29.606 26.506 29.642 ;
               RECT 26.454 30.806 26.506 30.842 ;
               RECT 26.454 32.006 26.506 32.042 ;
               RECT 26.454 33.206 26.506 33.242 ;
               RECT 26.454 34.406 26.506 34.442 ;
               RECT 26.454 35.606 26.506 35.642 ;
               RECT 26.454 36.806 26.506 36.842 ;
               RECT 26.454 38.006 26.506 38.042 ;
               RECT 26.454 39.206 26.506 39.242 ;
               RECT 26.454 40.406 26.506 40.442 ;
               RECT 26.454 41.606 26.506 41.642 ;
               RECT 26.454 42.806 26.506 42.842 ;
               RECT 26.454 44.006 26.506 44.042 ;
               RECT 26.454 45.206 26.506 45.242 ;
               RECT 26.454 46.406 26.506 46.442 ;
               RECT 26.454 47.606 26.506 47.642 ;
               RECT 26.454 49.422 26.506 49.458 ;
               RECT 26.454 49.662 26.506 49.698 ;
               RECT 26.454 51.102 26.506 51.138 ;
               RECT 26.454 51.582 26.506 51.618 ;
               RECT 26.454 53.502 26.506 53.538 ;
               RECT 26.454 53.982 26.506 54.018 ;
               RECT 26.454 55.422 26.506 55.458 ;
               RECT 26.454 55.662 26.506 55.698 ;
               RECT 26.454 56.726 26.506 56.762 ;
               RECT 26.454 57.926 26.506 57.962 ;
               RECT 26.454 59.126 26.506 59.162 ;
               RECT 26.454 60.326 26.506 60.362 ;
               RECT 26.454 61.526 26.506 61.562 ;
               RECT 26.454 62.726 26.506 62.762 ;
               RECT 26.454 63.926 26.506 63.962 ;
               RECT 26.454 65.126 26.506 65.162 ;
               RECT 26.454 66.326 26.506 66.362 ;
               RECT 26.454 67.526 26.506 67.562 ;
               RECT 26.454 68.726 26.506 68.762 ;
               RECT 26.454 69.926 26.506 69.962 ;
               RECT 26.454 71.126 26.506 71.162 ;
               RECT 26.454 72.326 26.506 72.362 ;
               RECT 26.454 73.526 26.506 73.562 ;
               RECT 26.454 74.726 26.506 74.762 ;
               RECT 26.454 75.926 26.506 75.962 ;
               RECT 26.454 77.126 26.506 77.162 ;
               RECT 26.454 78.326 26.506 78.362 ;
               RECT 26.454 79.526 26.506 79.562 ;
               RECT 26.454 80.726 26.506 80.762 ;
               RECT 26.454 81.926 26.506 81.962 ;
               RECT 26.454 83.126 26.506 83.162 ;
               RECT 26.454 84.326 26.506 84.362 ;
               RECT 26.454 85.526 26.506 85.562 ;
               RECT 26.454 86.726 26.506 86.762 ;
               RECT 26.454 87.926 26.506 87.962 ;
               RECT 26.454 89.126 26.506 89.162 ;
               RECT 26.454 90.326 26.506 90.362 ;
               RECT 26.454 91.526 26.506 91.562 ;
               RECT 26.454 92.726 26.506 92.762 ;
               RECT 26.454 93.926 26.506 93.962 ;
               RECT 26.454 95.126 26.506 95.162 ;
               RECT 26.454 96.326 26.506 96.362 ;
               RECT 26.454 97.526 26.506 97.562 ;
               RECT 26.454 98.726 26.506 98.762 ;
               RECT 26.454 99.926 26.506 99.962 ;
               RECT 26.454 101.126 26.506 101.162 ;
               RECT 26.454 102.326 26.506 102.362 ;
               RECT 26.454 103.526 26.506 103.562 ;
               RECT 26.534 1.558 26.586 1.594 ;
               RECT 26.534 2.758 26.586 2.794 ;
               RECT 26.534 3.958 26.586 3.994 ;
               RECT 26.534 5.158 26.586 5.194 ;
               RECT 26.534 6.358 26.586 6.394 ;
               RECT 26.534 7.558 26.586 7.594 ;
               RECT 26.534 8.758 26.586 8.794 ;
               RECT 26.534 9.958 26.586 9.994 ;
               RECT 26.534 11.158 26.586 11.194 ;
               RECT 26.534 12.358 26.586 12.394 ;
               RECT 26.534 13.558 26.586 13.594 ;
               RECT 26.534 14.758 26.586 14.794 ;
               RECT 26.534 15.958 26.586 15.994 ;
               RECT 26.534 17.158 26.586 17.194 ;
               RECT 26.534 18.358 26.586 18.394 ;
               RECT 26.534 19.558 26.586 19.594 ;
               RECT 26.534 20.758 26.586 20.794 ;
               RECT 26.534 21.958 26.586 21.994 ;
               RECT 26.534 23.158 26.586 23.194 ;
               RECT 26.534 24.358 26.586 24.394 ;
               RECT 26.534 25.558 26.586 25.594 ;
               RECT 26.534 26.758 26.586 26.794 ;
               RECT 26.534 27.958 26.586 27.994 ;
               RECT 26.534 29.158 26.586 29.194 ;
               RECT 26.534 30.358 26.586 30.394 ;
               RECT 26.534 31.558 26.586 31.594 ;
               RECT 26.534 32.758 26.586 32.794 ;
               RECT 26.534 33.958 26.586 33.994 ;
               RECT 26.534 35.158 26.586 35.194 ;
               RECT 26.534 36.358 26.586 36.394 ;
               RECT 26.534 37.558 26.586 37.594 ;
               RECT 26.534 38.758 26.586 38.794 ;
               RECT 26.534 39.958 26.586 39.994 ;
               RECT 26.534 41.158 26.586 41.194 ;
               RECT 26.534 42.358 26.586 42.394 ;
               RECT 26.534 43.558 26.586 43.594 ;
               RECT 26.534 44.758 26.586 44.794 ;
               RECT 26.534 45.958 26.586 45.994 ;
               RECT 26.534 47.158 26.586 47.194 ;
               RECT 26.534 48.358 26.586 48.394 ;
               RECT 26.534 50.142 26.586 50.178 ;
               RECT 26.534 50.382 26.586 50.418 ;
               RECT 26.534 54.702 26.586 54.738 ;
               RECT 26.534 54.942 26.586 54.978 ;
               RECT 26.534 57.478 26.586 57.514 ;
               RECT 26.534 58.678 26.586 58.714 ;
               RECT 26.534 59.878 26.586 59.914 ;
               RECT 26.534 61.078 26.586 61.114 ;
               RECT 26.534 62.278 26.586 62.314 ;
               RECT 26.534 63.478 26.586 63.514 ;
               RECT 26.534 64.678 26.586 64.714 ;
               RECT 26.534 65.878 26.586 65.914 ;
               RECT 26.534 67.078 26.586 67.114 ;
               RECT 26.534 68.278 26.586 68.314 ;
               RECT 26.534 69.478 26.586 69.514 ;
               RECT 26.534 70.678 26.586 70.714 ;
               RECT 26.534 71.878 26.586 71.914 ;
               RECT 26.534 73.078 26.586 73.114 ;
               RECT 26.534 74.278 26.586 74.314 ;
               RECT 26.534 75.478 26.586 75.514 ;
               RECT 26.534 76.678 26.586 76.714 ;
               RECT 26.534 77.878 26.586 77.914 ;
               RECT 26.534 79.078 26.586 79.114 ;
               RECT 26.534 80.278 26.586 80.314 ;
               RECT 26.534 81.478 26.586 81.514 ;
               RECT 26.534 82.678 26.586 82.714 ;
               RECT 26.534 83.878 26.586 83.914 ;
               RECT 26.534 85.078 26.586 85.114 ;
               RECT 26.534 86.278 26.586 86.314 ;
               RECT 26.534 87.478 26.586 87.514 ;
               RECT 26.534 88.678 26.586 88.714 ;
               RECT 26.534 89.878 26.586 89.914 ;
               RECT 26.534 91.078 26.586 91.114 ;
               RECT 26.534 92.278 26.586 92.314 ;
               RECT 26.534 93.478 26.586 93.514 ;
               RECT 26.534 94.678 26.586 94.714 ;
               RECT 26.534 95.878 26.586 95.914 ;
               RECT 26.534 97.078 26.586 97.114 ;
               RECT 26.534 98.278 26.586 98.314 ;
               RECT 26.534 99.478 26.586 99.514 ;
               RECT 26.534 100.678 26.586 100.714 ;
               RECT 26.534 101.878 26.586 101.914 ;
               RECT 26.534 103.078 26.586 103.114 ;
               RECT 26.534 104.278 26.586 104.314 ;
               RECT 26.614 0.806 26.666 0.842 ;
               RECT 26.614 2.006 26.666 2.042 ;
               RECT 26.614 3.206 26.666 3.242 ;
               RECT 26.614 4.406 26.666 4.442 ;
               RECT 26.614 5.606 26.666 5.642 ;
               RECT 26.614 6.806 26.666 6.842 ;
               RECT 26.614 8.006 26.666 8.042 ;
               RECT 26.614 9.206 26.666 9.242 ;
               RECT 26.614 10.406 26.666 10.442 ;
               RECT 26.614 11.606 26.666 11.642 ;
               RECT 26.614 12.806 26.666 12.842 ;
               RECT 26.614 14.006 26.666 14.042 ;
               RECT 26.614 15.206 26.666 15.242 ;
               RECT 26.614 16.406 26.666 16.442 ;
               RECT 26.614 17.606 26.666 17.642 ;
               RECT 26.614 18.806 26.666 18.842 ;
               RECT 26.614 20.006 26.666 20.042 ;
               RECT 26.614 21.206 26.666 21.242 ;
               RECT 26.614 22.406 26.666 22.442 ;
               RECT 26.614 23.606 26.666 23.642 ;
               RECT 26.614 24.806 26.666 24.842 ;
               RECT 26.614 26.006 26.666 26.042 ;
               RECT 26.614 27.206 26.666 27.242 ;
               RECT 26.614 28.406 26.666 28.442 ;
               RECT 26.614 29.606 26.666 29.642 ;
               RECT 26.614 30.806 26.666 30.842 ;
               RECT 26.614 32.006 26.666 32.042 ;
               RECT 26.614 33.206 26.666 33.242 ;
               RECT 26.614 34.406 26.666 34.442 ;
               RECT 26.614 35.606 26.666 35.642 ;
               RECT 26.614 36.806 26.666 36.842 ;
               RECT 26.614 38.006 26.666 38.042 ;
               RECT 26.614 39.206 26.666 39.242 ;
               RECT 26.614 40.406 26.666 40.442 ;
               RECT 26.614 41.606 26.666 41.642 ;
               RECT 26.614 42.806 26.666 42.842 ;
               RECT 26.614 44.006 26.666 44.042 ;
               RECT 26.614 45.206 26.666 45.242 ;
               RECT 26.614 46.406 26.666 46.442 ;
               RECT 26.614 47.606 26.666 47.642 ;
               RECT 26.614 49.422 26.666 49.458 ;
               RECT 26.614 49.662 26.666 49.698 ;
               RECT 26.614 55.422 26.666 55.458 ;
               RECT 26.614 55.662 26.666 55.698 ;
               RECT 26.614 56.726 26.666 56.762 ;
               RECT 26.614 57.926 26.666 57.962 ;
               RECT 26.614 59.126 26.666 59.162 ;
               RECT 26.614 60.326 26.666 60.362 ;
               RECT 26.614 61.526 26.666 61.562 ;
               RECT 26.614 62.726 26.666 62.762 ;
               RECT 26.614 63.926 26.666 63.962 ;
               RECT 26.614 65.126 26.666 65.162 ;
               RECT 26.614 66.326 26.666 66.362 ;
               RECT 26.614 67.526 26.666 67.562 ;
               RECT 26.614 68.726 26.666 68.762 ;
               RECT 26.614 69.926 26.666 69.962 ;
               RECT 26.614 71.126 26.666 71.162 ;
               RECT 26.614 72.326 26.666 72.362 ;
               RECT 26.614 73.526 26.666 73.562 ;
               RECT 26.614 74.726 26.666 74.762 ;
               RECT 26.614 75.926 26.666 75.962 ;
               RECT 26.614 77.126 26.666 77.162 ;
               RECT 26.614 78.326 26.666 78.362 ;
               RECT 26.614 79.526 26.666 79.562 ;
               RECT 26.614 80.726 26.666 80.762 ;
               RECT 26.614 81.926 26.666 81.962 ;
               RECT 26.614 83.126 26.666 83.162 ;
               RECT 26.614 84.326 26.666 84.362 ;
               RECT 26.614 85.526 26.666 85.562 ;
               RECT 26.614 86.726 26.666 86.762 ;
               RECT 26.614 87.926 26.666 87.962 ;
               RECT 26.614 89.126 26.666 89.162 ;
               RECT 26.614 90.326 26.666 90.362 ;
               RECT 26.614 91.526 26.666 91.562 ;
               RECT 26.614 92.726 26.666 92.762 ;
               RECT 26.614 93.926 26.666 93.962 ;
               RECT 26.614 95.126 26.666 95.162 ;
               RECT 26.614 96.326 26.666 96.362 ;
               RECT 26.614 97.526 26.666 97.562 ;
               RECT 26.614 98.726 26.666 98.762 ;
               RECT 26.614 99.926 26.666 99.962 ;
               RECT 26.614 101.126 26.666 101.162 ;
               RECT 26.614 102.326 26.666 102.362 ;
               RECT 26.614 103.526 26.666 103.562 ;
               RECT 26.694 1.558 26.746 1.594 ;
               RECT 26.694 2.758 26.746 2.794 ;
               RECT 26.694 3.958 26.746 3.994 ;
               RECT 26.694 5.158 26.746 5.194 ;
               RECT 26.694 6.358 26.746 6.394 ;
               RECT 26.694 7.558 26.746 7.594 ;
               RECT 26.694 8.758 26.746 8.794 ;
               RECT 26.694 9.958 26.746 9.994 ;
               RECT 26.694 11.158 26.746 11.194 ;
               RECT 26.694 12.358 26.746 12.394 ;
               RECT 26.694 13.558 26.746 13.594 ;
               RECT 26.694 14.758 26.746 14.794 ;
               RECT 26.694 15.958 26.746 15.994 ;
               RECT 26.694 17.158 26.746 17.194 ;
               RECT 26.694 18.358 26.746 18.394 ;
               RECT 26.694 19.558 26.746 19.594 ;
               RECT 26.694 20.758 26.746 20.794 ;
               RECT 26.694 21.958 26.746 21.994 ;
               RECT 26.694 23.158 26.746 23.194 ;
               RECT 26.694 24.358 26.746 24.394 ;
               RECT 26.694 25.558 26.746 25.594 ;
               RECT 26.694 26.758 26.746 26.794 ;
               RECT 26.694 27.958 26.746 27.994 ;
               RECT 26.694 29.158 26.746 29.194 ;
               RECT 26.694 30.358 26.746 30.394 ;
               RECT 26.694 31.558 26.746 31.594 ;
               RECT 26.694 32.758 26.746 32.794 ;
               RECT 26.694 33.958 26.746 33.994 ;
               RECT 26.694 35.158 26.746 35.194 ;
               RECT 26.694 36.358 26.746 36.394 ;
               RECT 26.694 37.558 26.746 37.594 ;
               RECT 26.694 38.758 26.746 38.794 ;
               RECT 26.694 39.958 26.746 39.994 ;
               RECT 26.694 41.158 26.746 41.194 ;
               RECT 26.694 42.358 26.746 42.394 ;
               RECT 26.694 43.558 26.746 43.594 ;
               RECT 26.694 44.758 26.746 44.794 ;
               RECT 26.694 45.958 26.746 45.994 ;
               RECT 26.694 47.158 26.746 47.194 ;
               RECT 26.694 48.358 26.746 48.394 ;
               RECT 26.694 50.142 26.746 50.178 ;
               RECT 26.694 50.382 26.746 50.418 ;
               RECT 26.694 54.702 26.746 54.738 ;
               RECT 26.694 54.942 26.746 54.978 ;
               RECT 26.694 57.478 26.746 57.514 ;
               RECT 26.694 58.678 26.746 58.714 ;
               RECT 26.694 59.878 26.746 59.914 ;
               RECT 26.694 61.078 26.746 61.114 ;
               RECT 26.694 62.278 26.746 62.314 ;
               RECT 26.694 63.478 26.746 63.514 ;
               RECT 26.694 64.678 26.746 64.714 ;
               RECT 26.694 65.878 26.746 65.914 ;
               RECT 26.694 67.078 26.746 67.114 ;
               RECT 26.694 68.278 26.746 68.314 ;
               RECT 26.694 69.478 26.746 69.514 ;
               RECT 26.694 70.678 26.746 70.714 ;
               RECT 26.694 71.878 26.746 71.914 ;
               RECT 26.694 73.078 26.746 73.114 ;
               RECT 26.694 74.278 26.746 74.314 ;
               RECT 26.694 75.478 26.746 75.514 ;
               RECT 26.694 76.678 26.746 76.714 ;
               RECT 26.694 77.878 26.746 77.914 ;
               RECT 26.694 79.078 26.746 79.114 ;
               RECT 26.694 80.278 26.746 80.314 ;
               RECT 26.694 81.478 26.746 81.514 ;
               RECT 26.694 82.678 26.746 82.714 ;
               RECT 26.694 83.878 26.746 83.914 ;
               RECT 26.694 85.078 26.746 85.114 ;
               RECT 26.694 86.278 26.746 86.314 ;
               RECT 26.694 87.478 26.746 87.514 ;
               RECT 26.694 88.678 26.746 88.714 ;
               RECT 26.694 89.878 26.746 89.914 ;
               RECT 26.694 91.078 26.746 91.114 ;
               RECT 26.694 92.278 26.746 92.314 ;
               RECT 26.694 93.478 26.746 93.514 ;
               RECT 26.694 94.678 26.746 94.714 ;
               RECT 26.694 95.878 26.746 95.914 ;
               RECT 26.694 97.078 26.746 97.114 ;
               RECT 26.694 98.278 26.746 98.314 ;
               RECT 26.694 99.478 26.746 99.514 ;
               RECT 26.694 100.678 26.746 100.714 ;
               RECT 26.694 101.878 26.746 101.914 ;
               RECT 26.694 103.078 26.746 103.114 ;
               RECT 26.694 104.278 26.746 104.314 ;
               RECT 26.774 0.281 26.826 0.317 ;
               RECT 26.774 104.803 26.826 104.839 ;
               RECT 26.854 0.806 26.906 0.842 ;
               RECT 26.854 2.006 26.906 2.042 ;
               RECT 26.854 3.206 26.906 3.242 ;
               RECT 26.854 4.406 26.906 4.442 ;
               RECT 26.854 5.606 26.906 5.642 ;
               RECT 26.854 6.806 26.906 6.842 ;
               RECT 26.854 8.006 26.906 8.042 ;
               RECT 26.854 9.206 26.906 9.242 ;
               RECT 26.854 10.406 26.906 10.442 ;
               RECT 26.854 11.606 26.906 11.642 ;
               RECT 26.854 12.806 26.906 12.842 ;
               RECT 26.854 14.006 26.906 14.042 ;
               RECT 26.854 15.206 26.906 15.242 ;
               RECT 26.854 16.406 26.906 16.442 ;
               RECT 26.854 17.606 26.906 17.642 ;
               RECT 26.854 18.806 26.906 18.842 ;
               RECT 26.854 20.006 26.906 20.042 ;
               RECT 26.854 21.206 26.906 21.242 ;
               RECT 26.854 22.406 26.906 22.442 ;
               RECT 26.854 23.606 26.906 23.642 ;
               RECT 26.854 24.806 26.906 24.842 ;
               RECT 26.854 26.006 26.906 26.042 ;
               RECT 26.854 27.206 26.906 27.242 ;
               RECT 26.854 28.406 26.906 28.442 ;
               RECT 26.854 29.606 26.906 29.642 ;
               RECT 26.854 30.806 26.906 30.842 ;
               RECT 26.854 32.006 26.906 32.042 ;
               RECT 26.854 33.206 26.906 33.242 ;
               RECT 26.854 34.406 26.906 34.442 ;
               RECT 26.854 35.606 26.906 35.642 ;
               RECT 26.854 36.806 26.906 36.842 ;
               RECT 26.854 38.006 26.906 38.042 ;
               RECT 26.854 39.206 26.906 39.242 ;
               RECT 26.854 40.406 26.906 40.442 ;
               RECT 26.854 41.606 26.906 41.642 ;
               RECT 26.854 42.806 26.906 42.842 ;
               RECT 26.854 44.006 26.906 44.042 ;
               RECT 26.854 45.206 26.906 45.242 ;
               RECT 26.854 46.406 26.906 46.442 ;
               RECT 26.854 47.606 26.906 47.642 ;
               RECT 26.854 49.422 26.906 49.458 ;
               RECT 26.854 49.662 26.906 49.698 ;
               RECT 26.854 55.422 26.906 55.458 ;
               RECT 26.854 55.662 26.906 55.698 ;
               RECT 26.854 56.726 26.906 56.762 ;
               RECT 26.854 57.926 26.906 57.962 ;
               RECT 26.854 59.126 26.906 59.162 ;
               RECT 26.854 60.326 26.906 60.362 ;
               RECT 26.854 61.526 26.906 61.562 ;
               RECT 26.854 62.726 26.906 62.762 ;
               RECT 26.854 63.926 26.906 63.962 ;
               RECT 26.854 65.126 26.906 65.162 ;
               RECT 26.854 66.326 26.906 66.362 ;
               RECT 26.854 67.526 26.906 67.562 ;
               RECT 26.854 68.726 26.906 68.762 ;
               RECT 26.854 69.926 26.906 69.962 ;
               RECT 26.854 71.126 26.906 71.162 ;
               RECT 26.854 72.326 26.906 72.362 ;
               RECT 26.854 73.526 26.906 73.562 ;
               RECT 26.854 74.726 26.906 74.762 ;
               RECT 26.854 75.926 26.906 75.962 ;
               RECT 26.854 77.126 26.906 77.162 ;
               RECT 26.854 78.326 26.906 78.362 ;
               RECT 26.854 79.526 26.906 79.562 ;
               RECT 26.854 80.726 26.906 80.762 ;
               RECT 26.854 81.926 26.906 81.962 ;
               RECT 26.854 83.126 26.906 83.162 ;
               RECT 26.854 84.326 26.906 84.362 ;
               RECT 26.854 85.526 26.906 85.562 ;
               RECT 26.854 86.726 26.906 86.762 ;
               RECT 26.854 87.926 26.906 87.962 ;
               RECT 26.854 89.126 26.906 89.162 ;
               RECT 26.854 90.326 26.906 90.362 ;
               RECT 26.854 91.526 26.906 91.562 ;
               RECT 26.854 92.726 26.906 92.762 ;
               RECT 26.854 93.926 26.906 93.962 ;
               RECT 26.854 95.126 26.906 95.162 ;
               RECT 26.854 96.326 26.906 96.362 ;
               RECT 26.854 97.526 26.906 97.562 ;
               RECT 26.854 98.726 26.906 98.762 ;
               RECT 26.854 99.926 26.906 99.962 ;
               RECT 26.854 101.126 26.906 101.162 ;
               RECT 26.854 102.326 26.906 102.362 ;
               RECT 26.854 103.526 26.906 103.562 ;
               RECT 26.934 1.558 26.986 1.594 ;
               RECT 26.934 2.758 26.986 2.794 ;
               RECT 26.934 3.958 26.986 3.994 ;
               RECT 26.934 5.158 26.986 5.194 ;
               RECT 26.934 6.358 26.986 6.394 ;
               RECT 26.934 7.558 26.986 7.594 ;
               RECT 26.934 8.758 26.986 8.794 ;
               RECT 26.934 9.958 26.986 9.994 ;
               RECT 26.934 11.158 26.986 11.194 ;
               RECT 26.934 12.358 26.986 12.394 ;
               RECT 26.934 13.558 26.986 13.594 ;
               RECT 26.934 14.758 26.986 14.794 ;
               RECT 26.934 15.958 26.986 15.994 ;
               RECT 26.934 17.158 26.986 17.194 ;
               RECT 26.934 18.358 26.986 18.394 ;
               RECT 26.934 19.558 26.986 19.594 ;
               RECT 26.934 20.758 26.986 20.794 ;
               RECT 26.934 21.958 26.986 21.994 ;
               RECT 26.934 23.158 26.986 23.194 ;
               RECT 26.934 24.358 26.986 24.394 ;
               RECT 26.934 25.558 26.986 25.594 ;
               RECT 26.934 26.758 26.986 26.794 ;
               RECT 26.934 27.958 26.986 27.994 ;
               RECT 26.934 29.158 26.986 29.194 ;
               RECT 26.934 30.358 26.986 30.394 ;
               RECT 26.934 31.558 26.986 31.594 ;
               RECT 26.934 32.758 26.986 32.794 ;
               RECT 26.934 33.958 26.986 33.994 ;
               RECT 26.934 35.158 26.986 35.194 ;
               RECT 26.934 36.358 26.986 36.394 ;
               RECT 26.934 37.558 26.986 37.594 ;
               RECT 26.934 38.758 26.986 38.794 ;
               RECT 26.934 39.958 26.986 39.994 ;
               RECT 26.934 41.158 26.986 41.194 ;
               RECT 26.934 42.358 26.986 42.394 ;
               RECT 26.934 43.558 26.986 43.594 ;
               RECT 26.934 44.758 26.986 44.794 ;
               RECT 26.934 45.958 26.986 45.994 ;
               RECT 26.934 47.158 26.986 47.194 ;
               RECT 26.934 48.358 26.986 48.394 ;
               RECT 26.934 50.142 26.986 50.178 ;
               RECT 26.934 50.382 26.986 50.418 ;
               RECT 26.934 54.702 26.986 54.738 ;
               RECT 26.934 54.942 26.986 54.978 ;
               RECT 26.934 57.478 26.986 57.514 ;
               RECT 26.934 58.678 26.986 58.714 ;
               RECT 26.934 59.878 26.986 59.914 ;
               RECT 26.934 61.078 26.986 61.114 ;
               RECT 26.934 62.278 26.986 62.314 ;
               RECT 26.934 63.478 26.986 63.514 ;
               RECT 26.934 64.678 26.986 64.714 ;
               RECT 26.934 65.878 26.986 65.914 ;
               RECT 26.934 67.078 26.986 67.114 ;
               RECT 26.934 68.278 26.986 68.314 ;
               RECT 26.934 69.478 26.986 69.514 ;
               RECT 26.934 70.678 26.986 70.714 ;
               RECT 26.934 71.878 26.986 71.914 ;
               RECT 26.934 73.078 26.986 73.114 ;
               RECT 26.934 74.278 26.986 74.314 ;
               RECT 26.934 75.478 26.986 75.514 ;
               RECT 26.934 76.678 26.986 76.714 ;
               RECT 26.934 77.878 26.986 77.914 ;
               RECT 26.934 79.078 26.986 79.114 ;
               RECT 26.934 80.278 26.986 80.314 ;
               RECT 26.934 81.478 26.986 81.514 ;
               RECT 26.934 82.678 26.986 82.714 ;
               RECT 26.934 83.878 26.986 83.914 ;
               RECT 26.934 85.078 26.986 85.114 ;
               RECT 26.934 86.278 26.986 86.314 ;
               RECT 26.934 87.478 26.986 87.514 ;
               RECT 26.934 88.678 26.986 88.714 ;
               RECT 26.934 89.878 26.986 89.914 ;
               RECT 26.934 91.078 26.986 91.114 ;
               RECT 26.934 92.278 26.986 92.314 ;
               RECT 26.934 93.478 26.986 93.514 ;
               RECT 26.934 94.678 26.986 94.714 ;
               RECT 26.934 95.878 26.986 95.914 ;
               RECT 26.934 97.078 26.986 97.114 ;
               RECT 26.934 98.278 26.986 98.314 ;
               RECT 26.934 99.478 26.986 99.514 ;
               RECT 26.934 100.678 26.986 100.714 ;
               RECT 26.934 101.878 26.986 101.914 ;
               RECT 26.934 103.078 26.986 103.114 ;
               RECT 26.934 104.278 26.986 104.314 ;
               RECT 27.014 0.806 27.066 0.842 ;
               RECT 27.014 2.006 27.066 2.042 ;
               RECT 27.014 3.206 27.066 3.242 ;
               RECT 27.014 4.406 27.066 4.442 ;
               RECT 27.014 5.606 27.066 5.642 ;
               RECT 27.014 6.806 27.066 6.842 ;
               RECT 27.014 8.006 27.066 8.042 ;
               RECT 27.014 9.206 27.066 9.242 ;
               RECT 27.014 10.406 27.066 10.442 ;
               RECT 27.014 11.606 27.066 11.642 ;
               RECT 27.014 12.806 27.066 12.842 ;
               RECT 27.014 14.006 27.066 14.042 ;
               RECT 27.014 15.206 27.066 15.242 ;
               RECT 27.014 16.406 27.066 16.442 ;
               RECT 27.014 17.606 27.066 17.642 ;
               RECT 27.014 18.806 27.066 18.842 ;
               RECT 27.014 20.006 27.066 20.042 ;
               RECT 27.014 21.206 27.066 21.242 ;
               RECT 27.014 22.406 27.066 22.442 ;
               RECT 27.014 23.606 27.066 23.642 ;
               RECT 27.014 24.806 27.066 24.842 ;
               RECT 27.014 26.006 27.066 26.042 ;
               RECT 27.014 27.206 27.066 27.242 ;
               RECT 27.014 28.406 27.066 28.442 ;
               RECT 27.014 29.606 27.066 29.642 ;
               RECT 27.014 30.806 27.066 30.842 ;
               RECT 27.014 32.006 27.066 32.042 ;
               RECT 27.014 33.206 27.066 33.242 ;
               RECT 27.014 34.406 27.066 34.442 ;
               RECT 27.014 35.606 27.066 35.642 ;
               RECT 27.014 36.806 27.066 36.842 ;
               RECT 27.014 38.006 27.066 38.042 ;
               RECT 27.014 39.206 27.066 39.242 ;
               RECT 27.014 40.406 27.066 40.442 ;
               RECT 27.014 41.606 27.066 41.642 ;
               RECT 27.014 42.806 27.066 42.842 ;
               RECT 27.014 44.006 27.066 44.042 ;
               RECT 27.014 45.206 27.066 45.242 ;
               RECT 27.014 46.406 27.066 46.442 ;
               RECT 27.014 47.606 27.066 47.642 ;
               RECT 27.014 49.422 27.066 49.458 ;
               RECT 27.014 49.662 27.066 49.698 ;
               RECT 27.014 55.422 27.066 55.458 ;
               RECT 27.014 55.662 27.066 55.698 ;
               RECT 27.014 56.726 27.066 56.762 ;
               RECT 27.014 57.926 27.066 57.962 ;
               RECT 27.014 59.126 27.066 59.162 ;
               RECT 27.014 60.326 27.066 60.362 ;
               RECT 27.014 61.526 27.066 61.562 ;
               RECT 27.014 62.726 27.066 62.762 ;
               RECT 27.014 63.926 27.066 63.962 ;
               RECT 27.014 65.126 27.066 65.162 ;
               RECT 27.014 66.326 27.066 66.362 ;
               RECT 27.014 67.526 27.066 67.562 ;
               RECT 27.014 68.726 27.066 68.762 ;
               RECT 27.014 69.926 27.066 69.962 ;
               RECT 27.014 71.126 27.066 71.162 ;
               RECT 27.014 72.326 27.066 72.362 ;
               RECT 27.014 73.526 27.066 73.562 ;
               RECT 27.014 74.726 27.066 74.762 ;
               RECT 27.014 75.926 27.066 75.962 ;
               RECT 27.014 77.126 27.066 77.162 ;
               RECT 27.014 78.326 27.066 78.362 ;
               RECT 27.014 79.526 27.066 79.562 ;
               RECT 27.014 80.726 27.066 80.762 ;
               RECT 27.014 81.926 27.066 81.962 ;
               RECT 27.014 83.126 27.066 83.162 ;
               RECT 27.014 84.326 27.066 84.362 ;
               RECT 27.014 85.526 27.066 85.562 ;
               RECT 27.014 86.726 27.066 86.762 ;
               RECT 27.014 87.926 27.066 87.962 ;
               RECT 27.014 89.126 27.066 89.162 ;
               RECT 27.014 90.326 27.066 90.362 ;
               RECT 27.014 91.526 27.066 91.562 ;
               RECT 27.014 92.726 27.066 92.762 ;
               RECT 27.014 93.926 27.066 93.962 ;
               RECT 27.014 95.126 27.066 95.162 ;
               RECT 27.014 96.326 27.066 96.362 ;
               RECT 27.014 97.526 27.066 97.562 ;
               RECT 27.014 98.726 27.066 98.762 ;
               RECT 27.014 99.926 27.066 99.962 ;
               RECT 27.014 101.126 27.066 101.162 ;
               RECT 27.014 102.326 27.066 102.362 ;
               RECT 27.014 103.526 27.066 103.562 ;
               RECT 27.094 1.558 27.146 1.594 ;
               RECT 27.094 2.758 27.146 2.794 ;
               RECT 27.094 3.958 27.146 3.994 ;
               RECT 27.094 5.158 27.146 5.194 ;
               RECT 27.094 6.358 27.146 6.394 ;
               RECT 27.094 7.558 27.146 7.594 ;
               RECT 27.094 8.758 27.146 8.794 ;
               RECT 27.094 9.958 27.146 9.994 ;
               RECT 27.094 11.158 27.146 11.194 ;
               RECT 27.094 12.358 27.146 12.394 ;
               RECT 27.094 13.558 27.146 13.594 ;
               RECT 27.094 14.758 27.146 14.794 ;
               RECT 27.094 15.958 27.146 15.994 ;
               RECT 27.094 17.158 27.146 17.194 ;
               RECT 27.094 18.358 27.146 18.394 ;
               RECT 27.094 19.558 27.146 19.594 ;
               RECT 27.094 20.758 27.146 20.794 ;
               RECT 27.094 21.958 27.146 21.994 ;
               RECT 27.094 23.158 27.146 23.194 ;
               RECT 27.094 24.358 27.146 24.394 ;
               RECT 27.094 25.558 27.146 25.594 ;
               RECT 27.094 26.758 27.146 26.794 ;
               RECT 27.094 27.958 27.146 27.994 ;
               RECT 27.094 29.158 27.146 29.194 ;
               RECT 27.094 30.358 27.146 30.394 ;
               RECT 27.094 31.558 27.146 31.594 ;
               RECT 27.094 32.758 27.146 32.794 ;
               RECT 27.094 33.958 27.146 33.994 ;
               RECT 27.094 35.158 27.146 35.194 ;
               RECT 27.094 36.358 27.146 36.394 ;
               RECT 27.094 37.558 27.146 37.594 ;
               RECT 27.094 38.758 27.146 38.794 ;
               RECT 27.094 39.958 27.146 39.994 ;
               RECT 27.094 41.158 27.146 41.194 ;
               RECT 27.094 42.358 27.146 42.394 ;
               RECT 27.094 43.558 27.146 43.594 ;
               RECT 27.094 44.758 27.146 44.794 ;
               RECT 27.094 45.958 27.146 45.994 ;
               RECT 27.094 47.158 27.146 47.194 ;
               RECT 27.094 48.358 27.146 48.394 ;
               RECT 27.094 50.142 27.146 50.178 ;
               RECT 27.094 50.382 27.146 50.418 ;
               RECT 27.094 54.702 27.146 54.738 ;
               RECT 27.094 54.942 27.146 54.978 ;
               RECT 27.094 57.478 27.146 57.514 ;
               RECT 27.094 58.678 27.146 58.714 ;
               RECT 27.094 59.878 27.146 59.914 ;
               RECT 27.094 61.078 27.146 61.114 ;
               RECT 27.094 62.278 27.146 62.314 ;
               RECT 27.094 63.478 27.146 63.514 ;
               RECT 27.094 64.678 27.146 64.714 ;
               RECT 27.094 65.878 27.146 65.914 ;
               RECT 27.094 67.078 27.146 67.114 ;
               RECT 27.094 68.278 27.146 68.314 ;
               RECT 27.094 69.478 27.146 69.514 ;
               RECT 27.094 70.678 27.146 70.714 ;
               RECT 27.094 71.878 27.146 71.914 ;
               RECT 27.094 73.078 27.146 73.114 ;
               RECT 27.094 74.278 27.146 74.314 ;
               RECT 27.094 75.478 27.146 75.514 ;
               RECT 27.094 76.678 27.146 76.714 ;
               RECT 27.094 77.878 27.146 77.914 ;
               RECT 27.094 79.078 27.146 79.114 ;
               RECT 27.094 80.278 27.146 80.314 ;
               RECT 27.094 81.478 27.146 81.514 ;
               RECT 27.094 82.678 27.146 82.714 ;
               RECT 27.094 83.878 27.146 83.914 ;
               RECT 27.094 85.078 27.146 85.114 ;
               RECT 27.094 86.278 27.146 86.314 ;
               RECT 27.094 87.478 27.146 87.514 ;
               RECT 27.094 88.678 27.146 88.714 ;
               RECT 27.094 89.878 27.146 89.914 ;
               RECT 27.094 91.078 27.146 91.114 ;
               RECT 27.094 92.278 27.146 92.314 ;
               RECT 27.094 93.478 27.146 93.514 ;
               RECT 27.094 94.678 27.146 94.714 ;
               RECT 27.094 95.878 27.146 95.914 ;
               RECT 27.094 97.078 27.146 97.114 ;
               RECT 27.094 98.278 27.146 98.314 ;
               RECT 27.094 99.478 27.146 99.514 ;
               RECT 27.094 100.678 27.146 100.714 ;
               RECT 27.094 101.878 27.146 101.914 ;
               RECT 27.094 103.078 27.146 103.114 ;
               RECT 27.094 104.278 27.146 104.314 ;
               RECT 27.174 0.281 27.226 0.317 ;
               RECT 27.174 104.803 27.226 104.839 ;
               RECT 27.254 0.806 27.306 0.842 ;
               RECT 27.254 2.006 27.306 2.042 ;
               RECT 27.254 3.206 27.306 3.242 ;
               RECT 27.254 4.406 27.306 4.442 ;
               RECT 27.254 5.606 27.306 5.642 ;
               RECT 27.254 6.806 27.306 6.842 ;
               RECT 27.254 8.006 27.306 8.042 ;
               RECT 27.254 9.206 27.306 9.242 ;
               RECT 27.254 10.406 27.306 10.442 ;
               RECT 27.254 11.606 27.306 11.642 ;
               RECT 27.254 12.806 27.306 12.842 ;
               RECT 27.254 14.006 27.306 14.042 ;
               RECT 27.254 15.206 27.306 15.242 ;
               RECT 27.254 16.406 27.306 16.442 ;
               RECT 27.254 17.606 27.306 17.642 ;
               RECT 27.254 18.806 27.306 18.842 ;
               RECT 27.254 20.006 27.306 20.042 ;
               RECT 27.254 21.206 27.306 21.242 ;
               RECT 27.254 22.406 27.306 22.442 ;
               RECT 27.254 23.606 27.306 23.642 ;
               RECT 27.254 24.806 27.306 24.842 ;
               RECT 27.254 26.006 27.306 26.042 ;
               RECT 27.254 27.206 27.306 27.242 ;
               RECT 27.254 28.406 27.306 28.442 ;
               RECT 27.254 29.606 27.306 29.642 ;
               RECT 27.254 30.806 27.306 30.842 ;
               RECT 27.254 32.006 27.306 32.042 ;
               RECT 27.254 33.206 27.306 33.242 ;
               RECT 27.254 34.406 27.306 34.442 ;
               RECT 27.254 35.606 27.306 35.642 ;
               RECT 27.254 36.806 27.306 36.842 ;
               RECT 27.254 38.006 27.306 38.042 ;
               RECT 27.254 39.206 27.306 39.242 ;
               RECT 27.254 40.406 27.306 40.442 ;
               RECT 27.254 41.606 27.306 41.642 ;
               RECT 27.254 42.806 27.306 42.842 ;
               RECT 27.254 44.006 27.306 44.042 ;
               RECT 27.254 45.206 27.306 45.242 ;
               RECT 27.254 46.406 27.306 46.442 ;
               RECT 27.254 47.606 27.306 47.642 ;
               RECT 27.254 49.422 27.306 49.458 ;
               RECT 27.254 49.662 27.306 49.698 ;
               RECT 27.254 51.102 27.306 51.138 ;
               RECT 27.254 51.582 27.306 51.618 ;
               RECT 27.254 53.502 27.306 53.538 ;
               RECT 27.254 53.982 27.306 54.018 ;
               RECT 27.254 55.422 27.306 55.458 ;
               RECT 27.254 55.662 27.306 55.698 ;
               RECT 27.254 56.726 27.306 56.762 ;
               RECT 27.254 57.926 27.306 57.962 ;
               RECT 27.254 59.126 27.306 59.162 ;
               RECT 27.254 60.326 27.306 60.362 ;
               RECT 27.254 61.526 27.306 61.562 ;
               RECT 27.254 62.726 27.306 62.762 ;
               RECT 27.254 63.926 27.306 63.962 ;
               RECT 27.254 65.126 27.306 65.162 ;
               RECT 27.254 66.326 27.306 66.362 ;
               RECT 27.254 67.526 27.306 67.562 ;
               RECT 27.254 68.726 27.306 68.762 ;
               RECT 27.254 69.926 27.306 69.962 ;
               RECT 27.254 71.126 27.306 71.162 ;
               RECT 27.254 72.326 27.306 72.362 ;
               RECT 27.254 73.526 27.306 73.562 ;
               RECT 27.254 74.726 27.306 74.762 ;
               RECT 27.254 75.926 27.306 75.962 ;
               RECT 27.254 77.126 27.306 77.162 ;
               RECT 27.254 78.326 27.306 78.362 ;
               RECT 27.254 79.526 27.306 79.562 ;
               RECT 27.254 80.726 27.306 80.762 ;
               RECT 27.254 81.926 27.306 81.962 ;
               RECT 27.254 83.126 27.306 83.162 ;
               RECT 27.254 84.326 27.306 84.362 ;
               RECT 27.254 85.526 27.306 85.562 ;
               RECT 27.254 86.726 27.306 86.762 ;
               RECT 27.254 87.926 27.306 87.962 ;
               RECT 27.254 89.126 27.306 89.162 ;
               RECT 27.254 90.326 27.306 90.362 ;
               RECT 27.254 91.526 27.306 91.562 ;
               RECT 27.254 92.726 27.306 92.762 ;
               RECT 27.254 93.926 27.306 93.962 ;
               RECT 27.254 95.126 27.306 95.162 ;
               RECT 27.254 96.326 27.306 96.362 ;
               RECT 27.254 97.526 27.306 97.562 ;
               RECT 27.254 98.726 27.306 98.762 ;
               RECT 27.254 99.926 27.306 99.962 ;
               RECT 27.254 101.126 27.306 101.162 ;
               RECT 27.254 102.326 27.306 102.362 ;
               RECT 27.254 103.526 27.306 103.562 ;
               RECT 27.334 1.558 27.386 1.594 ;
               RECT 27.334 2.758 27.386 2.794 ;
               RECT 27.334 3.958 27.386 3.994 ;
               RECT 27.334 5.158 27.386 5.194 ;
               RECT 27.334 6.358 27.386 6.394 ;
               RECT 27.334 7.558 27.386 7.594 ;
               RECT 27.334 8.758 27.386 8.794 ;
               RECT 27.334 9.958 27.386 9.994 ;
               RECT 27.334 11.158 27.386 11.194 ;
               RECT 27.334 12.358 27.386 12.394 ;
               RECT 27.334 13.558 27.386 13.594 ;
               RECT 27.334 14.758 27.386 14.794 ;
               RECT 27.334 15.958 27.386 15.994 ;
               RECT 27.334 17.158 27.386 17.194 ;
               RECT 27.334 18.358 27.386 18.394 ;
               RECT 27.334 19.558 27.386 19.594 ;
               RECT 27.334 20.758 27.386 20.794 ;
               RECT 27.334 21.958 27.386 21.994 ;
               RECT 27.334 23.158 27.386 23.194 ;
               RECT 27.334 24.358 27.386 24.394 ;
               RECT 27.334 25.558 27.386 25.594 ;
               RECT 27.334 26.758 27.386 26.794 ;
               RECT 27.334 27.958 27.386 27.994 ;
               RECT 27.334 29.158 27.386 29.194 ;
               RECT 27.334 30.358 27.386 30.394 ;
               RECT 27.334 31.558 27.386 31.594 ;
               RECT 27.334 32.758 27.386 32.794 ;
               RECT 27.334 33.958 27.386 33.994 ;
               RECT 27.334 35.158 27.386 35.194 ;
               RECT 27.334 36.358 27.386 36.394 ;
               RECT 27.334 37.558 27.386 37.594 ;
               RECT 27.334 38.758 27.386 38.794 ;
               RECT 27.334 39.958 27.386 39.994 ;
               RECT 27.334 41.158 27.386 41.194 ;
               RECT 27.334 42.358 27.386 42.394 ;
               RECT 27.334 43.558 27.386 43.594 ;
               RECT 27.334 44.758 27.386 44.794 ;
               RECT 27.334 45.958 27.386 45.994 ;
               RECT 27.334 47.158 27.386 47.194 ;
               RECT 27.334 48.358 27.386 48.394 ;
               RECT 27.334 50.142 27.386 50.178 ;
               RECT 27.334 50.382 27.386 50.418 ;
               RECT 27.334 54.702 27.386 54.738 ;
               RECT 27.334 54.942 27.386 54.978 ;
               RECT 27.334 57.478 27.386 57.514 ;
               RECT 27.334 58.678 27.386 58.714 ;
               RECT 27.334 59.878 27.386 59.914 ;
               RECT 27.334 61.078 27.386 61.114 ;
               RECT 27.334 62.278 27.386 62.314 ;
               RECT 27.334 63.478 27.386 63.514 ;
               RECT 27.334 64.678 27.386 64.714 ;
               RECT 27.334 65.878 27.386 65.914 ;
               RECT 27.334 67.078 27.386 67.114 ;
               RECT 27.334 68.278 27.386 68.314 ;
               RECT 27.334 69.478 27.386 69.514 ;
               RECT 27.334 70.678 27.386 70.714 ;
               RECT 27.334 71.878 27.386 71.914 ;
               RECT 27.334 73.078 27.386 73.114 ;
               RECT 27.334 74.278 27.386 74.314 ;
               RECT 27.334 75.478 27.386 75.514 ;
               RECT 27.334 76.678 27.386 76.714 ;
               RECT 27.334 77.878 27.386 77.914 ;
               RECT 27.334 79.078 27.386 79.114 ;
               RECT 27.334 80.278 27.386 80.314 ;
               RECT 27.334 81.478 27.386 81.514 ;
               RECT 27.334 82.678 27.386 82.714 ;
               RECT 27.334 83.878 27.386 83.914 ;
               RECT 27.334 85.078 27.386 85.114 ;
               RECT 27.334 86.278 27.386 86.314 ;
               RECT 27.334 87.478 27.386 87.514 ;
               RECT 27.334 88.678 27.386 88.714 ;
               RECT 27.334 89.878 27.386 89.914 ;
               RECT 27.334 91.078 27.386 91.114 ;
               RECT 27.334 92.278 27.386 92.314 ;
               RECT 27.334 93.478 27.386 93.514 ;
               RECT 27.334 94.678 27.386 94.714 ;
               RECT 27.334 95.878 27.386 95.914 ;
               RECT 27.334 97.078 27.386 97.114 ;
               RECT 27.334 98.278 27.386 98.314 ;
               RECT 27.334 99.478 27.386 99.514 ;
               RECT 27.334 100.678 27.386 100.714 ;
               RECT 27.334 101.878 27.386 101.914 ;
               RECT 27.334 103.078 27.386 103.114 ;
               RECT 27.334 104.278 27.386 104.314 ;
               RECT 27.414 0.806 27.466 0.842 ;
               RECT 27.414 2.006 27.466 2.042 ;
               RECT 27.414 3.206 27.466 3.242 ;
               RECT 27.414 4.406 27.466 4.442 ;
               RECT 27.414 5.606 27.466 5.642 ;
               RECT 27.414 6.806 27.466 6.842 ;
               RECT 27.414 8.006 27.466 8.042 ;
               RECT 27.414 9.206 27.466 9.242 ;
               RECT 27.414 10.406 27.466 10.442 ;
               RECT 27.414 11.606 27.466 11.642 ;
               RECT 27.414 12.806 27.466 12.842 ;
               RECT 27.414 14.006 27.466 14.042 ;
               RECT 27.414 15.206 27.466 15.242 ;
               RECT 27.414 16.406 27.466 16.442 ;
               RECT 27.414 17.606 27.466 17.642 ;
               RECT 27.414 18.806 27.466 18.842 ;
               RECT 27.414 20.006 27.466 20.042 ;
               RECT 27.414 21.206 27.466 21.242 ;
               RECT 27.414 22.406 27.466 22.442 ;
               RECT 27.414 23.606 27.466 23.642 ;
               RECT 27.414 24.806 27.466 24.842 ;
               RECT 27.414 26.006 27.466 26.042 ;
               RECT 27.414 27.206 27.466 27.242 ;
               RECT 27.414 28.406 27.466 28.442 ;
               RECT 27.414 29.606 27.466 29.642 ;
               RECT 27.414 30.806 27.466 30.842 ;
               RECT 27.414 32.006 27.466 32.042 ;
               RECT 27.414 33.206 27.466 33.242 ;
               RECT 27.414 34.406 27.466 34.442 ;
               RECT 27.414 35.606 27.466 35.642 ;
               RECT 27.414 36.806 27.466 36.842 ;
               RECT 27.414 38.006 27.466 38.042 ;
               RECT 27.414 39.206 27.466 39.242 ;
               RECT 27.414 40.406 27.466 40.442 ;
               RECT 27.414 41.606 27.466 41.642 ;
               RECT 27.414 42.806 27.466 42.842 ;
               RECT 27.414 44.006 27.466 44.042 ;
               RECT 27.414 45.206 27.466 45.242 ;
               RECT 27.414 46.406 27.466 46.442 ;
               RECT 27.414 47.606 27.466 47.642 ;
               RECT 27.414 49.422 27.466 49.458 ;
               RECT 27.414 49.662 27.466 49.698 ;
               RECT 27.414 55.422 27.466 55.458 ;
               RECT 27.414 55.662 27.466 55.698 ;
               RECT 27.414 56.726 27.466 56.762 ;
               RECT 27.414 57.926 27.466 57.962 ;
               RECT 27.414 59.126 27.466 59.162 ;
               RECT 27.414 60.326 27.466 60.362 ;
               RECT 27.414 61.526 27.466 61.562 ;
               RECT 27.414 62.726 27.466 62.762 ;
               RECT 27.414 63.926 27.466 63.962 ;
               RECT 27.414 65.126 27.466 65.162 ;
               RECT 27.414 66.326 27.466 66.362 ;
               RECT 27.414 67.526 27.466 67.562 ;
               RECT 27.414 68.726 27.466 68.762 ;
               RECT 27.414 69.926 27.466 69.962 ;
               RECT 27.414 71.126 27.466 71.162 ;
               RECT 27.414 72.326 27.466 72.362 ;
               RECT 27.414 73.526 27.466 73.562 ;
               RECT 27.414 74.726 27.466 74.762 ;
               RECT 27.414 75.926 27.466 75.962 ;
               RECT 27.414 77.126 27.466 77.162 ;
               RECT 27.414 78.326 27.466 78.362 ;
               RECT 27.414 79.526 27.466 79.562 ;
               RECT 27.414 80.726 27.466 80.762 ;
               RECT 27.414 81.926 27.466 81.962 ;
               RECT 27.414 83.126 27.466 83.162 ;
               RECT 27.414 84.326 27.466 84.362 ;
               RECT 27.414 85.526 27.466 85.562 ;
               RECT 27.414 86.726 27.466 86.762 ;
               RECT 27.414 87.926 27.466 87.962 ;
               RECT 27.414 89.126 27.466 89.162 ;
               RECT 27.414 90.326 27.466 90.362 ;
               RECT 27.414 91.526 27.466 91.562 ;
               RECT 27.414 92.726 27.466 92.762 ;
               RECT 27.414 93.926 27.466 93.962 ;
               RECT 27.414 95.126 27.466 95.162 ;
               RECT 27.414 96.326 27.466 96.362 ;
               RECT 27.414 97.526 27.466 97.562 ;
               RECT 27.414 98.726 27.466 98.762 ;
               RECT 27.414 99.926 27.466 99.962 ;
               RECT 27.414 101.126 27.466 101.162 ;
               RECT 27.414 102.326 27.466 102.362 ;
               RECT 27.414 103.526 27.466 103.562 ;
               RECT 27.494 1.558 27.546 1.594 ;
               RECT 27.494 2.758 27.546 2.794 ;
               RECT 27.494 3.958 27.546 3.994 ;
               RECT 27.494 5.158 27.546 5.194 ;
               RECT 27.494 6.358 27.546 6.394 ;
               RECT 27.494 7.558 27.546 7.594 ;
               RECT 27.494 8.758 27.546 8.794 ;
               RECT 27.494 9.958 27.546 9.994 ;
               RECT 27.494 11.158 27.546 11.194 ;
               RECT 27.494 12.358 27.546 12.394 ;
               RECT 27.494 13.558 27.546 13.594 ;
               RECT 27.494 14.758 27.546 14.794 ;
               RECT 27.494 15.958 27.546 15.994 ;
               RECT 27.494 17.158 27.546 17.194 ;
               RECT 27.494 18.358 27.546 18.394 ;
               RECT 27.494 19.558 27.546 19.594 ;
               RECT 27.494 20.758 27.546 20.794 ;
               RECT 27.494 21.958 27.546 21.994 ;
               RECT 27.494 23.158 27.546 23.194 ;
               RECT 27.494 24.358 27.546 24.394 ;
               RECT 27.494 25.558 27.546 25.594 ;
               RECT 27.494 26.758 27.546 26.794 ;
               RECT 27.494 27.958 27.546 27.994 ;
               RECT 27.494 29.158 27.546 29.194 ;
               RECT 27.494 30.358 27.546 30.394 ;
               RECT 27.494 31.558 27.546 31.594 ;
               RECT 27.494 32.758 27.546 32.794 ;
               RECT 27.494 33.958 27.546 33.994 ;
               RECT 27.494 35.158 27.546 35.194 ;
               RECT 27.494 36.358 27.546 36.394 ;
               RECT 27.494 37.558 27.546 37.594 ;
               RECT 27.494 38.758 27.546 38.794 ;
               RECT 27.494 39.958 27.546 39.994 ;
               RECT 27.494 41.158 27.546 41.194 ;
               RECT 27.494 42.358 27.546 42.394 ;
               RECT 27.494 43.558 27.546 43.594 ;
               RECT 27.494 44.758 27.546 44.794 ;
               RECT 27.494 45.958 27.546 45.994 ;
               RECT 27.494 47.158 27.546 47.194 ;
               RECT 27.494 48.358 27.546 48.394 ;
               RECT 27.494 50.142 27.546 50.178 ;
               RECT 27.494 50.382 27.546 50.418 ;
               RECT 27.494 54.702 27.546 54.738 ;
               RECT 27.494 54.942 27.546 54.978 ;
               RECT 27.494 57.478 27.546 57.514 ;
               RECT 27.494 58.678 27.546 58.714 ;
               RECT 27.494 59.878 27.546 59.914 ;
               RECT 27.494 61.078 27.546 61.114 ;
               RECT 27.494 62.278 27.546 62.314 ;
               RECT 27.494 63.478 27.546 63.514 ;
               RECT 27.494 64.678 27.546 64.714 ;
               RECT 27.494 65.878 27.546 65.914 ;
               RECT 27.494 67.078 27.546 67.114 ;
               RECT 27.494 68.278 27.546 68.314 ;
               RECT 27.494 69.478 27.546 69.514 ;
               RECT 27.494 70.678 27.546 70.714 ;
               RECT 27.494 71.878 27.546 71.914 ;
               RECT 27.494 73.078 27.546 73.114 ;
               RECT 27.494 74.278 27.546 74.314 ;
               RECT 27.494 75.478 27.546 75.514 ;
               RECT 27.494 76.678 27.546 76.714 ;
               RECT 27.494 77.878 27.546 77.914 ;
               RECT 27.494 79.078 27.546 79.114 ;
               RECT 27.494 80.278 27.546 80.314 ;
               RECT 27.494 81.478 27.546 81.514 ;
               RECT 27.494 82.678 27.546 82.714 ;
               RECT 27.494 83.878 27.546 83.914 ;
               RECT 27.494 85.078 27.546 85.114 ;
               RECT 27.494 86.278 27.546 86.314 ;
               RECT 27.494 87.478 27.546 87.514 ;
               RECT 27.494 88.678 27.546 88.714 ;
               RECT 27.494 89.878 27.546 89.914 ;
               RECT 27.494 91.078 27.546 91.114 ;
               RECT 27.494 92.278 27.546 92.314 ;
               RECT 27.494 93.478 27.546 93.514 ;
               RECT 27.494 94.678 27.546 94.714 ;
               RECT 27.494 95.878 27.546 95.914 ;
               RECT 27.494 97.078 27.546 97.114 ;
               RECT 27.494 98.278 27.546 98.314 ;
               RECT 27.494 99.478 27.546 99.514 ;
               RECT 27.494 100.678 27.546 100.714 ;
               RECT 27.494 101.878 27.546 101.914 ;
               RECT 27.494 103.078 27.546 103.114 ;
               RECT 27.494 104.278 27.546 104.314 ;
               RECT 27.574 0.281 27.626 0.317 ;
               RECT 27.574 104.803 27.626 104.839 ;
               RECT 27.654 0.806 27.706 0.842 ;
               RECT 27.654 2.006 27.706 2.042 ;
               RECT 27.654 3.206 27.706 3.242 ;
               RECT 27.654 4.406 27.706 4.442 ;
               RECT 27.654 5.606 27.706 5.642 ;
               RECT 27.654 6.806 27.706 6.842 ;
               RECT 27.654 8.006 27.706 8.042 ;
               RECT 27.654 9.206 27.706 9.242 ;
               RECT 27.654 10.406 27.706 10.442 ;
               RECT 27.654 11.606 27.706 11.642 ;
               RECT 27.654 12.806 27.706 12.842 ;
               RECT 27.654 14.006 27.706 14.042 ;
               RECT 27.654 15.206 27.706 15.242 ;
               RECT 27.654 16.406 27.706 16.442 ;
               RECT 27.654 17.606 27.706 17.642 ;
               RECT 27.654 18.806 27.706 18.842 ;
               RECT 27.654 20.006 27.706 20.042 ;
               RECT 27.654 21.206 27.706 21.242 ;
               RECT 27.654 22.406 27.706 22.442 ;
               RECT 27.654 23.606 27.706 23.642 ;
               RECT 27.654 24.806 27.706 24.842 ;
               RECT 27.654 26.006 27.706 26.042 ;
               RECT 27.654 27.206 27.706 27.242 ;
               RECT 27.654 28.406 27.706 28.442 ;
               RECT 27.654 29.606 27.706 29.642 ;
               RECT 27.654 30.806 27.706 30.842 ;
               RECT 27.654 32.006 27.706 32.042 ;
               RECT 27.654 33.206 27.706 33.242 ;
               RECT 27.654 34.406 27.706 34.442 ;
               RECT 27.654 35.606 27.706 35.642 ;
               RECT 27.654 36.806 27.706 36.842 ;
               RECT 27.654 38.006 27.706 38.042 ;
               RECT 27.654 39.206 27.706 39.242 ;
               RECT 27.654 40.406 27.706 40.442 ;
               RECT 27.654 41.606 27.706 41.642 ;
               RECT 27.654 42.806 27.706 42.842 ;
               RECT 27.654 44.006 27.706 44.042 ;
               RECT 27.654 45.206 27.706 45.242 ;
               RECT 27.654 46.406 27.706 46.442 ;
               RECT 27.654 47.606 27.706 47.642 ;
               RECT 27.654 49.422 27.706 49.458 ;
               RECT 27.654 49.662 27.706 49.698 ;
               RECT 27.654 55.422 27.706 55.458 ;
               RECT 27.654 55.662 27.706 55.698 ;
               RECT 27.654 56.726 27.706 56.762 ;
               RECT 27.654 57.926 27.706 57.962 ;
               RECT 27.654 59.126 27.706 59.162 ;
               RECT 27.654 60.326 27.706 60.362 ;
               RECT 27.654 61.526 27.706 61.562 ;
               RECT 27.654 62.726 27.706 62.762 ;
               RECT 27.654 63.926 27.706 63.962 ;
               RECT 27.654 65.126 27.706 65.162 ;
               RECT 27.654 66.326 27.706 66.362 ;
               RECT 27.654 67.526 27.706 67.562 ;
               RECT 27.654 68.726 27.706 68.762 ;
               RECT 27.654 69.926 27.706 69.962 ;
               RECT 27.654 71.126 27.706 71.162 ;
               RECT 27.654 72.326 27.706 72.362 ;
               RECT 27.654 73.526 27.706 73.562 ;
               RECT 27.654 74.726 27.706 74.762 ;
               RECT 27.654 75.926 27.706 75.962 ;
               RECT 27.654 77.126 27.706 77.162 ;
               RECT 27.654 78.326 27.706 78.362 ;
               RECT 27.654 79.526 27.706 79.562 ;
               RECT 27.654 80.726 27.706 80.762 ;
               RECT 27.654 81.926 27.706 81.962 ;
               RECT 27.654 83.126 27.706 83.162 ;
               RECT 27.654 84.326 27.706 84.362 ;
               RECT 27.654 85.526 27.706 85.562 ;
               RECT 27.654 86.726 27.706 86.762 ;
               RECT 27.654 87.926 27.706 87.962 ;
               RECT 27.654 89.126 27.706 89.162 ;
               RECT 27.654 90.326 27.706 90.362 ;
               RECT 27.654 91.526 27.706 91.562 ;
               RECT 27.654 92.726 27.706 92.762 ;
               RECT 27.654 93.926 27.706 93.962 ;
               RECT 27.654 95.126 27.706 95.162 ;
               RECT 27.654 96.326 27.706 96.362 ;
               RECT 27.654 97.526 27.706 97.562 ;
               RECT 27.654 98.726 27.706 98.762 ;
               RECT 27.654 99.926 27.706 99.962 ;
               RECT 27.654 101.126 27.706 101.162 ;
               RECT 27.654 102.326 27.706 102.362 ;
               RECT 27.654 103.526 27.706 103.562 ;
               RECT 27.734 1.558 27.786 1.594 ;
               RECT 27.734 2.758 27.786 2.794 ;
               RECT 27.734 3.958 27.786 3.994 ;
               RECT 27.734 5.158 27.786 5.194 ;
               RECT 27.734 6.358 27.786 6.394 ;
               RECT 27.734 7.558 27.786 7.594 ;
               RECT 27.734 8.758 27.786 8.794 ;
               RECT 27.734 9.958 27.786 9.994 ;
               RECT 27.734 11.158 27.786 11.194 ;
               RECT 27.734 12.358 27.786 12.394 ;
               RECT 27.734 13.558 27.786 13.594 ;
               RECT 27.734 14.758 27.786 14.794 ;
               RECT 27.734 15.958 27.786 15.994 ;
               RECT 27.734 17.158 27.786 17.194 ;
               RECT 27.734 18.358 27.786 18.394 ;
               RECT 27.734 19.558 27.786 19.594 ;
               RECT 27.734 20.758 27.786 20.794 ;
               RECT 27.734 21.958 27.786 21.994 ;
               RECT 27.734 23.158 27.786 23.194 ;
               RECT 27.734 24.358 27.786 24.394 ;
               RECT 27.734 25.558 27.786 25.594 ;
               RECT 27.734 26.758 27.786 26.794 ;
               RECT 27.734 27.958 27.786 27.994 ;
               RECT 27.734 29.158 27.786 29.194 ;
               RECT 27.734 30.358 27.786 30.394 ;
               RECT 27.734 31.558 27.786 31.594 ;
               RECT 27.734 32.758 27.786 32.794 ;
               RECT 27.734 33.958 27.786 33.994 ;
               RECT 27.734 35.158 27.786 35.194 ;
               RECT 27.734 36.358 27.786 36.394 ;
               RECT 27.734 37.558 27.786 37.594 ;
               RECT 27.734 38.758 27.786 38.794 ;
               RECT 27.734 39.958 27.786 39.994 ;
               RECT 27.734 41.158 27.786 41.194 ;
               RECT 27.734 42.358 27.786 42.394 ;
               RECT 27.734 43.558 27.786 43.594 ;
               RECT 27.734 44.758 27.786 44.794 ;
               RECT 27.734 45.958 27.786 45.994 ;
               RECT 27.734 47.158 27.786 47.194 ;
               RECT 27.734 48.358 27.786 48.394 ;
               RECT 27.734 50.142 27.786 50.178 ;
               RECT 27.734 50.382 27.786 50.418 ;
               RECT 27.734 54.702 27.786 54.738 ;
               RECT 27.734 54.942 27.786 54.978 ;
               RECT 27.734 57.478 27.786 57.514 ;
               RECT 27.734 58.678 27.786 58.714 ;
               RECT 27.734 59.878 27.786 59.914 ;
               RECT 27.734 61.078 27.786 61.114 ;
               RECT 27.734 62.278 27.786 62.314 ;
               RECT 27.734 63.478 27.786 63.514 ;
               RECT 27.734 64.678 27.786 64.714 ;
               RECT 27.734 65.878 27.786 65.914 ;
               RECT 27.734 67.078 27.786 67.114 ;
               RECT 27.734 68.278 27.786 68.314 ;
               RECT 27.734 69.478 27.786 69.514 ;
               RECT 27.734 70.678 27.786 70.714 ;
               RECT 27.734 71.878 27.786 71.914 ;
               RECT 27.734 73.078 27.786 73.114 ;
               RECT 27.734 74.278 27.786 74.314 ;
               RECT 27.734 75.478 27.786 75.514 ;
               RECT 27.734 76.678 27.786 76.714 ;
               RECT 27.734 77.878 27.786 77.914 ;
               RECT 27.734 79.078 27.786 79.114 ;
               RECT 27.734 80.278 27.786 80.314 ;
               RECT 27.734 81.478 27.786 81.514 ;
               RECT 27.734 82.678 27.786 82.714 ;
               RECT 27.734 83.878 27.786 83.914 ;
               RECT 27.734 85.078 27.786 85.114 ;
               RECT 27.734 86.278 27.786 86.314 ;
               RECT 27.734 87.478 27.786 87.514 ;
               RECT 27.734 88.678 27.786 88.714 ;
               RECT 27.734 89.878 27.786 89.914 ;
               RECT 27.734 91.078 27.786 91.114 ;
               RECT 27.734 92.278 27.786 92.314 ;
               RECT 27.734 93.478 27.786 93.514 ;
               RECT 27.734 94.678 27.786 94.714 ;
               RECT 27.734 95.878 27.786 95.914 ;
               RECT 27.734 97.078 27.786 97.114 ;
               RECT 27.734 98.278 27.786 98.314 ;
               RECT 27.734 99.478 27.786 99.514 ;
               RECT 27.734 100.678 27.786 100.714 ;
               RECT 27.734 101.878 27.786 101.914 ;
               RECT 27.734 103.078 27.786 103.114 ;
               RECT 27.734 104.278 27.786 104.314 ;
               RECT 27.814 0.806 27.866 0.842 ;
               RECT 27.814 2.006 27.866 2.042 ;
               RECT 27.814 3.206 27.866 3.242 ;
               RECT 27.814 4.406 27.866 4.442 ;
               RECT 27.814 5.606 27.866 5.642 ;
               RECT 27.814 6.806 27.866 6.842 ;
               RECT 27.814 8.006 27.866 8.042 ;
               RECT 27.814 9.206 27.866 9.242 ;
               RECT 27.814 10.406 27.866 10.442 ;
               RECT 27.814 11.606 27.866 11.642 ;
               RECT 27.814 12.806 27.866 12.842 ;
               RECT 27.814 14.006 27.866 14.042 ;
               RECT 27.814 15.206 27.866 15.242 ;
               RECT 27.814 16.406 27.866 16.442 ;
               RECT 27.814 17.606 27.866 17.642 ;
               RECT 27.814 18.806 27.866 18.842 ;
               RECT 27.814 20.006 27.866 20.042 ;
               RECT 27.814 21.206 27.866 21.242 ;
               RECT 27.814 22.406 27.866 22.442 ;
               RECT 27.814 23.606 27.866 23.642 ;
               RECT 27.814 24.806 27.866 24.842 ;
               RECT 27.814 26.006 27.866 26.042 ;
               RECT 27.814 27.206 27.866 27.242 ;
               RECT 27.814 28.406 27.866 28.442 ;
               RECT 27.814 29.606 27.866 29.642 ;
               RECT 27.814 30.806 27.866 30.842 ;
               RECT 27.814 32.006 27.866 32.042 ;
               RECT 27.814 33.206 27.866 33.242 ;
               RECT 27.814 34.406 27.866 34.442 ;
               RECT 27.814 35.606 27.866 35.642 ;
               RECT 27.814 36.806 27.866 36.842 ;
               RECT 27.814 38.006 27.866 38.042 ;
               RECT 27.814 39.206 27.866 39.242 ;
               RECT 27.814 40.406 27.866 40.442 ;
               RECT 27.814 41.606 27.866 41.642 ;
               RECT 27.814 42.806 27.866 42.842 ;
               RECT 27.814 44.006 27.866 44.042 ;
               RECT 27.814 45.206 27.866 45.242 ;
               RECT 27.814 46.406 27.866 46.442 ;
               RECT 27.814 47.606 27.866 47.642 ;
               RECT 27.814 49.422 27.866 49.458 ;
               RECT 27.814 49.662 27.866 49.698 ;
               RECT 27.814 55.422 27.866 55.458 ;
               RECT 27.814 55.662 27.866 55.698 ;
               RECT 27.814 56.726 27.866 56.762 ;
               RECT 27.814 57.926 27.866 57.962 ;
               RECT 27.814 59.126 27.866 59.162 ;
               RECT 27.814 60.326 27.866 60.362 ;
               RECT 27.814 61.526 27.866 61.562 ;
               RECT 27.814 62.726 27.866 62.762 ;
               RECT 27.814 63.926 27.866 63.962 ;
               RECT 27.814 65.126 27.866 65.162 ;
               RECT 27.814 66.326 27.866 66.362 ;
               RECT 27.814 67.526 27.866 67.562 ;
               RECT 27.814 68.726 27.866 68.762 ;
               RECT 27.814 69.926 27.866 69.962 ;
               RECT 27.814 71.126 27.866 71.162 ;
               RECT 27.814 72.326 27.866 72.362 ;
               RECT 27.814 73.526 27.866 73.562 ;
               RECT 27.814 74.726 27.866 74.762 ;
               RECT 27.814 75.926 27.866 75.962 ;
               RECT 27.814 77.126 27.866 77.162 ;
               RECT 27.814 78.326 27.866 78.362 ;
               RECT 27.814 79.526 27.866 79.562 ;
               RECT 27.814 80.726 27.866 80.762 ;
               RECT 27.814 81.926 27.866 81.962 ;
               RECT 27.814 83.126 27.866 83.162 ;
               RECT 27.814 84.326 27.866 84.362 ;
               RECT 27.814 85.526 27.866 85.562 ;
               RECT 27.814 86.726 27.866 86.762 ;
               RECT 27.814 87.926 27.866 87.962 ;
               RECT 27.814 89.126 27.866 89.162 ;
               RECT 27.814 90.326 27.866 90.362 ;
               RECT 27.814 91.526 27.866 91.562 ;
               RECT 27.814 92.726 27.866 92.762 ;
               RECT 27.814 93.926 27.866 93.962 ;
               RECT 27.814 95.126 27.866 95.162 ;
               RECT 27.814 96.326 27.866 96.362 ;
               RECT 27.814 97.526 27.866 97.562 ;
               RECT 27.814 98.726 27.866 98.762 ;
               RECT 27.814 99.926 27.866 99.962 ;
               RECT 27.814 101.126 27.866 101.162 ;
               RECT 27.814 102.326 27.866 102.362 ;
               RECT 27.814 103.526 27.866 103.562 ;
               RECT 27.894 1.558 27.946 1.594 ;
               RECT 27.894 2.758 27.946 2.794 ;
               RECT 27.894 3.958 27.946 3.994 ;
               RECT 27.894 5.158 27.946 5.194 ;
               RECT 27.894 6.358 27.946 6.394 ;
               RECT 27.894 7.558 27.946 7.594 ;
               RECT 27.894 8.758 27.946 8.794 ;
               RECT 27.894 9.958 27.946 9.994 ;
               RECT 27.894 11.158 27.946 11.194 ;
               RECT 27.894 12.358 27.946 12.394 ;
               RECT 27.894 13.558 27.946 13.594 ;
               RECT 27.894 14.758 27.946 14.794 ;
               RECT 27.894 15.958 27.946 15.994 ;
               RECT 27.894 17.158 27.946 17.194 ;
               RECT 27.894 18.358 27.946 18.394 ;
               RECT 27.894 19.558 27.946 19.594 ;
               RECT 27.894 20.758 27.946 20.794 ;
               RECT 27.894 21.958 27.946 21.994 ;
               RECT 27.894 23.158 27.946 23.194 ;
               RECT 27.894 24.358 27.946 24.394 ;
               RECT 27.894 25.558 27.946 25.594 ;
               RECT 27.894 26.758 27.946 26.794 ;
               RECT 27.894 27.958 27.946 27.994 ;
               RECT 27.894 29.158 27.946 29.194 ;
               RECT 27.894 30.358 27.946 30.394 ;
               RECT 27.894 31.558 27.946 31.594 ;
               RECT 27.894 32.758 27.946 32.794 ;
               RECT 27.894 33.958 27.946 33.994 ;
               RECT 27.894 35.158 27.946 35.194 ;
               RECT 27.894 36.358 27.946 36.394 ;
               RECT 27.894 37.558 27.946 37.594 ;
               RECT 27.894 38.758 27.946 38.794 ;
               RECT 27.894 39.958 27.946 39.994 ;
               RECT 27.894 41.158 27.946 41.194 ;
               RECT 27.894 42.358 27.946 42.394 ;
               RECT 27.894 43.558 27.946 43.594 ;
               RECT 27.894 44.758 27.946 44.794 ;
               RECT 27.894 45.958 27.946 45.994 ;
               RECT 27.894 47.158 27.946 47.194 ;
               RECT 27.894 48.358 27.946 48.394 ;
               RECT 27.894 50.142 27.946 50.178 ;
               RECT 27.894 50.382 27.946 50.418 ;
               RECT 27.894 54.702 27.946 54.738 ;
               RECT 27.894 54.942 27.946 54.978 ;
               RECT 27.894 57.478 27.946 57.514 ;
               RECT 27.894 58.678 27.946 58.714 ;
               RECT 27.894 59.878 27.946 59.914 ;
               RECT 27.894 61.078 27.946 61.114 ;
               RECT 27.894 62.278 27.946 62.314 ;
               RECT 27.894 63.478 27.946 63.514 ;
               RECT 27.894 64.678 27.946 64.714 ;
               RECT 27.894 65.878 27.946 65.914 ;
               RECT 27.894 67.078 27.946 67.114 ;
               RECT 27.894 68.278 27.946 68.314 ;
               RECT 27.894 69.478 27.946 69.514 ;
               RECT 27.894 70.678 27.946 70.714 ;
               RECT 27.894 71.878 27.946 71.914 ;
               RECT 27.894 73.078 27.946 73.114 ;
               RECT 27.894 74.278 27.946 74.314 ;
               RECT 27.894 75.478 27.946 75.514 ;
               RECT 27.894 76.678 27.946 76.714 ;
               RECT 27.894 77.878 27.946 77.914 ;
               RECT 27.894 79.078 27.946 79.114 ;
               RECT 27.894 80.278 27.946 80.314 ;
               RECT 27.894 81.478 27.946 81.514 ;
               RECT 27.894 82.678 27.946 82.714 ;
               RECT 27.894 83.878 27.946 83.914 ;
               RECT 27.894 85.078 27.946 85.114 ;
               RECT 27.894 86.278 27.946 86.314 ;
               RECT 27.894 87.478 27.946 87.514 ;
               RECT 27.894 88.678 27.946 88.714 ;
               RECT 27.894 89.878 27.946 89.914 ;
               RECT 27.894 91.078 27.946 91.114 ;
               RECT 27.894 92.278 27.946 92.314 ;
               RECT 27.894 93.478 27.946 93.514 ;
               RECT 27.894 94.678 27.946 94.714 ;
               RECT 27.894 95.878 27.946 95.914 ;
               RECT 27.894 97.078 27.946 97.114 ;
               RECT 27.894 98.278 27.946 98.314 ;
               RECT 27.894 99.478 27.946 99.514 ;
               RECT 27.894 100.678 27.946 100.714 ;
               RECT 27.894 101.878 27.946 101.914 ;
               RECT 27.894 103.078 27.946 103.114 ;
               RECT 27.894 104.278 27.946 104.314 ;
               RECT 27.974 0.281 28.026 0.317 ;
               RECT 27.974 104.803 28.026 104.839 ;
               RECT 28.054 0.806 28.106 0.842 ;
               RECT 28.054 2.006 28.106 2.042 ;
               RECT 28.054 3.206 28.106 3.242 ;
               RECT 28.054 4.406 28.106 4.442 ;
               RECT 28.054 5.606 28.106 5.642 ;
               RECT 28.054 6.806 28.106 6.842 ;
               RECT 28.054 8.006 28.106 8.042 ;
               RECT 28.054 9.206 28.106 9.242 ;
               RECT 28.054 10.406 28.106 10.442 ;
               RECT 28.054 11.606 28.106 11.642 ;
               RECT 28.054 12.806 28.106 12.842 ;
               RECT 28.054 14.006 28.106 14.042 ;
               RECT 28.054 15.206 28.106 15.242 ;
               RECT 28.054 16.406 28.106 16.442 ;
               RECT 28.054 17.606 28.106 17.642 ;
               RECT 28.054 18.806 28.106 18.842 ;
               RECT 28.054 20.006 28.106 20.042 ;
               RECT 28.054 21.206 28.106 21.242 ;
               RECT 28.054 22.406 28.106 22.442 ;
               RECT 28.054 23.606 28.106 23.642 ;
               RECT 28.054 24.806 28.106 24.842 ;
               RECT 28.054 26.006 28.106 26.042 ;
               RECT 28.054 27.206 28.106 27.242 ;
               RECT 28.054 28.406 28.106 28.442 ;
               RECT 28.054 29.606 28.106 29.642 ;
               RECT 28.054 30.806 28.106 30.842 ;
               RECT 28.054 32.006 28.106 32.042 ;
               RECT 28.054 33.206 28.106 33.242 ;
               RECT 28.054 34.406 28.106 34.442 ;
               RECT 28.054 35.606 28.106 35.642 ;
               RECT 28.054 36.806 28.106 36.842 ;
               RECT 28.054 38.006 28.106 38.042 ;
               RECT 28.054 39.206 28.106 39.242 ;
               RECT 28.054 40.406 28.106 40.442 ;
               RECT 28.054 41.606 28.106 41.642 ;
               RECT 28.054 42.806 28.106 42.842 ;
               RECT 28.054 44.006 28.106 44.042 ;
               RECT 28.054 45.206 28.106 45.242 ;
               RECT 28.054 46.406 28.106 46.442 ;
               RECT 28.054 47.606 28.106 47.642 ;
               RECT 28.054 49.422 28.106 49.458 ;
               RECT 28.054 49.662 28.106 49.698 ;
               RECT 28.054 51.102 28.106 51.138 ;
               RECT 28.054 51.582 28.106 51.618 ;
               RECT 28.054 53.502 28.106 53.538 ;
               RECT 28.054 53.982 28.106 54.018 ;
               RECT 28.054 55.422 28.106 55.458 ;
               RECT 28.054 55.662 28.106 55.698 ;
               RECT 28.054 56.726 28.106 56.762 ;
               RECT 28.054 57.926 28.106 57.962 ;
               RECT 28.054 59.126 28.106 59.162 ;
               RECT 28.054 60.326 28.106 60.362 ;
               RECT 28.054 61.526 28.106 61.562 ;
               RECT 28.054 62.726 28.106 62.762 ;
               RECT 28.054 63.926 28.106 63.962 ;
               RECT 28.054 65.126 28.106 65.162 ;
               RECT 28.054 66.326 28.106 66.362 ;
               RECT 28.054 67.526 28.106 67.562 ;
               RECT 28.054 68.726 28.106 68.762 ;
               RECT 28.054 69.926 28.106 69.962 ;
               RECT 28.054 71.126 28.106 71.162 ;
               RECT 28.054 72.326 28.106 72.362 ;
               RECT 28.054 73.526 28.106 73.562 ;
               RECT 28.054 74.726 28.106 74.762 ;
               RECT 28.054 75.926 28.106 75.962 ;
               RECT 28.054 77.126 28.106 77.162 ;
               RECT 28.054 78.326 28.106 78.362 ;
               RECT 28.054 79.526 28.106 79.562 ;
               RECT 28.054 80.726 28.106 80.762 ;
               RECT 28.054 81.926 28.106 81.962 ;
               RECT 28.054 83.126 28.106 83.162 ;
               RECT 28.054 84.326 28.106 84.362 ;
               RECT 28.054 85.526 28.106 85.562 ;
               RECT 28.054 86.726 28.106 86.762 ;
               RECT 28.054 87.926 28.106 87.962 ;
               RECT 28.054 89.126 28.106 89.162 ;
               RECT 28.054 90.326 28.106 90.362 ;
               RECT 28.054 91.526 28.106 91.562 ;
               RECT 28.054 92.726 28.106 92.762 ;
               RECT 28.054 93.926 28.106 93.962 ;
               RECT 28.054 95.126 28.106 95.162 ;
               RECT 28.054 96.326 28.106 96.362 ;
               RECT 28.054 97.526 28.106 97.562 ;
               RECT 28.054 98.726 28.106 98.762 ;
               RECT 28.054 99.926 28.106 99.962 ;
               RECT 28.054 101.126 28.106 101.162 ;
               RECT 28.054 102.326 28.106 102.362 ;
               RECT 28.054 103.526 28.106 103.562 ;
               RECT 28.134 1.558 28.186 1.594 ;
               RECT 28.134 2.758 28.186 2.794 ;
               RECT 28.134 3.958 28.186 3.994 ;
               RECT 28.134 5.158 28.186 5.194 ;
               RECT 28.134 6.358 28.186 6.394 ;
               RECT 28.134 7.558 28.186 7.594 ;
               RECT 28.134 8.758 28.186 8.794 ;
               RECT 28.134 9.958 28.186 9.994 ;
               RECT 28.134 11.158 28.186 11.194 ;
               RECT 28.134 12.358 28.186 12.394 ;
               RECT 28.134 13.558 28.186 13.594 ;
               RECT 28.134 14.758 28.186 14.794 ;
               RECT 28.134 15.958 28.186 15.994 ;
               RECT 28.134 17.158 28.186 17.194 ;
               RECT 28.134 18.358 28.186 18.394 ;
               RECT 28.134 19.558 28.186 19.594 ;
               RECT 28.134 20.758 28.186 20.794 ;
               RECT 28.134 21.958 28.186 21.994 ;
               RECT 28.134 23.158 28.186 23.194 ;
               RECT 28.134 24.358 28.186 24.394 ;
               RECT 28.134 25.558 28.186 25.594 ;
               RECT 28.134 26.758 28.186 26.794 ;
               RECT 28.134 27.958 28.186 27.994 ;
               RECT 28.134 29.158 28.186 29.194 ;
               RECT 28.134 30.358 28.186 30.394 ;
               RECT 28.134 31.558 28.186 31.594 ;
               RECT 28.134 32.758 28.186 32.794 ;
               RECT 28.134 33.958 28.186 33.994 ;
               RECT 28.134 35.158 28.186 35.194 ;
               RECT 28.134 36.358 28.186 36.394 ;
               RECT 28.134 37.558 28.186 37.594 ;
               RECT 28.134 38.758 28.186 38.794 ;
               RECT 28.134 39.958 28.186 39.994 ;
               RECT 28.134 41.158 28.186 41.194 ;
               RECT 28.134 42.358 28.186 42.394 ;
               RECT 28.134 43.558 28.186 43.594 ;
               RECT 28.134 44.758 28.186 44.794 ;
               RECT 28.134 45.958 28.186 45.994 ;
               RECT 28.134 47.158 28.186 47.194 ;
               RECT 28.134 48.358 28.186 48.394 ;
               RECT 28.134 50.142 28.186 50.178 ;
               RECT 28.134 50.382 28.186 50.418 ;
               RECT 28.134 54.702 28.186 54.738 ;
               RECT 28.134 54.942 28.186 54.978 ;
               RECT 28.134 57.478 28.186 57.514 ;
               RECT 28.134 58.678 28.186 58.714 ;
               RECT 28.134 59.878 28.186 59.914 ;
               RECT 28.134 61.078 28.186 61.114 ;
               RECT 28.134 62.278 28.186 62.314 ;
               RECT 28.134 63.478 28.186 63.514 ;
               RECT 28.134 64.678 28.186 64.714 ;
               RECT 28.134 65.878 28.186 65.914 ;
               RECT 28.134 67.078 28.186 67.114 ;
               RECT 28.134 68.278 28.186 68.314 ;
               RECT 28.134 69.478 28.186 69.514 ;
               RECT 28.134 70.678 28.186 70.714 ;
               RECT 28.134 71.878 28.186 71.914 ;
               RECT 28.134 73.078 28.186 73.114 ;
               RECT 28.134 74.278 28.186 74.314 ;
               RECT 28.134 75.478 28.186 75.514 ;
               RECT 28.134 76.678 28.186 76.714 ;
               RECT 28.134 77.878 28.186 77.914 ;
               RECT 28.134 79.078 28.186 79.114 ;
               RECT 28.134 80.278 28.186 80.314 ;
               RECT 28.134 81.478 28.186 81.514 ;
               RECT 28.134 82.678 28.186 82.714 ;
               RECT 28.134 83.878 28.186 83.914 ;
               RECT 28.134 85.078 28.186 85.114 ;
               RECT 28.134 86.278 28.186 86.314 ;
               RECT 28.134 87.478 28.186 87.514 ;
               RECT 28.134 88.678 28.186 88.714 ;
               RECT 28.134 89.878 28.186 89.914 ;
               RECT 28.134 91.078 28.186 91.114 ;
               RECT 28.134 92.278 28.186 92.314 ;
               RECT 28.134 93.478 28.186 93.514 ;
               RECT 28.134 94.678 28.186 94.714 ;
               RECT 28.134 95.878 28.186 95.914 ;
               RECT 28.134 97.078 28.186 97.114 ;
               RECT 28.134 98.278 28.186 98.314 ;
               RECT 28.134 99.478 28.186 99.514 ;
               RECT 28.134 100.678 28.186 100.714 ;
               RECT 28.134 101.878 28.186 101.914 ;
               RECT 28.134 103.078 28.186 103.114 ;
               RECT 28.134 104.278 28.186 104.314 ;
               RECT 28.214 0.806 28.266 0.842 ;
               RECT 28.214 2.006 28.266 2.042 ;
               RECT 28.214 3.206 28.266 3.242 ;
               RECT 28.214 4.406 28.266 4.442 ;
               RECT 28.214 5.606 28.266 5.642 ;
               RECT 28.214 6.806 28.266 6.842 ;
               RECT 28.214 8.006 28.266 8.042 ;
               RECT 28.214 9.206 28.266 9.242 ;
               RECT 28.214 10.406 28.266 10.442 ;
               RECT 28.214 11.606 28.266 11.642 ;
               RECT 28.214 12.806 28.266 12.842 ;
               RECT 28.214 14.006 28.266 14.042 ;
               RECT 28.214 15.206 28.266 15.242 ;
               RECT 28.214 16.406 28.266 16.442 ;
               RECT 28.214 17.606 28.266 17.642 ;
               RECT 28.214 18.806 28.266 18.842 ;
               RECT 28.214 20.006 28.266 20.042 ;
               RECT 28.214 21.206 28.266 21.242 ;
               RECT 28.214 22.406 28.266 22.442 ;
               RECT 28.214 23.606 28.266 23.642 ;
               RECT 28.214 24.806 28.266 24.842 ;
               RECT 28.214 26.006 28.266 26.042 ;
               RECT 28.214 27.206 28.266 27.242 ;
               RECT 28.214 28.406 28.266 28.442 ;
               RECT 28.214 29.606 28.266 29.642 ;
               RECT 28.214 30.806 28.266 30.842 ;
               RECT 28.214 32.006 28.266 32.042 ;
               RECT 28.214 33.206 28.266 33.242 ;
               RECT 28.214 34.406 28.266 34.442 ;
               RECT 28.214 35.606 28.266 35.642 ;
               RECT 28.214 36.806 28.266 36.842 ;
               RECT 28.214 38.006 28.266 38.042 ;
               RECT 28.214 39.206 28.266 39.242 ;
               RECT 28.214 40.406 28.266 40.442 ;
               RECT 28.214 41.606 28.266 41.642 ;
               RECT 28.214 42.806 28.266 42.842 ;
               RECT 28.214 44.006 28.266 44.042 ;
               RECT 28.214 45.206 28.266 45.242 ;
               RECT 28.214 46.406 28.266 46.442 ;
               RECT 28.214 47.606 28.266 47.642 ;
               RECT 28.214 49.422 28.266 49.458 ;
               RECT 28.214 49.662 28.266 49.698 ;
               RECT 28.214 55.422 28.266 55.458 ;
               RECT 28.214 55.662 28.266 55.698 ;
               RECT 28.214 56.726 28.266 56.762 ;
               RECT 28.214 57.926 28.266 57.962 ;
               RECT 28.214 59.126 28.266 59.162 ;
               RECT 28.214 60.326 28.266 60.362 ;
               RECT 28.214 61.526 28.266 61.562 ;
               RECT 28.214 62.726 28.266 62.762 ;
               RECT 28.214 63.926 28.266 63.962 ;
               RECT 28.214 65.126 28.266 65.162 ;
               RECT 28.214 66.326 28.266 66.362 ;
               RECT 28.214 67.526 28.266 67.562 ;
               RECT 28.214 68.726 28.266 68.762 ;
               RECT 28.214 69.926 28.266 69.962 ;
               RECT 28.214 71.126 28.266 71.162 ;
               RECT 28.214 72.326 28.266 72.362 ;
               RECT 28.214 73.526 28.266 73.562 ;
               RECT 28.214 74.726 28.266 74.762 ;
               RECT 28.214 75.926 28.266 75.962 ;
               RECT 28.214 77.126 28.266 77.162 ;
               RECT 28.214 78.326 28.266 78.362 ;
               RECT 28.214 79.526 28.266 79.562 ;
               RECT 28.214 80.726 28.266 80.762 ;
               RECT 28.214 81.926 28.266 81.962 ;
               RECT 28.214 83.126 28.266 83.162 ;
               RECT 28.214 84.326 28.266 84.362 ;
               RECT 28.214 85.526 28.266 85.562 ;
               RECT 28.214 86.726 28.266 86.762 ;
               RECT 28.214 87.926 28.266 87.962 ;
               RECT 28.214 89.126 28.266 89.162 ;
               RECT 28.214 90.326 28.266 90.362 ;
               RECT 28.214 91.526 28.266 91.562 ;
               RECT 28.214 92.726 28.266 92.762 ;
               RECT 28.214 93.926 28.266 93.962 ;
               RECT 28.214 95.126 28.266 95.162 ;
               RECT 28.214 96.326 28.266 96.362 ;
               RECT 28.214 97.526 28.266 97.562 ;
               RECT 28.214 98.726 28.266 98.762 ;
               RECT 28.214 99.926 28.266 99.962 ;
               RECT 28.214 101.126 28.266 101.162 ;
               RECT 28.214 102.326 28.266 102.362 ;
               RECT 28.214 103.526 28.266 103.562 ;
               RECT 28.294 1.558 28.346 1.594 ;
               RECT 28.294 2.758 28.346 2.794 ;
               RECT 28.294 3.958 28.346 3.994 ;
               RECT 28.294 5.158 28.346 5.194 ;
               RECT 28.294 6.358 28.346 6.394 ;
               RECT 28.294 7.558 28.346 7.594 ;
               RECT 28.294 8.758 28.346 8.794 ;
               RECT 28.294 9.958 28.346 9.994 ;
               RECT 28.294 11.158 28.346 11.194 ;
               RECT 28.294 12.358 28.346 12.394 ;
               RECT 28.294 13.558 28.346 13.594 ;
               RECT 28.294 14.758 28.346 14.794 ;
               RECT 28.294 15.958 28.346 15.994 ;
               RECT 28.294 17.158 28.346 17.194 ;
               RECT 28.294 18.358 28.346 18.394 ;
               RECT 28.294 19.558 28.346 19.594 ;
               RECT 28.294 20.758 28.346 20.794 ;
               RECT 28.294 21.958 28.346 21.994 ;
               RECT 28.294 23.158 28.346 23.194 ;
               RECT 28.294 24.358 28.346 24.394 ;
               RECT 28.294 25.558 28.346 25.594 ;
               RECT 28.294 26.758 28.346 26.794 ;
               RECT 28.294 27.958 28.346 27.994 ;
               RECT 28.294 29.158 28.346 29.194 ;
               RECT 28.294 30.358 28.346 30.394 ;
               RECT 28.294 31.558 28.346 31.594 ;
               RECT 28.294 32.758 28.346 32.794 ;
               RECT 28.294 33.958 28.346 33.994 ;
               RECT 28.294 35.158 28.346 35.194 ;
               RECT 28.294 36.358 28.346 36.394 ;
               RECT 28.294 37.558 28.346 37.594 ;
               RECT 28.294 38.758 28.346 38.794 ;
               RECT 28.294 39.958 28.346 39.994 ;
               RECT 28.294 41.158 28.346 41.194 ;
               RECT 28.294 42.358 28.346 42.394 ;
               RECT 28.294 43.558 28.346 43.594 ;
               RECT 28.294 44.758 28.346 44.794 ;
               RECT 28.294 45.958 28.346 45.994 ;
               RECT 28.294 47.158 28.346 47.194 ;
               RECT 28.294 48.358 28.346 48.394 ;
               RECT 28.294 50.142 28.346 50.178 ;
               RECT 28.294 50.382 28.346 50.418 ;
               RECT 28.294 54.702 28.346 54.738 ;
               RECT 28.294 54.942 28.346 54.978 ;
               RECT 28.294 57.478 28.346 57.514 ;
               RECT 28.294 58.678 28.346 58.714 ;
               RECT 28.294 59.878 28.346 59.914 ;
               RECT 28.294 61.078 28.346 61.114 ;
               RECT 28.294 62.278 28.346 62.314 ;
               RECT 28.294 63.478 28.346 63.514 ;
               RECT 28.294 64.678 28.346 64.714 ;
               RECT 28.294 65.878 28.346 65.914 ;
               RECT 28.294 67.078 28.346 67.114 ;
               RECT 28.294 68.278 28.346 68.314 ;
               RECT 28.294 69.478 28.346 69.514 ;
               RECT 28.294 70.678 28.346 70.714 ;
               RECT 28.294 71.878 28.346 71.914 ;
               RECT 28.294 73.078 28.346 73.114 ;
               RECT 28.294 74.278 28.346 74.314 ;
               RECT 28.294 75.478 28.346 75.514 ;
               RECT 28.294 76.678 28.346 76.714 ;
               RECT 28.294 77.878 28.346 77.914 ;
               RECT 28.294 79.078 28.346 79.114 ;
               RECT 28.294 80.278 28.346 80.314 ;
               RECT 28.294 81.478 28.346 81.514 ;
               RECT 28.294 82.678 28.346 82.714 ;
               RECT 28.294 83.878 28.346 83.914 ;
               RECT 28.294 85.078 28.346 85.114 ;
               RECT 28.294 86.278 28.346 86.314 ;
               RECT 28.294 87.478 28.346 87.514 ;
               RECT 28.294 88.678 28.346 88.714 ;
               RECT 28.294 89.878 28.346 89.914 ;
               RECT 28.294 91.078 28.346 91.114 ;
               RECT 28.294 92.278 28.346 92.314 ;
               RECT 28.294 93.478 28.346 93.514 ;
               RECT 28.294 94.678 28.346 94.714 ;
               RECT 28.294 95.878 28.346 95.914 ;
               RECT 28.294 97.078 28.346 97.114 ;
               RECT 28.294 98.278 28.346 98.314 ;
               RECT 28.294 99.478 28.346 99.514 ;
               RECT 28.294 100.678 28.346 100.714 ;
               RECT 28.294 101.878 28.346 101.914 ;
               RECT 28.294 103.078 28.346 103.114 ;
               RECT 28.294 104.278 28.346 104.314 ;
               RECT 28.374 0.281 28.426 0.317 ;
               RECT 28.374 104.803 28.426 104.839 ;
               RECT 28.454 0.806 28.506 0.842 ;
               RECT 28.454 2.006 28.506 2.042 ;
               RECT 28.454 3.206 28.506 3.242 ;
               RECT 28.454 4.406 28.506 4.442 ;
               RECT 28.454 5.606 28.506 5.642 ;
               RECT 28.454 6.806 28.506 6.842 ;
               RECT 28.454 8.006 28.506 8.042 ;
               RECT 28.454 9.206 28.506 9.242 ;
               RECT 28.454 10.406 28.506 10.442 ;
               RECT 28.454 11.606 28.506 11.642 ;
               RECT 28.454 12.806 28.506 12.842 ;
               RECT 28.454 14.006 28.506 14.042 ;
               RECT 28.454 15.206 28.506 15.242 ;
               RECT 28.454 16.406 28.506 16.442 ;
               RECT 28.454 17.606 28.506 17.642 ;
               RECT 28.454 18.806 28.506 18.842 ;
               RECT 28.454 20.006 28.506 20.042 ;
               RECT 28.454 21.206 28.506 21.242 ;
               RECT 28.454 22.406 28.506 22.442 ;
               RECT 28.454 23.606 28.506 23.642 ;
               RECT 28.454 24.806 28.506 24.842 ;
               RECT 28.454 26.006 28.506 26.042 ;
               RECT 28.454 27.206 28.506 27.242 ;
               RECT 28.454 28.406 28.506 28.442 ;
               RECT 28.454 29.606 28.506 29.642 ;
               RECT 28.454 30.806 28.506 30.842 ;
               RECT 28.454 32.006 28.506 32.042 ;
               RECT 28.454 33.206 28.506 33.242 ;
               RECT 28.454 34.406 28.506 34.442 ;
               RECT 28.454 35.606 28.506 35.642 ;
               RECT 28.454 36.806 28.506 36.842 ;
               RECT 28.454 38.006 28.506 38.042 ;
               RECT 28.454 39.206 28.506 39.242 ;
               RECT 28.454 40.406 28.506 40.442 ;
               RECT 28.454 41.606 28.506 41.642 ;
               RECT 28.454 42.806 28.506 42.842 ;
               RECT 28.454 44.006 28.506 44.042 ;
               RECT 28.454 45.206 28.506 45.242 ;
               RECT 28.454 46.406 28.506 46.442 ;
               RECT 28.454 47.606 28.506 47.642 ;
               RECT 28.454 49.422 28.506 49.458 ;
               RECT 28.454 49.662 28.506 49.698 ;
               RECT 28.454 55.422 28.506 55.458 ;
               RECT 28.454 55.662 28.506 55.698 ;
               RECT 28.454 56.726 28.506 56.762 ;
               RECT 28.454 57.926 28.506 57.962 ;
               RECT 28.454 59.126 28.506 59.162 ;
               RECT 28.454 60.326 28.506 60.362 ;
               RECT 28.454 61.526 28.506 61.562 ;
               RECT 28.454 62.726 28.506 62.762 ;
               RECT 28.454 63.926 28.506 63.962 ;
               RECT 28.454 65.126 28.506 65.162 ;
               RECT 28.454 66.326 28.506 66.362 ;
               RECT 28.454 67.526 28.506 67.562 ;
               RECT 28.454 68.726 28.506 68.762 ;
               RECT 28.454 69.926 28.506 69.962 ;
               RECT 28.454 71.126 28.506 71.162 ;
               RECT 28.454 72.326 28.506 72.362 ;
               RECT 28.454 73.526 28.506 73.562 ;
               RECT 28.454 74.726 28.506 74.762 ;
               RECT 28.454 75.926 28.506 75.962 ;
               RECT 28.454 77.126 28.506 77.162 ;
               RECT 28.454 78.326 28.506 78.362 ;
               RECT 28.454 79.526 28.506 79.562 ;
               RECT 28.454 80.726 28.506 80.762 ;
               RECT 28.454 81.926 28.506 81.962 ;
               RECT 28.454 83.126 28.506 83.162 ;
               RECT 28.454 84.326 28.506 84.362 ;
               RECT 28.454 85.526 28.506 85.562 ;
               RECT 28.454 86.726 28.506 86.762 ;
               RECT 28.454 87.926 28.506 87.962 ;
               RECT 28.454 89.126 28.506 89.162 ;
               RECT 28.454 90.326 28.506 90.362 ;
               RECT 28.454 91.526 28.506 91.562 ;
               RECT 28.454 92.726 28.506 92.762 ;
               RECT 28.454 93.926 28.506 93.962 ;
               RECT 28.454 95.126 28.506 95.162 ;
               RECT 28.454 96.326 28.506 96.362 ;
               RECT 28.454 97.526 28.506 97.562 ;
               RECT 28.454 98.726 28.506 98.762 ;
               RECT 28.454 99.926 28.506 99.962 ;
               RECT 28.454 101.126 28.506 101.162 ;
               RECT 28.454 102.326 28.506 102.362 ;
               RECT 28.454 103.526 28.506 103.562 ;
               RECT 28.534 1.558 28.586 1.594 ;
               RECT 28.534 2.758 28.586 2.794 ;
               RECT 28.534 3.958 28.586 3.994 ;
               RECT 28.534 5.158 28.586 5.194 ;
               RECT 28.534 6.358 28.586 6.394 ;
               RECT 28.534 7.558 28.586 7.594 ;
               RECT 28.534 8.758 28.586 8.794 ;
               RECT 28.534 9.958 28.586 9.994 ;
               RECT 28.534 11.158 28.586 11.194 ;
               RECT 28.534 12.358 28.586 12.394 ;
               RECT 28.534 13.558 28.586 13.594 ;
               RECT 28.534 14.758 28.586 14.794 ;
               RECT 28.534 15.958 28.586 15.994 ;
               RECT 28.534 17.158 28.586 17.194 ;
               RECT 28.534 18.358 28.586 18.394 ;
               RECT 28.534 19.558 28.586 19.594 ;
               RECT 28.534 20.758 28.586 20.794 ;
               RECT 28.534 21.958 28.586 21.994 ;
               RECT 28.534 23.158 28.586 23.194 ;
               RECT 28.534 24.358 28.586 24.394 ;
               RECT 28.534 25.558 28.586 25.594 ;
               RECT 28.534 26.758 28.586 26.794 ;
               RECT 28.534 27.958 28.586 27.994 ;
               RECT 28.534 29.158 28.586 29.194 ;
               RECT 28.534 30.358 28.586 30.394 ;
               RECT 28.534 31.558 28.586 31.594 ;
               RECT 28.534 32.758 28.586 32.794 ;
               RECT 28.534 33.958 28.586 33.994 ;
               RECT 28.534 35.158 28.586 35.194 ;
               RECT 28.534 36.358 28.586 36.394 ;
               RECT 28.534 37.558 28.586 37.594 ;
               RECT 28.534 38.758 28.586 38.794 ;
               RECT 28.534 39.958 28.586 39.994 ;
               RECT 28.534 41.158 28.586 41.194 ;
               RECT 28.534 42.358 28.586 42.394 ;
               RECT 28.534 43.558 28.586 43.594 ;
               RECT 28.534 44.758 28.586 44.794 ;
               RECT 28.534 45.958 28.586 45.994 ;
               RECT 28.534 47.158 28.586 47.194 ;
               RECT 28.534 48.358 28.586 48.394 ;
               RECT 28.534 50.142 28.586 50.178 ;
               RECT 28.534 50.382 28.586 50.418 ;
               RECT 28.534 54.702 28.586 54.738 ;
               RECT 28.534 54.942 28.586 54.978 ;
               RECT 28.534 57.478 28.586 57.514 ;
               RECT 28.534 58.678 28.586 58.714 ;
               RECT 28.534 59.878 28.586 59.914 ;
               RECT 28.534 61.078 28.586 61.114 ;
               RECT 28.534 62.278 28.586 62.314 ;
               RECT 28.534 63.478 28.586 63.514 ;
               RECT 28.534 64.678 28.586 64.714 ;
               RECT 28.534 65.878 28.586 65.914 ;
               RECT 28.534 67.078 28.586 67.114 ;
               RECT 28.534 68.278 28.586 68.314 ;
               RECT 28.534 69.478 28.586 69.514 ;
               RECT 28.534 70.678 28.586 70.714 ;
               RECT 28.534 71.878 28.586 71.914 ;
               RECT 28.534 73.078 28.586 73.114 ;
               RECT 28.534 74.278 28.586 74.314 ;
               RECT 28.534 75.478 28.586 75.514 ;
               RECT 28.534 76.678 28.586 76.714 ;
               RECT 28.534 77.878 28.586 77.914 ;
               RECT 28.534 79.078 28.586 79.114 ;
               RECT 28.534 80.278 28.586 80.314 ;
               RECT 28.534 81.478 28.586 81.514 ;
               RECT 28.534 82.678 28.586 82.714 ;
               RECT 28.534 83.878 28.586 83.914 ;
               RECT 28.534 85.078 28.586 85.114 ;
               RECT 28.534 86.278 28.586 86.314 ;
               RECT 28.534 87.478 28.586 87.514 ;
               RECT 28.534 88.678 28.586 88.714 ;
               RECT 28.534 89.878 28.586 89.914 ;
               RECT 28.534 91.078 28.586 91.114 ;
               RECT 28.534 92.278 28.586 92.314 ;
               RECT 28.534 93.478 28.586 93.514 ;
               RECT 28.534 94.678 28.586 94.714 ;
               RECT 28.534 95.878 28.586 95.914 ;
               RECT 28.534 97.078 28.586 97.114 ;
               RECT 28.534 98.278 28.586 98.314 ;
               RECT 28.534 99.478 28.586 99.514 ;
               RECT 28.534 100.678 28.586 100.714 ;
               RECT 28.534 101.878 28.586 101.914 ;
               RECT 28.534 103.078 28.586 103.114 ;
               RECT 28.534 104.278 28.586 104.314 ;
               RECT 28.614 0.806 28.666 0.842 ;
               RECT 28.614 2.006 28.666 2.042 ;
               RECT 28.614 3.206 28.666 3.242 ;
               RECT 28.614 4.406 28.666 4.442 ;
               RECT 28.614 5.606 28.666 5.642 ;
               RECT 28.614 6.806 28.666 6.842 ;
               RECT 28.614 8.006 28.666 8.042 ;
               RECT 28.614 9.206 28.666 9.242 ;
               RECT 28.614 10.406 28.666 10.442 ;
               RECT 28.614 11.606 28.666 11.642 ;
               RECT 28.614 12.806 28.666 12.842 ;
               RECT 28.614 14.006 28.666 14.042 ;
               RECT 28.614 15.206 28.666 15.242 ;
               RECT 28.614 16.406 28.666 16.442 ;
               RECT 28.614 17.606 28.666 17.642 ;
               RECT 28.614 18.806 28.666 18.842 ;
               RECT 28.614 20.006 28.666 20.042 ;
               RECT 28.614 21.206 28.666 21.242 ;
               RECT 28.614 22.406 28.666 22.442 ;
               RECT 28.614 23.606 28.666 23.642 ;
               RECT 28.614 24.806 28.666 24.842 ;
               RECT 28.614 26.006 28.666 26.042 ;
               RECT 28.614 27.206 28.666 27.242 ;
               RECT 28.614 28.406 28.666 28.442 ;
               RECT 28.614 29.606 28.666 29.642 ;
               RECT 28.614 30.806 28.666 30.842 ;
               RECT 28.614 32.006 28.666 32.042 ;
               RECT 28.614 33.206 28.666 33.242 ;
               RECT 28.614 34.406 28.666 34.442 ;
               RECT 28.614 35.606 28.666 35.642 ;
               RECT 28.614 36.806 28.666 36.842 ;
               RECT 28.614 38.006 28.666 38.042 ;
               RECT 28.614 39.206 28.666 39.242 ;
               RECT 28.614 40.406 28.666 40.442 ;
               RECT 28.614 41.606 28.666 41.642 ;
               RECT 28.614 42.806 28.666 42.842 ;
               RECT 28.614 44.006 28.666 44.042 ;
               RECT 28.614 45.206 28.666 45.242 ;
               RECT 28.614 46.406 28.666 46.442 ;
               RECT 28.614 47.606 28.666 47.642 ;
               RECT 28.614 49.422 28.666 49.458 ;
               RECT 28.614 49.662 28.666 49.698 ;
               RECT 28.614 55.422 28.666 55.458 ;
               RECT 28.614 55.662 28.666 55.698 ;
               RECT 28.614 56.726 28.666 56.762 ;
               RECT 28.614 57.926 28.666 57.962 ;
               RECT 28.614 59.126 28.666 59.162 ;
               RECT 28.614 60.326 28.666 60.362 ;
               RECT 28.614 61.526 28.666 61.562 ;
               RECT 28.614 62.726 28.666 62.762 ;
               RECT 28.614 63.926 28.666 63.962 ;
               RECT 28.614 65.126 28.666 65.162 ;
               RECT 28.614 66.326 28.666 66.362 ;
               RECT 28.614 67.526 28.666 67.562 ;
               RECT 28.614 68.726 28.666 68.762 ;
               RECT 28.614 69.926 28.666 69.962 ;
               RECT 28.614 71.126 28.666 71.162 ;
               RECT 28.614 72.326 28.666 72.362 ;
               RECT 28.614 73.526 28.666 73.562 ;
               RECT 28.614 74.726 28.666 74.762 ;
               RECT 28.614 75.926 28.666 75.962 ;
               RECT 28.614 77.126 28.666 77.162 ;
               RECT 28.614 78.326 28.666 78.362 ;
               RECT 28.614 79.526 28.666 79.562 ;
               RECT 28.614 80.726 28.666 80.762 ;
               RECT 28.614 81.926 28.666 81.962 ;
               RECT 28.614 83.126 28.666 83.162 ;
               RECT 28.614 84.326 28.666 84.362 ;
               RECT 28.614 85.526 28.666 85.562 ;
               RECT 28.614 86.726 28.666 86.762 ;
               RECT 28.614 87.926 28.666 87.962 ;
               RECT 28.614 89.126 28.666 89.162 ;
               RECT 28.614 90.326 28.666 90.362 ;
               RECT 28.614 91.526 28.666 91.562 ;
               RECT 28.614 92.726 28.666 92.762 ;
               RECT 28.614 93.926 28.666 93.962 ;
               RECT 28.614 95.126 28.666 95.162 ;
               RECT 28.614 96.326 28.666 96.362 ;
               RECT 28.614 97.526 28.666 97.562 ;
               RECT 28.614 98.726 28.666 98.762 ;
               RECT 28.614 99.926 28.666 99.962 ;
               RECT 28.614 101.126 28.666 101.162 ;
               RECT 28.614 102.326 28.666 102.362 ;
               RECT 28.614 103.526 28.666 103.562 ;
               RECT 28.694 1.558 28.746 1.594 ;
               RECT 28.694 2.758 28.746 2.794 ;
               RECT 28.694 3.958 28.746 3.994 ;
               RECT 28.694 5.158 28.746 5.194 ;
               RECT 28.694 6.358 28.746 6.394 ;
               RECT 28.694 7.558 28.746 7.594 ;
               RECT 28.694 8.758 28.746 8.794 ;
               RECT 28.694 9.958 28.746 9.994 ;
               RECT 28.694 11.158 28.746 11.194 ;
               RECT 28.694 12.358 28.746 12.394 ;
               RECT 28.694 13.558 28.746 13.594 ;
               RECT 28.694 14.758 28.746 14.794 ;
               RECT 28.694 15.958 28.746 15.994 ;
               RECT 28.694 17.158 28.746 17.194 ;
               RECT 28.694 18.358 28.746 18.394 ;
               RECT 28.694 19.558 28.746 19.594 ;
               RECT 28.694 20.758 28.746 20.794 ;
               RECT 28.694 21.958 28.746 21.994 ;
               RECT 28.694 23.158 28.746 23.194 ;
               RECT 28.694 24.358 28.746 24.394 ;
               RECT 28.694 25.558 28.746 25.594 ;
               RECT 28.694 26.758 28.746 26.794 ;
               RECT 28.694 27.958 28.746 27.994 ;
               RECT 28.694 29.158 28.746 29.194 ;
               RECT 28.694 30.358 28.746 30.394 ;
               RECT 28.694 31.558 28.746 31.594 ;
               RECT 28.694 32.758 28.746 32.794 ;
               RECT 28.694 33.958 28.746 33.994 ;
               RECT 28.694 35.158 28.746 35.194 ;
               RECT 28.694 36.358 28.746 36.394 ;
               RECT 28.694 37.558 28.746 37.594 ;
               RECT 28.694 38.758 28.746 38.794 ;
               RECT 28.694 39.958 28.746 39.994 ;
               RECT 28.694 41.158 28.746 41.194 ;
               RECT 28.694 42.358 28.746 42.394 ;
               RECT 28.694 43.558 28.746 43.594 ;
               RECT 28.694 44.758 28.746 44.794 ;
               RECT 28.694 45.958 28.746 45.994 ;
               RECT 28.694 47.158 28.746 47.194 ;
               RECT 28.694 48.358 28.746 48.394 ;
               RECT 28.694 50.142 28.746 50.178 ;
               RECT 28.694 50.382 28.746 50.418 ;
               RECT 28.694 54.702 28.746 54.738 ;
               RECT 28.694 54.942 28.746 54.978 ;
               RECT 28.694 57.478 28.746 57.514 ;
               RECT 28.694 58.678 28.746 58.714 ;
               RECT 28.694 59.878 28.746 59.914 ;
               RECT 28.694 61.078 28.746 61.114 ;
               RECT 28.694 62.278 28.746 62.314 ;
               RECT 28.694 63.478 28.746 63.514 ;
               RECT 28.694 64.678 28.746 64.714 ;
               RECT 28.694 65.878 28.746 65.914 ;
               RECT 28.694 67.078 28.746 67.114 ;
               RECT 28.694 68.278 28.746 68.314 ;
               RECT 28.694 69.478 28.746 69.514 ;
               RECT 28.694 70.678 28.746 70.714 ;
               RECT 28.694 71.878 28.746 71.914 ;
               RECT 28.694 73.078 28.746 73.114 ;
               RECT 28.694 74.278 28.746 74.314 ;
               RECT 28.694 75.478 28.746 75.514 ;
               RECT 28.694 76.678 28.746 76.714 ;
               RECT 28.694 77.878 28.746 77.914 ;
               RECT 28.694 79.078 28.746 79.114 ;
               RECT 28.694 80.278 28.746 80.314 ;
               RECT 28.694 81.478 28.746 81.514 ;
               RECT 28.694 82.678 28.746 82.714 ;
               RECT 28.694 83.878 28.746 83.914 ;
               RECT 28.694 85.078 28.746 85.114 ;
               RECT 28.694 86.278 28.746 86.314 ;
               RECT 28.694 87.478 28.746 87.514 ;
               RECT 28.694 88.678 28.746 88.714 ;
               RECT 28.694 89.878 28.746 89.914 ;
               RECT 28.694 91.078 28.746 91.114 ;
               RECT 28.694 92.278 28.746 92.314 ;
               RECT 28.694 93.478 28.746 93.514 ;
               RECT 28.694 94.678 28.746 94.714 ;
               RECT 28.694 95.878 28.746 95.914 ;
               RECT 28.694 97.078 28.746 97.114 ;
               RECT 28.694 98.278 28.746 98.314 ;
               RECT 28.694 99.478 28.746 99.514 ;
               RECT 28.694 100.678 28.746 100.714 ;
               RECT 28.694 101.878 28.746 101.914 ;
               RECT 28.694 103.078 28.746 103.114 ;
               RECT 28.694 104.278 28.746 104.314 ;
               RECT 28.774 0.281 28.826 0.317 ;
               RECT 28.774 104.803 28.826 104.839 ;
               RECT 28.854 0.806 28.906 0.842 ;
               RECT 28.854 2.006 28.906 2.042 ;
               RECT 28.854 3.206 28.906 3.242 ;
               RECT 28.854 4.406 28.906 4.442 ;
               RECT 28.854 5.606 28.906 5.642 ;
               RECT 28.854 6.806 28.906 6.842 ;
               RECT 28.854 8.006 28.906 8.042 ;
               RECT 28.854 9.206 28.906 9.242 ;
               RECT 28.854 10.406 28.906 10.442 ;
               RECT 28.854 11.606 28.906 11.642 ;
               RECT 28.854 12.806 28.906 12.842 ;
               RECT 28.854 14.006 28.906 14.042 ;
               RECT 28.854 15.206 28.906 15.242 ;
               RECT 28.854 16.406 28.906 16.442 ;
               RECT 28.854 17.606 28.906 17.642 ;
               RECT 28.854 18.806 28.906 18.842 ;
               RECT 28.854 20.006 28.906 20.042 ;
               RECT 28.854 21.206 28.906 21.242 ;
               RECT 28.854 22.406 28.906 22.442 ;
               RECT 28.854 23.606 28.906 23.642 ;
               RECT 28.854 24.806 28.906 24.842 ;
               RECT 28.854 26.006 28.906 26.042 ;
               RECT 28.854 27.206 28.906 27.242 ;
               RECT 28.854 28.406 28.906 28.442 ;
               RECT 28.854 29.606 28.906 29.642 ;
               RECT 28.854 30.806 28.906 30.842 ;
               RECT 28.854 32.006 28.906 32.042 ;
               RECT 28.854 33.206 28.906 33.242 ;
               RECT 28.854 34.406 28.906 34.442 ;
               RECT 28.854 35.606 28.906 35.642 ;
               RECT 28.854 36.806 28.906 36.842 ;
               RECT 28.854 38.006 28.906 38.042 ;
               RECT 28.854 39.206 28.906 39.242 ;
               RECT 28.854 40.406 28.906 40.442 ;
               RECT 28.854 41.606 28.906 41.642 ;
               RECT 28.854 42.806 28.906 42.842 ;
               RECT 28.854 44.006 28.906 44.042 ;
               RECT 28.854 45.206 28.906 45.242 ;
               RECT 28.854 46.406 28.906 46.442 ;
               RECT 28.854 47.606 28.906 47.642 ;
               RECT 28.854 49.422 28.906 49.458 ;
               RECT 28.854 49.662 28.906 49.698 ;
               RECT 28.854 51.102 28.906 51.138 ;
               RECT 28.854 51.582 28.906 51.618 ;
               RECT 28.854 53.502 28.906 53.538 ;
               RECT 28.854 53.982 28.906 54.018 ;
               RECT 28.854 55.422 28.906 55.458 ;
               RECT 28.854 55.662 28.906 55.698 ;
               RECT 28.854 56.726 28.906 56.762 ;
               RECT 28.854 57.926 28.906 57.962 ;
               RECT 28.854 59.126 28.906 59.162 ;
               RECT 28.854 60.326 28.906 60.362 ;
               RECT 28.854 61.526 28.906 61.562 ;
               RECT 28.854 62.726 28.906 62.762 ;
               RECT 28.854 63.926 28.906 63.962 ;
               RECT 28.854 65.126 28.906 65.162 ;
               RECT 28.854 66.326 28.906 66.362 ;
               RECT 28.854 67.526 28.906 67.562 ;
               RECT 28.854 68.726 28.906 68.762 ;
               RECT 28.854 69.926 28.906 69.962 ;
               RECT 28.854 71.126 28.906 71.162 ;
               RECT 28.854 72.326 28.906 72.362 ;
               RECT 28.854 73.526 28.906 73.562 ;
               RECT 28.854 74.726 28.906 74.762 ;
               RECT 28.854 75.926 28.906 75.962 ;
               RECT 28.854 77.126 28.906 77.162 ;
               RECT 28.854 78.326 28.906 78.362 ;
               RECT 28.854 79.526 28.906 79.562 ;
               RECT 28.854 80.726 28.906 80.762 ;
               RECT 28.854 81.926 28.906 81.962 ;
               RECT 28.854 83.126 28.906 83.162 ;
               RECT 28.854 84.326 28.906 84.362 ;
               RECT 28.854 85.526 28.906 85.562 ;
               RECT 28.854 86.726 28.906 86.762 ;
               RECT 28.854 87.926 28.906 87.962 ;
               RECT 28.854 89.126 28.906 89.162 ;
               RECT 28.854 90.326 28.906 90.362 ;
               RECT 28.854 91.526 28.906 91.562 ;
               RECT 28.854 92.726 28.906 92.762 ;
               RECT 28.854 93.926 28.906 93.962 ;
               RECT 28.854 95.126 28.906 95.162 ;
               RECT 28.854 96.326 28.906 96.362 ;
               RECT 28.854 97.526 28.906 97.562 ;
               RECT 28.854 98.726 28.906 98.762 ;
               RECT 28.854 99.926 28.906 99.962 ;
               RECT 28.854 101.126 28.906 101.162 ;
               RECT 28.854 102.326 28.906 102.362 ;
               RECT 28.854 103.526 28.906 103.562 ;
               RECT 28.934 1.558 28.986 1.594 ;
               RECT 28.934 2.758 28.986 2.794 ;
               RECT 28.934 3.958 28.986 3.994 ;
               RECT 28.934 5.158 28.986 5.194 ;
               RECT 28.934 6.358 28.986 6.394 ;
               RECT 28.934 7.558 28.986 7.594 ;
               RECT 28.934 8.758 28.986 8.794 ;
               RECT 28.934 9.958 28.986 9.994 ;
               RECT 28.934 11.158 28.986 11.194 ;
               RECT 28.934 12.358 28.986 12.394 ;
               RECT 28.934 13.558 28.986 13.594 ;
               RECT 28.934 14.758 28.986 14.794 ;
               RECT 28.934 15.958 28.986 15.994 ;
               RECT 28.934 17.158 28.986 17.194 ;
               RECT 28.934 18.358 28.986 18.394 ;
               RECT 28.934 19.558 28.986 19.594 ;
               RECT 28.934 20.758 28.986 20.794 ;
               RECT 28.934 21.958 28.986 21.994 ;
               RECT 28.934 23.158 28.986 23.194 ;
               RECT 28.934 24.358 28.986 24.394 ;
               RECT 28.934 25.558 28.986 25.594 ;
               RECT 28.934 26.758 28.986 26.794 ;
               RECT 28.934 27.958 28.986 27.994 ;
               RECT 28.934 29.158 28.986 29.194 ;
               RECT 28.934 30.358 28.986 30.394 ;
               RECT 28.934 31.558 28.986 31.594 ;
               RECT 28.934 32.758 28.986 32.794 ;
               RECT 28.934 33.958 28.986 33.994 ;
               RECT 28.934 35.158 28.986 35.194 ;
               RECT 28.934 36.358 28.986 36.394 ;
               RECT 28.934 37.558 28.986 37.594 ;
               RECT 28.934 38.758 28.986 38.794 ;
               RECT 28.934 39.958 28.986 39.994 ;
               RECT 28.934 41.158 28.986 41.194 ;
               RECT 28.934 42.358 28.986 42.394 ;
               RECT 28.934 43.558 28.986 43.594 ;
               RECT 28.934 44.758 28.986 44.794 ;
               RECT 28.934 45.958 28.986 45.994 ;
               RECT 28.934 47.158 28.986 47.194 ;
               RECT 28.934 48.358 28.986 48.394 ;
               RECT 28.934 50.142 28.986 50.178 ;
               RECT 28.934 50.382 28.986 50.418 ;
               RECT 28.934 54.702 28.986 54.738 ;
               RECT 28.934 54.942 28.986 54.978 ;
               RECT 28.934 57.478 28.986 57.514 ;
               RECT 28.934 58.678 28.986 58.714 ;
               RECT 28.934 59.878 28.986 59.914 ;
               RECT 28.934 61.078 28.986 61.114 ;
               RECT 28.934 62.278 28.986 62.314 ;
               RECT 28.934 63.478 28.986 63.514 ;
               RECT 28.934 64.678 28.986 64.714 ;
               RECT 28.934 65.878 28.986 65.914 ;
               RECT 28.934 67.078 28.986 67.114 ;
               RECT 28.934 68.278 28.986 68.314 ;
               RECT 28.934 69.478 28.986 69.514 ;
               RECT 28.934 70.678 28.986 70.714 ;
               RECT 28.934 71.878 28.986 71.914 ;
               RECT 28.934 73.078 28.986 73.114 ;
               RECT 28.934 74.278 28.986 74.314 ;
               RECT 28.934 75.478 28.986 75.514 ;
               RECT 28.934 76.678 28.986 76.714 ;
               RECT 28.934 77.878 28.986 77.914 ;
               RECT 28.934 79.078 28.986 79.114 ;
               RECT 28.934 80.278 28.986 80.314 ;
               RECT 28.934 81.478 28.986 81.514 ;
               RECT 28.934 82.678 28.986 82.714 ;
               RECT 28.934 83.878 28.986 83.914 ;
               RECT 28.934 85.078 28.986 85.114 ;
               RECT 28.934 86.278 28.986 86.314 ;
               RECT 28.934 87.478 28.986 87.514 ;
               RECT 28.934 88.678 28.986 88.714 ;
               RECT 28.934 89.878 28.986 89.914 ;
               RECT 28.934 91.078 28.986 91.114 ;
               RECT 28.934 92.278 28.986 92.314 ;
               RECT 28.934 93.478 28.986 93.514 ;
               RECT 28.934 94.678 28.986 94.714 ;
               RECT 28.934 95.878 28.986 95.914 ;
               RECT 28.934 97.078 28.986 97.114 ;
               RECT 28.934 98.278 28.986 98.314 ;
               RECT 28.934 99.478 28.986 99.514 ;
               RECT 28.934 100.678 28.986 100.714 ;
               RECT 28.934 101.878 28.986 101.914 ;
               RECT 28.934 103.078 28.986 103.114 ;
               RECT 28.934 104.278 28.986 104.314 ;
               RECT 29.014 0.806 29.066 0.842 ;
               RECT 29.014 2.006 29.066 2.042 ;
               RECT 29.014 3.206 29.066 3.242 ;
               RECT 29.014 4.406 29.066 4.442 ;
               RECT 29.014 5.606 29.066 5.642 ;
               RECT 29.014 6.806 29.066 6.842 ;
               RECT 29.014 8.006 29.066 8.042 ;
               RECT 29.014 9.206 29.066 9.242 ;
               RECT 29.014 10.406 29.066 10.442 ;
               RECT 29.014 11.606 29.066 11.642 ;
               RECT 29.014 12.806 29.066 12.842 ;
               RECT 29.014 14.006 29.066 14.042 ;
               RECT 29.014 15.206 29.066 15.242 ;
               RECT 29.014 16.406 29.066 16.442 ;
               RECT 29.014 17.606 29.066 17.642 ;
               RECT 29.014 18.806 29.066 18.842 ;
               RECT 29.014 20.006 29.066 20.042 ;
               RECT 29.014 21.206 29.066 21.242 ;
               RECT 29.014 22.406 29.066 22.442 ;
               RECT 29.014 23.606 29.066 23.642 ;
               RECT 29.014 24.806 29.066 24.842 ;
               RECT 29.014 26.006 29.066 26.042 ;
               RECT 29.014 27.206 29.066 27.242 ;
               RECT 29.014 28.406 29.066 28.442 ;
               RECT 29.014 29.606 29.066 29.642 ;
               RECT 29.014 30.806 29.066 30.842 ;
               RECT 29.014 32.006 29.066 32.042 ;
               RECT 29.014 33.206 29.066 33.242 ;
               RECT 29.014 34.406 29.066 34.442 ;
               RECT 29.014 35.606 29.066 35.642 ;
               RECT 29.014 36.806 29.066 36.842 ;
               RECT 29.014 38.006 29.066 38.042 ;
               RECT 29.014 39.206 29.066 39.242 ;
               RECT 29.014 40.406 29.066 40.442 ;
               RECT 29.014 41.606 29.066 41.642 ;
               RECT 29.014 42.806 29.066 42.842 ;
               RECT 29.014 44.006 29.066 44.042 ;
               RECT 29.014 45.206 29.066 45.242 ;
               RECT 29.014 46.406 29.066 46.442 ;
               RECT 29.014 47.606 29.066 47.642 ;
               RECT 29.014 49.422 29.066 49.458 ;
               RECT 29.014 49.662 29.066 49.698 ;
               RECT 29.014 55.422 29.066 55.458 ;
               RECT 29.014 55.662 29.066 55.698 ;
               RECT 29.014 56.726 29.066 56.762 ;
               RECT 29.014 57.926 29.066 57.962 ;
               RECT 29.014 59.126 29.066 59.162 ;
               RECT 29.014 60.326 29.066 60.362 ;
               RECT 29.014 61.526 29.066 61.562 ;
               RECT 29.014 62.726 29.066 62.762 ;
               RECT 29.014 63.926 29.066 63.962 ;
               RECT 29.014 65.126 29.066 65.162 ;
               RECT 29.014 66.326 29.066 66.362 ;
               RECT 29.014 67.526 29.066 67.562 ;
               RECT 29.014 68.726 29.066 68.762 ;
               RECT 29.014 69.926 29.066 69.962 ;
               RECT 29.014 71.126 29.066 71.162 ;
               RECT 29.014 72.326 29.066 72.362 ;
               RECT 29.014 73.526 29.066 73.562 ;
               RECT 29.014 74.726 29.066 74.762 ;
               RECT 29.014 75.926 29.066 75.962 ;
               RECT 29.014 77.126 29.066 77.162 ;
               RECT 29.014 78.326 29.066 78.362 ;
               RECT 29.014 79.526 29.066 79.562 ;
               RECT 29.014 80.726 29.066 80.762 ;
               RECT 29.014 81.926 29.066 81.962 ;
               RECT 29.014 83.126 29.066 83.162 ;
               RECT 29.014 84.326 29.066 84.362 ;
               RECT 29.014 85.526 29.066 85.562 ;
               RECT 29.014 86.726 29.066 86.762 ;
               RECT 29.014 87.926 29.066 87.962 ;
               RECT 29.014 89.126 29.066 89.162 ;
               RECT 29.014 90.326 29.066 90.362 ;
               RECT 29.014 91.526 29.066 91.562 ;
               RECT 29.014 92.726 29.066 92.762 ;
               RECT 29.014 93.926 29.066 93.962 ;
               RECT 29.014 95.126 29.066 95.162 ;
               RECT 29.014 96.326 29.066 96.362 ;
               RECT 29.014 97.526 29.066 97.562 ;
               RECT 29.014 98.726 29.066 98.762 ;
               RECT 29.014 99.926 29.066 99.962 ;
               RECT 29.014 101.126 29.066 101.162 ;
               RECT 29.014 102.326 29.066 102.362 ;
               RECT 29.014 103.526 29.066 103.562 ;
               RECT 29.094 1.558 29.146 1.594 ;
               RECT 29.094 2.758 29.146 2.794 ;
               RECT 29.094 3.958 29.146 3.994 ;
               RECT 29.094 5.158 29.146 5.194 ;
               RECT 29.094 6.358 29.146 6.394 ;
               RECT 29.094 7.558 29.146 7.594 ;
               RECT 29.094 8.758 29.146 8.794 ;
               RECT 29.094 9.958 29.146 9.994 ;
               RECT 29.094 11.158 29.146 11.194 ;
               RECT 29.094 12.358 29.146 12.394 ;
               RECT 29.094 13.558 29.146 13.594 ;
               RECT 29.094 14.758 29.146 14.794 ;
               RECT 29.094 15.958 29.146 15.994 ;
               RECT 29.094 17.158 29.146 17.194 ;
               RECT 29.094 18.358 29.146 18.394 ;
               RECT 29.094 19.558 29.146 19.594 ;
               RECT 29.094 20.758 29.146 20.794 ;
               RECT 29.094 21.958 29.146 21.994 ;
               RECT 29.094 23.158 29.146 23.194 ;
               RECT 29.094 24.358 29.146 24.394 ;
               RECT 29.094 25.558 29.146 25.594 ;
               RECT 29.094 26.758 29.146 26.794 ;
               RECT 29.094 27.958 29.146 27.994 ;
               RECT 29.094 29.158 29.146 29.194 ;
               RECT 29.094 30.358 29.146 30.394 ;
               RECT 29.094 31.558 29.146 31.594 ;
               RECT 29.094 32.758 29.146 32.794 ;
               RECT 29.094 33.958 29.146 33.994 ;
               RECT 29.094 35.158 29.146 35.194 ;
               RECT 29.094 36.358 29.146 36.394 ;
               RECT 29.094 37.558 29.146 37.594 ;
               RECT 29.094 38.758 29.146 38.794 ;
               RECT 29.094 39.958 29.146 39.994 ;
               RECT 29.094 41.158 29.146 41.194 ;
               RECT 29.094 42.358 29.146 42.394 ;
               RECT 29.094 43.558 29.146 43.594 ;
               RECT 29.094 44.758 29.146 44.794 ;
               RECT 29.094 45.958 29.146 45.994 ;
               RECT 29.094 47.158 29.146 47.194 ;
               RECT 29.094 48.358 29.146 48.394 ;
               RECT 29.094 50.142 29.146 50.178 ;
               RECT 29.094 50.382 29.146 50.418 ;
               RECT 29.094 54.702 29.146 54.738 ;
               RECT 29.094 54.942 29.146 54.978 ;
               RECT 29.094 57.478 29.146 57.514 ;
               RECT 29.094 58.678 29.146 58.714 ;
               RECT 29.094 59.878 29.146 59.914 ;
               RECT 29.094 61.078 29.146 61.114 ;
               RECT 29.094 62.278 29.146 62.314 ;
               RECT 29.094 63.478 29.146 63.514 ;
               RECT 29.094 64.678 29.146 64.714 ;
               RECT 29.094 65.878 29.146 65.914 ;
               RECT 29.094 67.078 29.146 67.114 ;
               RECT 29.094 68.278 29.146 68.314 ;
               RECT 29.094 69.478 29.146 69.514 ;
               RECT 29.094 70.678 29.146 70.714 ;
               RECT 29.094 71.878 29.146 71.914 ;
               RECT 29.094 73.078 29.146 73.114 ;
               RECT 29.094 74.278 29.146 74.314 ;
               RECT 29.094 75.478 29.146 75.514 ;
               RECT 29.094 76.678 29.146 76.714 ;
               RECT 29.094 77.878 29.146 77.914 ;
               RECT 29.094 79.078 29.146 79.114 ;
               RECT 29.094 80.278 29.146 80.314 ;
               RECT 29.094 81.478 29.146 81.514 ;
               RECT 29.094 82.678 29.146 82.714 ;
               RECT 29.094 83.878 29.146 83.914 ;
               RECT 29.094 85.078 29.146 85.114 ;
               RECT 29.094 86.278 29.146 86.314 ;
               RECT 29.094 87.478 29.146 87.514 ;
               RECT 29.094 88.678 29.146 88.714 ;
               RECT 29.094 89.878 29.146 89.914 ;
               RECT 29.094 91.078 29.146 91.114 ;
               RECT 29.094 92.278 29.146 92.314 ;
               RECT 29.094 93.478 29.146 93.514 ;
               RECT 29.094 94.678 29.146 94.714 ;
               RECT 29.094 95.878 29.146 95.914 ;
               RECT 29.094 97.078 29.146 97.114 ;
               RECT 29.094 98.278 29.146 98.314 ;
               RECT 29.094 99.478 29.146 99.514 ;
               RECT 29.094 100.678 29.146 100.714 ;
               RECT 29.094 101.878 29.146 101.914 ;
               RECT 29.094 103.078 29.146 103.114 ;
               RECT 29.094 104.278 29.146 104.314 ;
               RECT 29.174 0.281 29.226 0.317 ;
               RECT 29.174 104.803 29.226 104.839 ;
               RECT 29.254 0.806 29.306 0.842 ;
               RECT 29.254 2.006 29.306 2.042 ;
               RECT 29.254 3.206 29.306 3.242 ;
               RECT 29.254 4.406 29.306 4.442 ;
               RECT 29.254 5.606 29.306 5.642 ;
               RECT 29.254 6.806 29.306 6.842 ;
               RECT 29.254 8.006 29.306 8.042 ;
               RECT 29.254 9.206 29.306 9.242 ;
               RECT 29.254 10.406 29.306 10.442 ;
               RECT 29.254 11.606 29.306 11.642 ;
               RECT 29.254 12.806 29.306 12.842 ;
               RECT 29.254 14.006 29.306 14.042 ;
               RECT 29.254 15.206 29.306 15.242 ;
               RECT 29.254 16.406 29.306 16.442 ;
               RECT 29.254 17.606 29.306 17.642 ;
               RECT 29.254 18.806 29.306 18.842 ;
               RECT 29.254 20.006 29.306 20.042 ;
               RECT 29.254 21.206 29.306 21.242 ;
               RECT 29.254 22.406 29.306 22.442 ;
               RECT 29.254 23.606 29.306 23.642 ;
               RECT 29.254 24.806 29.306 24.842 ;
               RECT 29.254 26.006 29.306 26.042 ;
               RECT 29.254 27.206 29.306 27.242 ;
               RECT 29.254 28.406 29.306 28.442 ;
               RECT 29.254 29.606 29.306 29.642 ;
               RECT 29.254 30.806 29.306 30.842 ;
               RECT 29.254 32.006 29.306 32.042 ;
               RECT 29.254 33.206 29.306 33.242 ;
               RECT 29.254 34.406 29.306 34.442 ;
               RECT 29.254 35.606 29.306 35.642 ;
               RECT 29.254 36.806 29.306 36.842 ;
               RECT 29.254 38.006 29.306 38.042 ;
               RECT 29.254 39.206 29.306 39.242 ;
               RECT 29.254 40.406 29.306 40.442 ;
               RECT 29.254 41.606 29.306 41.642 ;
               RECT 29.254 42.806 29.306 42.842 ;
               RECT 29.254 44.006 29.306 44.042 ;
               RECT 29.254 45.206 29.306 45.242 ;
               RECT 29.254 46.406 29.306 46.442 ;
               RECT 29.254 47.606 29.306 47.642 ;
               RECT 29.254 49.422 29.306 49.458 ;
               RECT 29.254 49.662 29.306 49.698 ;
               RECT 29.254 55.422 29.306 55.458 ;
               RECT 29.254 55.662 29.306 55.698 ;
               RECT 29.254 56.726 29.306 56.762 ;
               RECT 29.254 57.926 29.306 57.962 ;
               RECT 29.254 59.126 29.306 59.162 ;
               RECT 29.254 60.326 29.306 60.362 ;
               RECT 29.254 61.526 29.306 61.562 ;
               RECT 29.254 62.726 29.306 62.762 ;
               RECT 29.254 63.926 29.306 63.962 ;
               RECT 29.254 65.126 29.306 65.162 ;
               RECT 29.254 66.326 29.306 66.362 ;
               RECT 29.254 67.526 29.306 67.562 ;
               RECT 29.254 68.726 29.306 68.762 ;
               RECT 29.254 69.926 29.306 69.962 ;
               RECT 29.254 71.126 29.306 71.162 ;
               RECT 29.254 72.326 29.306 72.362 ;
               RECT 29.254 73.526 29.306 73.562 ;
               RECT 29.254 74.726 29.306 74.762 ;
               RECT 29.254 75.926 29.306 75.962 ;
               RECT 29.254 77.126 29.306 77.162 ;
               RECT 29.254 78.326 29.306 78.362 ;
               RECT 29.254 79.526 29.306 79.562 ;
               RECT 29.254 80.726 29.306 80.762 ;
               RECT 29.254 81.926 29.306 81.962 ;
               RECT 29.254 83.126 29.306 83.162 ;
               RECT 29.254 84.326 29.306 84.362 ;
               RECT 29.254 85.526 29.306 85.562 ;
               RECT 29.254 86.726 29.306 86.762 ;
               RECT 29.254 87.926 29.306 87.962 ;
               RECT 29.254 89.126 29.306 89.162 ;
               RECT 29.254 90.326 29.306 90.362 ;
               RECT 29.254 91.526 29.306 91.562 ;
               RECT 29.254 92.726 29.306 92.762 ;
               RECT 29.254 93.926 29.306 93.962 ;
               RECT 29.254 95.126 29.306 95.162 ;
               RECT 29.254 96.326 29.306 96.362 ;
               RECT 29.254 97.526 29.306 97.562 ;
               RECT 29.254 98.726 29.306 98.762 ;
               RECT 29.254 99.926 29.306 99.962 ;
               RECT 29.254 101.126 29.306 101.162 ;
               RECT 29.254 102.326 29.306 102.362 ;
               RECT 29.254 103.526 29.306 103.562 ;
               RECT 29.334 1.558 29.386 1.594 ;
               RECT 29.334 2.758 29.386 2.794 ;
               RECT 29.334 3.958 29.386 3.994 ;
               RECT 29.334 5.158 29.386 5.194 ;
               RECT 29.334 6.358 29.386 6.394 ;
               RECT 29.334 7.558 29.386 7.594 ;
               RECT 29.334 8.758 29.386 8.794 ;
               RECT 29.334 9.958 29.386 9.994 ;
               RECT 29.334 11.158 29.386 11.194 ;
               RECT 29.334 12.358 29.386 12.394 ;
               RECT 29.334 13.558 29.386 13.594 ;
               RECT 29.334 14.758 29.386 14.794 ;
               RECT 29.334 15.958 29.386 15.994 ;
               RECT 29.334 17.158 29.386 17.194 ;
               RECT 29.334 18.358 29.386 18.394 ;
               RECT 29.334 19.558 29.386 19.594 ;
               RECT 29.334 20.758 29.386 20.794 ;
               RECT 29.334 21.958 29.386 21.994 ;
               RECT 29.334 23.158 29.386 23.194 ;
               RECT 29.334 24.358 29.386 24.394 ;
               RECT 29.334 25.558 29.386 25.594 ;
               RECT 29.334 26.758 29.386 26.794 ;
               RECT 29.334 27.958 29.386 27.994 ;
               RECT 29.334 29.158 29.386 29.194 ;
               RECT 29.334 30.358 29.386 30.394 ;
               RECT 29.334 31.558 29.386 31.594 ;
               RECT 29.334 32.758 29.386 32.794 ;
               RECT 29.334 33.958 29.386 33.994 ;
               RECT 29.334 35.158 29.386 35.194 ;
               RECT 29.334 36.358 29.386 36.394 ;
               RECT 29.334 37.558 29.386 37.594 ;
               RECT 29.334 38.758 29.386 38.794 ;
               RECT 29.334 39.958 29.386 39.994 ;
               RECT 29.334 41.158 29.386 41.194 ;
               RECT 29.334 42.358 29.386 42.394 ;
               RECT 29.334 43.558 29.386 43.594 ;
               RECT 29.334 44.758 29.386 44.794 ;
               RECT 29.334 45.958 29.386 45.994 ;
               RECT 29.334 47.158 29.386 47.194 ;
               RECT 29.334 48.358 29.386 48.394 ;
               RECT 29.334 50.142 29.386 50.178 ;
               RECT 29.334 50.382 29.386 50.418 ;
               RECT 29.334 54.702 29.386 54.738 ;
               RECT 29.334 54.942 29.386 54.978 ;
               RECT 29.334 57.478 29.386 57.514 ;
               RECT 29.334 58.678 29.386 58.714 ;
               RECT 29.334 59.878 29.386 59.914 ;
               RECT 29.334 61.078 29.386 61.114 ;
               RECT 29.334 62.278 29.386 62.314 ;
               RECT 29.334 63.478 29.386 63.514 ;
               RECT 29.334 64.678 29.386 64.714 ;
               RECT 29.334 65.878 29.386 65.914 ;
               RECT 29.334 67.078 29.386 67.114 ;
               RECT 29.334 68.278 29.386 68.314 ;
               RECT 29.334 69.478 29.386 69.514 ;
               RECT 29.334 70.678 29.386 70.714 ;
               RECT 29.334 71.878 29.386 71.914 ;
               RECT 29.334 73.078 29.386 73.114 ;
               RECT 29.334 74.278 29.386 74.314 ;
               RECT 29.334 75.478 29.386 75.514 ;
               RECT 29.334 76.678 29.386 76.714 ;
               RECT 29.334 77.878 29.386 77.914 ;
               RECT 29.334 79.078 29.386 79.114 ;
               RECT 29.334 80.278 29.386 80.314 ;
               RECT 29.334 81.478 29.386 81.514 ;
               RECT 29.334 82.678 29.386 82.714 ;
               RECT 29.334 83.878 29.386 83.914 ;
               RECT 29.334 85.078 29.386 85.114 ;
               RECT 29.334 86.278 29.386 86.314 ;
               RECT 29.334 87.478 29.386 87.514 ;
               RECT 29.334 88.678 29.386 88.714 ;
               RECT 29.334 89.878 29.386 89.914 ;
               RECT 29.334 91.078 29.386 91.114 ;
               RECT 29.334 92.278 29.386 92.314 ;
               RECT 29.334 93.478 29.386 93.514 ;
               RECT 29.334 94.678 29.386 94.714 ;
               RECT 29.334 95.878 29.386 95.914 ;
               RECT 29.334 97.078 29.386 97.114 ;
               RECT 29.334 98.278 29.386 98.314 ;
               RECT 29.334 99.478 29.386 99.514 ;
               RECT 29.334 100.678 29.386 100.714 ;
               RECT 29.334 101.878 29.386 101.914 ;
               RECT 29.334 103.078 29.386 103.114 ;
               RECT 29.334 104.278 29.386 104.314 ;
               RECT 29.414 0.806 29.466 0.842 ;
               RECT 29.414 2.006 29.466 2.042 ;
               RECT 29.414 3.206 29.466 3.242 ;
               RECT 29.414 4.406 29.466 4.442 ;
               RECT 29.414 5.606 29.466 5.642 ;
               RECT 29.414 6.806 29.466 6.842 ;
               RECT 29.414 8.006 29.466 8.042 ;
               RECT 29.414 9.206 29.466 9.242 ;
               RECT 29.414 10.406 29.466 10.442 ;
               RECT 29.414 11.606 29.466 11.642 ;
               RECT 29.414 12.806 29.466 12.842 ;
               RECT 29.414 14.006 29.466 14.042 ;
               RECT 29.414 15.206 29.466 15.242 ;
               RECT 29.414 16.406 29.466 16.442 ;
               RECT 29.414 17.606 29.466 17.642 ;
               RECT 29.414 18.806 29.466 18.842 ;
               RECT 29.414 20.006 29.466 20.042 ;
               RECT 29.414 21.206 29.466 21.242 ;
               RECT 29.414 22.406 29.466 22.442 ;
               RECT 29.414 23.606 29.466 23.642 ;
               RECT 29.414 24.806 29.466 24.842 ;
               RECT 29.414 26.006 29.466 26.042 ;
               RECT 29.414 27.206 29.466 27.242 ;
               RECT 29.414 28.406 29.466 28.442 ;
               RECT 29.414 29.606 29.466 29.642 ;
               RECT 29.414 30.806 29.466 30.842 ;
               RECT 29.414 32.006 29.466 32.042 ;
               RECT 29.414 33.206 29.466 33.242 ;
               RECT 29.414 34.406 29.466 34.442 ;
               RECT 29.414 35.606 29.466 35.642 ;
               RECT 29.414 36.806 29.466 36.842 ;
               RECT 29.414 38.006 29.466 38.042 ;
               RECT 29.414 39.206 29.466 39.242 ;
               RECT 29.414 40.406 29.466 40.442 ;
               RECT 29.414 41.606 29.466 41.642 ;
               RECT 29.414 42.806 29.466 42.842 ;
               RECT 29.414 44.006 29.466 44.042 ;
               RECT 29.414 45.206 29.466 45.242 ;
               RECT 29.414 46.406 29.466 46.442 ;
               RECT 29.414 47.606 29.466 47.642 ;
               RECT 29.414 49.422 29.466 49.458 ;
               RECT 29.414 49.662 29.466 49.698 ;
               RECT 29.414 55.422 29.466 55.458 ;
               RECT 29.414 55.662 29.466 55.698 ;
               RECT 29.414 56.726 29.466 56.762 ;
               RECT 29.414 57.926 29.466 57.962 ;
               RECT 29.414 59.126 29.466 59.162 ;
               RECT 29.414 60.326 29.466 60.362 ;
               RECT 29.414 61.526 29.466 61.562 ;
               RECT 29.414 62.726 29.466 62.762 ;
               RECT 29.414 63.926 29.466 63.962 ;
               RECT 29.414 65.126 29.466 65.162 ;
               RECT 29.414 66.326 29.466 66.362 ;
               RECT 29.414 67.526 29.466 67.562 ;
               RECT 29.414 68.726 29.466 68.762 ;
               RECT 29.414 69.926 29.466 69.962 ;
               RECT 29.414 71.126 29.466 71.162 ;
               RECT 29.414 72.326 29.466 72.362 ;
               RECT 29.414 73.526 29.466 73.562 ;
               RECT 29.414 74.726 29.466 74.762 ;
               RECT 29.414 75.926 29.466 75.962 ;
               RECT 29.414 77.126 29.466 77.162 ;
               RECT 29.414 78.326 29.466 78.362 ;
               RECT 29.414 79.526 29.466 79.562 ;
               RECT 29.414 80.726 29.466 80.762 ;
               RECT 29.414 81.926 29.466 81.962 ;
               RECT 29.414 83.126 29.466 83.162 ;
               RECT 29.414 84.326 29.466 84.362 ;
               RECT 29.414 85.526 29.466 85.562 ;
               RECT 29.414 86.726 29.466 86.762 ;
               RECT 29.414 87.926 29.466 87.962 ;
               RECT 29.414 89.126 29.466 89.162 ;
               RECT 29.414 90.326 29.466 90.362 ;
               RECT 29.414 91.526 29.466 91.562 ;
               RECT 29.414 92.726 29.466 92.762 ;
               RECT 29.414 93.926 29.466 93.962 ;
               RECT 29.414 95.126 29.466 95.162 ;
               RECT 29.414 96.326 29.466 96.362 ;
               RECT 29.414 97.526 29.466 97.562 ;
               RECT 29.414 98.726 29.466 98.762 ;
               RECT 29.414 99.926 29.466 99.962 ;
               RECT 29.414 101.126 29.466 101.162 ;
               RECT 29.414 102.326 29.466 102.362 ;
               RECT 29.414 103.526 29.466 103.562 ;
               RECT 29.494 1.558 29.546 1.594 ;
               RECT 29.494 2.758 29.546 2.794 ;
               RECT 29.494 3.958 29.546 3.994 ;
               RECT 29.494 5.158 29.546 5.194 ;
               RECT 29.494 6.358 29.546 6.394 ;
               RECT 29.494 7.558 29.546 7.594 ;
               RECT 29.494 8.758 29.546 8.794 ;
               RECT 29.494 9.958 29.546 9.994 ;
               RECT 29.494 11.158 29.546 11.194 ;
               RECT 29.494 12.358 29.546 12.394 ;
               RECT 29.494 13.558 29.546 13.594 ;
               RECT 29.494 14.758 29.546 14.794 ;
               RECT 29.494 15.958 29.546 15.994 ;
               RECT 29.494 17.158 29.546 17.194 ;
               RECT 29.494 18.358 29.546 18.394 ;
               RECT 29.494 19.558 29.546 19.594 ;
               RECT 29.494 20.758 29.546 20.794 ;
               RECT 29.494 21.958 29.546 21.994 ;
               RECT 29.494 23.158 29.546 23.194 ;
               RECT 29.494 24.358 29.546 24.394 ;
               RECT 29.494 25.558 29.546 25.594 ;
               RECT 29.494 26.758 29.546 26.794 ;
               RECT 29.494 27.958 29.546 27.994 ;
               RECT 29.494 29.158 29.546 29.194 ;
               RECT 29.494 30.358 29.546 30.394 ;
               RECT 29.494 31.558 29.546 31.594 ;
               RECT 29.494 32.758 29.546 32.794 ;
               RECT 29.494 33.958 29.546 33.994 ;
               RECT 29.494 35.158 29.546 35.194 ;
               RECT 29.494 36.358 29.546 36.394 ;
               RECT 29.494 37.558 29.546 37.594 ;
               RECT 29.494 38.758 29.546 38.794 ;
               RECT 29.494 39.958 29.546 39.994 ;
               RECT 29.494 41.158 29.546 41.194 ;
               RECT 29.494 42.358 29.546 42.394 ;
               RECT 29.494 43.558 29.546 43.594 ;
               RECT 29.494 44.758 29.546 44.794 ;
               RECT 29.494 45.958 29.546 45.994 ;
               RECT 29.494 47.158 29.546 47.194 ;
               RECT 29.494 48.358 29.546 48.394 ;
               RECT 29.494 50.142 29.546 50.178 ;
               RECT 29.494 50.382 29.546 50.418 ;
               RECT 29.494 54.702 29.546 54.738 ;
               RECT 29.494 54.942 29.546 54.978 ;
               RECT 29.494 57.478 29.546 57.514 ;
               RECT 29.494 58.678 29.546 58.714 ;
               RECT 29.494 59.878 29.546 59.914 ;
               RECT 29.494 61.078 29.546 61.114 ;
               RECT 29.494 62.278 29.546 62.314 ;
               RECT 29.494 63.478 29.546 63.514 ;
               RECT 29.494 64.678 29.546 64.714 ;
               RECT 29.494 65.878 29.546 65.914 ;
               RECT 29.494 67.078 29.546 67.114 ;
               RECT 29.494 68.278 29.546 68.314 ;
               RECT 29.494 69.478 29.546 69.514 ;
               RECT 29.494 70.678 29.546 70.714 ;
               RECT 29.494 71.878 29.546 71.914 ;
               RECT 29.494 73.078 29.546 73.114 ;
               RECT 29.494 74.278 29.546 74.314 ;
               RECT 29.494 75.478 29.546 75.514 ;
               RECT 29.494 76.678 29.546 76.714 ;
               RECT 29.494 77.878 29.546 77.914 ;
               RECT 29.494 79.078 29.546 79.114 ;
               RECT 29.494 80.278 29.546 80.314 ;
               RECT 29.494 81.478 29.546 81.514 ;
               RECT 29.494 82.678 29.546 82.714 ;
               RECT 29.494 83.878 29.546 83.914 ;
               RECT 29.494 85.078 29.546 85.114 ;
               RECT 29.494 86.278 29.546 86.314 ;
               RECT 29.494 87.478 29.546 87.514 ;
               RECT 29.494 88.678 29.546 88.714 ;
               RECT 29.494 89.878 29.546 89.914 ;
               RECT 29.494 91.078 29.546 91.114 ;
               RECT 29.494 92.278 29.546 92.314 ;
               RECT 29.494 93.478 29.546 93.514 ;
               RECT 29.494 94.678 29.546 94.714 ;
               RECT 29.494 95.878 29.546 95.914 ;
               RECT 29.494 97.078 29.546 97.114 ;
               RECT 29.494 98.278 29.546 98.314 ;
               RECT 29.494 99.478 29.546 99.514 ;
               RECT 29.494 100.678 29.546 100.714 ;
               RECT 29.494 101.878 29.546 101.914 ;
               RECT 29.494 103.078 29.546 103.114 ;
               RECT 29.494 104.278 29.546 104.314 ;
               RECT 29.574 0.281 29.626 0.317 ;
               RECT 29.574 104.803 29.626 104.839 ;
               RECT 29.654 0.806 29.706 0.842 ;
               RECT 29.654 2.006 29.706 2.042 ;
               RECT 29.654 3.206 29.706 3.242 ;
               RECT 29.654 4.406 29.706 4.442 ;
               RECT 29.654 5.606 29.706 5.642 ;
               RECT 29.654 6.806 29.706 6.842 ;
               RECT 29.654 8.006 29.706 8.042 ;
               RECT 29.654 9.206 29.706 9.242 ;
               RECT 29.654 10.406 29.706 10.442 ;
               RECT 29.654 11.606 29.706 11.642 ;
               RECT 29.654 12.806 29.706 12.842 ;
               RECT 29.654 14.006 29.706 14.042 ;
               RECT 29.654 15.206 29.706 15.242 ;
               RECT 29.654 16.406 29.706 16.442 ;
               RECT 29.654 17.606 29.706 17.642 ;
               RECT 29.654 18.806 29.706 18.842 ;
               RECT 29.654 20.006 29.706 20.042 ;
               RECT 29.654 21.206 29.706 21.242 ;
               RECT 29.654 22.406 29.706 22.442 ;
               RECT 29.654 23.606 29.706 23.642 ;
               RECT 29.654 24.806 29.706 24.842 ;
               RECT 29.654 26.006 29.706 26.042 ;
               RECT 29.654 27.206 29.706 27.242 ;
               RECT 29.654 28.406 29.706 28.442 ;
               RECT 29.654 29.606 29.706 29.642 ;
               RECT 29.654 30.806 29.706 30.842 ;
               RECT 29.654 32.006 29.706 32.042 ;
               RECT 29.654 33.206 29.706 33.242 ;
               RECT 29.654 34.406 29.706 34.442 ;
               RECT 29.654 35.606 29.706 35.642 ;
               RECT 29.654 36.806 29.706 36.842 ;
               RECT 29.654 38.006 29.706 38.042 ;
               RECT 29.654 39.206 29.706 39.242 ;
               RECT 29.654 40.406 29.706 40.442 ;
               RECT 29.654 41.606 29.706 41.642 ;
               RECT 29.654 42.806 29.706 42.842 ;
               RECT 29.654 44.006 29.706 44.042 ;
               RECT 29.654 45.206 29.706 45.242 ;
               RECT 29.654 46.406 29.706 46.442 ;
               RECT 29.654 47.606 29.706 47.642 ;
               RECT 29.654 49.422 29.706 49.458 ;
               RECT 29.654 49.662 29.706 49.698 ;
               RECT 29.654 51.102 29.706 51.138 ;
               RECT 29.654 51.582 29.706 51.618 ;
               RECT 29.654 53.502 29.706 53.538 ;
               RECT 29.654 53.982 29.706 54.018 ;
               RECT 29.654 55.422 29.706 55.458 ;
               RECT 29.654 55.662 29.706 55.698 ;
               RECT 29.654 56.726 29.706 56.762 ;
               RECT 29.654 57.926 29.706 57.962 ;
               RECT 29.654 59.126 29.706 59.162 ;
               RECT 29.654 60.326 29.706 60.362 ;
               RECT 29.654 61.526 29.706 61.562 ;
               RECT 29.654 62.726 29.706 62.762 ;
               RECT 29.654 63.926 29.706 63.962 ;
               RECT 29.654 65.126 29.706 65.162 ;
               RECT 29.654 66.326 29.706 66.362 ;
               RECT 29.654 67.526 29.706 67.562 ;
               RECT 29.654 68.726 29.706 68.762 ;
               RECT 29.654 69.926 29.706 69.962 ;
               RECT 29.654 71.126 29.706 71.162 ;
               RECT 29.654 72.326 29.706 72.362 ;
               RECT 29.654 73.526 29.706 73.562 ;
               RECT 29.654 74.726 29.706 74.762 ;
               RECT 29.654 75.926 29.706 75.962 ;
               RECT 29.654 77.126 29.706 77.162 ;
               RECT 29.654 78.326 29.706 78.362 ;
               RECT 29.654 79.526 29.706 79.562 ;
               RECT 29.654 80.726 29.706 80.762 ;
               RECT 29.654 81.926 29.706 81.962 ;
               RECT 29.654 83.126 29.706 83.162 ;
               RECT 29.654 84.326 29.706 84.362 ;
               RECT 29.654 85.526 29.706 85.562 ;
               RECT 29.654 86.726 29.706 86.762 ;
               RECT 29.654 87.926 29.706 87.962 ;
               RECT 29.654 89.126 29.706 89.162 ;
               RECT 29.654 90.326 29.706 90.362 ;
               RECT 29.654 91.526 29.706 91.562 ;
               RECT 29.654 92.726 29.706 92.762 ;
               RECT 29.654 93.926 29.706 93.962 ;
               RECT 29.654 95.126 29.706 95.162 ;
               RECT 29.654 96.326 29.706 96.362 ;
               RECT 29.654 97.526 29.706 97.562 ;
               RECT 29.654 98.726 29.706 98.762 ;
               RECT 29.654 99.926 29.706 99.962 ;
               RECT 29.654 101.126 29.706 101.162 ;
               RECT 29.654 102.326 29.706 102.362 ;
               RECT 29.654 103.526 29.706 103.562 ;
               RECT 29.734 1.558 29.786 1.594 ;
               RECT 29.734 2.758 29.786 2.794 ;
               RECT 29.734 3.958 29.786 3.994 ;
               RECT 29.734 5.158 29.786 5.194 ;
               RECT 29.734 6.358 29.786 6.394 ;
               RECT 29.734 7.558 29.786 7.594 ;
               RECT 29.734 8.758 29.786 8.794 ;
               RECT 29.734 9.958 29.786 9.994 ;
               RECT 29.734 11.158 29.786 11.194 ;
               RECT 29.734 12.358 29.786 12.394 ;
               RECT 29.734 13.558 29.786 13.594 ;
               RECT 29.734 14.758 29.786 14.794 ;
               RECT 29.734 15.958 29.786 15.994 ;
               RECT 29.734 17.158 29.786 17.194 ;
               RECT 29.734 18.358 29.786 18.394 ;
               RECT 29.734 19.558 29.786 19.594 ;
               RECT 29.734 20.758 29.786 20.794 ;
               RECT 29.734 21.958 29.786 21.994 ;
               RECT 29.734 23.158 29.786 23.194 ;
               RECT 29.734 24.358 29.786 24.394 ;
               RECT 29.734 25.558 29.786 25.594 ;
               RECT 29.734 26.758 29.786 26.794 ;
               RECT 29.734 27.958 29.786 27.994 ;
               RECT 29.734 29.158 29.786 29.194 ;
               RECT 29.734 30.358 29.786 30.394 ;
               RECT 29.734 31.558 29.786 31.594 ;
               RECT 29.734 32.758 29.786 32.794 ;
               RECT 29.734 33.958 29.786 33.994 ;
               RECT 29.734 35.158 29.786 35.194 ;
               RECT 29.734 36.358 29.786 36.394 ;
               RECT 29.734 37.558 29.786 37.594 ;
               RECT 29.734 38.758 29.786 38.794 ;
               RECT 29.734 39.958 29.786 39.994 ;
               RECT 29.734 41.158 29.786 41.194 ;
               RECT 29.734 42.358 29.786 42.394 ;
               RECT 29.734 43.558 29.786 43.594 ;
               RECT 29.734 44.758 29.786 44.794 ;
               RECT 29.734 45.958 29.786 45.994 ;
               RECT 29.734 47.158 29.786 47.194 ;
               RECT 29.734 48.358 29.786 48.394 ;
               RECT 29.734 50.142 29.786 50.178 ;
               RECT 29.734 50.382 29.786 50.418 ;
               RECT 29.734 54.702 29.786 54.738 ;
               RECT 29.734 54.942 29.786 54.978 ;
               RECT 29.734 57.478 29.786 57.514 ;
               RECT 29.734 58.678 29.786 58.714 ;
               RECT 29.734 59.878 29.786 59.914 ;
               RECT 29.734 61.078 29.786 61.114 ;
               RECT 29.734 62.278 29.786 62.314 ;
               RECT 29.734 63.478 29.786 63.514 ;
               RECT 29.734 64.678 29.786 64.714 ;
               RECT 29.734 65.878 29.786 65.914 ;
               RECT 29.734 67.078 29.786 67.114 ;
               RECT 29.734 68.278 29.786 68.314 ;
               RECT 29.734 69.478 29.786 69.514 ;
               RECT 29.734 70.678 29.786 70.714 ;
               RECT 29.734 71.878 29.786 71.914 ;
               RECT 29.734 73.078 29.786 73.114 ;
               RECT 29.734 74.278 29.786 74.314 ;
               RECT 29.734 75.478 29.786 75.514 ;
               RECT 29.734 76.678 29.786 76.714 ;
               RECT 29.734 77.878 29.786 77.914 ;
               RECT 29.734 79.078 29.786 79.114 ;
               RECT 29.734 80.278 29.786 80.314 ;
               RECT 29.734 81.478 29.786 81.514 ;
               RECT 29.734 82.678 29.786 82.714 ;
               RECT 29.734 83.878 29.786 83.914 ;
               RECT 29.734 85.078 29.786 85.114 ;
               RECT 29.734 86.278 29.786 86.314 ;
               RECT 29.734 87.478 29.786 87.514 ;
               RECT 29.734 88.678 29.786 88.714 ;
               RECT 29.734 89.878 29.786 89.914 ;
               RECT 29.734 91.078 29.786 91.114 ;
               RECT 29.734 92.278 29.786 92.314 ;
               RECT 29.734 93.478 29.786 93.514 ;
               RECT 29.734 94.678 29.786 94.714 ;
               RECT 29.734 95.878 29.786 95.914 ;
               RECT 29.734 97.078 29.786 97.114 ;
               RECT 29.734 98.278 29.786 98.314 ;
               RECT 29.734 99.478 29.786 99.514 ;
               RECT 29.734 100.678 29.786 100.714 ;
               RECT 29.734 101.878 29.786 101.914 ;
               RECT 29.734 103.078 29.786 103.114 ;
               RECT 29.734 104.278 29.786 104.314 ;
               RECT 29.814 0.806 29.866 0.842 ;
               RECT 29.814 2.006 29.866 2.042 ;
               RECT 29.814 3.206 29.866 3.242 ;
               RECT 29.814 4.406 29.866 4.442 ;
               RECT 29.814 5.606 29.866 5.642 ;
               RECT 29.814 6.806 29.866 6.842 ;
               RECT 29.814 8.006 29.866 8.042 ;
               RECT 29.814 9.206 29.866 9.242 ;
               RECT 29.814 10.406 29.866 10.442 ;
               RECT 29.814 11.606 29.866 11.642 ;
               RECT 29.814 12.806 29.866 12.842 ;
               RECT 29.814 14.006 29.866 14.042 ;
               RECT 29.814 15.206 29.866 15.242 ;
               RECT 29.814 16.406 29.866 16.442 ;
               RECT 29.814 17.606 29.866 17.642 ;
               RECT 29.814 18.806 29.866 18.842 ;
               RECT 29.814 20.006 29.866 20.042 ;
               RECT 29.814 21.206 29.866 21.242 ;
               RECT 29.814 22.406 29.866 22.442 ;
               RECT 29.814 23.606 29.866 23.642 ;
               RECT 29.814 24.806 29.866 24.842 ;
               RECT 29.814 26.006 29.866 26.042 ;
               RECT 29.814 27.206 29.866 27.242 ;
               RECT 29.814 28.406 29.866 28.442 ;
               RECT 29.814 29.606 29.866 29.642 ;
               RECT 29.814 30.806 29.866 30.842 ;
               RECT 29.814 32.006 29.866 32.042 ;
               RECT 29.814 33.206 29.866 33.242 ;
               RECT 29.814 34.406 29.866 34.442 ;
               RECT 29.814 35.606 29.866 35.642 ;
               RECT 29.814 36.806 29.866 36.842 ;
               RECT 29.814 38.006 29.866 38.042 ;
               RECT 29.814 39.206 29.866 39.242 ;
               RECT 29.814 40.406 29.866 40.442 ;
               RECT 29.814 41.606 29.866 41.642 ;
               RECT 29.814 42.806 29.866 42.842 ;
               RECT 29.814 44.006 29.866 44.042 ;
               RECT 29.814 45.206 29.866 45.242 ;
               RECT 29.814 46.406 29.866 46.442 ;
               RECT 29.814 47.606 29.866 47.642 ;
               RECT 29.814 49.422 29.866 49.458 ;
               RECT 29.814 49.662 29.866 49.698 ;
               RECT 29.814 55.422 29.866 55.458 ;
               RECT 29.814 55.662 29.866 55.698 ;
               RECT 29.814 56.726 29.866 56.762 ;
               RECT 29.814 57.926 29.866 57.962 ;
               RECT 29.814 59.126 29.866 59.162 ;
               RECT 29.814 60.326 29.866 60.362 ;
               RECT 29.814 61.526 29.866 61.562 ;
               RECT 29.814 62.726 29.866 62.762 ;
               RECT 29.814 63.926 29.866 63.962 ;
               RECT 29.814 65.126 29.866 65.162 ;
               RECT 29.814 66.326 29.866 66.362 ;
               RECT 29.814 67.526 29.866 67.562 ;
               RECT 29.814 68.726 29.866 68.762 ;
               RECT 29.814 69.926 29.866 69.962 ;
               RECT 29.814 71.126 29.866 71.162 ;
               RECT 29.814 72.326 29.866 72.362 ;
               RECT 29.814 73.526 29.866 73.562 ;
               RECT 29.814 74.726 29.866 74.762 ;
               RECT 29.814 75.926 29.866 75.962 ;
               RECT 29.814 77.126 29.866 77.162 ;
               RECT 29.814 78.326 29.866 78.362 ;
               RECT 29.814 79.526 29.866 79.562 ;
               RECT 29.814 80.726 29.866 80.762 ;
               RECT 29.814 81.926 29.866 81.962 ;
               RECT 29.814 83.126 29.866 83.162 ;
               RECT 29.814 84.326 29.866 84.362 ;
               RECT 29.814 85.526 29.866 85.562 ;
               RECT 29.814 86.726 29.866 86.762 ;
               RECT 29.814 87.926 29.866 87.962 ;
               RECT 29.814 89.126 29.866 89.162 ;
               RECT 29.814 90.326 29.866 90.362 ;
               RECT 29.814 91.526 29.866 91.562 ;
               RECT 29.814 92.726 29.866 92.762 ;
               RECT 29.814 93.926 29.866 93.962 ;
               RECT 29.814 95.126 29.866 95.162 ;
               RECT 29.814 96.326 29.866 96.362 ;
               RECT 29.814 97.526 29.866 97.562 ;
               RECT 29.814 98.726 29.866 98.762 ;
               RECT 29.814 99.926 29.866 99.962 ;
               RECT 29.814 101.126 29.866 101.162 ;
               RECT 29.814 102.326 29.866 102.362 ;
               RECT 29.814 103.526 29.866 103.562 ;
               RECT 29.894 1.558 29.946 1.594 ;
               RECT 29.894 2.758 29.946 2.794 ;
               RECT 29.894 3.958 29.946 3.994 ;
               RECT 29.894 5.158 29.946 5.194 ;
               RECT 29.894 6.358 29.946 6.394 ;
               RECT 29.894 7.558 29.946 7.594 ;
               RECT 29.894 8.758 29.946 8.794 ;
               RECT 29.894 9.958 29.946 9.994 ;
               RECT 29.894 11.158 29.946 11.194 ;
               RECT 29.894 12.358 29.946 12.394 ;
               RECT 29.894 13.558 29.946 13.594 ;
               RECT 29.894 14.758 29.946 14.794 ;
               RECT 29.894 15.958 29.946 15.994 ;
               RECT 29.894 17.158 29.946 17.194 ;
               RECT 29.894 18.358 29.946 18.394 ;
               RECT 29.894 19.558 29.946 19.594 ;
               RECT 29.894 20.758 29.946 20.794 ;
               RECT 29.894 21.958 29.946 21.994 ;
               RECT 29.894 23.158 29.946 23.194 ;
               RECT 29.894 24.358 29.946 24.394 ;
               RECT 29.894 25.558 29.946 25.594 ;
               RECT 29.894 26.758 29.946 26.794 ;
               RECT 29.894 27.958 29.946 27.994 ;
               RECT 29.894 29.158 29.946 29.194 ;
               RECT 29.894 30.358 29.946 30.394 ;
               RECT 29.894 31.558 29.946 31.594 ;
               RECT 29.894 32.758 29.946 32.794 ;
               RECT 29.894 33.958 29.946 33.994 ;
               RECT 29.894 35.158 29.946 35.194 ;
               RECT 29.894 36.358 29.946 36.394 ;
               RECT 29.894 37.558 29.946 37.594 ;
               RECT 29.894 38.758 29.946 38.794 ;
               RECT 29.894 39.958 29.946 39.994 ;
               RECT 29.894 41.158 29.946 41.194 ;
               RECT 29.894 42.358 29.946 42.394 ;
               RECT 29.894 43.558 29.946 43.594 ;
               RECT 29.894 44.758 29.946 44.794 ;
               RECT 29.894 45.958 29.946 45.994 ;
               RECT 29.894 47.158 29.946 47.194 ;
               RECT 29.894 48.358 29.946 48.394 ;
               RECT 29.894 50.142 29.946 50.178 ;
               RECT 29.894 50.382 29.946 50.418 ;
               RECT 29.894 54.702 29.946 54.738 ;
               RECT 29.894 54.942 29.946 54.978 ;
               RECT 29.894 57.478 29.946 57.514 ;
               RECT 29.894 58.678 29.946 58.714 ;
               RECT 29.894 59.878 29.946 59.914 ;
               RECT 29.894 61.078 29.946 61.114 ;
               RECT 29.894 62.278 29.946 62.314 ;
               RECT 29.894 63.478 29.946 63.514 ;
               RECT 29.894 64.678 29.946 64.714 ;
               RECT 29.894 65.878 29.946 65.914 ;
               RECT 29.894 67.078 29.946 67.114 ;
               RECT 29.894 68.278 29.946 68.314 ;
               RECT 29.894 69.478 29.946 69.514 ;
               RECT 29.894 70.678 29.946 70.714 ;
               RECT 29.894 71.878 29.946 71.914 ;
               RECT 29.894 73.078 29.946 73.114 ;
               RECT 29.894 74.278 29.946 74.314 ;
               RECT 29.894 75.478 29.946 75.514 ;
               RECT 29.894 76.678 29.946 76.714 ;
               RECT 29.894 77.878 29.946 77.914 ;
               RECT 29.894 79.078 29.946 79.114 ;
               RECT 29.894 80.278 29.946 80.314 ;
               RECT 29.894 81.478 29.946 81.514 ;
               RECT 29.894 82.678 29.946 82.714 ;
               RECT 29.894 83.878 29.946 83.914 ;
               RECT 29.894 85.078 29.946 85.114 ;
               RECT 29.894 86.278 29.946 86.314 ;
               RECT 29.894 87.478 29.946 87.514 ;
               RECT 29.894 88.678 29.946 88.714 ;
               RECT 29.894 89.878 29.946 89.914 ;
               RECT 29.894 91.078 29.946 91.114 ;
               RECT 29.894 92.278 29.946 92.314 ;
               RECT 29.894 93.478 29.946 93.514 ;
               RECT 29.894 94.678 29.946 94.714 ;
               RECT 29.894 95.878 29.946 95.914 ;
               RECT 29.894 97.078 29.946 97.114 ;
               RECT 29.894 98.278 29.946 98.314 ;
               RECT 29.894 99.478 29.946 99.514 ;
               RECT 29.894 100.678 29.946 100.714 ;
               RECT 29.894 101.878 29.946 101.914 ;
               RECT 29.894 103.078 29.946 103.114 ;
               RECT 29.894 104.278 29.946 104.314 ;
               RECT 29.974 0.281 30.026 0.317 ;
               RECT 29.974 104.803 30.026 104.839 ;
               RECT 30.054 0.806 30.106 0.842 ;
               RECT 30.054 2.006 30.106 2.042 ;
               RECT 30.054 3.206 30.106 3.242 ;
               RECT 30.054 4.406 30.106 4.442 ;
               RECT 30.054 5.606 30.106 5.642 ;
               RECT 30.054 6.806 30.106 6.842 ;
               RECT 30.054 8.006 30.106 8.042 ;
               RECT 30.054 9.206 30.106 9.242 ;
               RECT 30.054 10.406 30.106 10.442 ;
               RECT 30.054 11.606 30.106 11.642 ;
               RECT 30.054 12.806 30.106 12.842 ;
               RECT 30.054 14.006 30.106 14.042 ;
               RECT 30.054 15.206 30.106 15.242 ;
               RECT 30.054 16.406 30.106 16.442 ;
               RECT 30.054 17.606 30.106 17.642 ;
               RECT 30.054 18.806 30.106 18.842 ;
               RECT 30.054 20.006 30.106 20.042 ;
               RECT 30.054 21.206 30.106 21.242 ;
               RECT 30.054 22.406 30.106 22.442 ;
               RECT 30.054 23.606 30.106 23.642 ;
               RECT 30.054 24.806 30.106 24.842 ;
               RECT 30.054 26.006 30.106 26.042 ;
               RECT 30.054 27.206 30.106 27.242 ;
               RECT 30.054 28.406 30.106 28.442 ;
               RECT 30.054 29.606 30.106 29.642 ;
               RECT 30.054 30.806 30.106 30.842 ;
               RECT 30.054 32.006 30.106 32.042 ;
               RECT 30.054 33.206 30.106 33.242 ;
               RECT 30.054 34.406 30.106 34.442 ;
               RECT 30.054 35.606 30.106 35.642 ;
               RECT 30.054 36.806 30.106 36.842 ;
               RECT 30.054 38.006 30.106 38.042 ;
               RECT 30.054 39.206 30.106 39.242 ;
               RECT 30.054 40.406 30.106 40.442 ;
               RECT 30.054 41.606 30.106 41.642 ;
               RECT 30.054 42.806 30.106 42.842 ;
               RECT 30.054 44.006 30.106 44.042 ;
               RECT 30.054 45.206 30.106 45.242 ;
               RECT 30.054 46.406 30.106 46.442 ;
               RECT 30.054 47.606 30.106 47.642 ;
               RECT 30.054 49.422 30.106 49.458 ;
               RECT 30.054 49.662 30.106 49.698 ;
               RECT 30.054 55.422 30.106 55.458 ;
               RECT 30.054 55.662 30.106 55.698 ;
               RECT 30.054 56.726 30.106 56.762 ;
               RECT 30.054 57.926 30.106 57.962 ;
               RECT 30.054 59.126 30.106 59.162 ;
               RECT 30.054 60.326 30.106 60.362 ;
               RECT 30.054 61.526 30.106 61.562 ;
               RECT 30.054 62.726 30.106 62.762 ;
               RECT 30.054 63.926 30.106 63.962 ;
               RECT 30.054 65.126 30.106 65.162 ;
               RECT 30.054 66.326 30.106 66.362 ;
               RECT 30.054 67.526 30.106 67.562 ;
               RECT 30.054 68.726 30.106 68.762 ;
               RECT 30.054 69.926 30.106 69.962 ;
               RECT 30.054 71.126 30.106 71.162 ;
               RECT 30.054 72.326 30.106 72.362 ;
               RECT 30.054 73.526 30.106 73.562 ;
               RECT 30.054 74.726 30.106 74.762 ;
               RECT 30.054 75.926 30.106 75.962 ;
               RECT 30.054 77.126 30.106 77.162 ;
               RECT 30.054 78.326 30.106 78.362 ;
               RECT 30.054 79.526 30.106 79.562 ;
               RECT 30.054 80.726 30.106 80.762 ;
               RECT 30.054 81.926 30.106 81.962 ;
               RECT 30.054 83.126 30.106 83.162 ;
               RECT 30.054 84.326 30.106 84.362 ;
               RECT 30.054 85.526 30.106 85.562 ;
               RECT 30.054 86.726 30.106 86.762 ;
               RECT 30.054 87.926 30.106 87.962 ;
               RECT 30.054 89.126 30.106 89.162 ;
               RECT 30.054 90.326 30.106 90.362 ;
               RECT 30.054 91.526 30.106 91.562 ;
               RECT 30.054 92.726 30.106 92.762 ;
               RECT 30.054 93.926 30.106 93.962 ;
               RECT 30.054 95.126 30.106 95.162 ;
               RECT 30.054 96.326 30.106 96.362 ;
               RECT 30.054 97.526 30.106 97.562 ;
               RECT 30.054 98.726 30.106 98.762 ;
               RECT 30.054 99.926 30.106 99.962 ;
               RECT 30.054 101.126 30.106 101.162 ;
               RECT 30.054 102.326 30.106 102.362 ;
               RECT 30.054 103.526 30.106 103.562 ;
               RECT 30.134 1.558 30.186 1.594 ;
               RECT 30.134 2.758 30.186 2.794 ;
               RECT 30.134 3.958 30.186 3.994 ;
               RECT 30.134 5.158 30.186 5.194 ;
               RECT 30.134 6.358 30.186 6.394 ;
               RECT 30.134 7.558 30.186 7.594 ;
               RECT 30.134 8.758 30.186 8.794 ;
               RECT 30.134 9.958 30.186 9.994 ;
               RECT 30.134 11.158 30.186 11.194 ;
               RECT 30.134 12.358 30.186 12.394 ;
               RECT 30.134 13.558 30.186 13.594 ;
               RECT 30.134 14.758 30.186 14.794 ;
               RECT 30.134 15.958 30.186 15.994 ;
               RECT 30.134 17.158 30.186 17.194 ;
               RECT 30.134 18.358 30.186 18.394 ;
               RECT 30.134 19.558 30.186 19.594 ;
               RECT 30.134 20.758 30.186 20.794 ;
               RECT 30.134 21.958 30.186 21.994 ;
               RECT 30.134 23.158 30.186 23.194 ;
               RECT 30.134 24.358 30.186 24.394 ;
               RECT 30.134 25.558 30.186 25.594 ;
               RECT 30.134 26.758 30.186 26.794 ;
               RECT 30.134 27.958 30.186 27.994 ;
               RECT 30.134 29.158 30.186 29.194 ;
               RECT 30.134 30.358 30.186 30.394 ;
               RECT 30.134 31.558 30.186 31.594 ;
               RECT 30.134 32.758 30.186 32.794 ;
               RECT 30.134 33.958 30.186 33.994 ;
               RECT 30.134 35.158 30.186 35.194 ;
               RECT 30.134 36.358 30.186 36.394 ;
               RECT 30.134 37.558 30.186 37.594 ;
               RECT 30.134 38.758 30.186 38.794 ;
               RECT 30.134 39.958 30.186 39.994 ;
               RECT 30.134 41.158 30.186 41.194 ;
               RECT 30.134 42.358 30.186 42.394 ;
               RECT 30.134 43.558 30.186 43.594 ;
               RECT 30.134 44.758 30.186 44.794 ;
               RECT 30.134 45.958 30.186 45.994 ;
               RECT 30.134 47.158 30.186 47.194 ;
               RECT 30.134 48.358 30.186 48.394 ;
               RECT 30.134 50.142 30.186 50.178 ;
               RECT 30.134 50.382 30.186 50.418 ;
               RECT 30.134 54.702 30.186 54.738 ;
               RECT 30.134 54.942 30.186 54.978 ;
               RECT 30.134 57.478 30.186 57.514 ;
               RECT 30.134 58.678 30.186 58.714 ;
               RECT 30.134 59.878 30.186 59.914 ;
               RECT 30.134 61.078 30.186 61.114 ;
               RECT 30.134 62.278 30.186 62.314 ;
               RECT 30.134 63.478 30.186 63.514 ;
               RECT 30.134 64.678 30.186 64.714 ;
               RECT 30.134 65.878 30.186 65.914 ;
               RECT 30.134 67.078 30.186 67.114 ;
               RECT 30.134 68.278 30.186 68.314 ;
               RECT 30.134 69.478 30.186 69.514 ;
               RECT 30.134 70.678 30.186 70.714 ;
               RECT 30.134 71.878 30.186 71.914 ;
               RECT 30.134 73.078 30.186 73.114 ;
               RECT 30.134 74.278 30.186 74.314 ;
               RECT 30.134 75.478 30.186 75.514 ;
               RECT 30.134 76.678 30.186 76.714 ;
               RECT 30.134 77.878 30.186 77.914 ;
               RECT 30.134 79.078 30.186 79.114 ;
               RECT 30.134 80.278 30.186 80.314 ;
               RECT 30.134 81.478 30.186 81.514 ;
               RECT 30.134 82.678 30.186 82.714 ;
               RECT 30.134 83.878 30.186 83.914 ;
               RECT 30.134 85.078 30.186 85.114 ;
               RECT 30.134 86.278 30.186 86.314 ;
               RECT 30.134 87.478 30.186 87.514 ;
               RECT 30.134 88.678 30.186 88.714 ;
               RECT 30.134 89.878 30.186 89.914 ;
               RECT 30.134 91.078 30.186 91.114 ;
               RECT 30.134 92.278 30.186 92.314 ;
               RECT 30.134 93.478 30.186 93.514 ;
               RECT 30.134 94.678 30.186 94.714 ;
               RECT 30.134 95.878 30.186 95.914 ;
               RECT 30.134 97.078 30.186 97.114 ;
               RECT 30.134 98.278 30.186 98.314 ;
               RECT 30.134 99.478 30.186 99.514 ;
               RECT 30.134 100.678 30.186 100.714 ;
               RECT 30.134 101.878 30.186 101.914 ;
               RECT 30.134 103.078 30.186 103.114 ;
               RECT 30.134 104.278 30.186 104.314 ;
               RECT 30.214 0.806 30.266 0.842 ;
               RECT 30.214 2.006 30.266 2.042 ;
               RECT 30.214 3.206 30.266 3.242 ;
               RECT 30.214 4.406 30.266 4.442 ;
               RECT 30.214 5.606 30.266 5.642 ;
               RECT 30.214 6.806 30.266 6.842 ;
               RECT 30.214 8.006 30.266 8.042 ;
               RECT 30.214 9.206 30.266 9.242 ;
               RECT 30.214 10.406 30.266 10.442 ;
               RECT 30.214 11.606 30.266 11.642 ;
               RECT 30.214 12.806 30.266 12.842 ;
               RECT 30.214 14.006 30.266 14.042 ;
               RECT 30.214 15.206 30.266 15.242 ;
               RECT 30.214 16.406 30.266 16.442 ;
               RECT 30.214 17.606 30.266 17.642 ;
               RECT 30.214 18.806 30.266 18.842 ;
               RECT 30.214 20.006 30.266 20.042 ;
               RECT 30.214 21.206 30.266 21.242 ;
               RECT 30.214 22.406 30.266 22.442 ;
               RECT 30.214 23.606 30.266 23.642 ;
               RECT 30.214 24.806 30.266 24.842 ;
               RECT 30.214 26.006 30.266 26.042 ;
               RECT 30.214 27.206 30.266 27.242 ;
               RECT 30.214 28.406 30.266 28.442 ;
               RECT 30.214 29.606 30.266 29.642 ;
               RECT 30.214 30.806 30.266 30.842 ;
               RECT 30.214 32.006 30.266 32.042 ;
               RECT 30.214 33.206 30.266 33.242 ;
               RECT 30.214 34.406 30.266 34.442 ;
               RECT 30.214 35.606 30.266 35.642 ;
               RECT 30.214 36.806 30.266 36.842 ;
               RECT 30.214 38.006 30.266 38.042 ;
               RECT 30.214 39.206 30.266 39.242 ;
               RECT 30.214 40.406 30.266 40.442 ;
               RECT 30.214 41.606 30.266 41.642 ;
               RECT 30.214 42.806 30.266 42.842 ;
               RECT 30.214 44.006 30.266 44.042 ;
               RECT 30.214 45.206 30.266 45.242 ;
               RECT 30.214 46.406 30.266 46.442 ;
               RECT 30.214 47.606 30.266 47.642 ;
               RECT 30.214 49.422 30.266 49.458 ;
               RECT 30.214 49.662 30.266 49.698 ;
               RECT 30.214 55.422 30.266 55.458 ;
               RECT 30.214 55.662 30.266 55.698 ;
               RECT 30.214 56.726 30.266 56.762 ;
               RECT 30.214 57.926 30.266 57.962 ;
               RECT 30.214 59.126 30.266 59.162 ;
               RECT 30.214 60.326 30.266 60.362 ;
               RECT 30.214 61.526 30.266 61.562 ;
               RECT 30.214 62.726 30.266 62.762 ;
               RECT 30.214 63.926 30.266 63.962 ;
               RECT 30.214 65.126 30.266 65.162 ;
               RECT 30.214 66.326 30.266 66.362 ;
               RECT 30.214 67.526 30.266 67.562 ;
               RECT 30.214 68.726 30.266 68.762 ;
               RECT 30.214 69.926 30.266 69.962 ;
               RECT 30.214 71.126 30.266 71.162 ;
               RECT 30.214 72.326 30.266 72.362 ;
               RECT 30.214 73.526 30.266 73.562 ;
               RECT 30.214 74.726 30.266 74.762 ;
               RECT 30.214 75.926 30.266 75.962 ;
               RECT 30.214 77.126 30.266 77.162 ;
               RECT 30.214 78.326 30.266 78.362 ;
               RECT 30.214 79.526 30.266 79.562 ;
               RECT 30.214 80.726 30.266 80.762 ;
               RECT 30.214 81.926 30.266 81.962 ;
               RECT 30.214 83.126 30.266 83.162 ;
               RECT 30.214 84.326 30.266 84.362 ;
               RECT 30.214 85.526 30.266 85.562 ;
               RECT 30.214 86.726 30.266 86.762 ;
               RECT 30.214 87.926 30.266 87.962 ;
               RECT 30.214 89.126 30.266 89.162 ;
               RECT 30.214 90.326 30.266 90.362 ;
               RECT 30.214 91.526 30.266 91.562 ;
               RECT 30.214 92.726 30.266 92.762 ;
               RECT 30.214 93.926 30.266 93.962 ;
               RECT 30.214 95.126 30.266 95.162 ;
               RECT 30.214 96.326 30.266 96.362 ;
               RECT 30.214 97.526 30.266 97.562 ;
               RECT 30.214 98.726 30.266 98.762 ;
               RECT 30.214 99.926 30.266 99.962 ;
               RECT 30.214 101.126 30.266 101.162 ;
               RECT 30.214 102.326 30.266 102.362 ;
               RECT 30.214 103.526 30.266 103.562 ;
               RECT 30.294 1.558 30.346 1.594 ;
               RECT 30.294 2.758 30.346 2.794 ;
               RECT 30.294 3.958 30.346 3.994 ;
               RECT 30.294 5.158 30.346 5.194 ;
               RECT 30.294 6.358 30.346 6.394 ;
               RECT 30.294 7.558 30.346 7.594 ;
               RECT 30.294 8.758 30.346 8.794 ;
               RECT 30.294 9.958 30.346 9.994 ;
               RECT 30.294 11.158 30.346 11.194 ;
               RECT 30.294 12.358 30.346 12.394 ;
               RECT 30.294 13.558 30.346 13.594 ;
               RECT 30.294 14.758 30.346 14.794 ;
               RECT 30.294 15.958 30.346 15.994 ;
               RECT 30.294 17.158 30.346 17.194 ;
               RECT 30.294 18.358 30.346 18.394 ;
               RECT 30.294 19.558 30.346 19.594 ;
               RECT 30.294 20.758 30.346 20.794 ;
               RECT 30.294 21.958 30.346 21.994 ;
               RECT 30.294 23.158 30.346 23.194 ;
               RECT 30.294 24.358 30.346 24.394 ;
               RECT 30.294 25.558 30.346 25.594 ;
               RECT 30.294 26.758 30.346 26.794 ;
               RECT 30.294 27.958 30.346 27.994 ;
               RECT 30.294 29.158 30.346 29.194 ;
               RECT 30.294 30.358 30.346 30.394 ;
               RECT 30.294 31.558 30.346 31.594 ;
               RECT 30.294 32.758 30.346 32.794 ;
               RECT 30.294 33.958 30.346 33.994 ;
               RECT 30.294 35.158 30.346 35.194 ;
               RECT 30.294 36.358 30.346 36.394 ;
               RECT 30.294 37.558 30.346 37.594 ;
               RECT 30.294 38.758 30.346 38.794 ;
               RECT 30.294 39.958 30.346 39.994 ;
               RECT 30.294 41.158 30.346 41.194 ;
               RECT 30.294 42.358 30.346 42.394 ;
               RECT 30.294 43.558 30.346 43.594 ;
               RECT 30.294 44.758 30.346 44.794 ;
               RECT 30.294 45.958 30.346 45.994 ;
               RECT 30.294 47.158 30.346 47.194 ;
               RECT 30.294 48.358 30.346 48.394 ;
               RECT 30.294 50.142 30.346 50.178 ;
               RECT 30.294 50.382 30.346 50.418 ;
               RECT 30.294 54.702 30.346 54.738 ;
               RECT 30.294 54.942 30.346 54.978 ;
               RECT 30.294 57.478 30.346 57.514 ;
               RECT 30.294 58.678 30.346 58.714 ;
               RECT 30.294 59.878 30.346 59.914 ;
               RECT 30.294 61.078 30.346 61.114 ;
               RECT 30.294 62.278 30.346 62.314 ;
               RECT 30.294 63.478 30.346 63.514 ;
               RECT 30.294 64.678 30.346 64.714 ;
               RECT 30.294 65.878 30.346 65.914 ;
               RECT 30.294 67.078 30.346 67.114 ;
               RECT 30.294 68.278 30.346 68.314 ;
               RECT 30.294 69.478 30.346 69.514 ;
               RECT 30.294 70.678 30.346 70.714 ;
               RECT 30.294 71.878 30.346 71.914 ;
               RECT 30.294 73.078 30.346 73.114 ;
               RECT 30.294 74.278 30.346 74.314 ;
               RECT 30.294 75.478 30.346 75.514 ;
               RECT 30.294 76.678 30.346 76.714 ;
               RECT 30.294 77.878 30.346 77.914 ;
               RECT 30.294 79.078 30.346 79.114 ;
               RECT 30.294 80.278 30.346 80.314 ;
               RECT 30.294 81.478 30.346 81.514 ;
               RECT 30.294 82.678 30.346 82.714 ;
               RECT 30.294 83.878 30.346 83.914 ;
               RECT 30.294 85.078 30.346 85.114 ;
               RECT 30.294 86.278 30.346 86.314 ;
               RECT 30.294 87.478 30.346 87.514 ;
               RECT 30.294 88.678 30.346 88.714 ;
               RECT 30.294 89.878 30.346 89.914 ;
               RECT 30.294 91.078 30.346 91.114 ;
               RECT 30.294 92.278 30.346 92.314 ;
               RECT 30.294 93.478 30.346 93.514 ;
               RECT 30.294 94.678 30.346 94.714 ;
               RECT 30.294 95.878 30.346 95.914 ;
               RECT 30.294 97.078 30.346 97.114 ;
               RECT 30.294 98.278 30.346 98.314 ;
               RECT 30.294 99.478 30.346 99.514 ;
               RECT 30.294 100.678 30.346 100.714 ;
               RECT 30.294 101.878 30.346 101.914 ;
               RECT 30.294 103.078 30.346 103.114 ;
               RECT 30.294 104.278 30.346 104.314 ;
               RECT 30.374 0.281 30.426 0.317 ;
               RECT 30.374 104.803 30.426 104.839 ;
               RECT 30.454 0.806 30.506 0.842 ;
               RECT 30.454 2.006 30.506 2.042 ;
               RECT 30.454 3.206 30.506 3.242 ;
               RECT 30.454 4.406 30.506 4.442 ;
               RECT 30.454 5.606 30.506 5.642 ;
               RECT 30.454 6.806 30.506 6.842 ;
               RECT 30.454 8.006 30.506 8.042 ;
               RECT 30.454 9.206 30.506 9.242 ;
               RECT 30.454 10.406 30.506 10.442 ;
               RECT 30.454 11.606 30.506 11.642 ;
               RECT 30.454 12.806 30.506 12.842 ;
               RECT 30.454 14.006 30.506 14.042 ;
               RECT 30.454 15.206 30.506 15.242 ;
               RECT 30.454 16.406 30.506 16.442 ;
               RECT 30.454 17.606 30.506 17.642 ;
               RECT 30.454 18.806 30.506 18.842 ;
               RECT 30.454 20.006 30.506 20.042 ;
               RECT 30.454 21.206 30.506 21.242 ;
               RECT 30.454 22.406 30.506 22.442 ;
               RECT 30.454 23.606 30.506 23.642 ;
               RECT 30.454 24.806 30.506 24.842 ;
               RECT 30.454 26.006 30.506 26.042 ;
               RECT 30.454 27.206 30.506 27.242 ;
               RECT 30.454 28.406 30.506 28.442 ;
               RECT 30.454 29.606 30.506 29.642 ;
               RECT 30.454 30.806 30.506 30.842 ;
               RECT 30.454 32.006 30.506 32.042 ;
               RECT 30.454 33.206 30.506 33.242 ;
               RECT 30.454 34.406 30.506 34.442 ;
               RECT 30.454 35.606 30.506 35.642 ;
               RECT 30.454 36.806 30.506 36.842 ;
               RECT 30.454 38.006 30.506 38.042 ;
               RECT 30.454 39.206 30.506 39.242 ;
               RECT 30.454 40.406 30.506 40.442 ;
               RECT 30.454 41.606 30.506 41.642 ;
               RECT 30.454 42.806 30.506 42.842 ;
               RECT 30.454 44.006 30.506 44.042 ;
               RECT 30.454 45.206 30.506 45.242 ;
               RECT 30.454 46.406 30.506 46.442 ;
               RECT 30.454 47.606 30.506 47.642 ;
               RECT 30.454 49.422 30.506 49.458 ;
               RECT 30.454 49.662 30.506 49.698 ;
               RECT 30.454 51.102 30.506 51.138 ;
               RECT 30.454 51.582 30.506 51.618 ;
               RECT 30.454 53.502 30.506 53.538 ;
               RECT 30.454 53.982 30.506 54.018 ;
               RECT 30.454 55.422 30.506 55.458 ;
               RECT 30.454 55.662 30.506 55.698 ;
               RECT 30.454 56.726 30.506 56.762 ;
               RECT 30.454 57.926 30.506 57.962 ;
               RECT 30.454 59.126 30.506 59.162 ;
               RECT 30.454 60.326 30.506 60.362 ;
               RECT 30.454 61.526 30.506 61.562 ;
               RECT 30.454 62.726 30.506 62.762 ;
               RECT 30.454 63.926 30.506 63.962 ;
               RECT 30.454 65.126 30.506 65.162 ;
               RECT 30.454 66.326 30.506 66.362 ;
               RECT 30.454 67.526 30.506 67.562 ;
               RECT 30.454 68.726 30.506 68.762 ;
               RECT 30.454 69.926 30.506 69.962 ;
               RECT 30.454 71.126 30.506 71.162 ;
               RECT 30.454 72.326 30.506 72.362 ;
               RECT 30.454 73.526 30.506 73.562 ;
               RECT 30.454 74.726 30.506 74.762 ;
               RECT 30.454 75.926 30.506 75.962 ;
               RECT 30.454 77.126 30.506 77.162 ;
               RECT 30.454 78.326 30.506 78.362 ;
               RECT 30.454 79.526 30.506 79.562 ;
               RECT 30.454 80.726 30.506 80.762 ;
               RECT 30.454 81.926 30.506 81.962 ;
               RECT 30.454 83.126 30.506 83.162 ;
               RECT 30.454 84.326 30.506 84.362 ;
               RECT 30.454 85.526 30.506 85.562 ;
               RECT 30.454 86.726 30.506 86.762 ;
               RECT 30.454 87.926 30.506 87.962 ;
               RECT 30.454 89.126 30.506 89.162 ;
               RECT 30.454 90.326 30.506 90.362 ;
               RECT 30.454 91.526 30.506 91.562 ;
               RECT 30.454 92.726 30.506 92.762 ;
               RECT 30.454 93.926 30.506 93.962 ;
               RECT 30.454 95.126 30.506 95.162 ;
               RECT 30.454 96.326 30.506 96.362 ;
               RECT 30.454 97.526 30.506 97.562 ;
               RECT 30.454 98.726 30.506 98.762 ;
               RECT 30.454 99.926 30.506 99.962 ;
               RECT 30.454 101.126 30.506 101.162 ;
               RECT 30.454 102.326 30.506 102.362 ;
               RECT 30.454 103.526 30.506 103.562 ;
               RECT 30.534 1.558 30.586 1.594 ;
               RECT 30.534 2.758 30.586 2.794 ;
               RECT 30.534 3.958 30.586 3.994 ;
               RECT 30.534 5.158 30.586 5.194 ;
               RECT 30.534 6.358 30.586 6.394 ;
               RECT 30.534 7.558 30.586 7.594 ;
               RECT 30.534 8.758 30.586 8.794 ;
               RECT 30.534 9.958 30.586 9.994 ;
               RECT 30.534 11.158 30.586 11.194 ;
               RECT 30.534 12.358 30.586 12.394 ;
               RECT 30.534 13.558 30.586 13.594 ;
               RECT 30.534 14.758 30.586 14.794 ;
               RECT 30.534 15.958 30.586 15.994 ;
               RECT 30.534 17.158 30.586 17.194 ;
               RECT 30.534 18.358 30.586 18.394 ;
               RECT 30.534 19.558 30.586 19.594 ;
               RECT 30.534 20.758 30.586 20.794 ;
               RECT 30.534 21.958 30.586 21.994 ;
               RECT 30.534 23.158 30.586 23.194 ;
               RECT 30.534 24.358 30.586 24.394 ;
               RECT 30.534 25.558 30.586 25.594 ;
               RECT 30.534 26.758 30.586 26.794 ;
               RECT 30.534 27.958 30.586 27.994 ;
               RECT 30.534 29.158 30.586 29.194 ;
               RECT 30.534 30.358 30.586 30.394 ;
               RECT 30.534 31.558 30.586 31.594 ;
               RECT 30.534 32.758 30.586 32.794 ;
               RECT 30.534 33.958 30.586 33.994 ;
               RECT 30.534 35.158 30.586 35.194 ;
               RECT 30.534 36.358 30.586 36.394 ;
               RECT 30.534 37.558 30.586 37.594 ;
               RECT 30.534 38.758 30.586 38.794 ;
               RECT 30.534 39.958 30.586 39.994 ;
               RECT 30.534 41.158 30.586 41.194 ;
               RECT 30.534 42.358 30.586 42.394 ;
               RECT 30.534 43.558 30.586 43.594 ;
               RECT 30.534 44.758 30.586 44.794 ;
               RECT 30.534 45.958 30.586 45.994 ;
               RECT 30.534 47.158 30.586 47.194 ;
               RECT 30.534 48.358 30.586 48.394 ;
               RECT 30.534 50.142 30.586 50.178 ;
               RECT 30.534 50.382 30.586 50.418 ;
               RECT 30.534 54.702 30.586 54.738 ;
               RECT 30.534 54.942 30.586 54.978 ;
               RECT 30.534 57.478 30.586 57.514 ;
               RECT 30.534 58.678 30.586 58.714 ;
               RECT 30.534 59.878 30.586 59.914 ;
               RECT 30.534 61.078 30.586 61.114 ;
               RECT 30.534 62.278 30.586 62.314 ;
               RECT 30.534 63.478 30.586 63.514 ;
               RECT 30.534 64.678 30.586 64.714 ;
               RECT 30.534 65.878 30.586 65.914 ;
               RECT 30.534 67.078 30.586 67.114 ;
               RECT 30.534 68.278 30.586 68.314 ;
               RECT 30.534 69.478 30.586 69.514 ;
               RECT 30.534 70.678 30.586 70.714 ;
               RECT 30.534 71.878 30.586 71.914 ;
               RECT 30.534 73.078 30.586 73.114 ;
               RECT 30.534 74.278 30.586 74.314 ;
               RECT 30.534 75.478 30.586 75.514 ;
               RECT 30.534 76.678 30.586 76.714 ;
               RECT 30.534 77.878 30.586 77.914 ;
               RECT 30.534 79.078 30.586 79.114 ;
               RECT 30.534 80.278 30.586 80.314 ;
               RECT 30.534 81.478 30.586 81.514 ;
               RECT 30.534 82.678 30.586 82.714 ;
               RECT 30.534 83.878 30.586 83.914 ;
               RECT 30.534 85.078 30.586 85.114 ;
               RECT 30.534 86.278 30.586 86.314 ;
               RECT 30.534 87.478 30.586 87.514 ;
               RECT 30.534 88.678 30.586 88.714 ;
               RECT 30.534 89.878 30.586 89.914 ;
               RECT 30.534 91.078 30.586 91.114 ;
               RECT 30.534 92.278 30.586 92.314 ;
               RECT 30.534 93.478 30.586 93.514 ;
               RECT 30.534 94.678 30.586 94.714 ;
               RECT 30.534 95.878 30.586 95.914 ;
               RECT 30.534 97.078 30.586 97.114 ;
               RECT 30.534 98.278 30.586 98.314 ;
               RECT 30.534 99.478 30.586 99.514 ;
               RECT 30.534 100.678 30.586 100.714 ;
               RECT 30.534 101.878 30.586 101.914 ;
               RECT 30.534 103.078 30.586 103.114 ;
               RECT 30.534 104.278 30.586 104.314 ;
               RECT 30.614 0.806 30.666 0.842 ;
               RECT 30.614 2.006 30.666 2.042 ;
               RECT 30.614 3.206 30.666 3.242 ;
               RECT 30.614 4.406 30.666 4.442 ;
               RECT 30.614 5.606 30.666 5.642 ;
               RECT 30.614 6.806 30.666 6.842 ;
               RECT 30.614 8.006 30.666 8.042 ;
               RECT 30.614 9.206 30.666 9.242 ;
               RECT 30.614 10.406 30.666 10.442 ;
               RECT 30.614 11.606 30.666 11.642 ;
               RECT 30.614 12.806 30.666 12.842 ;
               RECT 30.614 14.006 30.666 14.042 ;
               RECT 30.614 15.206 30.666 15.242 ;
               RECT 30.614 16.406 30.666 16.442 ;
               RECT 30.614 17.606 30.666 17.642 ;
               RECT 30.614 18.806 30.666 18.842 ;
               RECT 30.614 20.006 30.666 20.042 ;
               RECT 30.614 21.206 30.666 21.242 ;
               RECT 30.614 22.406 30.666 22.442 ;
               RECT 30.614 23.606 30.666 23.642 ;
               RECT 30.614 24.806 30.666 24.842 ;
               RECT 30.614 26.006 30.666 26.042 ;
               RECT 30.614 27.206 30.666 27.242 ;
               RECT 30.614 28.406 30.666 28.442 ;
               RECT 30.614 29.606 30.666 29.642 ;
               RECT 30.614 30.806 30.666 30.842 ;
               RECT 30.614 32.006 30.666 32.042 ;
               RECT 30.614 33.206 30.666 33.242 ;
               RECT 30.614 34.406 30.666 34.442 ;
               RECT 30.614 35.606 30.666 35.642 ;
               RECT 30.614 36.806 30.666 36.842 ;
               RECT 30.614 38.006 30.666 38.042 ;
               RECT 30.614 39.206 30.666 39.242 ;
               RECT 30.614 40.406 30.666 40.442 ;
               RECT 30.614 41.606 30.666 41.642 ;
               RECT 30.614 42.806 30.666 42.842 ;
               RECT 30.614 44.006 30.666 44.042 ;
               RECT 30.614 45.206 30.666 45.242 ;
               RECT 30.614 46.406 30.666 46.442 ;
               RECT 30.614 47.606 30.666 47.642 ;
               RECT 30.614 49.422 30.666 49.458 ;
               RECT 30.614 49.662 30.666 49.698 ;
               RECT 30.614 55.422 30.666 55.458 ;
               RECT 30.614 55.662 30.666 55.698 ;
               RECT 30.614 56.726 30.666 56.762 ;
               RECT 30.614 57.926 30.666 57.962 ;
               RECT 30.614 59.126 30.666 59.162 ;
               RECT 30.614 60.326 30.666 60.362 ;
               RECT 30.614 61.526 30.666 61.562 ;
               RECT 30.614 62.726 30.666 62.762 ;
               RECT 30.614 63.926 30.666 63.962 ;
               RECT 30.614 65.126 30.666 65.162 ;
               RECT 30.614 66.326 30.666 66.362 ;
               RECT 30.614 67.526 30.666 67.562 ;
               RECT 30.614 68.726 30.666 68.762 ;
               RECT 30.614 69.926 30.666 69.962 ;
               RECT 30.614 71.126 30.666 71.162 ;
               RECT 30.614 72.326 30.666 72.362 ;
               RECT 30.614 73.526 30.666 73.562 ;
               RECT 30.614 74.726 30.666 74.762 ;
               RECT 30.614 75.926 30.666 75.962 ;
               RECT 30.614 77.126 30.666 77.162 ;
               RECT 30.614 78.326 30.666 78.362 ;
               RECT 30.614 79.526 30.666 79.562 ;
               RECT 30.614 80.726 30.666 80.762 ;
               RECT 30.614 81.926 30.666 81.962 ;
               RECT 30.614 83.126 30.666 83.162 ;
               RECT 30.614 84.326 30.666 84.362 ;
               RECT 30.614 85.526 30.666 85.562 ;
               RECT 30.614 86.726 30.666 86.762 ;
               RECT 30.614 87.926 30.666 87.962 ;
               RECT 30.614 89.126 30.666 89.162 ;
               RECT 30.614 90.326 30.666 90.362 ;
               RECT 30.614 91.526 30.666 91.562 ;
               RECT 30.614 92.726 30.666 92.762 ;
               RECT 30.614 93.926 30.666 93.962 ;
               RECT 30.614 95.126 30.666 95.162 ;
               RECT 30.614 96.326 30.666 96.362 ;
               RECT 30.614 97.526 30.666 97.562 ;
               RECT 30.614 98.726 30.666 98.762 ;
               RECT 30.614 99.926 30.666 99.962 ;
               RECT 30.614 101.126 30.666 101.162 ;
               RECT 30.614 102.326 30.666 102.362 ;
               RECT 30.614 103.526 30.666 103.562 ;
               RECT 30.694 1.558 30.746 1.594 ;
               RECT 30.694 2.758 30.746 2.794 ;
               RECT 30.694 3.958 30.746 3.994 ;
               RECT 30.694 5.158 30.746 5.194 ;
               RECT 30.694 6.358 30.746 6.394 ;
               RECT 30.694 7.558 30.746 7.594 ;
               RECT 30.694 8.758 30.746 8.794 ;
               RECT 30.694 9.958 30.746 9.994 ;
               RECT 30.694 11.158 30.746 11.194 ;
               RECT 30.694 12.358 30.746 12.394 ;
               RECT 30.694 13.558 30.746 13.594 ;
               RECT 30.694 14.758 30.746 14.794 ;
               RECT 30.694 15.958 30.746 15.994 ;
               RECT 30.694 17.158 30.746 17.194 ;
               RECT 30.694 18.358 30.746 18.394 ;
               RECT 30.694 19.558 30.746 19.594 ;
               RECT 30.694 20.758 30.746 20.794 ;
               RECT 30.694 21.958 30.746 21.994 ;
               RECT 30.694 23.158 30.746 23.194 ;
               RECT 30.694 24.358 30.746 24.394 ;
               RECT 30.694 25.558 30.746 25.594 ;
               RECT 30.694 26.758 30.746 26.794 ;
               RECT 30.694 27.958 30.746 27.994 ;
               RECT 30.694 29.158 30.746 29.194 ;
               RECT 30.694 30.358 30.746 30.394 ;
               RECT 30.694 31.558 30.746 31.594 ;
               RECT 30.694 32.758 30.746 32.794 ;
               RECT 30.694 33.958 30.746 33.994 ;
               RECT 30.694 35.158 30.746 35.194 ;
               RECT 30.694 36.358 30.746 36.394 ;
               RECT 30.694 37.558 30.746 37.594 ;
               RECT 30.694 38.758 30.746 38.794 ;
               RECT 30.694 39.958 30.746 39.994 ;
               RECT 30.694 41.158 30.746 41.194 ;
               RECT 30.694 42.358 30.746 42.394 ;
               RECT 30.694 43.558 30.746 43.594 ;
               RECT 30.694 44.758 30.746 44.794 ;
               RECT 30.694 45.958 30.746 45.994 ;
               RECT 30.694 47.158 30.746 47.194 ;
               RECT 30.694 48.358 30.746 48.394 ;
               RECT 30.694 50.142 30.746 50.178 ;
               RECT 30.694 50.382 30.746 50.418 ;
               RECT 30.694 54.702 30.746 54.738 ;
               RECT 30.694 54.942 30.746 54.978 ;
               RECT 30.694 57.478 30.746 57.514 ;
               RECT 30.694 58.678 30.746 58.714 ;
               RECT 30.694 59.878 30.746 59.914 ;
               RECT 30.694 61.078 30.746 61.114 ;
               RECT 30.694 62.278 30.746 62.314 ;
               RECT 30.694 63.478 30.746 63.514 ;
               RECT 30.694 64.678 30.746 64.714 ;
               RECT 30.694 65.878 30.746 65.914 ;
               RECT 30.694 67.078 30.746 67.114 ;
               RECT 30.694 68.278 30.746 68.314 ;
               RECT 30.694 69.478 30.746 69.514 ;
               RECT 30.694 70.678 30.746 70.714 ;
               RECT 30.694 71.878 30.746 71.914 ;
               RECT 30.694 73.078 30.746 73.114 ;
               RECT 30.694 74.278 30.746 74.314 ;
               RECT 30.694 75.478 30.746 75.514 ;
               RECT 30.694 76.678 30.746 76.714 ;
               RECT 30.694 77.878 30.746 77.914 ;
               RECT 30.694 79.078 30.746 79.114 ;
               RECT 30.694 80.278 30.746 80.314 ;
               RECT 30.694 81.478 30.746 81.514 ;
               RECT 30.694 82.678 30.746 82.714 ;
               RECT 30.694 83.878 30.746 83.914 ;
               RECT 30.694 85.078 30.746 85.114 ;
               RECT 30.694 86.278 30.746 86.314 ;
               RECT 30.694 87.478 30.746 87.514 ;
               RECT 30.694 88.678 30.746 88.714 ;
               RECT 30.694 89.878 30.746 89.914 ;
               RECT 30.694 91.078 30.746 91.114 ;
               RECT 30.694 92.278 30.746 92.314 ;
               RECT 30.694 93.478 30.746 93.514 ;
               RECT 30.694 94.678 30.746 94.714 ;
               RECT 30.694 95.878 30.746 95.914 ;
               RECT 30.694 97.078 30.746 97.114 ;
               RECT 30.694 98.278 30.746 98.314 ;
               RECT 30.694 99.478 30.746 99.514 ;
               RECT 30.694 100.678 30.746 100.714 ;
               RECT 30.694 101.878 30.746 101.914 ;
               RECT 30.694 103.078 30.746 103.114 ;
               RECT 30.694 104.278 30.746 104.314 ;
               RECT 30.774 0.281 30.826 0.317 ;
               RECT 30.774 104.803 30.826 104.839 ;
               RECT 30.854 0.806 30.906 0.842 ;
               RECT 30.854 2.006 30.906 2.042 ;
               RECT 30.854 3.206 30.906 3.242 ;
               RECT 30.854 4.406 30.906 4.442 ;
               RECT 30.854 5.606 30.906 5.642 ;
               RECT 30.854 6.806 30.906 6.842 ;
               RECT 30.854 8.006 30.906 8.042 ;
               RECT 30.854 9.206 30.906 9.242 ;
               RECT 30.854 10.406 30.906 10.442 ;
               RECT 30.854 11.606 30.906 11.642 ;
               RECT 30.854 12.806 30.906 12.842 ;
               RECT 30.854 14.006 30.906 14.042 ;
               RECT 30.854 15.206 30.906 15.242 ;
               RECT 30.854 16.406 30.906 16.442 ;
               RECT 30.854 17.606 30.906 17.642 ;
               RECT 30.854 18.806 30.906 18.842 ;
               RECT 30.854 20.006 30.906 20.042 ;
               RECT 30.854 21.206 30.906 21.242 ;
               RECT 30.854 22.406 30.906 22.442 ;
               RECT 30.854 23.606 30.906 23.642 ;
               RECT 30.854 24.806 30.906 24.842 ;
               RECT 30.854 26.006 30.906 26.042 ;
               RECT 30.854 27.206 30.906 27.242 ;
               RECT 30.854 28.406 30.906 28.442 ;
               RECT 30.854 29.606 30.906 29.642 ;
               RECT 30.854 30.806 30.906 30.842 ;
               RECT 30.854 32.006 30.906 32.042 ;
               RECT 30.854 33.206 30.906 33.242 ;
               RECT 30.854 34.406 30.906 34.442 ;
               RECT 30.854 35.606 30.906 35.642 ;
               RECT 30.854 36.806 30.906 36.842 ;
               RECT 30.854 38.006 30.906 38.042 ;
               RECT 30.854 39.206 30.906 39.242 ;
               RECT 30.854 40.406 30.906 40.442 ;
               RECT 30.854 41.606 30.906 41.642 ;
               RECT 30.854 42.806 30.906 42.842 ;
               RECT 30.854 44.006 30.906 44.042 ;
               RECT 30.854 45.206 30.906 45.242 ;
               RECT 30.854 46.406 30.906 46.442 ;
               RECT 30.854 47.606 30.906 47.642 ;
               RECT 30.854 49.422 30.906 49.458 ;
               RECT 30.854 49.662 30.906 49.698 ;
               RECT 30.854 55.422 30.906 55.458 ;
               RECT 30.854 55.662 30.906 55.698 ;
               RECT 30.854 56.726 30.906 56.762 ;
               RECT 30.854 57.926 30.906 57.962 ;
               RECT 30.854 59.126 30.906 59.162 ;
               RECT 30.854 60.326 30.906 60.362 ;
               RECT 30.854 61.526 30.906 61.562 ;
               RECT 30.854 62.726 30.906 62.762 ;
               RECT 30.854 63.926 30.906 63.962 ;
               RECT 30.854 65.126 30.906 65.162 ;
               RECT 30.854 66.326 30.906 66.362 ;
               RECT 30.854 67.526 30.906 67.562 ;
               RECT 30.854 68.726 30.906 68.762 ;
               RECT 30.854 69.926 30.906 69.962 ;
               RECT 30.854 71.126 30.906 71.162 ;
               RECT 30.854 72.326 30.906 72.362 ;
               RECT 30.854 73.526 30.906 73.562 ;
               RECT 30.854 74.726 30.906 74.762 ;
               RECT 30.854 75.926 30.906 75.962 ;
               RECT 30.854 77.126 30.906 77.162 ;
               RECT 30.854 78.326 30.906 78.362 ;
               RECT 30.854 79.526 30.906 79.562 ;
               RECT 30.854 80.726 30.906 80.762 ;
               RECT 30.854 81.926 30.906 81.962 ;
               RECT 30.854 83.126 30.906 83.162 ;
               RECT 30.854 84.326 30.906 84.362 ;
               RECT 30.854 85.526 30.906 85.562 ;
               RECT 30.854 86.726 30.906 86.762 ;
               RECT 30.854 87.926 30.906 87.962 ;
               RECT 30.854 89.126 30.906 89.162 ;
               RECT 30.854 90.326 30.906 90.362 ;
               RECT 30.854 91.526 30.906 91.562 ;
               RECT 30.854 92.726 30.906 92.762 ;
               RECT 30.854 93.926 30.906 93.962 ;
               RECT 30.854 95.126 30.906 95.162 ;
               RECT 30.854 96.326 30.906 96.362 ;
               RECT 30.854 97.526 30.906 97.562 ;
               RECT 30.854 98.726 30.906 98.762 ;
               RECT 30.854 99.926 30.906 99.962 ;
               RECT 30.854 101.126 30.906 101.162 ;
               RECT 30.854 102.326 30.906 102.362 ;
               RECT 30.854 103.526 30.906 103.562 ;
               RECT 30.934 1.558 30.986 1.594 ;
               RECT 30.934 2.758 30.986 2.794 ;
               RECT 30.934 3.958 30.986 3.994 ;
               RECT 30.934 5.158 30.986 5.194 ;
               RECT 30.934 6.358 30.986 6.394 ;
               RECT 30.934 7.558 30.986 7.594 ;
               RECT 30.934 8.758 30.986 8.794 ;
               RECT 30.934 9.958 30.986 9.994 ;
               RECT 30.934 11.158 30.986 11.194 ;
               RECT 30.934 12.358 30.986 12.394 ;
               RECT 30.934 13.558 30.986 13.594 ;
               RECT 30.934 14.758 30.986 14.794 ;
               RECT 30.934 15.958 30.986 15.994 ;
               RECT 30.934 17.158 30.986 17.194 ;
               RECT 30.934 18.358 30.986 18.394 ;
               RECT 30.934 19.558 30.986 19.594 ;
               RECT 30.934 20.758 30.986 20.794 ;
               RECT 30.934 21.958 30.986 21.994 ;
               RECT 30.934 23.158 30.986 23.194 ;
               RECT 30.934 24.358 30.986 24.394 ;
               RECT 30.934 25.558 30.986 25.594 ;
               RECT 30.934 26.758 30.986 26.794 ;
               RECT 30.934 27.958 30.986 27.994 ;
               RECT 30.934 29.158 30.986 29.194 ;
               RECT 30.934 30.358 30.986 30.394 ;
               RECT 30.934 31.558 30.986 31.594 ;
               RECT 30.934 32.758 30.986 32.794 ;
               RECT 30.934 33.958 30.986 33.994 ;
               RECT 30.934 35.158 30.986 35.194 ;
               RECT 30.934 36.358 30.986 36.394 ;
               RECT 30.934 37.558 30.986 37.594 ;
               RECT 30.934 38.758 30.986 38.794 ;
               RECT 30.934 39.958 30.986 39.994 ;
               RECT 30.934 41.158 30.986 41.194 ;
               RECT 30.934 42.358 30.986 42.394 ;
               RECT 30.934 43.558 30.986 43.594 ;
               RECT 30.934 44.758 30.986 44.794 ;
               RECT 30.934 45.958 30.986 45.994 ;
               RECT 30.934 47.158 30.986 47.194 ;
               RECT 30.934 48.358 30.986 48.394 ;
               RECT 30.934 50.142 30.986 50.178 ;
               RECT 30.934 50.382 30.986 50.418 ;
               RECT 30.934 54.702 30.986 54.738 ;
               RECT 30.934 54.942 30.986 54.978 ;
               RECT 30.934 57.478 30.986 57.514 ;
               RECT 30.934 58.678 30.986 58.714 ;
               RECT 30.934 59.878 30.986 59.914 ;
               RECT 30.934 61.078 30.986 61.114 ;
               RECT 30.934 62.278 30.986 62.314 ;
               RECT 30.934 63.478 30.986 63.514 ;
               RECT 30.934 64.678 30.986 64.714 ;
               RECT 30.934 65.878 30.986 65.914 ;
               RECT 30.934 67.078 30.986 67.114 ;
               RECT 30.934 68.278 30.986 68.314 ;
               RECT 30.934 69.478 30.986 69.514 ;
               RECT 30.934 70.678 30.986 70.714 ;
               RECT 30.934 71.878 30.986 71.914 ;
               RECT 30.934 73.078 30.986 73.114 ;
               RECT 30.934 74.278 30.986 74.314 ;
               RECT 30.934 75.478 30.986 75.514 ;
               RECT 30.934 76.678 30.986 76.714 ;
               RECT 30.934 77.878 30.986 77.914 ;
               RECT 30.934 79.078 30.986 79.114 ;
               RECT 30.934 80.278 30.986 80.314 ;
               RECT 30.934 81.478 30.986 81.514 ;
               RECT 30.934 82.678 30.986 82.714 ;
               RECT 30.934 83.878 30.986 83.914 ;
               RECT 30.934 85.078 30.986 85.114 ;
               RECT 30.934 86.278 30.986 86.314 ;
               RECT 30.934 87.478 30.986 87.514 ;
               RECT 30.934 88.678 30.986 88.714 ;
               RECT 30.934 89.878 30.986 89.914 ;
               RECT 30.934 91.078 30.986 91.114 ;
               RECT 30.934 92.278 30.986 92.314 ;
               RECT 30.934 93.478 30.986 93.514 ;
               RECT 30.934 94.678 30.986 94.714 ;
               RECT 30.934 95.878 30.986 95.914 ;
               RECT 30.934 97.078 30.986 97.114 ;
               RECT 30.934 98.278 30.986 98.314 ;
               RECT 30.934 99.478 30.986 99.514 ;
               RECT 30.934 100.678 30.986 100.714 ;
               RECT 30.934 101.878 30.986 101.914 ;
               RECT 30.934 103.078 30.986 103.114 ;
               RECT 30.934 104.278 30.986 104.314 ;
               RECT 31.014 0.806 31.066 0.842 ;
               RECT 31.014 2.006 31.066 2.042 ;
               RECT 31.014 3.206 31.066 3.242 ;
               RECT 31.014 4.406 31.066 4.442 ;
               RECT 31.014 5.606 31.066 5.642 ;
               RECT 31.014 6.806 31.066 6.842 ;
               RECT 31.014 8.006 31.066 8.042 ;
               RECT 31.014 9.206 31.066 9.242 ;
               RECT 31.014 10.406 31.066 10.442 ;
               RECT 31.014 11.606 31.066 11.642 ;
               RECT 31.014 12.806 31.066 12.842 ;
               RECT 31.014 14.006 31.066 14.042 ;
               RECT 31.014 15.206 31.066 15.242 ;
               RECT 31.014 16.406 31.066 16.442 ;
               RECT 31.014 17.606 31.066 17.642 ;
               RECT 31.014 18.806 31.066 18.842 ;
               RECT 31.014 20.006 31.066 20.042 ;
               RECT 31.014 21.206 31.066 21.242 ;
               RECT 31.014 22.406 31.066 22.442 ;
               RECT 31.014 23.606 31.066 23.642 ;
               RECT 31.014 24.806 31.066 24.842 ;
               RECT 31.014 26.006 31.066 26.042 ;
               RECT 31.014 27.206 31.066 27.242 ;
               RECT 31.014 28.406 31.066 28.442 ;
               RECT 31.014 29.606 31.066 29.642 ;
               RECT 31.014 30.806 31.066 30.842 ;
               RECT 31.014 32.006 31.066 32.042 ;
               RECT 31.014 33.206 31.066 33.242 ;
               RECT 31.014 34.406 31.066 34.442 ;
               RECT 31.014 35.606 31.066 35.642 ;
               RECT 31.014 36.806 31.066 36.842 ;
               RECT 31.014 38.006 31.066 38.042 ;
               RECT 31.014 39.206 31.066 39.242 ;
               RECT 31.014 40.406 31.066 40.442 ;
               RECT 31.014 41.606 31.066 41.642 ;
               RECT 31.014 42.806 31.066 42.842 ;
               RECT 31.014 44.006 31.066 44.042 ;
               RECT 31.014 45.206 31.066 45.242 ;
               RECT 31.014 46.406 31.066 46.442 ;
               RECT 31.014 47.606 31.066 47.642 ;
               RECT 31.014 49.422 31.066 49.458 ;
               RECT 31.014 49.662 31.066 49.698 ;
               RECT 31.014 55.422 31.066 55.458 ;
               RECT 31.014 55.662 31.066 55.698 ;
               RECT 31.014 56.726 31.066 56.762 ;
               RECT 31.014 57.926 31.066 57.962 ;
               RECT 31.014 59.126 31.066 59.162 ;
               RECT 31.014 60.326 31.066 60.362 ;
               RECT 31.014 61.526 31.066 61.562 ;
               RECT 31.014 62.726 31.066 62.762 ;
               RECT 31.014 63.926 31.066 63.962 ;
               RECT 31.014 65.126 31.066 65.162 ;
               RECT 31.014 66.326 31.066 66.362 ;
               RECT 31.014 67.526 31.066 67.562 ;
               RECT 31.014 68.726 31.066 68.762 ;
               RECT 31.014 69.926 31.066 69.962 ;
               RECT 31.014 71.126 31.066 71.162 ;
               RECT 31.014 72.326 31.066 72.362 ;
               RECT 31.014 73.526 31.066 73.562 ;
               RECT 31.014 74.726 31.066 74.762 ;
               RECT 31.014 75.926 31.066 75.962 ;
               RECT 31.014 77.126 31.066 77.162 ;
               RECT 31.014 78.326 31.066 78.362 ;
               RECT 31.014 79.526 31.066 79.562 ;
               RECT 31.014 80.726 31.066 80.762 ;
               RECT 31.014 81.926 31.066 81.962 ;
               RECT 31.014 83.126 31.066 83.162 ;
               RECT 31.014 84.326 31.066 84.362 ;
               RECT 31.014 85.526 31.066 85.562 ;
               RECT 31.014 86.726 31.066 86.762 ;
               RECT 31.014 87.926 31.066 87.962 ;
               RECT 31.014 89.126 31.066 89.162 ;
               RECT 31.014 90.326 31.066 90.362 ;
               RECT 31.014 91.526 31.066 91.562 ;
               RECT 31.014 92.726 31.066 92.762 ;
               RECT 31.014 93.926 31.066 93.962 ;
               RECT 31.014 95.126 31.066 95.162 ;
               RECT 31.014 96.326 31.066 96.362 ;
               RECT 31.014 97.526 31.066 97.562 ;
               RECT 31.014 98.726 31.066 98.762 ;
               RECT 31.014 99.926 31.066 99.962 ;
               RECT 31.014 101.126 31.066 101.162 ;
               RECT 31.014 102.326 31.066 102.362 ;
               RECT 31.014 103.526 31.066 103.562 ;
               RECT 31.094 1.558 31.146 1.594 ;
               RECT 31.094 2.758 31.146 2.794 ;
               RECT 31.094 3.958 31.146 3.994 ;
               RECT 31.094 5.158 31.146 5.194 ;
               RECT 31.094 6.358 31.146 6.394 ;
               RECT 31.094 7.558 31.146 7.594 ;
               RECT 31.094 8.758 31.146 8.794 ;
               RECT 31.094 9.958 31.146 9.994 ;
               RECT 31.094 11.158 31.146 11.194 ;
               RECT 31.094 12.358 31.146 12.394 ;
               RECT 31.094 13.558 31.146 13.594 ;
               RECT 31.094 14.758 31.146 14.794 ;
               RECT 31.094 15.958 31.146 15.994 ;
               RECT 31.094 17.158 31.146 17.194 ;
               RECT 31.094 18.358 31.146 18.394 ;
               RECT 31.094 19.558 31.146 19.594 ;
               RECT 31.094 20.758 31.146 20.794 ;
               RECT 31.094 21.958 31.146 21.994 ;
               RECT 31.094 23.158 31.146 23.194 ;
               RECT 31.094 24.358 31.146 24.394 ;
               RECT 31.094 25.558 31.146 25.594 ;
               RECT 31.094 26.758 31.146 26.794 ;
               RECT 31.094 27.958 31.146 27.994 ;
               RECT 31.094 29.158 31.146 29.194 ;
               RECT 31.094 30.358 31.146 30.394 ;
               RECT 31.094 31.558 31.146 31.594 ;
               RECT 31.094 32.758 31.146 32.794 ;
               RECT 31.094 33.958 31.146 33.994 ;
               RECT 31.094 35.158 31.146 35.194 ;
               RECT 31.094 36.358 31.146 36.394 ;
               RECT 31.094 37.558 31.146 37.594 ;
               RECT 31.094 38.758 31.146 38.794 ;
               RECT 31.094 39.958 31.146 39.994 ;
               RECT 31.094 41.158 31.146 41.194 ;
               RECT 31.094 42.358 31.146 42.394 ;
               RECT 31.094 43.558 31.146 43.594 ;
               RECT 31.094 44.758 31.146 44.794 ;
               RECT 31.094 45.958 31.146 45.994 ;
               RECT 31.094 47.158 31.146 47.194 ;
               RECT 31.094 48.358 31.146 48.394 ;
               RECT 31.094 50.142 31.146 50.178 ;
               RECT 31.094 50.382 31.146 50.418 ;
               RECT 31.094 54.702 31.146 54.738 ;
               RECT 31.094 54.942 31.146 54.978 ;
               RECT 31.094 57.478 31.146 57.514 ;
               RECT 31.094 58.678 31.146 58.714 ;
               RECT 31.094 59.878 31.146 59.914 ;
               RECT 31.094 61.078 31.146 61.114 ;
               RECT 31.094 62.278 31.146 62.314 ;
               RECT 31.094 63.478 31.146 63.514 ;
               RECT 31.094 64.678 31.146 64.714 ;
               RECT 31.094 65.878 31.146 65.914 ;
               RECT 31.094 67.078 31.146 67.114 ;
               RECT 31.094 68.278 31.146 68.314 ;
               RECT 31.094 69.478 31.146 69.514 ;
               RECT 31.094 70.678 31.146 70.714 ;
               RECT 31.094 71.878 31.146 71.914 ;
               RECT 31.094 73.078 31.146 73.114 ;
               RECT 31.094 74.278 31.146 74.314 ;
               RECT 31.094 75.478 31.146 75.514 ;
               RECT 31.094 76.678 31.146 76.714 ;
               RECT 31.094 77.878 31.146 77.914 ;
               RECT 31.094 79.078 31.146 79.114 ;
               RECT 31.094 80.278 31.146 80.314 ;
               RECT 31.094 81.478 31.146 81.514 ;
               RECT 31.094 82.678 31.146 82.714 ;
               RECT 31.094 83.878 31.146 83.914 ;
               RECT 31.094 85.078 31.146 85.114 ;
               RECT 31.094 86.278 31.146 86.314 ;
               RECT 31.094 87.478 31.146 87.514 ;
               RECT 31.094 88.678 31.146 88.714 ;
               RECT 31.094 89.878 31.146 89.914 ;
               RECT 31.094 91.078 31.146 91.114 ;
               RECT 31.094 92.278 31.146 92.314 ;
               RECT 31.094 93.478 31.146 93.514 ;
               RECT 31.094 94.678 31.146 94.714 ;
               RECT 31.094 95.878 31.146 95.914 ;
               RECT 31.094 97.078 31.146 97.114 ;
               RECT 31.094 98.278 31.146 98.314 ;
               RECT 31.094 99.478 31.146 99.514 ;
               RECT 31.094 100.678 31.146 100.714 ;
               RECT 31.094 101.878 31.146 101.914 ;
               RECT 31.094 103.078 31.146 103.114 ;
               RECT 31.094 104.278 31.146 104.314 ;
               RECT 31.174 0.281 31.226 0.317 ;
               RECT 31.174 104.803 31.226 104.839 ;
               RECT 31.254 0.806 31.306 0.842 ;
               RECT 31.254 2.006 31.306 2.042 ;
               RECT 31.254 3.206 31.306 3.242 ;
               RECT 31.254 4.406 31.306 4.442 ;
               RECT 31.254 5.606 31.306 5.642 ;
               RECT 31.254 6.806 31.306 6.842 ;
               RECT 31.254 8.006 31.306 8.042 ;
               RECT 31.254 9.206 31.306 9.242 ;
               RECT 31.254 10.406 31.306 10.442 ;
               RECT 31.254 11.606 31.306 11.642 ;
               RECT 31.254 12.806 31.306 12.842 ;
               RECT 31.254 14.006 31.306 14.042 ;
               RECT 31.254 15.206 31.306 15.242 ;
               RECT 31.254 16.406 31.306 16.442 ;
               RECT 31.254 17.606 31.306 17.642 ;
               RECT 31.254 18.806 31.306 18.842 ;
               RECT 31.254 20.006 31.306 20.042 ;
               RECT 31.254 21.206 31.306 21.242 ;
               RECT 31.254 22.406 31.306 22.442 ;
               RECT 31.254 23.606 31.306 23.642 ;
               RECT 31.254 24.806 31.306 24.842 ;
               RECT 31.254 26.006 31.306 26.042 ;
               RECT 31.254 27.206 31.306 27.242 ;
               RECT 31.254 28.406 31.306 28.442 ;
               RECT 31.254 29.606 31.306 29.642 ;
               RECT 31.254 30.806 31.306 30.842 ;
               RECT 31.254 32.006 31.306 32.042 ;
               RECT 31.254 33.206 31.306 33.242 ;
               RECT 31.254 34.406 31.306 34.442 ;
               RECT 31.254 35.606 31.306 35.642 ;
               RECT 31.254 36.806 31.306 36.842 ;
               RECT 31.254 38.006 31.306 38.042 ;
               RECT 31.254 39.206 31.306 39.242 ;
               RECT 31.254 40.406 31.306 40.442 ;
               RECT 31.254 41.606 31.306 41.642 ;
               RECT 31.254 42.806 31.306 42.842 ;
               RECT 31.254 44.006 31.306 44.042 ;
               RECT 31.254 45.206 31.306 45.242 ;
               RECT 31.254 46.406 31.306 46.442 ;
               RECT 31.254 47.606 31.306 47.642 ;
               RECT 31.254 49.422 31.306 49.458 ;
               RECT 31.254 49.662 31.306 49.698 ;
               RECT 31.254 51.102 31.306 51.138 ;
               RECT 31.254 51.582 31.306 51.618 ;
               RECT 31.254 53.502 31.306 53.538 ;
               RECT 31.254 53.982 31.306 54.018 ;
               RECT 31.254 55.422 31.306 55.458 ;
               RECT 31.254 55.662 31.306 55.698 ;
               RECT 31.254 56.726 31.306 56.762 ;
               RECT 31.254 57.926 31.306 57.962 ;
               RECT 31.254 59.126 31.306 59.162 ;
               RECT 31.254 60.326 31.306 60.362 ;
               RECT 31.254 61.526 31.306 61.562 ;
               RECT 31.254 62.726 31.306 62.762 ;
               RECT 31.254 63.926 31.306 63.962 ;
               RECT 31.254 65.126 31.306 65.162 ;
               RECT 31.254 66.326 31.306 66.362 ;
               RECT 31.254 67.526 31.306 67.562 ;
               RECT 31.254 68.726 31.306 68.762 ;
               RECT 31.254 69.926 31.306 69.962 ;
               RECT 31.254 71.126 31.306 71.162 ;
               RECT 31.254 72.326 31.306 72.362 ;
               RECT 31.254 73.526 31.306 73.562 ;
               RECT 31.254 74.726 31.306 74.762 ;
               RECT 31.254 75.926 31.306 75.962 ;
               RECT 31.254 77.126 31.306 77.162 ;
               RECT 31.254 78.326 31.306 78.362 ;
               RECT 31.254 79.526 31.306 79.562 ;
               RECT 31.254 80.726 31.306 80.762 ;
               RECT 31.254 81.926 31.306 81.962 ;
               RECT 31.254 83.126 31.306 83.162 ;
               RECT 31.254 84.326 31.306 84.362 ;
               RECT 31.254 85.526 31.306 85.562 ;
               RECT 31.254 86.726 31.306 86.762 ;
               RECT 31.254 87.926 31.306 87.962 ;
               RECT 31.254 89.126 31.306 89.162 ;
               RECT 31.254 90.326 31.306 90.362 ;
               RECT 31.254 91.526 31.306 91.562 ;
               RECT 31.254 92.726 31.306 92.762 ;
               RECT 31.254 93.926 31.306 93.962 ;
               RECT 31.254 95.126 31.306 95.162 ;
               RECT 31.254 96.326 31.306 96.362 ;
               RECT 31.254 97.526 31.306 97.562 ;
               RECT 31.254 98.726 31.306 98.762 ;
               RECT 31.254 99.926 31.306 99.962 ;
               RECT 31.254 101.126 31.306 101.162 ;
               RECT 31.254 102.326 31.306 102.362 ;
               RECT 31.254 103.526 31.306 103.562 ;
               RECT 31.334 1.558 31.386 1.594 ;
               RECT 31.334 2.758 31.386 2.794 ;
               RECT 31.334 3.958 31.386 3.994 ;
               RECT 31.334 5.158 31.386 5.194 ;
               RECT 31.334 6.358 31.386 6.394 ;
               RECT 31.334 7.558 31.386 7.594 ;
               RECT 31.334 8.758 31.386 8.794 ;
               RECT 31.334 9.958 31.386 9.994 ;
               RECT 31.334 11.158 31.386 11.194 ;
               RECT 31.334 12.358 31.386 12.394 ;
               RECT 31.334 13.558 31.386 13.594 ;
               RECT 31.334 14.758 31.386 14.794 ;
               RECT 31.334 15.958 31.386 15.994 ;
               RECT 31.334 17.158 31.386 17.194 ;
               RECT 31.334 18.358 31.386 18.394 ;
               RECT 31.334 19.558 31.386 19.594 ;
               RECT 31.334 20.758 31.386 20.794 ;
               RECT 31.334 21.958 31.386 21.994 ;
               RECT 31.334 23.158 31.386 23.194 ;
               RECT 31.334 24.358 31.386 24.394 ;
               RECT 31.334 25.558 31.386 25.594 ;
               RECT 31.334 26.758 31.386 26.794 ;
               RECT 31.334 27.958 31.386 27.994 ;
               RECT 31.334 29.158 31.386 29.194 ;
               RECT 31.334 30.358 31.386 30.394 ;
               RECT 31.334 31.558 31.386 31.594 ;
               RECT 31.334 32.758 31.386 32.794 ;
               RECT 31.334 33.958 31.386 33.994 ;
               RECT 31.334 35.158 31.386 35.194 ;
               RECT 31.334 36.358 31.386 36.394 ;
               RECT 31.334 37.558 31.386 37.594 ;
               RECT 31.334 38.758 31.386 38.794 ;
               RECT 31.334 39.958 31.386 39.994 ;
               RECT 31.334 41.158 31.386 41.194 ;
               RECT 31.334 42.358 31.386 42.394 ;
               RECT 31.334 43.558 31.386 43.594 ;
               RECT 31.334 44.758 31.386 44.794 ;
               RECT 31.334 45.958 31.386 45.994 ;
               RECT 31.334 47.158 31.386 47.194 ;
               RECT 31.334 48.358 31.386 48.394 ;
               RECT 31.334 50.142 31.386 50.178 ;
               RECT 31.334 50.382 31.386 50.418 ;
               RECT 31.334 54.702 31.386 54.738 ;
               RECT 31.334 54.942 31.386 54.978 ;
               RECT 31.334 57.478 31.386 57.514 ;
               RECT 31.334 58.678 31.386 58.714 ;
               RECT 31.334 59.878 31.386 59.914 ;
               RECT 31.334 61.078 31.386 61.114 ;
               RECT 31.334 62.278 31.386 62.314 ;
               RECT 31.334 63.478 31.386 63.514 ;
               RECT 31.334 64.678 31.386 64.714 ;
               RECT 31.334 65.878 31.386 65.914 ;
               RECT 31.334 67.078 31.386 67.114 ;
               RECT 31.334 68.278 31.386 68.314 ;
               RECT 31.334 69.478 31.386 69.514 ;
               RECT 31.334 70.678 31.386 70.714 ;
               RECT 31.334 71.878 31.386 71.914 ;
               RECT 31.334 73.078 31.386 73.114 ;
               RECT 31.334 74.278 31.386 74.314 ;
               RECT 31.334 75.478 31.386 75.514 ;
               RECT 31.334 76.678 31.386 76.714 ;
               RECT 31.334 77.878 31.386 77.914 ;
               RECT 31.334 79.078 31.386 79.114 ;
               RECT 31.334 80.278 31.386 80.314 ;
               RECT 31.334 81.478 31.386 81.514 ;
               RECT 31.334 82.678 31.386 82.714 ;
               RECT 31.334 83.878 31.386 83.914 ;
               RECT 31.334 85.078 31.386 85.114 ;
               RECT 31.334 86.278 31.386 86.314 ;
               RECT 31.334 87.478 31.386 87.514 ;
               RECT 31.334 88.678 31.386 88.714 ;
               RECT 31.334 89.878 31.386 89.914 ;
               RECT 31.334 91.078 31.386 91.114 ;
               RECT 31.334 92.278 31.386 92.314 ;
               RECT 31.334 93.478 31.386 93.514 ;
               RECT 31.334 94.678 31.386 94.714 ;
               RECT 31.334 95.878 31.386 95.914 ;
               RECT 31.334 97.078 31.386 97.114 ;
               RECT 31.334 98.278 31.386 98.314 ;
               RECT 31.334 99.478 31.386 99.514 ;
               RECT 31.334 100.678 31.386 100.714 ;
               RECT 31.334 101.878 31.386 101.914 ;
               RECT 31.334 103.078 31.386 103.114 ;
               RECT 31.334 104.278 31.386 104.314 ;
               RECT 31.414 0.806 31.466 0.842 ;
               RECT 31.414 2.006 31.466 2.042 ;
               RECT 31.414 3.206 31.466 3.242 ;
               RECT 31.414 4.406 31.466 4.442 ;
               RECT 31.414 5.606 31.466 5.642 ;
               RECT 31.414 6.806 31.466 6.842 ;
               RECT 31.414 8.006 31.466 8.042 ;
               RECT 31.414 9.206 31.466 9.242 ;
               RECT 31.414 10.406 31.466 10.442 ;
               RECT 31.414 11.606 31.466 11.642 ;
               RECT 31.414 12.806 31.466 12.842 ;
               RECT 31.414 14.006 31.466 14.042 ;
               RECT 31.414 15.206 31.466 15.242 ;
               RECT 31.414 16.406 31.466 16.442 ;
               RECT 31.414 17.606 31.466 17.642 ;
               RECT 31.414 18.806 31.466 18.842 ;
               RECT 31.414 20.006 31.466 20.042 ;
               RECT 31.414 21.206 31.466 21.242 ;
               RECT 31.414 22.406 31.466 22.442 ;
               RECT 31.414 23.606 31.466 23.642 ;
               RECT 31.414 24.806 31.466 24.842 ;
               RECT 31.414 26.006 31.466 26.042 ;
               RECT 31.414 27.206 31.466 27.242 ;
               RECT 31.414 28.406 31.466 28.442 ;
               RECT 31.414 29.606 31.466 29.642 ;
               RECT 31.414 30.806 31.466 30.842 ;
               RECT 31.414 32.006 31.466 32.042 ;
               RECT 31.414 33.206 31.466 33.242 ;
               RECT 31.414 34.406 31.466 34.442 ;
               RECT 31.414 35.606 31.466 35.642 ;
               RECT 31.414 36.806 31.466 36.842 ;
               RECT 31.414 38.006 31.466 38.042 ;
               RECT 31.414 39.206 31.466 39.242 ;
               RECT 31.414 40.406 31.466 40.442 ;
               RECT 31.414 41.606 31.466 41.642 ;
               RECT 31.414 42.806 31.466 42.842 ;
               RECT 31.414 44.006 31.466 44.042 ;
               RECT 31.414 45.206 31.466 45.242 ;
               RECT 31.414 46.406 31.466 46.442 ;
               RECT 31.414 47.606 31.466 47.642 ;
               RECT 31.414 49.422 31.466 49.458 ;
               RECT 31.414 49.662 31.466 49.698 ;
               RECT 31.414 55.422 31.466 55.458 ;
               RECT 31.414 55.662 31.466 55.698 ;
               RECT 31.414 56.726 31.466 56.762 ;
               RECT 31.414 57.926 31.466 57.962 ;
               RECT 31.414 59.126 31.466 59.162 ;
               RECT 31.414 60.326 31.466 60.362 ;
               RECT 31.414 61.526 31.466 61.562 ;
               RECT 31.414 62.726 31.466 62.762 ;
               RECT 31.414 63.926 31.466 63.962 ;
               RECT 31.414 65.126 31.466 65.162 ;
               RECT 31.414 66.326 31.466 66.362 ;
               RECT 31.414 67.526 31.466 67.562 ;
               RECT 31.414 68.726 31.466 68.762 ;
               RECT 31.414 69.926 31.466 69.962 ;
               RECT 31.414 71.126 31.466 71.162 ;
               RECT 31.414 72.326 31.466 72.362 ;
               RECT 31.414 73.526 31.466 73.562 ;
               RECT 31.414 74.726 31.466 74.762 ;
               RECT 31.414 75.926 31.466 75.962 ;
               RECT 31.414 77.126 31.466 77.162 ;
               RECT 31.414 78.326 31.466 78.362 ;
               RECT 31.414 79.526 31.466 79.562 ;
               RECT 31.414 80.726 31.466 80.762 ;
               RECT 31.414 81.926 31.466 81.962 ;
               RECT 31.414 83.126 31.466 83.162 ;
               RECT 31.414 84.326 31.466 84.362 ;
               RECT 31.414 85.526 31.466 85.562 ;
               RECT 31.414 86.726 31.466 86.762 ;
               RECT 31.414 87.926 31.466 87.962 ;
               RECT 31.414 89.126 31.466 89.162 ;
               RECT 31.414 90.326 31.466 90.362 ;
               RECT 31.414 91.526 31.466 91.562 ;
               RECT 31.414 92.726 31.466 92.762 ;
               RECT 31.414 93.926 31.466 93.962 ;
               RECT 31.414 95.126 31.466 95.162 ;
               RECT 31.414 96.326 31.466 96.362 ;
               RECT 31.414 97.526 31.466 97.562 ;
               RECT 31.414 98.726 31.466 98.762 ;
               RECT 31.414 99.926 31.466 99.962 ;
               RECT 31.414 101.126 31.466 101.162 ;
               RECT 31.414 102.326 31.466 102.362 ;
               RECT 31.414 103.526 31.466 103.562 ;
               RECT 31.494 1.558 31.546 1.594 ;
               RECT 31.494 2.758 31.546 2.794 ;
               RECT 31.494 3.958 31.546 3.994 ;
               RECT 31.494 5.158 31.546 5.194 ;
               RECT 31.494 6.358 31.546 6.394 ;
               RECT 31.494 7.558 31.546 7.594 ;
               RECT 31.494 8.758 31.546 8.794 ;
               RECT 31.494 9.958 31.546 9.994 ;
               RECT 31.494 11.158 31.546 11.194 ;
               RECT 31.494 12.358 31.546 12.394 ;
               RECT 31.494 13.558 31.546 13.594 ;
               RECT 31.494 14.758 31.546 14.794 ;
               RECT 31.494 15.958 31.546 15.994 ;
               RECT 31.494 17.158 31.546 17.194 ;
               RECT 31.494 18.358 31.546 18.394 ;
               RECT 31.494 19.558 31.546 19.594 ;
               RECT 31.494 20.758 31.546 20.794 ;
               RECT 31.494 21.958 31.546 21.994 ;
               RECT 31.494 23.158 31.546 23.194 ;
               RECT 31.494 24.358 31.546 24.394 ;
               RECT 31.494 25.558 31.546 25.594 ;
               RECT 31.494 26.758 31.546 26.794 ;
               RECT 31.494 27.958 31.546 27.994 ;
               RECT 31.494 29.158 31.546 29.194 ;
               RECT 31.494 30.358 31.546 30.394 ;
               RECT 31.494 31.558 31.546 31.594 ;
               RECT 31.494 32.758 31.546 32.794 ;
               RECT 31.494 33.958 31.546 33.994 ;
               RECT 31.494 35.158 31.546 35.194 ;
               RECT 31.494 36.358 31.546 36.394 ;
               RECT 31.494 37.558 31.546 37.594 ;
               RECT 31.494 38.758 31.546 38.794 ;
               RECT 31.494 39.958 31.546 39.994 ;
               RECT 31.494 41.158 31.546 41.194 ;
               RECT 31.494 42.358 31.546 42.394 ;
               RECT 31.494 43.558 31.546 43.594 ;
               RECT 31.494 44.758 31.546 44.794 ;
               RECT 31.494 45.958 31.546 45.994 ;
               RECT 31.494 47.158 31.546 47.194 ;
               RECT 31.494 48.358 31.546 48.394 ;
               RECT 31.494 50.142 31.546 50.178 ;
               RECT 31.494 50.382 31.546 50.418 ;
               RECT 31.494 54.702 31.546 54.738 ;
               RECT 31.494 54.942 31.546 54.978 ;
               RECT 31.494 57.478 31.546 57.514 ;
               RECT 31.494 58.678 31.546 58.714 ;
               RECT 31.494 59.878 31.546 59.914 ;
               RECT 31.494 61.078 31.546 61.114 ;
               RECT 31.494 62.278 31.546 62.314 ;
               RECT 31.494 63.478 31.546 63.514 ;
               RECT 31.494 64.678 31.546 64.714 ;
               RECT 31.494 65.878 31.546 65.914 ;
               RECT 31.494 67.078 31.546 67.114 ;
               RECT 31.494 68.278 31.546 68.314 ;
               RECT 31.494 69.478 31.546 69.514 ;
               RECT 31.494 70.678 31.546 70.714 ;
               RECT 31.494 71.878 31.546 71.914 ;
               RECT 31.494 73.078 31.546 73.114 ;
               RECT 31.494 74.278 31.546 74.314 ;
               RECT 31.494 75.478 31.546 75.514 ;
               RECT 31.494 76.678 31.546 76.714 ;
               RECT 31.494 77.878 31.546 77.914 ;
               RECT 31.494 79.078 31.546 79.114 ;
               RECT 31.494 80.278 31.546 80.314 ;
               RECT 31.494 81.478 31.546 81.514 ;
               RECT 31.494 82.678 31.546 82.714 ;
               RECT 31.494 83.878 31.546 83.914 ;
               RECT 31.494 85.078 31.546 85.114 ;
               RECT 31.494 86.278 31.546 86.314 ;
               RECT 31.494 87.478 31.546 87.514 ;
               RECT 31.494 88.678 31.546 88.714 ;
               RECT 31.494 89.878 31.546 89.914 ;
               RECT 31.494 91.078 31.546 91.114 ;
               RECT 31.494 92.278 31.546 92.314 ;
               RECT 31.494 93.478 31.546 93.514 ;
               RECT 31.494 94.678 31.546 94.714 ;
               RECT 31.494 95.878 31.546 95.914 ;
               RECT 31.494 97.078 31.546 97.114 ;
               RECT 31.494 98.278 31.546 98.314 ;
               RECT 31.494 99.478 31.546 99.514 ;
               RECT 31.494 100.678 31.546 100.714 ;
               RECT 31.494 101.878 31.546 101.914 ;
               RECT 31.494 103.078 31.546 103.114 ;
               RECT 31.494 104.278 31.546 104.314 ;
               RECT 31.574 0.281 31.626 0.317 ;
               RECT 31.574 104.803 31.626 104.839 ;
               RECT 31.654 0.806 31.706 0.842 ;
               RECT 31.654 2.006 31.706 2.042 ;
               RECT 31.654 3.206 31.706 3.242 ;
               RECT 31.654 4.406 31.706 4.442 ;
               RECT 31.654 5.606 31.706 5.642 ;
               RECT 31.654 6.806 31.706 6.842 ;
               RECT 31.654 8.006 31.706 8.042 ;
               RECT 31.654 9.206 31.706 9.242 ;
               RECT 31.654 10.406 31.706 10.442 ;
               RECT 31.654 11.606 31.706 11.642 ;
               RECT 31.654 12.806 31.706 12.842 ;
               RECT 31.654 14.006 31.706 14.042 ;
               RECT 31.654 15.206 31.706 15.242 ;
               RECT 31.654 16.406 31.706 16.442 ;
               RECT 31.654 17.606 31.706 17.642 ;
               RECT 31.654 18.806 31.706 18.842 ;
               RECT 31.654 20.006 31.706 20.042 ;
               RECT 31.654 21.206 31.706 21.242 ;
               RECT 31.654 22.406 31.706 22.442 ;
               RECT 31.654 23.606 31.706 23.642 ;
               RECT 31.654 24.806 31.706 24.842 ;
               RECT 31.654 26.006 31.706 26.042 ;
               RECT 31.654 27.206 31.706 27.242 ;
               RECT 31.654 28.406 31.706 28.442 ;
               RECT 31.654 29.606 31.706 29.642 ;
               RECT 31.654 30.806 31.706 30.842 ;
               RECT 31.654 32.006 31.706 32.042 ;
               RECT 31.654 33.206 31.706 33.242 ;
               RECT 31.654 34.406 31.706 34.442 ;
               RECT 31.654 35.606 31.706 35.642 ;
               RECT 31.654 36.806 31.706 36.842 ;
               RECT 31.654 38.006 31.706 38.042 ;
               RECT 31.654 39.206 31.706 39.242 ;
               RECT 31.654 40.406 31.706 40.442 ;
               RECT 31.654 41.606 31.706 41.642 ;
               RECT 31.654 42.806 31.706 42.842 ;
               RECT 31.654 44.006 31.706 44.042 ;
               RECT 31.654 45.206 31.706 45.242 ;
               RECT 31.654 46.406 31.706 46.442 ;
               RECT 31.654 47.606 31.706 47.642 ;
               RECT 31.654 49.422 31.706 49.458 ;
               RECT 31.654 49.662 31.706 49.698 ;
               RECT 31.654 55.422 31.706 55.458 ;
               RECT 31.654 55.662 31.706 55.698 ;
               RECT 31.654 56.726 31.706 56.762 ;
               RECT 31.654 57.926 31.706 57.962 ;
               RECT 31.654 59.126 31.706 59.162 ;
               RECT 31.654 60.326 31.706 60.362 ;
               RECT 31.654 61.526 31.706 61.562 ;
               RECT 31.654 62.726 31.706 62.762 ;
               RECT 31.654 63.926 31.706 63.962 ;
               RECT 31.654 65.126 31.706 65.162 ;
               RECT 31.654 66.326 31.706 66.362 ;
               RECT 31.654 67.526 31.706 67.562 ;
               RECT 31.654 68.726 31.706 68.762 ;
               RECT 31.654 69.926 31.706 69.962 ;
               RECT 31.654 71.126 31.706 71.162 ;
               RECT 31.654 72.326 31.706 72.362 ;
               RECT 31.654 73.526 31.706 73.562 ;
               RECT 31.654 74.726 31.706 74.762 ;
               RECT 31.654 75.926 31.706 75.962 ;
               RECT 31.654 77.126 31.706 77.162 ;
               RECT 31.654 78.326 31.706 78.362 ;
               RECT 31.654 79.526 31.706 79.562 ;
               RECT 31.654 80.726 31.706 80.762 ;
               RECT 31.654 81.926 31.706 81.962 ;
               RECT 31.654 83.126 31.706 83.162 ;
               RECT 31.654 84.326 31.706 84.362 ;
               RECT 31.654 85.526 31.706 85.562 ;
               RECT 31.654 86.726 31.706 86.762 ;
               RECT 31.654 87.926 31.706 87.962 ;
               RECT 31.654 89.126 31.706 89.162 ;
               RECT 31.654 90.326 31.706 90.362 ;
               RECT 31.654 91.526 31.706 91.562 ;
               RECT 31.654 92.726 31.706 92.762 ;
               RECT 31.654 93.926 31.706 93.962 ;
               RECT 31.654 95.126 31.706 95.162 ;
               RECT 31.654 96.326 31.706 96.362 ;
               RECT 31.654 97.526 31.706 97.562 ;
               RECT 31.654 98.726 31.706 98.762 ;
               RECT 31.654 99.926 31.706 99.962 ;
               RECT 31.654 101.126 31.706 101.162 ;
               RECT 31.654 102.326 31.706 102.362 ;
               RECT 31.654 103.526 31.706 103.562 ;
               RECT 31.734 1.558 31.786 1.594 ;
               RECT 31.734 2.758 31.786 2.794 ;
               RECT 31.734 3.958 31.786 3.994 ;
               RECT 31.734 5.158 31.786 5.194 ;
               RECT 31.734 6.358 31.786 6.394 ;
               RECT 31.734 7.558 31.786 7.594 ;
               RECT 31.734 8.758 31.786 8.794 ;
               RECT 31.734 9.958 31.786 9.994 ;
               RECT 31.734 11.158 31.786 11.194 ;
               RECT 31.734 12.358 31.786 12.394 ;
               RECT 31.734 13.558 31.786 13.594 ;
               RECT 31.734 14.758 31.786 14.794 ;
               RECT 31.734 15.958 31.786 15.994 ;
               RECT 31.734 17.158 31.786 17.194 ;
               RECT 31.734 18.358 31.786 18.394 ;
               RECT 31.734 19.558 31.786 19.594 ;
               RECT 31.734 20.758 31.786 20.794 ;
               RECT 31.734 21.958 31.786 21.994 ;
               RECT 31.734 23.158 31.786 23.194 ;
               RECT 31.734 24.358 31.786 24.394 ;
               RECT 31.734 25.558 31.786 25.594 ;
               RECT 31.734 26.758 31.786 26.794 ;
               RECT 31.734 27.958 31.786 27.994 ;
               RECT 31.734 29.158 31.786 29.194 ;
               RECT 31.734 30.358 31.786 30.394 ;
               RECT 31.734 31.558 31.786 31.594 ;
               RECT 31.734 32.758 31.786 32.794 ;
               RECT 31.734 33.958 31.786 33.994 ;
               RECT 31.734 35.158 31.786 35.194 ;
               RECT 31.734 36.358 31.786 36.394 ;
               RECT 31.734 37.558 31.786 37.594 ;
               RECT 31.734 38.758 31.786 38.794 ;
               RECT 31.734 39.958 31.786 39.994 ;
               RECT 31.734 41.158 31.786 41.194 ;
               RECT 31.734 42.358 31.786 42.394 ;
               RECT 31.734 43.558 31.786 43.594 ;
               RECT 31.734 44.758 31.786 44.794 ;
               RECT 31.734 45.958 31.786 45.994 ;
               RECT 31.734 47.158 31.786 47.194 ;
               RECT 31.734 48.358 31.786 48.394 ;
               RECT 31.734 50.142 31.786 50.178 ;
               RECT 31.734 50.382 31.786 50.418 ;
               RECT 31.734 54.702 31.786 54.738 ;
               RECT 31.734 54.942 31.786 54.978 ;
               RECT 31.734 57.478 31.786 57.514 ;
               RECT 31.734 58.678 31.786 58.714 ;
               RECT 31.734 59.878 31.786 59.914 ;
               RECT 31.734 61.078 31.786 61.114 ;
               RECT 31.734 62.278 31.786 62.314 ;
               RECT 31.734 63.478 31.786 63.514 ;
               RECT 31.734 64.678 31.786 64.714 ;
               RECT 31.734 65.878 31.786 65.914 ;
               RECT 31.734 67.078 31.786 67.114 ;
               RECT 31.734 68.278 31.786 68.314 ;
               RECT 31.734 69.478 31.786 69.514 ;
               RECT 31.734 70.678 31.786 70.714 ;
               RECT 31.734 71.878 31.786 71.914 ;
               RECT 31.734 73.078 31.786 73.114 ;
               RECT 31.734 74.278 31.786 74.314 ;
               RECT 31.734 75.478 31.786 75.514 ;
               RECT 31.734 76.678 31.786 76.714 ;
               RECT 31.734 77.878 31.786 77.914 ;
               RECT 31.734 79.078 31.786 79.114 ;
               RECT 31.734 80.278 31.786 80.314 ;
               RECT 31.734 81.478 31.786 81.514 ;
               RECT 31.734 82.678 31.786 82.714 ;
               RECT 31.734 83.878 31.786 83.914 ;
               RECT 31.734 85.078 31.786 85.114 ;
               RECT 31.734 86.278 31.786 86.314 ;
               RECT 31.734 87.478 31.786 87.514 ;
               RECT 31.734 88.678 31.786 88.714 ;
               RECT 31.734 89.878 31.786 89.914 ;
               RECT 31.734 91.078 31.786 91.114 ;
               RECT 31.734 92.278 31.786 92.314 ;
               RECT 31.734 93.478 31.786 93.514 ;
               RECT 31.734 94.678 31.786 94.714 ;
               RECT 31.734 95.878 31.786 95.914 ;
               RECT 31.734 97.078 31.786 97.114 ;
               RECT 31.734 98.278 31.786 98.314 ;
               RECT 31.734 99.478 31.786 99.514 ;
               RECT 31.734 100.678 31.786 100.714 ;
               RECT 31.734 101.878 31.786 101.914 ;
               RECT 31.734 103.078 31.786 103.114 ;
               RECT 31.734 104.278 31.786 104.314 ;
               RECT 31.814 0.806 31.866 0.842 ;
               RECT 31.814 2.006 31.866 2.042 ;
               RECT 31.814 3.206 31.866 3.242 ;
               RECT 31.814 4.406 31.866 4.442 ;
               RECT 31.814 5.606 31.866 5.642 ;
               RECT 31.814 6.806 31.866 6.842 ;
               RECT 31.814 8.006 31.866 8.042 ;
               RECT 31.814 9.206 31.866 9.242 ;
               RECT 31.814 10.406 31.866 10.442 ;
               RECT 31.814 11.606 31.866 11.642 ;
               RECT 31.814 12.806 31.866 12.842 ;
               RECT 31.814 14.006 31.866 14.042 ;
               RECT 31.814 15.206 31.866 15.242 ;
               RECT 31.814 16.406 31.866 16.442 ;
               RECT 31.814 17.606 31.866 17.642 ;
               RECT 31.814 18.806 31.866 18.842 ;
               RECT 31.814 20.006 31.866 20.042 ;
               RECT 31.814 21.206 31.866 21.242 ;
               RECT 31.814 22.406 31.866 22.442 ;
               RECT 31.814 23.606 31.866 23.642 ;
               RECT 31.814 24.806 31.866 24.842 ;
               RECT 31.814 26.006 31.866 26.042 ;
               RECT 31.814 27.206 31.866 27.242 ;
               RECT 31.814 28.406 31.866 28.442 ;
               RECT 31.814 29.606 31.866 29.642 ;
               RECT 31.814 30.806 31.866 30.842 ;
               RECT 31.814 32.006 31.866 32.042 ;
               RECT 31.814 33.206 31.866 33.242 ;
               RECT 31.814 34.406 31.866 34.442 ;
               RECT 31.814 35.606 31.866 35.642 ;
               RECT 31.814 36.806 31.866 36.842 ;
               RECT 31.814 38.006 31.866 38.042 ;
               RECT 31.814 39.206 31.866 39.242 ;
               RECT 31.814 40.406 31.866 40.442 ;
               RECT 31.814 41.606 31.866 41.642 ;
               RECT 31.814 42.806 31.866 42.842 ;
               RECT 31.814 44.006 31.866 44.042 ;
               RECT 31.814 45.206 31.866 45.242 ;
               RECT 31.814 46.406 31.866 46.442 ;
               RECT 31.814 47.606 31.866 47.642 ;
               RECT 31.814 49.422 31.866 49.458 ;
               RECT 31.814 49.662 31.866 49.698 ;
               RECT 31.814 55.422 31.866 55.458 ;
               RECT 31.814 55.662 31.866 55.698 ;
               RECT 31.814 56.726 31.866 56.762 ;
               RECT 31.814 57.926 31.866 57.962 ;
               RECT 31.814 59.126 31.866 59.162 ;
               RECT 31.814 60.326 31.866 60.362 ;
               RECT 31.814 61.526 31.866 61.562 ;
               RECT 31.814 62.726 31.866 62.762 ;
               RECT 31.814 63.926 31.866 63.962 ;
               RECT 31.814 65.126 31.866 65.162 ;
               RECT 31.814 66.326 31.866 66.362 ;
               RECT 31.814 67.526 31.866 67.562 ;
               RECT 31.814 68.726 31.866 68.762 ;
               RECT 31.814 69.926 31.866 69.962 ;
               RECT 31.814 71.126 31.866 71.162 ;
               RECT 31.814 72.326 31.866 72.362 ;
               RECT 31.814 73.526 31.866 73.562 ;
               RECT 31.814 74.726 31.866 74.762 ;
               RECT 31.814 75.926 31.866 75.962 ;
               RECT 31.814 77.126 31.866 77.162 ;
               RECT 31.814 78.326 31.866 78.362 ;
               RECT 31.814 79.526 31.866 79.562 ;
               RECT 31.814 80.726 31.866 80.762 ;
               RECT 31.814 81.926 31.866 81.962 ;
               RECT 31.814 83.126 31.866 83.162 ;
               RECT 31.814 84.326 31.866 84.362 ;
               RECT 31.814 85.526 31.866 85.562 ;
               RECT 31.814 86.726 31.866 86.762 ;
               RECT 31.814 87.926 31.866 87.962 ;
               RECT 31.814 89.126 31.866 89.162 ;
               RECT 31.814 90.326 31.866 90.362 ;
               RECT 31.814 91.526 31.866 91.562 ;
               RECT 31.814 92.726 31.866 92.762 ;
               RECT 31.814 93.926 31.866 93.962 ;
               RECT 31.814 95.126 31.866 95.162 ;
               RECT 31.814 96.326 31.866 96.362 ;
               RECT 31.814 97.526 31.866 97.562 ;
               RECT 31.814 98.726 31.866 98.762 ;
               RECT 31.814 99.926 31.866 99.962 ;
               RECT 31.814 101.126 31.866 101.162 ;
               RECT 31.814 102.326 31.866 102.362 ;
               RECT 31.814 103.526 31.866 103.562 ;
               RECT 31.894 1.558 31.946 1.594 ;
               RECT 31.894 2.758 31.946 2.794 ;
               RECT 31.894 3.958 31.946 3.994 ;
               RECT 31.894 5.158 31.946 5.194 ;
               RECT 31.894 6.358 31.946 6.394 ;
               RECT 31.894 7.558 31.946 7.594 ;
               RECT 31.894 8.758 31.946 8.794 ;
               RECT 31.894 9.958 31.946 9.994 ;
               RECT 31.894 11.158 31.946 11.194 ;
               RECT 31.894 12.358 31.946 12.394 ;
               RECT 31.894 13.558 31.946 13.594 ;
               RECT 31.894 14.758 31.946 14.794 ;
               RECT 31.894 15.958 31.946 15.994 ;
               RECT 31.894 17.158 31.946 17.194 ;
               RECT 31.894 18.358 31.946 18.394 ;
               RECT 31.894 19.558 31.946 19.594 ;
               RECT 31.894 20.758 31.946 20.794 ;
               RECT 31.894 21.958 31.946 21.994 ;
               RECT 31.894 23.158 31.946 23.194 ;
               RECT 31.894 24.358 31.946 24.394 ;
               RECT 31.894 25.558 31.946 25.594 ;
               RECT 31.894 26.758 31.946 26.794 ;
               RECT 31.894 27.958 31.946 27.994 ;
               RECT 31.894 29.158 31.946 29.194 ;
               RECT 31.894 30.358 31.946 30.394 ;
               RECT 31.894 31.558 31.946 31.594 ;
               RECT 31.894 32.758 31.946 32.794 ;
               RECT 31.894 33.958 31.946 33.994 ;
               RECT 31.894 35.158 31.946 35.194 ;
               RECT 31.894 36.358 31.946 36.394 ;
               RECT 31.894 37.558 31.946 37.594 ;
               RECT 31.894 38.758 31.946 38.794 ;
               RECT 31.894 39.958 31.946 39.994 ;
               RECT 31.894 41.158 31.946 41.194 ;
               RECT 31.894 42.358 31.946 42.394 ;
               RECT 31.894 43.558 31.946 43.594 ;
               RECT 31.894 44.758 31.946 44.794 ;
               RECT 31.894 45.958 31.946 45.994 ;
               RECT 31.894 47.158 31.946 47.194 ;
               RECT 31.894 48.358 31.946 48.394 ;
               RECT 31.894 50.142 31.946 50.178 ;
               RECT 31.894 50.382 31.946 50.418 ;
               RECT 31.894 54.702 31.946 54.738 ;
               RECT 31.894 54.942 31.946 54.978 ;
               RECT 31.894 57.478 31.946 57.514 ;
               RECT 31.894 58.678 31.946 58.714 ;
               RECT 31.894 59.878 31.946 59.914 ;
               RECT 31.894 61.078 31.946 61.114 ;
               RECT 31.894 62.278 31.946 62.314 ;
               RECT 31.894 63.478 31.946 63.514 ;
               RECT 31.894 64.678 31.946 64.714 ;
               RECT 31.894 65.878 31.946 65.914 ;
               RECT 31.894 67.078 31.946 67.114 ;
               RECT 31.894 68.278 31.946 68.314 ;
               RECT 31.894 69.478 31.946 69.514 ;
               RECT 31.894 70.678 31.946 70.714 ;
               RECT 31.894 71.878 31.946 71.914 ;
               RECT 31.894 73.078 31.946 73.114 ;
               RECT 31.894 74.278 31.946 74.314 ;
               RECT 31.894 75.478 31.946 75.514 ;
               RECT 31.894 76.678 31.946 76.714 ;
               RECT 31.894 77.878 31.946 77.914 ;
               RECT 31.894 79.078 31.946 79.114 ;
               RECT 31.894 80.278 31.946 80.314 ;
               RECT 31.894 81.478 31.946 81.514 ;
               RECT 31.894 82.678 31.946 82.714 ;
               RECT 31.894 83.878 31.946 83.914 ;
               RECT 31.894 85.078 31.946 85.114 ;
               RECT 31.894 86.278 31.946 86.314 ;
               RECT 31.894 87.478 31.946 87.514 ;
               RECT 31.894 88.678 31.946 88.714 ;
               RECT 31.894 89.878 31.946 89.914 ;
               RECT 31.894 91.078 31.946 91.114 ;
               RECT 31.894 92.278 31.946 92.314 ;
               RECT 31.894 93.478 31.946 93.514 ;
               RECT 31.894 94.678 31.946 94.714 ;
               RECT 31.894 95.878 31.946 95.914 ;
               RECT 31.894 97.078 31.946 97.114 ;
               RECT 31.894 98.278 31.946 98.314 ;
               RECT 31.894 99.478 31.946 99.514 ;
               RECT 31.894 100.678 31.946 100.714 ;
               RECT 31.894 101.878 31.946 101.914 ;
               RECT 31.894 103.078 31.946 103.114 ;
               RECT 31.894 104.278 31.946 104.314 ;
               RECT 31.974 0.281 32.026 0.317 ;
               RECT 31.974 104.803 32.026 104.839 ;
               RECT 32.054 0.806 32.106 0.842 ;
               RECT 32.054 2.006 32.106 2.042 ;
               RECT 32.054 3.206 32.106 3.242 ;
               RECT 32.054 4.406 32.106 4.442 ;
               RECT 32.054 5.606 32.106 5.642 ;
               RECT 32.054 6.806 32.106 6.842 ;
               RECT 32.054 8.006 32.106 8.042 ;
               RECT 32.054 9.206 32.106 9.242 ;
               RECT 32.054 10.406 32.106 10.442 ;
               RECT 32.054 11.606 32.106 11.642 ;
               RECT 32.054 12.806 32.106 12.842 ;
               RECT 32.054 14.006 32.106 14.042 ;
               RECT 32.054 15.206 32.106 15.242 ;
               RECT 32.054 16.406 32.106 16.442 ;
               RECT 32.054 17.606 32.106 17.642 ;
               RECT 32.054 18.806 32.106 18.842 ;
               RECT 32.054 20.006 32.106 20.042 ;
               RECT 32.054 21.206 32.106 21.242 ;
               RECT 32.054 22.406 32.106 22.442 ;
               RECT 32.054 23.606 32.106 23.642 ;
               RECT 32.054 24.806 32.106 24.842 ;
               RECT 32.054 26.006 32.106 26.042 ;
               RECT 32.054 27.206 32.106 27.242 ;
               RECT 32.054 28.406 32.106 28.442 ;
               RECT 32.054 29.606 32.106 29.642 ;
               RECT 32.054 30.806 32.106 30.842 ;
               RECT 32.054 32.006 32.106 32.042 ;
               RECT 32.054 33.206 32.106 33.242 ;
               RECT 32.054 34.406 32.106 34.442 ;
               RECT 32.054 35.606 32.106 35.642 ;
               RECT 32.054 36.806 32.106 36.842 ;
               RECT 32.054 38.006 32.106 38.042 ;
               RECT 32.054 39.206 32.106 39.242 ;
               RECT 32.054 40.406 32.106 40.442 ;
               RECT 32.054 41.606 32.106 41.642 ;
               RECT 32.054 42.806 32.106 42.842 ;
               RECT 32.054 44.006 32.106 44.042 ;
               RECT 32.054 45.206 32.106 45.242 ;
               RECT 32.054 46.406 32.106 46.442 ;
               RECT 32.054 47.606 32.106 47.642 ;
               RECT 32.054 49.422 32.106 49.458 ;
               RECT 32.054 49.662 32.106 49.698 ;
               RECT 32.054 51.102 32.106 51.138 ;
               RECT 32.054 51.582 32.106 51.618 ;
               RECT 32.054 53.502 32.106 53.538 ;
               RECT 32.054 53.982 32.106 54.018 ;
               RECT 32.054 55.422 32.106 55.458 ;
               RECT 32.054 55.662 32.106 55.698 ;
               RECT 32.054 56.726 32.106 56.762 ;
               RECT 32.054 57.926 32.106 57.962 ;
               RECT 32.054 59.126 32.106 59.162 ;
               RECT 32.054 60.326 32.106 60.362 ;
               RECT 32.054 61.526 32.106 61.562 ;
               RECT 32.054 62.726 32.106 62.762 ;
               RECT 32.054 63.926 32.106 63.962 ;
               RECT 32.054 65.126 32.106 65.162 ;
               RECT 32.054 66.326 32.106 66.362 ;
               RECT 32.054 67.526 32.106 67.562 ;
               RECT 32.054 68.726 32.106 68.762 ;
               RECT 32.054 69.926 32.106 69.962 ;
               RECT 32.054 71.126 32.106 71.162 ;
               RECT 32.054 72.326 32.106 72.362 ;
               RECT 32.054 73.526 32.106 73.562 ;
               RECT 32.054 74.726 32.106 74.762 ;
               RECT 32.054 75.926 32.106 75.962 ;
               RECT 32.054 77.126 32.106 77.162 ;
               RECT 32.054 78.326 32.106 78.362 ;
               RECT 32.054 79.526 32.106 79.562 ;
               RECT 32.054 80.726 32.106 80.762 ;
               RECT 32.054 81.926 32.106 81.962 ;
               RECT 32.054 83.126 32.106 83.162 ;
               RECT 32.054 84.326 32.106 84.362 ;
               RECT 32.054 85.526 32.106 85.562 ;
               RECT 32.054 86.726 32.106 86.762 ;
               RECT 32.054 87.926 32.106 87.962 ;
               RECT 32.054 89.126 32.106 89.162 ;
               RECT 32.054 90.326 32.106 90.362 ;
               RECT 32.054 91.526 32.106 91.562 ;
               RECT 32.054 92.726 32.106 92.762 ;
               RECT 32.054 93.926 32.106 93.962 ;
               RECT 32.054 95.126 32.106 95.162 ;
               RECT 32.054 96.326 32.106 96.362 ;
               RECT 32.054 97.526 32.106 97.562 ;
               RECT 32.054 98.726 32.106 98.762 ;
               RECT 32.054 99.926 32.106 99.962 ;
               RECT 32.054 101.126 32.106 101.162 ;
               RECT 32.054 102.326 32.106 102.362 ;
               RECT 32.054 103.526 32.106 103.562 ;
               RECT 32.134 1.558 32.186 1.594 ;
               RECT 32.134 2.758 32.186 2.794 ;
               RECT 32.134 3.958 32.186 3.994 ;
               RECT 32.134 5.158 32.186 5.194 ;
               RECT 32.134 6.358 32.186 6.394 ;
               RECT 32.134 7.558 32.186 7.594 ;
               RECT 32.134 8.758 32.186 8.794 ;
               RECT 32.134 9.958 32.186 9.994 ;
               RECT 32.134 11.158 32.186 11.194 ;
               RECT 32.134 12.358 32.186 12.394 ;
               RECT 32.134 13.558 32.186 13.594 ;
               RECT 32.134 14.758 32.186 14.794 ;
               RECT 32.134 15.958 32.186 15.994 ;
               RECT 32.134 17.158 32.186 17.194 ;
               RECT 32.134 18.358 32.186 18.394 ;
               RECT 32.134 19.558 32.186 19.594 ;
               RECT 32.134 20.758 32.186 20.794 ;
               RECT 32.134 21.958 32.186 21.994 ;
               RECT 32.134 23.158 32.186 23.194 ;
               RECT 32.134 24.358 32.186 24.394 ;
               RECT 32.134 25.558 32.186 25.594 ;
               RECT 32.134 26.758 32.186 26.794 ;
               RECT 32.134 27.958 32.186 27.994 ;
               RECT 32.134 29.158 32.186 29.194 ;
               RECT 32.134 30.358 32.186 30.394 ;
               RECT 32.134 31.558 32.186 31.594 ;
               RECT 32.134 32.758 32.186 32.794 ;
               RECT 32.134 33.958 32.186 33.994 ;
               RECT 32.134 35.158 32.186 35.194 ;
               RECT 32.134 36.358 32.186 36.394 ;
               RECT 32.134 37.558 32.186 37.594 ;
               RECT 32.134 38.758 32.186 38.794 ;
               RECT 32.134 39.958 32.186 39.994 ;
               RECT 32.134 41.158 32.186 41.194 ;
               RECT 32.134 42.358 32.186 42.394 ;
               RECT 32.134 43.558 32.186 43.594 ;
               RECT 32.134 44.758 32.186 44.794 ;
               RECT 32.134 45.958 32.186 45.994 ;
               RECT 32.134 47.158 32.186 47.194 ;
               RECT 32.134 48.358 32.186 48.394 ;
               RECT 32.134 50.142 32.186 50.178 ;
               RECT 32.134 50.382 32.186 50.418 ;
               RECT 32.134 54.702 32.186 54.738 ;
               RECT 32.134 54.942 32.186 54.978 ;
               RECT 32.134 57.478 32.186 57.514 ;
               RECT 32.134 58.678 32.186 58.714 ;
               RECT 32.134 59.878 32.186 59.914 ;
               RECT 32.134 61.078 32.186 61.114 ;
               RECT 32.134 62.278 32.186 62.314 ;
               RECT 32.134 63.478 32.186 63.514 ;
               RECT 32.134 64.678 32.186 64.714 ;
               RECT 32.134 65.878 32.186 65.914 ;
               RECT 32.134 67.078 32.186 67.114 ;
               RECT 32.134 68.278 32.186 68.314 ;
               RECT 32.134 69.478 32.186 69.514 ;
               RECT 32.134 70.678 32.186 70.714 ;
               RECT 32.134 71.878 32.186 71.914 ;
               RECT 32.134 73.078 32.186 73.114 ;
               RECT 32.134 74.278 32.186 74.314 ;
               RECT 32.134 75.478 32.186 75.514 ;
               RECT 32.134 76.678 32.186 76.714 ;
               RECT 32.134 77.878 32.186 77.914 ;
               RECT 32.134 79.078 32.186 79.114 ;
               RECT 32.134 80.278 32.186 80.314 ;
               RECT 32.134 81.478 32.186 81.514 ;
               RECT 32.134 82.678 32.186 82.714 ;
               RECT 32.134 83.878 32.186 83.914 ;
               RECT 32.134 85.078 32.186 85.114 ;
               RECT 32.134 86.278 32.186 86.314 ;
               RECT 32.134 87.478 32.186 87.514 ;
               RECT 32.134 88.678 32.186 88.714 ;
               RECT 32.134 89.878 32.186 89.914 ;
               RECT 32.134 91.078 32.186 91.114 ;
               RECT 32.134 92.278 32.186 92.314 ;
               RECT 32.134 93.478 32.186 93.514 ;
               RECT 32.134 94.678 32.186 94.714 ;
               RECT 32.134 95.878 32.186 95.914 ;
               RECT 32.134 97.078 32.186 97.114 ;
               RECT 32.134 98.278 32.186 98.314 ;
               RECT 32.134 99.478 32.186 99.514 ;
               RECT 32.134 100.678 32.186 100.714 ;
               RECT 32.134 101.878 32.186 101.914 ;
               RECT 32.134 103.078 32.186 103.114 ;
               RECT 32.134 104.278 32.186 104.314 ;
               RECT 32.214 0.806 32.266 0.842 ;
               RECT 32.214 2.006 32.266 2.042 ;
               RECT 32.214 3.206 32.266 3.242 ;
               RECT 32.214 4.406 32.266 4.442 ;
               RECT 32.214 5.606 32.266 5.642 ;
               RECT 32.214 6.806 32.266 6.842 ;
               RECT 32.214 8.006 32.266 8.042 ;
               RECT 32.214 9.206 32.266 9.242 ;
               RECT 32.214 10.406 32.266 10.442 ;
               RECT 32.214 11.606 32.266 11.642 ;
               RECT 32.214 12.806 32.266 12.842 ;
               RECT 32.214 14.006 32.266 14.042 ;
               RECT 32.214 15.206 32.266 15.242 ;
               RECT 32.214 16.406 32.266 16.442 ;
               RECT 32.214 17.606 32.266 17.642 ;
               RECT 32.214 18.806 32.266 18.842 ;
               RECT 32.214 20.006 32.266 20.042 ;
               RECT 32.214 21.206 32.266 21.242 ;
               RECT 32.214 22.406 32.266 22.442 ;
               RECT 32.214 23.606 32.266 23.642 ;
               RECT 32.214 24.806 32.266 24.842 ;
               RECT 32.214 26.006 32.266 26.042 ;
               RECT 32.214 27.206 32.266 27.242 ;
               RECT 32.214 28.406 32.266 28.442 ;
               RECT 32.214 29.606 32.266 29.642 ;
               RECT 32.214 30.806 32.266 30.842 ;
               RECT 32.214 32.006 32.266 32.042 ;
               RECT 32.214 33.206 32.266 33.242 ;
               RECT 32.214 34.406 32.266 34.442 ;
               RECT 32.214 35.606 32.266 35.642 ;
               RECT 32.214 36.806 32.266 36.842 ;
               RECT 32.214 38.006 32.266 38.042 ;
               RECT 32.214 39.206 32.266 39.242 ;
               RECT 32.214 40.406 32.266 40.442 ;
               RECT 32.214 41.606 32.266 41.642 ;
               RECT 32.214 42.806 32.266 42.842 ;
               RECT 32.214 44.006 32.266 44.042 ;
               RECT 32.214 45.206 32.266 45.242 ;
               RECT 32.214 46.406 32.266 46.442 ;
               RECT 32.214 47.606 32.266 47.642 ;
               RECT 32.214 49.422 32.266 49.458 ;
               RECT 32.214 49.662 32.266 49.698 ;
               RECT 32.214 55.422 32.266 55.458 ;
               RECT 32.214 55.662 32.266 55.698 ;
               RECT 32.214 56.726 32.266 56.762 ;
               RECT 32.214 57.926 32.266 57.962 ;
               RECT 32.214 59.126 32.266 59.162 ;
               RECT 32.214 60.326 32.266 60.362 ;
               RECT 32.214 61.526 32.266 61.562 ;
               RECT 32.214 62.726 32.266 62.762 ;
               RECT 32.214 63.926 32.266 63.962 ;
               RECT 32.214 65.126 32.266 65.162 ;
               RECT 32.214 66.326 32.266 66.362 ;
               RECT 32.214 67.526 32.266 67.562 ;
               RECT 32.214 68.726 32.266 68.762 ;
               RECT 32.214 69.926 32.266 69.962 ;
               RECT 32.214 71.126 32.266 71.162 ;
               RECT 32.214 72.326 32.266 72.362 ;
               RECT 32.214 73.526 32.266 73.562 ;
               RECT 32.214 74.726 32.266 74.762 ;
               RECT 32.214 75.926 32.266 75.962 ;
               RECT 32.214 77.126 32.266 77.162 ;
               RECT 32.214 78.326 32.266 78.362 ;
               RECT 32.214 79.526 32.266 79.562 ;
               RECT 32.214 80.726 32.266 80.762 ;
               RECT 32.214 81.926 32.266 81.962 ;
               RECT 32.214 83.126 32.266 83.162 ;
               RECT 32.214 84.326 32.266 84.362 ;
               RECT 32.214 85.526 32.266 85.562 ;
               RECT 32.214 86.726 32.266 86.762 ;
               RECT 32.214 87.926 32.266 87.962 ;
               RECT 32.214 89.126 32.266 89.162 ;
               RECT 32.214 90.326 32.266 90.362 ;
               RECT 32.214 91.526 32.266 91.562 ;
               RECT 32.214 92.726 32.266 92.762 ;
               RECT 32.214 93.926 32.266 93.962 ;
               RECT 32.214 95.126 32.266 95.162 ;
               RECT 32.214 96.326 32.266 96.362 ;
               RECT 32.214 97.526 32.266 97.562 ;
               RECT 32.214 98.726 32.266 98.762 ;
               RECT 32.214 99.926 32.266 99.962 ;
               RECT 32.214 101.126 32.266 101.162 ;
               RECT 32.214 102.326 32.266 102.362 ;
               RECT 32.214 103.526 32.266 103.562 ;
               RECT 32.294 1.558 32.346 1.594 ;
               RECT 32.294 2.758 32.346 2.794 ;
               RECT 32.294 3.958 32.346 3.994 ;
               RECT 32.294 5.158 32.346 5.194 ;
               RECT 32.294 6.358 32.346 6.394 ;
               RECT 32.294 7.558 32.346 7.594 ;
               RECT 32.294 8.758 32.346 8.794 ;
               RECT 32.294 9.958 32.346 9.994 ;
               RECT 32.294 11.158 32.346 11.194 ;
               RECT 32.294 12.358 32.346 12.394 ;
               RECT 32.294 13.558 32.346 13.594 ;
               RECT 32.294 14.758 32.346 14.794 ;
               RECT 32.294 15.958 32.346 15.994 ;
               RECT 32.294 17.158 32.346 17.194 ;
               RECT 32.294 18.358 32.346 18.394 ;
               RECT 32.294 19.558 32.346 19.594 ;
               RECT 32.294 20.758 32.346 20.794 ;
               RECT 32.294 21.958 32.346 21.994 ;
               RECT 32.294 23.158 32.346 23.194 ;
               RECT 32.294 24.358 32.346 24.394 ;
               RECT 32.294 25.558 32.346 25.594 ;
               RECT 32.294 26.758 32.346 26.794 ;
               RECT 32.294 27.958 32.346 27.994 ;
               RECT 32.294 29.158 32.346 29.194 ;
               RECT 32.294 30.358 32.346 30.394 ;
               RECT 32.294 31.558 32.346 31.594 ;
               RECT 32.294 32.758 32.346 32.794 ;
               RECT 32.294 33.958 32.346 33.994 ;
               RECT 32.294 35.158 32.346 35.194 ;
               RECT 32.294 36.358 32.346 36.394 ;
               RECT 32.294 37.558 32.346 37.594 ;
               RECT 32.294 38.758 32.346 38.794 ;
               RECT 32.294 39.958 32.346 39.994 ;
               RECT 32.294 41.158 32.346 41.194 ;
               RECT 32.294 42.358 32.346 42.394 ;
               RECT 32.294 43.558 32.346 43.594 ;
               RECT 32.294 44.758 32.346 44.794 ;
               RECT 32.294 45.958 32.346 45.994 ;
               RECT 32.294 47.158 32.346 47.194 ;
               RECT 32.294 48.358 32.346 48.394 ;
               RECT 32.294 50.142 32.346 50.178 ;
               RECT 32.294 50.382 32.346 50.418 ;
               RECT 32.294 54.702 32.346 54.738 ;
               RECT 32.294 54.942 32.346 54.978 ;
               RECT 32.294 57.478 32.346 57.514 ;
               RECT 32.294 58.678 32.346 58.714 ;
               RECT 32.294 59.878 32.346 59.914 ;
               RECT 32.294 61.078 32.346 61.114 ;
               RECT 32.294 62.278 32.346 62.314 ;
               RECT 32.294 63.478 32.346 63.514 ;
               RECT 32.294 64.678 32.346 64.714 ;
               RECT 32.294 65.878 32.346 65.914 ;
               RECT 32.294 67.078 32.346 67.114 ;
               RECT 32.294 68.278 32.346 68.314 ;
               RECT 32.294 69.478 32.346 69.514 ;
               RECT 32.294 70.678 32.346 70.714 ;
               RECT 32.294 71.878 32.346 71.914 ;
               RECT 32.294 73.078 32.346 73.114 ;
               RECT 32.294 74.278 32.346 74.314 ;
               RECT 32.294 75.478 32.346 75.514 ;
               RECT 32.294 76.678 32.346 76.714 ;
               RECT 32.294 77.878 32.346 77.914 ;
               RECT 32.294 79.078 32.346 79.114 ;
               RECT 32.294 80.278 32.346 80.314 ;
               RECT 32.294 81.478 32.346 81.514 ;
               RECT 32.294 82.678 32.346 82.714 ;
               RECT 32.294 83.878 32.346 83.914 ;
               RECT 32.294 85.078 32.346 85.114 ;
               RECT 32.294 86.278 32.346 86.314 ;
               RECT 32.294 87.478 32.346 87.514 ;
               RECT 32.294 88.678 32.346 88.714 ;
               RECT 32.294 89.878 32.346 89.914 ;
               RECT 32.294 91.078 32.346 91.114 ;
               RECT 32.294 92.278 32.346 92.314 ;
               RECT 32.294 93.478 32.346 93.514 ;
               RECT 32.294 94.678 32.346 94.714 ;
               RECT 32.294 95.878 32.346 95.914 ;
               RECT 32.294 97.078 32.346 97.114 ;
               RECT 32.294 98.278 32.346 98.314 ;
               RECT 32.294 99.478 32.346 99.514 ;
               RECT 32.294 100.678 32.346 100.714 ;
               RECT 32.294 101.878 32.346 101.914 ;
               RECT 32.294 103.078 32.346 103.114 ;
               RECT 32.294 104.278 32.346 104.314 ;
               RECT 32.374 0.281 32.426 0.317 ;
               RECT 32.374 104.803 32.426 104.839 ;
               RECT 32.454 0.806 32.506 0.842 ;
               RECT 32.454 2.006 32.506 2.042 ;
               RECT 32.454 3.206 32.506 3.242 ;
               RECT 32.454 4.406 32.506 4.442 ;
               RECT 32.454 5.606 32.506 5.642 ;
               RECT 32.454 6.806 32.506 6.842 ;
               RECT 32.454 8.006 32.506 8.042 ;
               RECT 32.454 9.206 32.506 9.242 ;
               RECT 32.454 10.406 32.506 10.442 ;
               RECT 32.454 11.606 32.506 11.642 ;
               RECT 32.454 12.806 32.506 12.842 ;
               RECT 32.454 14.006 32.506 14.042 ;
               RECT 32.454 15.206 32.506 15.242 ;
               RECT 32.454 16.406 32.506 16.442 ;
               RECT 32.454 17.606 32.506 17.642 ;
               RECT 32.454 18.806 32.506 18.842 ;
               RECT 32.454 20.006 32.506 20.042 ;
               RECT 32.454 21.206 32.506 21.242 ;
               RECT 32.454 22.406 32.506 22.442 ;
               RECT 32.454 23.606 32.506 23.642 ;
               RECT 32.454 24.806 32.506 24.842 ;
               RECT 32.454 26.006 32.506 26.042 ;
               RECT 32.454 27.206 32.506 27.242 ;
               RECT 32.454 28.406 32.506 28.442 ;
               RECT 32.454 29.606 32.506 29.642 ;
               RECT 32.454 30.806 32.506 30.842 ;
               RECT 32.454 32.006 32.506 32.042 ;
               RECT 32.454 33.206 32.506 33.242 ;
               RECT 32.454 34.406 32.506 34.442 ;
               RECT 32.454 35.606 32.506 35.642 ;
               RECT 32.454 36.806 32.506 36.842 ;
               RECT 32.454 38.006 32.506 38.042 ;
               RECT 32.454 39.206 32.506 39.242 ;
               RECT 32.454 40.406 32.506 40.442 ;
               RECT 32.454 41.606 32.506 41.642 ;
               RECT 32.454 42.806 32.506 42.842 ;
               RECT 32.454 44.006 32.506 44.042 ;
               RECT 32.454 45.206 32.506 45.242 ;
               RECT 32.454 46.406 32.506 46.442 ;
               RECT 32.454 47.606 32.506 47.642 ;
               RECT 32.454 49.422 32.506 49.458 ;
               RECT 32.454 49.662 32.506 49.698 ;
               RECT 32.454 55.422 32.506 55.458 ;
               RECT 32.454 55.662 32.506 55.698 ;
               RECT 32.454 56.726 32.506 56.762 ;
               RECT 32.454 57.926 32.506 57.962 ;
               RECT 32.454 59.126 32.506 59.162 ;
               RECT 32.454 60.326 32.506 60.362 ;
               RECT 32.454 61.526 32.506 61.562 ;
               RECT 32.454 62.726 32.506 62.762 ;
               RECT 32.454 63.926 32.506 63.962 ;
               RECT 32.454 65.126 32.506 65.162 ;
               RECT 32.454 66.326 32.506 66.362 ;
               RECT 32.454 67.526 32.506 67.562 ;
               RECT 32.454 68.726 32.506 68.762 ;
               RECT 32.454 69.926 32.506 69.962 ;
               RECT 32.454 71.126 32.506 71.162 ;
               RECT 32.454 72.326 32.506 72.362 ;
               RECT 32.454 73.526 32.506 73.562 ;
               RECT 32.454 74.726 32.506 74.762 ;
               RECT 32.454 75.926 32.506 75.962 ;
               RECT 32.454 77.126 32.506 77.162 ;
               RECT 32.454 78.326 32.506 78.362 ;
               RECT 32.454 79.526 32.506 79.562 ;
               RECT 32.454 80.726 32.506 80.762 ;
               RECT 32.454 81.926 32.506 81.962 ;
               RECT 32.454 83.126 32.506 83.162 ;
               RECT 32.454 84.326 32.506 84.362 ;
               RECT 32.454 85.526 32.506 85.562 ;
               RECT 32.454 86.726 32.506 86.762 ;
               RECT 32.454 87.926 32.506 87.962 ;
               RECT 32.454 89.126 32.506 89.162 ;
               RECT 32.454 90.326 32.506 90.362 ;
               RECT 32.454 91.526 32.506 91.562 ;
               RECT 32.454 92.726 32.506 92.762 ;
               RECT 32.454 93.926 32.506 93.962 ;
               RECT 32.454 95.126 32.506 95.162 ;
               RECT 32.454 96.326 32.506 96.362 ;
               RECT 32.454 97.526 32.506 97.562 ;
               RECT 32.454 98.726 32.506 98.762 ;
               RECT 32.454 99.926 32.506 99.962 ;
               RECT 32.454 101.126 32.506 101.162 ;
               RECT 32.454 102.326 32.506 102.362 ;
               RECT 32.454 103.526 32.506 103.562 ;
               RECT 32.534 1.558 32.586 1.594 ;
               RECT 32.534 2.758 32.586 2.794 ;
               RECT 32.534 3.958 32.586 3.994 ;
               RECT 32.534 5.158 32.586 5.194 ;
               RECT 32.534 6.358 32.586 6.394 ;
               RECT 32.534 7.558 32.586 7.594 ;
               RECT 32.534 8.758 32.586 8.794 ;
               RECT 32.534 9.958 32.586 9.994 ;
               RECT 32.534 11.158 32.586 11.194 ;
               RECT 32.534 12.358 32.586 12.394 ;
               RECT 32.534 13.558 32.586 13.594 ;
               RECT 32.534 14.758 32.586 14.794 ;
               RECT 32.534 15.958 32.586 15.994 ;
               RECT 32.534 17.158 32.586 17.194 ;
               RECT 32.534 18.358 32.586 18.394 ;
               RECT 32.534 19.558 32.586 19.594 ;
               RECT 32.534 20.758 32.586 20.794 ;
               RECT 32.534 21.958 32.586 21.994 ;
               RECT 32.534 23.158 32.586 23.194 ;
               RECT 32.534 24.358 32.586 24.394 ;
               RECT 32.534 25.558 32.586 25.594 ;
               RECT 32.534 26.758 32.586 26.794 ;
               RECT 32.534 27.958 32.586 27.994 ;
               RECT 32.534 29.158 32.586 29.194 ;
               RECT 32.534 30.358 32.586 30.394 ;
               RECT 32.534 31.558 32.586 31.594 ;
               RECT 32.534 32.758 32.586 32.794 ;
               RECT 32.534 33.958 32.586 33.994 ;
               RECT 32.534 35.158 32.586 35.194 ;
               RECT 32.534 36.358 32.586 36.394 ;
               RECT 32.534 37.558 32.586 37.594 ;
               RECT 32.534 38.758 32.586 38.794 ;
               RECT 32.534 39.958 32.586 39.994 ;
               RECT 32.534 41.158 32.586 41.194 ;
               RECT 32.534 42.358 32.586 42.394 ;
               RECT 32.534 43.558 32.586 43.594 ;
               RECT 32.534 44.758 32.586 44.794 ;
               RECT 32.534 45.958 32.586 45.994 ;
               RECT 32.534 47.158 32.586 47.194 ;
               RECT 32.534 48.358 32.586 48.394 ;
               RECT 32.534 50.142 32.586 50.178 ;
               RECT 32.534 50.382 32.586 50.418 ;
               RECT 32.534 54.702 32.586 54.738 ;
               RECT 32.534 54.942 32.586 54.978 ;
               RECT 32.534 57.478 32.586 57.514 ;
               RECT 32.534 58.678 32.586 58.714 ;
               RECT 32.534 59.878 32.586 59.914 ;
               RECT 32.534 61.078 32.586 61.114 ;
               RECT 32.534 62.278 32.586 62.314 ;
               RECT 32.534 63.478 32.586 63.514 ;
               RECT 32.534 64.678 32.586 64.714 ;
               RECT 32.534 65.878 32.586 65.914 ;
               RECT 32.534 67.078 32.586 67.114 ;
               RECT 32.534 68.278 32.586 68.314 ;
               RECT 32.534 69.478 32.586 69.514 ;
               RECT 32.534 70.678 32.586 70.714 ;
               RECT 32.534 71.878 32.586 71.914 ;
               RECT 32.534 73.078 32.586 73.114 ;
               RECT 32.534 74.278 32.586 74.314 ;
               RECT 32.534 75.478 32.586 75.514 ;
               RECT 32.534 76.678 32.586 76.714 ;
               RECT 32.534 77.878 32.586 77.914 ;
               RECT 32.534 79.078 32.586 79.114 ;
               RECT 32.534 80.278 32.586 80.314 ;
               RECT 32.534 81.478 32.586 81.514 ;
               RECT 32.534 82.678 32.586 82.714 ;
               RECT 32.534 83.878 32.586 83.914 ;
               RECT 32.534 85.078 32.586 85.114 ;
               RECT 32.534 86.278 32.586 86.314 ;
               RECT 32.534 87.478 32.586 87.514 ;
               RECT 32.534 88.678 32.586 88.714 ;
               RECT 32.534 89.878 32.586 89.914 ;
               RECT 32.534 91.078 32.586 91.114 ;
               RECT 32.534 92.278 32.586 92.314 ;
               RECT 32.534 93.478 32.586 93.514 ;
               RECT 32.534 94.678 32.586 94.714 ;
               RECT 32.534 95.878 32.586 95.914 ;
               RECT 32.534 97.078 32.586 97.114 ;
               RECT 32.534 98.278 32.586 98.314 ;
               RECT 32.534 99.478 32.586 99.514 ;
               RECT 32.534 100.678 32.586 100.714 ;
               RECT 32.534 101.878 32.586 101.914 ;
               RECT 32.534 103.078 32.586 103.114 ;
               RECT 32.534 104.278 32.586 104.314 ;
               RECT 32.614 0.806 32.666 0.842 ;
               RECT 32.614 2.006 32.666 2.042 ;
               RECT 32.614 3.206 32.666 3.242 ;
               RECT 32.614 4.406 32.666 4.442 ;
               RECT 32.614 5.606 32.666 5.642 ;
               RECT 32.614 6.806 32.666 6.842 ;
               RECT 32.614 8.006 32.666 8.042 ;
               RECT 32.614 9.206 32.666 9.242 ;
               RECT 32.614 10.406 32.666 10.442 ;
               RECT 32.614 11.606 32.666 11.642 ;
               RECT 32.614 12.806 32.666 12.842 ;
               RECT 32.614 14.006 32.666 14.042 ;
               RECT 32.614 15.206 32.666 15.242 ;
               RECT 32.614 16.406 32.666 16.442 ;
               RECT 32.614 17.606 32.666 17.642 ;
               RECT 32.614 18.806 32.666 18.842 ;
               RECT 32.614 20.006 32.666 20.042 ;
               RECT 32.614 21.206 32.666 21.242 ;
               RECT 32.614 22.406 32.666 22.442 ;
               RECT 32.614 23.606 32.666 23.642 ;
               RECT 32.614 24.806 32.666 24.842 ;
               RECT 32.614 26.006 32.666 26.042 ;
               RECT 32.614 27.206 32.666 27.242 ;
               RECT 32.614 28.406 32.666 28.442 ;
               RECT 32.614 29.606 32.666 29.642 ;
               RECT 32.614 30.806 32.666 30.842 ;
               RECT 32.614 32.006 32.666 32.042 ;
               RECT 32.614 33.206 32.666 33.242 ;
               RECT 32.614 34.406 32.666 34.442 ;
               RECT 32.614 35.606 32.666 35.642 ;
               RECT 32.614 36.806 32.666 36.842 ;
               RECT 32.614 38.006 32.666 38.042 ;
               RECT 32.614 39.206 32.666 39.242 ;
               RECT 32.614 40.406 32.666 40.442 ;
               RECT 32.614 41.606 32.666 41.642 ;
               RECT 32.614 42.806 32.666 42.842 ;
               RECT 32.614 44.006 32.666 44.042 ;
               RECT 32.614 45.206 32.666 45.242 ;
               RECT 32.614 46.406 32.666 46.442 ;
               RECT 32.614 47.606 32.666 47.642 ;
               RECT 32.614 49.422 32.666 49.458 ;
               RECT 32.614 49.662 32.666 49.698 ;
               RECT 32.614 55.422 32.666 55.458 ;
               RECT 32.614 55.662 32.666 55.698 ;
               RECT 32.614 56.726 32.666 56.762 ;
               RECT 32.614 57.926 32.666 57.962 ;
               RECT 32.614 59.126 32.666 59.162 ;
               RECT 32.614 60.326 32.666 60.362 ;
               RECT 32.614 61.526 32.666 61.562 ;
               RECT 32.614 62.726 32.666 62.762 ;
               RECT 32.614 63.926 32.666 63.962 ;
               RECT 32.614 65.126 32.666 65.162 ;
               RECT 32.614 66.326 32.666 66.362 ;
               RECT 32.614 67.526 32.666 67.562 ;
               RECT 32.614 68.726 32.666 68.762 ;
               RECT 32.614 69.926 32.666 69.962 ;
               RECT 32.614 71.126 32.666 71.162 ;
               RECT 32.614 72.326 32.666 72.362 ;
               RECT 32.614 73.526 32.666 73.562 ;
               RECT 32.614 74.726 32.666 74.762 ;
               RECT 32.614 75.926 32.666 75.962 ;
               RECT 32.614 77.126 32.666 77.162 ;
               RECT 32.614 78.326 32.666 78.362 ;
               RECT 32.614 79.526 32.666 79.562 ;
               RECT 32.614 80.726 32.666 80.762 ;
               RECT 32.614 81.926 32.666 81.962 ;
               RECT 32.614 83.126 32.666 83.162 ;
               RECT 32.614 84.326 32.666 84.362 ;
               RECT 32.614 85.526 32.666 85.562 ;
               RECT 32.614 86.726 32.666 86.762 ;
               RECT 32.614 87.926 32.666 87.962 ;
               RECT 32.614 89.126 32.666 89.162 ;
               RECT 32.614 90.326 32.666 90.362 ;
               RECT 32.614 91.526 32.666 91.562 ;
               RECT 32.614 92.726 32.666 92.762 ;
               RECT 32.614 93.926 32.666 93.962 ;
               RECT 32.614 95.126 32.666 95.162 ;
               RECT 32.614 96.326 32.666 96.362 ;
               RECT 32.614 97.526 32.666 97.562 ;
               RECT 32.614 98.726 32.666 98.762 ;
               RECT 32.614 99.926 32.666 99.962 ;
               RECT 32.614 101.126 32.666 101.162 ;
               RECT 32.614 102.326 32.666 102.362 ;
               RECT 32.614 103.526 32.666 103.562 ;
               RECT 32.694 1.558 32.746 1.594 ;
               RECT 32.694 2.758 32.746 2.794 ;
               RECT 32.694 3.958 32.746 3.994 ;
               RECT 32.694 5.158 32.746 5.194 ;
               RECT 32.694 6.358 32.746 6.394 ;
               RECT 32.694 7.558 32.746 7.594 ;
               RECT 32.694 8.758 32.746 8.794 ;
               RECT 32.694 9.958 32.746 9.994 ;
               RECT 32.694 11.158 32.746 11.194 ;
               RECT 32.694 12.358 32.746 12.394 ;
               RECT 32.694 13.558 32.746 13.594 ;
               RECT 32.694 14.758 32.746 14.794 ;
               RECT 32.694 15.958 32.746 15.994 ;
               RECT 32.694 17.158 32.746 17.194 ;
               RECT 32.694 18.358 32.746 18.394 ;
               RECT 32.694 19.558 32.746 19.594 ;
               RECT 32.694 20.758 32.746 20.794 ;
               RECT 32.694 21.958 32.746 21.994 ;
               RECT 32.694 23.158 32.746 23.194 ;
               RECT 32.694 24.358 32.746 24.394 ;
               RECT 32.694 25.558 32.746 25.594 ;
               RECT 32.694 26.758 32.746 26.794 ;
               RECT 32.694 27.958 32.746 27.994 ;
               RECT 32.694 29.158 32.746 29.194 ;
               RECT 32.694 30.358 32.746 30.394 ;
               RECT 32.694 31.558 32.746 31.594 ;
               RECT 32.694 32.758 32.746 32.794 ;
               RECT 32.694 33.958 32.746 33.994 ;
               RECT 32.694 35.158 32.746 35.194 ;
               RECT 32.694 36.358 32.746 36.394 ;
               RECT 32.694 37.558 32.746 37.594 ;
               RECT 32.694 38.758 32.746 38.794 ;
               RECT 32.694 39.958 32.746 39.994 ;
               RECT 32.694 41.158 32.746 41.194 ;
               RECT 32.694 42.358 32.746 42.394 ;
               RECT 32.694 43.558 32.746 43.594 ;
               RECT 32.694 44.758 32.746 44.794 ;
               RECT 32.694 45.958 32.746 45.994 ;
               RECT 32.694 47.158 32.746 47.194 ;
               RECT 32.694 48.358 32.746 48.394 ;
               RECT 32.694 50.142 32.746 50.178 ;
               RECT 32.694 50.382 32.746 50.418 ;
               RECT 32.694 54.702 32.746 54.738 ;
               RECT 32.694 54.942 32.746 54.978 ;
               RECT 32.694 57.478 32.746 57.514 ;
               RECT 32.694 58.678 32.746 58.714 ;
               RECT 32.694 59.878 32.746 59.914 ;
               RECT 32.694 61.078 32.746 61.114 ;
               RECT 32.694 62.278 32.746 62.314 ;
               RECT 32.694 63.478 32.746 63.514 ;
               RECT 32.694 64.678 32.746 64.714 ;
               RECT 32.694 65.878 32.746 65.914 ;
               RECT 32.694 67.078 32.746 67.114 ;
               RECT 32.694 68.278 32.746 68.314 ;
               RECT 32.694 69.478 32.746 69.514 ;
               RECT 32.694 70.678 32.746 70.714 ;
               RECT 32.694 71.878 32.746 71.914 ;
               RECT 32.694 73.078 32.746 73.114 ;
               RECT 32.694 74.278 32.746 74.314 ;
               RECT 32.694 75.478 32.746 75.514 ;
               RECT 32.694 76.678 32.746 76.714 ;
               RECT 32.694 77.878 32.746 77.914 ;
               RECT 32.694 79.078 32.746 79.114 ;
               RECT 32.694 80.278 32.746 80.314 ;
               RECT 32.694 81.478 32.746 81.514 ;
               RECT 32.694 82.678 32.746 82.714 ;
               RECT 32.694 83.878 32.746 83.914 ;
               RECT 32.694 85.078 32.746 85.114 ;
               RECT 32.694 86.278 32.746 86.314 ;
               RECT 32.694 87.478 32.746 87.514 ;
               RECT 32.694 88.678 32.746 88.714 ;
               RECT 32.694 89.878 32.746 89.914 ;
               RECT 32.694 91.078 32.746 91.114 ;
               RECT 32.694 92.278 32.746 92.314 ;
               RECT 32.694 93.478 32.746 93.514 ;
               RECT 32.694 94.678 32.746 94.714 ;
               RECT 32.694 95.878 32.746 95.914 ;
               RECT 32.694 97.078 32.746 97.114 ;
               RECT 32.694 98.278 32.746 98.314 ;
               RECT 32.694 99.478 32.746 99.514 ;
               RECT 32.694 100.678 32.746 100.714 ;
               RECT 32.694 101.878 32.746 101.914 ;
               RECT 32.694 103.078 32.746 103.114 ;
               RECT 32.694 104.278 32.746 104.314 ;
               RECT 32.774 0.281 32.826 0.317 ;
               RECT 32.774 104.803 32.826 104.839 ;
               RECT 32.854 0.806 32.906 0.842 ;
               RECT 32.854 2.006 32.906 2.042 ;
               RECT 32.854 3.206 32.906 3.242 ;
               RECT 32.854 4.406 32.906 4.442 ;
               RECT 32.854 5.606 32.906 5.642 ;
               RECT 32.854 6.806 32.906 6.842 ;
               RECT 32.854 8.006 32.906 8.042 ;
               RECT 32.854 9.206 32.906 9.242 ;
               RECT 32.854 10.406 32.906 10.442 ;
               RECT 32.854 11.606 32.906 11.642 ;
               RECT 32.854 12.806 32.906 12.842 ;
               RECT 32.854 14.006 32.906 14.042 ;
               RECT 32.854 15.206 32.906 15.242 ;
               RECT 32.854 16.406 32.906 16.442 ;
               RECT 32.854 17.606 32.906 17.642 ;
               RECT 32.854 18.806 32.906 18.842 ;
               RECT 32.854 20.006 32.906 20.042 ;
               RECT 32.854 21.206 32.906 21.242 ;
               RECT 32.854 22.406 32.906 22.442 ;
               RECT 32.854 23.606 32.906 23.642 ;
               RECT 32.854 24.806 32.906 24.842 ;
               RECT 32.854 26.006 32.906 26.042 ;
               RECT 32.854 27.206 32.906 27.242 ;
               RECT 32.854 28.406 32.906 28.442 ;
               RECT 32.854 29.606 32.906 29.642 ;
               RECT 32.854 30.806 32.906 30.842 ;
               RECT 32.854 32.006 32.906 32.042 ;
               RECT 32.854 33.206 32.906 33.242 ;
               RECT 32.854 34.406 32.906 34.442 ;
               RECT 32.854 35.606 32.906 35.642 ;
               RECT 32.854 36.806 32.906 36.842 ;
               RECT 32.854 38.006 32.906 38.042 ;
               RECT 32.854 39.206 32.906 39.242 ;
               RECT 32.854 40.406 32.906 40.442 ;
               RECT 32.854 41.606 32.906 41.642 ;
               RECT 32.854 42.806 32.906 42.842 ;
               RECT 32.854 44.006 32.906 44.042 ;
               RECT 32.854 45.206 32.906 45.242 ;
               RECT 32.854 46.406 32.906 46.442 ;
               RECT 32.854 47.606 32.906 47.642 ;
               RECT 32.854 49.422 32.906 49.458 ;
               RECT 32.854 49.662 32.906 49.698 ;
               RECT 32.854 51.102 32.906 51.138 ;
               RECT 32.854 51.582 32.906 51.618 ;
               RECT 32.854 53.502 32.906 53.538 ;
               RECT 32.854 53.982 32.906 54.018 ;
               RECT 32.854 55.422 32.906 55.458 ;
               RECT 32.854 55.662 32.906 55.698 ;
               RECT 32.854 56.726 32.906 56.762 ;
               RECT 32.854 57.926 32.906 57.962 ;
               RECT 32.854 59.126 32.906 59.162 ;
               RECT 32.854 60.326 32.906 60.362 ;
               RECT 32.854 61.526 32.906 61.562 ;
               RECT 32.854 62.726 32.906 62.762 ;
               RECT 32.854 63.926 32.906 63.962 ;
               RECT 32.854 65.126 32.906 65.162 ;
               RECT 32.854 66.326 32.906 66.362 ;
               RECT 32.854 67.526 32.906 67.562 ;
               RECT 32.854 68.726 32.906 68.762 ;
               RECT 32.854 69.926 32.906 69.962 ;
               RECT 32.854 71.126 32.906 71.162 ;
               RECT 32.854 72.326 32.906 72.362 ;
               RECT 32.854 73.526 32.906 73.562 ;
               RECT 32.854 74.726 32.906 74.762 ;
               RECT 32.854 75.926 32.906 75.962 ;
               RECT 32.854 77.126 32.906 77.162 ;
               RECT 32.854 78.326 32.906 78.362 ;
               RECT 32.854 79.526 32.906 79.562 ;
               RECT 32.854 80.726 32.906 80.762 ;
               RECT 32.854 81.926 32.906 81.962 ;
               RECT 32.854 83.126 32.906 83.162 ;
               RECT 32.854 84.326 32.906 84.362 ;
               RECT 32.854 85.526 32.906 85.562 ;
               RECT 32.854 86.726 32.906 86.762 ;
               RECT 32.854 87.926 32.906 87.962 ;
               RECT 32.854 89.126 32.906 89.162 ;
               RECT 32.854 90.326 32.906 90.362 ;
               RECT 32.854 91.526 32.906 91.562 ;
               RECT 32.854 92.726 32.906 92.762 ;
               RECT 32.854 93.926 32.906 93.962 ;
               RECT 32.854 95.126 32.906 95.162 ;
               RECT 32.854 96.326 32.906 96.362 ;
               RECT 32.854 97.526 32.906 97.562 ;
               RECT 32.854 98.726 32.906 98.762 ;
               RECT 32.854 99.926 32.906 99.962 ;
               RECT 32.854 101.126 32.906 101.162 ;
               RECT 32.854 102.326 32.906 102.362 ;
               RECT 32.854 103.526 32.906 103.562 ;
               RECT 32.934 1.558 32.986 1.594 ;
               RECT 32.934 2.758 32.986 2.794 ;
               RECT 32.934 3.958 32.986 3.994 ;
               RECT 32.934 5.158 32.986 5.194 ;
               RECT 32.934 6.358 32.986 6.394 ;
               RECT 32.934 7.558 32.986 7.594 ;
               RECT 32.934 8.758 32.986 8.794 ;
               RECT 32.934 9.958 32.986 9.994 ;
               RECT 32.934 11.158 32.986 11.194 ;
               RECT 32.934 12.358 32.986 12.394 ;
               RECT 32.934 13.558 32.986 13.594 ;
               RECT 32.934 14.758 32.986 14.794 ;
               RECT 32.934 15.958 32.986 15.994 ;
               RECT 32.934 17.158 32.986 17.194 ;
               RECT 32.934 18.358 32.986 18.394 ;
               RECT 32.934 19.558 32.986 19.594 ;
               RECT 32.934 20.758 32.986 20.794 ;
               RECT 32.934 21.958 32.986 21.994 ;
               RECT 32.934 23.158 32.986 23.194 ;
               RECT 32.934 24.358 32.986 24.394 ;
               RECT 32.934 25.558 32.986 25.594 ;
               RECT 32.934 26.758 32.986 26.794 ;
               RECT 32.934 27.958 32.986 27.994 ;
               RECT 32.934 29.158 32.986 29.194 ;
               RECT 32.934 30.358 32.986 30.394 ;
               RECT 32.934 31.558 32.986 31.594 ;
               RECT 32.934 32.758 32.986 32.794 ;
               RECT 32.934 33.958 32.986 33.994 ;
               RECT 32.934 35.158 32.986 35.194 ;
               RECT 32.934 36.358 32.986 36.394 ;
               RECT 32.934 37.558 32.986 37.594 ;
               RECT 32.934 38.758 32.986 38.794 ;
               RECT 32.934 39.958 32.986 39.994 ;
               RECT 32.934 41.158 32.986 41.194 ;
               RECT 32.934 42.358 32.986 42.394 ;
               RECT 32.934 43.558 32.986 43.594 ;
               RECT 32.934 44.758 32.986 44.794 ;
               RECT 32.934 45.958 32.986 45.994 ;
               RECT 32.934 47.158 32.986 47.194 ;
               RECT 32.934 48.358 32.986 48.394 ;
               RECT 32.934 50.142 32.986 50.178 ;
               RECT 32.934 50.382 32.986 50.418 ;
               RECT 32.934 54.702 32.986 54.738 ;
               RECT 32.934 54.942 32.986 54.978 ;
               RECT 32.934 57.478 32.986 57.514 ;
               RECT 32.934 58.678 32.986 58.714 ;
               RECT 32.934 59.878 32.986 59.914 ;
               RECT 32.934 61.078 32.986 61.114 ;
               RECT 32.934 62.278 32.986 62.314 ;
               RECT 32.934 63.478 32.986 63.514 ;
               RECT 32.934 64.678 32.986 64.714 ;
               RECT 32.934 65.878 32.986 65.914 ;
               RECT 32.934 67.078 32.986 67.114 ;
               RECT 32.934 68.278 32.986 68.314 ;
               RECT 32.934 69.478 32.986 69.514 ;
               RECT 32.934 70.678 32.986 70.714 ;
               RECT 32.934 71.878 32.986 71.914 ;
               RECT 32.934 73.078 32.986 73.114 ;
               RECT 32.934 74.278 32.986 74.314 ;
               RECT 32.934 75.478 32.986 75.514 ;
               RECT 32.934 76.678 32.986 76.714 ;
               RECT 32.934 77.878 32.986 77.914 ;
               RECT 32.934 79.078 32.986 79.114 ;
               RECT 32.934 80.278 32.986 80.314 ;
               RECT 32.934 81.478 32.986 81.514 ;
               RECT 32.934 82.678 32.986 82.714 ;
               RECT 32.934 83.878 32.986 83.914 ;
               RECT 32.934 85.078 32.986 85.114 ;
               RECT 32.934 86.278 32.986 86.314 ;
               RECT 32.934 87.478 32.986 87.514 ;
               RECT 32.934 88.678 32.986 88.714 ;
               RECT 32.934 89.878 32.986 89.914 ;
               RECT 32.934 91.078 32.986 91.114 ;
               RECT 32.934 92.278 32.986 92.314 ;
               RECT 32.934 93.478 32.986 93.514 ;
               RECT 32.934 94.678 32.986 94.714 ;
               RECT 32.934 95.878 32.986 95.914 ;
               RECT 32.934 97.078 32.986 97.114 ;
               RECT 32.934 98.278 32.986 98.314 ;
               RECT 32.934 99.478 32.986 99.514 ;
               RECT 32.934 100.678 32.986 100.714 ;
               RECT 32.934 101.878 32.986 101.914 ;
               RECT 32.934 103.078 32.986 103.114 ;
               RECT 32.934 104.278 32.986 104.314 ;
               RECT 33.014 0.806 33.066 0.842 ;
               RECT 33.014 2.006 33.066 2.042 ;
               RECT 33.014 3.206 33.066 3.242 ;
               RECT 33.014 4.406 33.066 4.442 ;
               RECT 33.014 5.606 33.066 5.642 ;
               RECT 33.014 6.806 33.066 6.842 ;
               RECT 33.014 8.006 33.066 8.042 ;
               RECT 33.014 9.206 33.066 9.242 ;
               RECT 33.014 10.406 33.066 10.442 ;
               RECT 33.014 11.606 33.066 11.642 ;
               RECT 33.014 12.806 33.066 12.842 ;
               RECT 33.014 14.006 33.066 14.042 ;
               RECT 33.014 15.206 33.066 15.242 ;
               RECT 33.014 16.406 33.066 16.442 ;
               RECT 33.014 17.606 33.066 17.642 ;
               RECT 33.014 18.806 33.066 18.842 ;
               RECT 33.014 20.006 33.066 20.042 ;
               RECT 33.014 21.206 33.066 21.242 ;
               RECT 33.014 22.406 33.066 22.442 ;
               RECT 33.014 23.606 33.066 23.642 ;
               RECT 33.014 24.806 33.066 24.842 ;
               RECT 33.014 26.006 33.066 26.042 ;
               RECT 33.014 27.206 33.066 27.242 ;
               RECT 33.014 28.406 33.066 28.442 ;
               RECT 33.014 29.606 33.066 29.642 ;
               RECT 33.014 30.806 33.066 30.842 ;
               RECT 33.014 32.006 33.066 32.042 ;
               RECT 33.014 33.206 33.066 33.242 ;
               RECT 33.014 34.406 33.066 34.442 ;
               RECT 33.014 35.606 33.066 35.642 ;
               RECT 33.014 36.806 33.066 36.842 ;
               RECT 33.014 38.006 33.066 38.042 ;
               RECT 33.014 39.206 33.066 39.242 ;
               RECT 33.014 40.406 33.066 40.442 ;
               RECT 33.014 41.606 33.066 41.642 ;
               RECT 33.014 42.806 33.066 42.842 ;
               RECT 33.014 44.006 33.066 44.042 ;
               RECT 33.014 45.206 33.066 45.242 ;
               RECT 33.014 46.406 33.066 46.442 ;
               RECT 33.014 47.606 33.066 47.642 ;
               RECT 33.014 49.422 33.066 49.458 ;
               RECT 33.014 49.662 33.066 49.698 ;
               RECT 33.014 55.422 33.066 55.458 ;
               RECT 33.014 55.662 33.066 55.698 ;
               RECT 33.014 56.726 33.066 56.762 ;
               RECT 33.014 57.926 33.066 57.962 ;
               RECT 33.014 59.126 33.066 59.162 ;
               RECT 33.014 60.326 33.066 60.362 ;
               RECT 33.014 61.526 33.066 61.562 ;
               RECT 33.014 62.726 33.066 62.762 ;
               RECT 33.014 63.926 33.066 63.962 ;
               RECT 33.014 65.126 33.066 65.162 ;
               RECT 33.014 66.326 33.066 66.362 ;
               RECT 33.014 67.526 33.066 67.562 ;
               RECT 33.014 68.726 33.066 68.762 ;
               RECT 33.014 69.926 33.066 69.962 ;
               RECT 33.014 71.126 33.066 71.162 ;
               RECT 33.014 72.326 33.066 72.362 ;
               RECT 33.014 73.526 33.066 73.562 ;
               RECT 33.014 74.726 33.066 74.762 ;
               RECT 33.014 75.926 33.066 75.962 ;
               RECT 33.014 77.126 33.066 77.162 ;
               RECT 33.014 78.326 33.066 78.362 ;
               RECT 33.014 79.526 33.066 79.562 ;
               RECT 33.014 80.726 33.066 80.762 ;
               RECT 33.014 81.926 33.066 81.962 ;
               RECT 33.014 83.126 33.066 83.162 ;
               RECT 33.014 84.326 33.066 84.362 ;
               RECT 33.014 85.526 33.066 85.562 ;
               RECT 33.014 86.726 33.066 86.762 ;
               RECT 33.014 87.926 33.066 87.962 ;
               RECT 33.014 89.126 33.066 89.162 ;
               RECT 33.014 90.326 33.066 90.362 ;
               RECT 33.014 91.526 33.066 91.562 ;
               RECT 33.014 92.726 33.066 92.762 ;
               RECT 33.014 93.926 33.066 93.962 ;
               RECT 33.014 95.126 33.066 95.162 ;
               RECT 33.014 96.326 33.066 96.362 ;
               RECT 33.014 97.526 33.066 97.562 ;
               RECT 33.014 98.726 33.066 98.762 ;
               RECT 33.014 99.926 33.066 99.962 ;
               RECT 33.014 101.126 33.066 101.162 ;
               RECT 33.014 102.326 33.066 102.362 ;
               RECT 33.014 103.526 33.066 103.562 ;
               RECT 33.094 1.558 33.146 1.594 ;
               RECT 33.094 2.758 33.146 2.794 ;
               RECT 33.094 3.958 33.146 3.994 ;
               RECT 33.094 5.158 33.146 5.194 ;
               RECT 33.094 6.358 33.146 6.394 ;
               RECT 33.094 7.558 33.146 7.594 ;
               RECT 33.094 8.758 33.146 8.794 ;
               RECT 33.094 9.958 33.146 9.994 ;
               RECT 33.094 11.158 33.146 11.194 ;
               RECT 33.094 12.358 33.146 12.394 ;
               RECT 33.094 13.558 33.146 13.594 ;
               RECT 33.094 14.758 33.146 14.794 ;
               RECT 33.094 15.958 33.146 15.994 ;
               RECT 33.094 17.158 33.146 17.194 ;
               RECT 33.094 18.358 33.146 18.394 ;
               RECT 33.094 19.558 33.146 19.594 ;
               RECT 33.094 20.758 33.146 20.794 ;
               RECT 33.094 21.958 33.146 21.994 ;
               RECT 33.094 23.158 33.146 23.194 ;
               RECT 33.094 24.358 33.146 24.394 ;
               RECT 33.094 25.558 33.146 25.594 ;
               RECT 33.094 26.758 33.146 26.794 ;
               RECT 33.094 27.958 33.146 27.994 ;
               RECT 33.094 29.158 33.146 29.194 ;
               RECT 33.094 30.358 33.146 30.394 ;
               RECT 33.094 31.558 33.146 31.594 ;
               RECT 33.094 32.758 33.146 32.794 ;
               RECT 33.094 33.958 33.146 33.994 ;
               RECT 33.094 35.158 33.146 35.194 ;
               RECT 33.094 36.358 33.146 36.394 ;
               RECT 33.094 37.558 33.146 37.594 ;
               RECT 33.094 38.758 33.146 38.794 ;
               RECT 33.094 39.958 33.146 39.994 ;
               RECT 33.094 41.158 33.146 41.194 ;
               RECT 33.094 42.358 33.146 42.394 ;
               RECT 33.094 43.558 33.146 43.594 ;
               RECT 33.094 44.758 33.146 44.794 ;
               RECT 33.094 45.958 33.146 45.994 ;
               RECT 33.094 47.158 33.146 47.194 ;
               RECT 33.094 48.358 33.146 48.394 ;
               RECT 33.094 50.142 33.146 50.178 ;
               RECT 33.094 50.382 33.146 50.418 ;
               RECT 33.094 54.702 33.146 54.738 ;
               RECT 33.094 54.942 33.146 54.978 ;
               RECT 33.094 57.478 33.146 57.514 ;
               RECT 33.094 58.678 33.146 58.714 ;
               RECT 33.094 59.878 33.146 59.914 ;
               RECT 33.094 61.078 33.146 61.114 ;
               RECT 33.094 62.278 33.146 62.314 ;
               RECT 33.094 63.478 33.146 63.514 ;
               RECT 33.094 64.678 33.146 64.714 ;
               RECT 33.094 65.878 33.146 65.914 ;
               RECT 33.094 67.078 33.146 67.114 ;
               RECT 33.094 68.278 33.146 68.314 ;
               RECT 33.094 69.478 33.146 69.514 ;
               RECT 33.094 70.678 33.146 70.714 ;
               RECT 33.094 71.878 33.146 71.914 ;
               RECT 33.094 73.078 33.146 73.114 ;
               RECT 33.094 74.278 33.146 74.314 ;
               RECT 33.094 75.478 33.146 75.514 ;
               RECT 33.094 76.678 33.146 76.714 ;
               RECT 33.094 77.878 33.146 77.914 ;
               RECT 33.094 79.078 33.146 79.114 ;
               RECT 33.094 80.278 33.146 80.314 ;
               RECT 33.094 81.478 33.146 81.514 ;
               RECT 33.094 82.678 33.146 82.714 ;
               RECT 33.094 83.878 33.146 83.914 ;
               RECT 33.094 85.078 33.146 85.114 ;
               RECT 33.094 86.278 33.146 86.314 ;
               RECT 33.094 87.478 33.146 87.514 ;
               RECT 33.094 88.678 33.146 88.714 ;
               RECT 33.094 89.878 33.146 89.914 ;
               RECT 33.094 91.078 33.146 91.114 ;
               RECT 33.094 92.278 33.146 92.314 ;
               RECT 33.094 93.478 33.146 93.514 ;
               RECT 33.094 94.678 33.146 94.714 ;
               RECT 33.094 95.878 33.146 95.914 ;
               RECT 33.094 97.078 33.146 97.114 ;
               RECT 33.094 98.278 33.146 98.314 ;
               RECT 33.094 99.478 33.146 99.514 ;
               RECT 33.094 100.678 33.146 100.714 ;
               RECT 33.094 101.878 33.146 101.914 ;
               RECT 33.094 103.078 33.146 103.114 ;
               RECT 33.094 104.278 33.146 104.314 ;
               RECT 33.174 0.281 33.226 0.317 ;
               RECT 33.174 104.803 33.226 104.839 ;
               RECT 33.254 0.806 33.306 0.842 ;
               RECT 33.254 2.006 33.306 2.042 ;
               RECT 33.254 3.206 33.306 3.242 ;
               RECT 33.254 4.406 33.306 4.442 ;
               RECT 33.254 5.606 33.306 5.642 ;
               RECT 33.254 6.806 33.306 6.842 ;
               RECT 33.254 8.006 33.306 8.042 ;
               RECT 33.254 9.206 33.306 9.242 ;
               RECT 33.254 10.406 33.306 10.442 ;
               RECT 33.254 11.606 33.306 11.642 ;
               RECT 33.254 12.806 33.306 12.842 ;
               RECT 33.254 14.006 33.306 14.042 ;
               RECT 33.254 15.206 33.306 15.242 ;
               RECT 33.254 16.406 33.306 16.442 ;
               RECT 33.254 17.606 33.306 17.642 ;
               RECT 33.254 18.806 33.306 18.842 ;
               RECT 33.254 20.006 33.306 20.042 ;
               RECT 33.254 21.206 33.306 21.242 ;
               RECT 33.254 22.406 33.306 22.442 ;
               RECT 33.254 23.606 33.306 23.642 ;
               RECT 33.254 24.806 33.306 24.842 ;
               RECT 33.254 26.006 33.306 26.042 ;
               RECT 33.254 27.206 33.306 27.242 ;
               RECT 33.254 28.406 33.306 28.442 ;
               RECT 33.254 29.606 33.306 29.642 ;
               RECT 33.254 30.806 33.306 30.842 ;
               RECT 33.254 32.006 33.306 32.042 ;
               RECT 33.254 33.206 33.306 33.242 ;
               RECT 33.254 34.406 33.306 34.442 ;
               RECT 33.254 35.606 33.306 35.642 ;
               RECT 33.254 36.806 33.306 36.842 ;
               RECT 33.254 38.006 33.306 38.042 ;
               RECT 33.254 39.206 33.306 39.242 ;
               RECT 33.254 40.406 33.306 40.442 ;
               RECT 33.254 41.606 33.306 41.642 ;
               RECT 33.254 42.806 33.306 42.842 ;
               RECT 33.254 44.006 33.306 44.042 ;
               RECT 33.254 45.206 33.306 45.242 ;
               RECT 33.254 46.406 33.306 46.442 ;
               RECT 33.254 47.606 33.306 47.642 ;
               RECT 33.254 49.422 33.306 49.458 ;
               RECT 33.254 49.662 33.306 49.698 ;
               RECT 33.254 55.422 33.306 55.458 ;
               RECT 33.254 55.662 33.306 55.698 ;
               RECT 33.254 56.726 33.306 56.762 ;
               RECT 33.254 57.926 33.306 57.962 ;
               RECT 33.254 59.126 33.306 59.162 ;
               RECT 33.254 60.326 33.306 60.362 ;
               RECT 33.254 61.526 33.306 61.562 ;
               RECT 33.254 62.726 33.306 62.762 ;
               RECT 33.254 63.926 33.306 63.962 ;
               RECT 33.254 65.126 33.306 65.162 ;
               RECT 33.254 66.326 33.306 66.362 ;
               RECT 33.254 67.526 33.306 67.562 ;
               RECT 33.254 68.726 33.306 68.762 ;
               RECT 33.254 69.926 33.306 69.962 ;
               RECT 33.254 71.126 33.306 71.162 ;
               RECT 33.254 72.326 33.306 72.362 ;
               RECT 33.254 73.526 33.306 73.562 ;
               RECT 33.254 74.726 33.306 74.762 ;
               RECT 33.254 75.926 33.306 75.962 ;
               RECT 33.254 77.126 33.306 77.162 ;
               RECT 33.254 78.326 33.306 78.362 ;
               RECT 33.254 79.526 33.306 79.562 ;
               RECT 33.254 80.726 33.306 80.762 ;
               RECT 33.254 81.926 33.306 81.962 ;
               RECT 33.254 83.126 33.306 83.162 ;
               RECT 33.254 84.326 33.306 84.362 ;
               RECT 33.254 85.526 33.306 85.562 ;
               RECT 33.254 86.726 33.306 86.762 ;
               RECT 33.254 87.926 33.306 87.962 ;
               RECT 33.254 89.126 33.306 89.162 ;
               RECT 33.254 90.326 33.306 90.362 ;
               RECT 33.254 91.526 33.306 91.562 ;
               RECT 33.254 92.726 33.306 92.762 ;
               RECT 33.254 93.926 33.306 93.962 ;
               RECT 33.254 95.126 33.306 95.162 ;
               RECT 33.254 96.326 33.306 96.362 ;
               RECT 33.254 97.526 33.306 97.562 ;
               RECT 33.254 98.726 33.306 98.762 ;
               RECT 33.254 99.926 33.306 99.962 ;
               RECT 33.254 101.126 33.306 101.162 ;
               RECT 33.254 102.326 33.306 102.362 ;
               RECT 33.254 103.526 33.306 103.562 ;
               RECT 33.334 1.558 33.386 1.594 ;
               RECT 33.334 2.758 33.386 2.794 ;
               RECT 33.334 3.958 33.386 3.994 ;
               RECT 33.334 5.158 33.386 5.194 ;
               RECT 33.334 6.358 33.386 6.394 ;
               RECT 33.334 7.558 33.386 7.594 ;
               RECT 33.334 8.758 33.386 8.794 ;
               RECT 33.334 9.958 33.386 9.994 ;
               RECT 33.334 11.158 33.386 11.194 ;
               RECT 33.334 12.358 33.386 12.394 ;
               RECT 33.334 13.558 33.386 13.594 ;
               RECT 33.334 14.758 33.386 14.794 ;
               RECT 33.334 15.958 33.386 15.994 ;
               RECT 33.334 17.158 33.386 17.194 ;
               RECT 33.334 18.358 33.386 18.394 ;
               RECT 33.334 19.558 33.386 19.594 ;
               RECT 33.334 20.758 33.386 20.794 ;
               RECT 33.334 21.958 33.386 21.994 ;
               RECT 33.334 23.158 33.386 23.194 ;
               RECT 33.334 24.358 33.386 24.394 ;
               RECT 33.334 25.558 33.386 25.594 ;
               RECT 33.334 26.758 33.386 26.794 ;
               RECT 33.334 27.958 33.386 27.994 ;
               RECT 33.334 29.158 33.386 29.194 ;
               RECT 33.334 30.358 33.386 30.394 ;
               RECT 33.334 31.558 33.386 31.594 ;
               RECT 33.334 32.758 33.386 32.794 ;
               RECT 33.334 33.958 33.386 33.994 ;
               RECT 33.334 35.158 33.386 35.194 ;
               RECT 33.334 36.358 33.386 36.394 ;
               RECT 33.334 37.558 33.386 37.594 ;
               RECT 33.334 38.758 33.386 38.794 ;
               RECT 33.334 39.958 33.386 39.994 ;
               RECT 33.334 41.158 33.386 41.194 ;
               RECT 33.334 42.358 33.386 42.394 ;
               RECT 33.334 43.558 33.386 43.594 ;
               RECT 33.334 44.758 33.386 44.794 ;
               RECT 33.334 45.958 33.386 45.994 ;
               RECT 33.334 47.158 33.386 47.194 ;
               RECT 33.334 48.358 33.386 48.394 ;
               RECT 33.334 50.142 33.386 50.178 ;
               RECT 33.334 50.382 33.386 50.418 ;
               RECT 33.334 54.702 33.386 54.738 ;
               RECT 33.334 54.942 33.386 54.978 ;
               RECT 33.334 57.478 33.386 57.514 ;
               RECT 33.334 58.678 33.386 58.714 ;
               RECT 33.334 59.878 33.386 59.914 ;
               RECT 33.334 61.078 33.386 61.114 ;
               RECT 33.334 62.278 33.386 62.314 ;
               RECT 33.334 63.478 33.386 63.514 ;
               RECT 33.334 64.678 33.386 64.714 ;
               RECT 33.334 65.878 33.386 65.914 ;
               RECT 33.334 67.078 33.386 67.114 ;
               RECT 33.334 68.278 33.386 68.314 ;
               RECT 33.334 69.478 33.386 69.514 ;
               RECT 33.334 70.678 33.386 70.714 ;
               RECT 33.334 71.878 33.386 71.914 ;
               RECT 33.334 73.078 33.386 73.114 ;
               RECT 33.334 74.278 33.386 74.314 ;
               RECT 33.334 75.478 33.386 75.514 ;
               RECT 33.334 76.678 33.386 76.714 ;
               RECT 33.334 77.878 33.386 77.914 ;
               RECT 33.334 79.078 33.386 79.114 ;
               RECT 33.334 80.278 33.386 80.314 ;
               RECT 33.334 81.478 33.386 81.514 ;
               RECT 33.334 82.678 33.386 82.714 ;
               RECT 33.334 83.878 33.386 83.914 ;
               RECT 33.334 85.078 33.386 85.114 ;
               RECT 33.334 86.278 33.386 86.314 ;
               RECT 33.334 87.478 33.386 87.514 ;
               RECT 33.334 88.678 33.386 88.714 ;
               RECT 33.334 89.878 33.386 89.914 ;
               RECT 33.334 91.078 33.386 91.114 ;
               RECT 33.334 92.278 33.386 92.314 ;
               RECT 33.334 93.478 33.386 93.514 ;
               RECT 33.334 94.678 33.386 94.714 ;
               RECT 33.334 95.878 33.386 95.914 ;
               RECT 33.334 97.078 33.386 97.114 ;
               RECT 33.334 98.278 33.386 98.314 ;
               RECT 33.334 99.478 33.386 99.514 ;
               RECT 33.334 100.678 33.386 100.714 ;
               RECT 33.334 101.878 33.386 101.914 ;
               RECT 33.334 103.078 33.386 103.114 ;
               RECT 33.334 104.278 33.386 104.314 ;
               RECT 33.414 0.806 33.466 0.842 ;
               RECT 33.414 2.006 33.466 2.042 ;
               RECT 33.414 3.206 33.466 3.242 ;
               RECT 33.414 4.406 33.466 4.442 ;
               RECT 33.414 5.606 33.466 5.642 ;
               RECT 33.414 6.806 33.466 6.842 ;
               RECT 33.414 8.006 33.466 8.042 ;
               RECT 33.414 9.206 33.466 9.242 ;
               RECT 33.414 10.406 33.466 10.442 ;
               RECT 33.414 11.606 33.466 11.642 ;
               RECT 33.414 12.806 33.466 12.842 ;
               RECT 33.414 14.006 33.466 14.042 ;
               RECT 33.414 15.206 33.466 15.242 ;
               RECT 33.414 16.406 33.466 16.442 ;
               RECT 33.414 17.606 33.466 17.642 ;
               RECT 33.414 18.806 33.466 18.842 ;
               RECT 33.414 20.006 33.466 20.042 ;
               RECT 33.414 21.206 33.466 21.242 ;
               RECT 33.414 22.406 33.466 22.442 ;
               RECT 33.414 23.606 33.466 23.642 ;
               RECT 33.414 24.806 33.466 24.842 ;
               RECT 33.414 26.006 33.466 26.042 ;
               RECT 33.414 27.206 33.466 27.242 ;
               RECT 33.414 28.406 33.466 28.442 ;
               RECT 33.414 29.606 33.466 29.642 ;
               RECT 33.414 30.806 33.466 30.842 ;
               RECT 33.414 32.006 33.466 32.042 ;
               RECT 33.414 33.206 33.466 33.242 ;
               RECT 33.414 34.406 33.466 34.442 ;
               RECT 33.414 35.606 33.466 35.642 ;
               RECT 33.414 36.806 33.466 36.842 ;
               RECT 33.414 38.006 33.466 38.042 ;
               RECT 33.414 39.206 33.466 39.242 ;
               RECT 33.414 40.406 33.466 40.442 ;
               RECT 33.414 41.606 33.466 41.642 ;
               RECT 33.414 42.806 33.466 42.842 ;
               RECT 33.414 44.006 33.466 44.042 ;
               RECT 33.414 45.206 33.466 45.242 ;
               RECT 33.414 46.406 33.466 46.442 ;
               RECT 33.414 47.606 33.466 47.642 ;
               RECT 33.414 49.422 33.466 49.458 ;
               RECT 33.414 49.662 33.466 49.698 ;
               RECT 33.414 55.422 33.466 55.458 ;
               RECT 33.414 55.662 33.466 55.698 ;
               RECT 33.414 56.726 33.466 56.762 ;
               RECT 33.414 57.926 33.466 57.962 ;
               RECT 33.414 59.126 33.466 59.162 ;
               RECT 33.414 60.326 33.466 60.362 ;
               RECT 33.414 61.526 33.466 61.562 ;
               RECT 33.414 62.726 33.466 62.762 ;
               RECT 33.414 63.926 33.466 63.962 ;
               RECT 33.414 65.126 33.466 65.162 ;
               RECT 33.414 66.326 33.466 66.362 ;
               RECT 33.414 67.526 33.466 67.562 ;
               RECT 33.414 68.726 33.466 68.762 ;
               RECT 33.414 69.926 33.466 69.962 ;
               RECT 33.414 71.126 33.466 71.162 ;
               RECT 33.414 72.326 33.466 72.362 ;
               RECT 33.414 73.526 33.466 73.562 ;
               RECT 33.414 74.726 33.466 74.762 ;
               RECT 33.414 75.926 33.466 75.962 ;
               RECT 33.414 77.126 33.466 77.162 ;
               RECT 33.414 78.326 33.466 78.362 ;
               RECT 33.414 79.526 33.466 79.562 ;
               RECT 33.414 80.726 33.466 80.762 ;
               RECT 33.414 81.926 33.466 81.962 ;
               RECT 33.414 83.126 33.466 83.162 ;
               RECT 33.414 84.326 33.466 84.362 ;
               RECT 33.414 85.526 33.466 85.562 ;
               RECT 33.414 86.726 33.466 86.762 ;
               RECT 33.414 87.926 33.466 87.962 ;
               RECT 33.414 89.126 33.466 89.162 ;
               RECT 33.414 90.326 33.466 90.362 ;
               RECT 33.414 91.526 33.466 91.562 ;
               RECT 33.414 92.726 33.466 92.762 ;
               RECT 33.414 93.926 33.466 93.962 ;
               RECT 33.414 95.126 33.466 95.162 ;
               RECT 33.414 96.326 33.466 96.362 ;
               RECT 33.414 97.526 33.466 97.562 ;
               RECT 33.414 98.726 33.466 98.762 ;
               RECT 33.414 99.926 33.466 99.962 ;
               RECT 33.414 101.126 33.466 101.162 ;
               RECT 33.414 102.326 33.466 102.362 ;
               RECT 33.414 103.526 33.466 103.562 ;
               RECT 33.494 1.558 33.546 1.594 ;
               RECT 33.494 2.758 33.546 2.794 ;
               RECT 33.494 3.958 33.546 3.994 ;
               RECT 33.494 5.158 33.546 5.194 ;
               RECT 33.494 6.358 33.546 6.394 ;
               RECT 33.494 7.558 33.546 7.594 ;
               RECT 33.494 8.758 33.546 8.794 ;
               RECT 33.494 9.958 33.546 9.994 ;
               RECT 33.494 11.158 33.546 11.194 ;
               RECT 33.494 12.358 33.546 12.394 ;
               RECT 33.494 13.558 33.546 13.594 ;
               RECT 33.494 14.758 33.546 14.794 ;
               RECT 33.494 15.958 33.546 15.994 ;
               RECT 33.494 17.158 33.546 17.194 ;
               RECT 33.494 18.358 33.546 18.394 ;
               RECT 33.494 19.558 33.546 19.594 ;
               RECT 33.494 20.758 33.546 20.794 ;
               RECT 33.494 21.958 33.546 21.994 ;
               RECT 33.494 23.158 33.546 23.194 ;
               RECT 33.494 24.358 33.546 24.394 ;
               RECT 33.494 25.558 33.546 25.594 ;
               RECT 33.494 26.758 33.546 26.794 ;
               RECT 33.494 27.958 33.546 27.994 ;
               RECT 33.494 29.158 33.546 29.194 ;
               RECT 33.494 30.358 33.546 30.394 ;
               RECT 33.494 31.558 33.546 31.594 ;
               RECT 33.494 32.758 33.546 32.794 ;
               RECT 33.494 33.958 33.546 33.994 ;
               RECT 33.494 35.158 33.546 35.194 ;
               RECT 33.494 36.358 33.546 36.394 ;
               RECT 33.494 37.558 33.546 37.594 ;
               RECT 33.494 38.758 33.546 38.794 ;
               RECT 33.494 39.958 33.546 39.994 ;
               RECT 33.494 41.158 33.546 41.194 ;
               RECT 33.494 42.358 33.546 42.394 ;
               RECT 33.494 43.558 33.546 43.594 ;
               RECT 33.494 44.758 33.546 44.794 ;
               RECT 33.494 45.958 33.546 45.994 ;
               RECT 33.494 47.158 33.546 47.194 ;
               RECT 33.494 48.358 33.546 48.394 ;
               RECT 33.494 50.142 33.546 50.178 ;
               RECT 33.494 50.382 33.546 50.418 ;
               RECT 33.494 54.702 33.546 54.738 ;
               RECT 33.494 54.942 33.546 54.978 ;
               RECT 33.494 57.478 33.546 57.514 ;
               RECT 33.494 58.678 33.546 58.714 ;
               RECT 33.494 59.878 33.546 59.914 ;
               RECT 33.494 61.078 33.546 61.114 ;
               RECT 33.494 62.278 33.546 62.314 ;
               RECT 33.494 63.478 33.546 63.514 ;
               RECT 33.494 64.678 33.546 64.714 ;
               RECT 33.494 65.878 33.546 65.914 ;
               RECT 33.494 67.078 33.546 67.114 ;
               RECT 33.494 68.278 33.546 68.314 ;
               RECT 33.494 69.478 33.546 69.514 ;
               RECT 33.494 70.678 33.546 70.714 ;
               RECT 33.494 71.878 33.546 71.914 ;
               RECT 33.494 73.078 33.546 73.114 ;
               RECT 33.494 74.278 33.546 74.314 ;
               RECT 33.494 75.478 33.546 75.514 ;
               RECT 33.494 76.678 33.546 76.714 ;
               RECT 33.494 77.878 33.546 77.914 ;
               RECT 33.494 79.078 33.546 79.114 ;
               RECT 33.494 80.278 33.546 80.314 ;
               RECT 33.494 81.478 33.546 81.514 ;
               RECT 33.494 82.678 33.546 82.714 ;
               RECT 33.494 83.878 33.546 83.914 ;
               RECT 33.494 85.078 33.546 85.114 ;
               RECT 33.494 86.278 33.546 86.314 ;
               RECT 33.494 87.478 33.546 87.514 ;
               RECT 33.494 88.678 33.546 88.714 ;
               RECT 33.494 89.878 33.546 89.914 ;
               RECT 33.494 91.078 33.546 91.114 ;
               RECT 33.494 92.278 33.546 92.314 ;
               RECT 33.494 93.478 33.546 93.514 ;
               RECT 33.494 94.678 33.546 94.714 ;
               RECT 33.494 95.878 33.546 95.914 ;
               RECT 33.494 97.078 33.546 97.114 ;
               RECT 33.494 98.278 33.546 98.314 ;
               RECT 33.494 99.478 33.546 99.514 ;
               RECT 33.494 100.678 33.546 100.714 ;
               RECT 33.494 101.878 33.546 101.914 ;
               RECT 33.494 103.078 33.546 103.114 ;
               RECT 33.494 104.278 33.546 104.314 ;
               RECT 33.574 0.281 33.626 0.317 ;
               RECT 33.574 104.803 33.626 104.839 ;
               RECT 33.654 0.806 33.706 0.842 ;
               RECT 33.654 2.006 33.706 2.042 ;
               RECT 33.654 3.206 33.706 3.242 ;
               RECT 33.654 4.406 33.706 4.442 ;
               RECT 33.654 5.606 33.706 5.642 ;
               RECT 33.654 6.806 33.706 6.842 ;
               RECT 33.654 8.006 33.706 8.042 ;
               RECT 33.654 9.206 33.706 9.242 ;
               RECT 33.654 10.406 33.706 10.442 ;
               RECT 33.654 11.606 33.706 11.642 ;
               RECT 33.654 12.806 33.706 12.842 ;
               RECT 33.654 14.006 33.706 14.042 ;
               RECT 33.654 15.206 33.706 15.242 ;
               RECT 33.654 16.406 33.706 16.442 ;
               RECT 33.654 17.606 33.706 17.642 ;
               RECT 33.654 18.806 33.706 18.842 ;
               RECT 33.654 20.006 33.706 20.042 ;
               RECT 33.654 21.206 33.706 21.242 ;
               RECT 33.654 22.406 33.706 22.442 ;
               RECT 33.654 23.606 33.706 23.642 ;
               RECT 33.654 24.806 33.706 24.842 ;
               RECT 33.654 26.006 33.706 26.042 ;
               RECT 33.654 27.206 33.706 27.242 ;
               RECT 33.654 28.406 33.706 28.442 ;
               RECT 33.654 29.606 33.706 29.642 ;
               RECT 33.654 30.806 33.706 30.842 ;
               RECT 33.654 32.006 33.706 32.042 ;
               RECT 33.654 33.206 33.706 33.242 ;
               RECT 33.654 34.406 33.706 34.442 ;
               RECT 33.654 35.606 33.706 35.642 ;
               RECT 33.654 36.806 33.706 36.842 ;
               RECT 33.654 38.006 33.706 38.042 ;
               RECT 33.654 39.206 33.706 39.242 ;
               RECT 33.654 40.406 33.706 40.442 ;
               RECT 33.654 41.606 33.706 41.642 ;
               RECT 33.654 42.806 33.706 42.842 ;
               RECT 33.654 44.006 33.706 44.042 ;
               RECT 33.654 45.206 33.706 45.242 ;
               RECT 33.654 46.406 33.706 46.442 ;
               RECT 33.654 47.606 33.706 47.642 ;
               RECT 33.654 49.422 33.706 49.458 ;
               RECT 33.654 49.662 33.706 49.698 ;
               RECT 33.654 51.102 33.706 51.138 ;
               RECT 33.654 51.582 33.706 51.618 ;
               RECT 33.654 53.502 33.706 53.538 ;
               RECT 33.654 53.982 33.706 54.018 ;
               RECT 33.654 55.422 33.706 55.458 ;
               RECT 33.654 55.662 33.706 55.698 ;
               RECT 33.654 56.726 33.706 56.762 ;
               RECT 33.654 57.926 33.706 57.962 ;
               RECT 33.654 59.126 33.706 59.162 ;
               RECT 33.654 60.326 33.706 60.362 ;
               RECT 33.654 61.526 33.706 61.562 ;
               RECT 33.654 62.726 33.706 62.762 ;
               RECT 33.654 63.926 33.706 63.962 ;
               RECT 33.654 65.126 33.706 65.162 ;
               RECT 33.654 66.326 33.706 66.362 ;
               RECT 33.654 67.526 33.706 67.562 ;
               RECT 33.654 68.726 33.706 68.762 ;
               RECT 33.654 69.926 33.706 69.962 ;
               RECT 33.654 71.126 33.706 71.162 ;
               RECT 33.654 72.326 33.706 72.362 ;
               RECT 33.654 73.526 33.706 73.562 ;
               RECT 33.654 74.726 33.706 74.762 ;
               RECT 33.654 75.926 33.706 75.962 ;
               RECT 33.654 77.126 33.706 77.162 ;
               RECT 33.654 78.326 33.706 78.362 ;
               RECT 33.654 79.526 33.706 79.562 ;
               RECT 33.654 80.726 33.706 80.762 ;
               RECT 33.654 81.926 33.706 81.962 ;
               RECT 33.654 83.126 33.706 83.162 ;
               RECT 33.654 84.326 33.706 84.362 ;
               RECT 33.654 85.526 33.706 85.562 ;
               RECT 33.654 86.726 33.706 86.762 ;
               RECT 33.654 87.926 33.706 87.962 ;
               RECT 33.654 89.126 33.706 89.162 ;
               RECT 33.654 90.326 33.706 90.362 ;
               RECT 33.654 91.526 33.706 91.562 ;
               RECT 33.654 92.726 33.706 92.762 ;
               RECT 33.654 93.926 33.706 93.962 ;
               RECT 33.654 95.126 33.706 95.162 ;
               RECT 33.654 96.326 33.706 96.362 ;
               RECT 33.654 97.526 33.706 97.562 ;
               RECT 33.654 98.726 33.706 98.762 ;
               RECT 33.654 99.926 33.706 99.962 ;
               RECT 33.654 101.126 33.706 101.162 ;
               RECT 33.654 102.326 33.706 102.362 ;
               RECT 33.654 103.526 33.706 103.562 ;
               RECT 33.734 1.558 33.786 1.594 ;
               RECT 33.734 2.758 33.786 2.794 ;
               RECT 33.734 3.958 33.786 3.994 ;
               RECT 33.734 5.158 33.786 5.194 ;
               RECT 33.734 6.358 33.786 6.394 ;
               RECT 33.734 7.558 33.786 7.594 ;
               RECT 33.734 8.758 33.786 8.794 ;
               RECT 33.734 9.958 33.786 9.994 ;
               RECT 33.734 11.158 33.786 11.194 ;
               RECT 33.734 12.358 33.786 12.394 ;
               RECT 33.734 13.558 33.786 13.594 ;
               RECT 33.734 14.758 33.786 14.794 ;
               RECT 33.734 15.958 33.786 15.994 ;
               RECT 33.734 17.158 33.786 17.194 ;
               RECT 33.734 18.358 33.786 18.394 ;
               RECT 33.734 19.558 33.786 19.594 ;
               RECT 33.734 20.758 33.786 20.794 ;
               RECT 33.734 21.958 33.786 21.994 ;
               RECT 33.734 23.158 33.786 23.194 ;
               RECT 33.734 24.358 33.786 24.394 ;
               RECT 33.734 25.558 33.786 25.594 ;
               RECT 33.734 26.758 33.786 26.794 ;
               RECT 33.734 27.958 33.786 27.994 ;
               RECT 33.734 29.158 33.786 29.194 ;
               RECT 33.734 30.358 33.786 30.394 ;
               RECT 33.734 31.558 33.786 31.594 ;
               RECT 33.734 32.758 33.786 32.794 ;
               RECT 33.734 33.958 33.786 33.994 ;
               RECT 33.734 35.158 33.786 35.194 ;
               RECT 33.734 36.358 33.786 36.394 ;
               RECT 33.734 37.558 33.786 37.594 ;
               RECT 33.734 38.758 33.786 38.794 ;
               RECT 33.734 39.958 33.786 39.994 ;
               RECT 33.734 41.158 33.786 41.194 ;
               RECT 33.734 42.358 33.786 42.394 ;
               RECT 33.734 43.558 33.786 43.594 ;
               RECT 33.734 44.758 33.786 44.794 ;
               RECT 33.734 45.958 33.786 45.994 ;
               RECT 33.734 47.158 33.786 47.194 ;
               RECT 33.734 48.358 33.786 48.394 ;
               RECT 33.734 50.142 33.786 50.178 ;
               RECT 33.734 50.382 33.786 50.418 ;
               RECT 33.734 54.702 33.786 54.738 ;
               RECT 33.734 54.942 33.786 54.978 ;
               RECT 33.734 57.478 33.786 57.514 ;
               RECT 33.734 58.678 33.786 58.714 ;
               RECT 33.734 59.878 33.786 59.914 ;
               RECT 33.734 61.078 33.786 61.114 ;
               RECT 33.734 62.278 33.786 62.314 ;
               RECT 33.734 63.478 33.786 63.514 ;
               RECT 33.734 64.678 33.786 64.714 ;
               RECT 33.734 65.878 33.786 65.914 ;
               RECT 33.734 67.078 33.786 67.114 ;
               RECT 33.734 68.278 33.786 68.314 ;
               RECT 33.734 69.478 33.786 69.514 ;
               RECT 33.734 70.678 33.786 70.714 ;
               RECT 33.734 71.878 33.786 71.914 ;
               RECT 33.734 73.078 33.786 73.114 ;
               RECT 33.734 74.278 33.786 74.314 ;
               RECT 33.734 75.478 33.786 75.514 ;
               RECT 33.734 76.678 33.786 76.714 ;
               RECT 33.734 77.878 33.786 77.914 ;
               RECT 33.734 79.078 33.786 79.114 ;
               RECT 33.734 80.278 33.786 80.314 ;
               RECT 33.734 81.478 33.786 81.514 ;
               RECT 33.734 82.678 33.786 82.714 ;
               RECT 33.734 83.878 33.786 83.914 ;
               RECT 33.734 85.078 33.786 85.114 ;
               RECT 33.734 86.278 33.786 86.314 ;
               RECT 33.734 87.478 33.786 87.514 ;
               RECT 33.734 88.678 33.786 88.714 ;
               RECT 33.734 89.878 33.786 89.914 ;
               RECT 33.734 91.078 33.786 91.114 ;
               RECT 33.734 92.278 33.786 92.314 ;
               RECT 33.734 93.478 33.786 93.514 ;
               RECT 33.734 94.678 33.786 94.714 ;
               RECT 33.734 95.878 33.786 95.914 ;
               RECT 33.734 97.078 33.786 97.114 ;
               RECT 33.734 98.278 33.786 98.314 ;
               RECT 33.734 99.478 33.786 99.514 ;
               RECT 33.734 100.678 33.786 100.714 ;
               RECT 33.734 101.878 33.786 101.914 ;
               RECT 33.734 103.078 33.786 103.114 ;
               RECT 33.734 104.278 33.786 104.314 ;
               RECT 33.814 0.806 33.866 0.842 ;
               RECT 33.814 2.006 33.866 2.042 ;
               RECT 33.814 3.206 33.866 3.242 ;
               RECT 33.814 4.406 33.866 4.442 ;
               RECT 33.814 5.606 33.866 5.642 ;
               RECT 33.814 6.806 33.866 6.842 ;
               RECT 33.814 8.006 33.866 8.042 ;
               RECT 33.814 9.206 33.866 9.242 ;
               RECT 33.814 10.406 33.866 10.442 ;
               RECT 33.814 11.606 33.866 11.642 ;
               RECT 33.814 12.806 33.866 12.842 ;
               RECT 33.814 14.006 33.866 14.042 ;
               RECT 33.814 15.206 33.866 15.242 ;
               RECT 33.814 16.406 33.866 16.442 ;
               RECT 33.814 17.606 33.866 17.642 ;
               RECT 33.814 18.806 33.866 18.842 ;
               RECT 33.814 20.006 33.866 20.042 ;
               RECT 33.814 21.206 33.866 21.242 ;
               RECT 33.814 22.406 33.866 22.442 ;
               RECT 33.814 23.606 33.866 23.642 ;
               RECT 33.814 24.806 33.866 24.842 ;
               RECT 33.814 26.006 33.866 26.042 ;
               RECT 33.814 27.206 33.866 27.242 ;
               RECT 33.814 28.406 33.866 28.442 ;
               RECT 33.814 29.606 33.866 29.642 ;
               RECT 33.814 30.806 33.866 30.842 ;
               RECT 33.814 32.006 33.866 32.042 ;
               RECT 33.814 33.206 33.866 33.242 ;
               RECT 33.814 34.406 33.866 34.442 ;
               RECT 33.814 35.606 33.866 35.642 ;
               RECT 33.814 36.806 33.866 36.842 ;
               RECT 33.814 38.006 33.866 38.042 ;
               RECT 33.814 39.206 33.866 39.242 ;
               RECT 33.814 40.406 33.866 40.442 ;
               RECT 33.814 41.606 33.866 41.642 ;
               RECT 33.814 42.806 33.866 42.842 ;
               RECT 33.814 44.006 33.866 44.042 ;
               RECT 33.814 45.206 33.866 45.242 ;
               RECT 33.814 46.406 33.866 46.442 ;
               RECT 33.814 47.606 33.866 47.642 ;
               RECT 33.814 49.422 33.866 49.458 ;
               RECT 33.814 49.662 33.866 49.698 ;
               RECT 33.814 55.422 33.866 55.458 ;
               RECT 33.814 55.662 33.866 55.698 ;
               RECT 33.814 56.726 33.866 56.762 ;
               RECT 33.814 57.926 33.866 57.962 ;
               RECT 33.814 59.126 33.866 59.162 ;
               RECT 33.814 60.326 33.866 60.362 ;
               RECT 33.814 61.526 33.866 61.562 ;
               RECT 33.814 62.726 33.866 62.762 ;
               RECT 33.814 63.926 33.866 63.962 ;
               RECT 33.814 65.126 33.866 65.162 ;
               RECT 33.814 66.326 33.866 66.362 ;
               RECT 33.814 67.526 33.866 67.562 ;
               RECT 33.814 68.726 33.866 68.762 ;
               RECT 33.814 69.926 33.866 69.962 ;
               RECT 33.814 71.126 33.866 71.162 ;
               RECT 33.814 72.326 33.866 72.362 ;
               RECT 33.814 73.526 33.866 73.562 ;
               RECT 33.814 74.726 33.866 74.762 ;
               RECT 33.814 75.926 33.866 75.962 ;
               RECT 33.814 77.126 33.866 77.162 ;
               RECT 33.814 78.326 33.866 78.362 ;
               RECT 33.814 79.526 33.866 79.562 ;
               RECT 33.814 80.726 33.866 80.762 ;
               RECT 33.814 81.926 33.866 81.962 ;
               RECT 33.814 83.126 33.866 83.162 ;
               RECT 33.814 84.326 33.866 84.362 ;
               RECT 33.814 85.526 33.866 85.562 ;
               RECT 33.814 86.726 33.866 86.762 ;
               RECT 33.814 87.926 33.866 87.962 ;
               RECT 33.814 89.126 33.866 89.162 ;
               RECT 33.814 90.326 33.866 90.362 ;
               RECT 33.814 91.526 33.866 91.562 ;
               RECT 33.814 92.726 33.866 92.762 ;
               RECT 33.814 93.926 33.866 93.962 ;
               RECT 33.814 95.126 33.866 95.162 ;
               RECT 33.814 96.326 33.866 96.362 ;
               RECT 33.814 97.526 33.866 97.562 ;
               RECT 33.814 98.726 33.866 98.762 ;
               RECT 33.814 99.926 33.866 99.962 ;
               RECT 33.814 101.126 33.866 101.162 ;
               RECT 33.814 102.326 33.866 102.362 ;
               RECT 33.814 103.526 33.866 103.562 ;
               RECT 33.894 1.558 33.946 1.594 ;
               RECT 33.894 2.758 33.946 2.794 ;
               RECT 33.894 3.958 33.946 3.994 ;
               RECT 33.894 5.158 33.946 5.194 ;
               RECT 33.894 6.358 33.946 6.394 ;
               RECT 33.894 7.558 33.946 7.594 ;
               RECT 33.894 8.758 33.946 8.794 ;
               RECT 33.894 9.958 33.946 9.994 ;
               RECT 33.894 11.158 33.946 11.194 ;
               RECT 33.894 12.358 33.946 12.394 ;
               RECT 33.894 13.558 33.946 13.594 ;
               RECT 33.894 14.758 33.946 14.794 ;
               RECT 33.894 15.958 33.946 15.994 ;
               RECT 33.894 17.158 33.946 17.194 ;
               RECT 33.894 18.358 33.946 18.394 ;
               RECT 33.894 19.558 33.946 19.594 ;
               RECT 33.894 20.758 33.946 20.794 ;
               RECT 33.894 21.958 33.946 21.994 ;
               RECT 33.894 23.158 33.946 23.194 ;
               RECT 33.894 24.358 33.946 24.394 ;
               RECT 33.894 25.558 33.946 25.594 ;
               RECT 33.894 26.758 33.946 26.794 ;
               RECT 33.894 27.958 33.946 27.994 ;
               RECT 33.894 29.158 33.946 29.194 ;
               RECT 33.894 30.358 33.946 30.394 ;
               RECT 33.894 31.558 33.946 31.594 ;
               RECT 33.894 32.758 33.946 32.794 ;
               RECT 33.894 33.958 33.946 33.994 ;
               RECT 33.894 35.158 33.946 35.194 ;
               RECT 33.894 36.358 33.946 36.394 ;
               RECT 33.894 37.558 33.946 37.594 ;
               RECT 33.894 38.758 33.946 38.794 ;
               RECT 33.894 39.958 33.946 39.994 ;
               RECT 33.894 41.158 33.946 41.194 ;
               RECT 33.894 42.358 33.946 42.394 ;
               RECT 33.894 43.558 33.946 43.594 ;
               RECT 33.894 44.758 33.946 44.794 ;
               RECT 33.894 45.958 33.946 45.994 ;
               RECT 33.894 47.158 33.946 47.194 ;
               RECT 33.894 48.358 33.946 48.394 ;
               RECT 33.894 50.142 33.946 50.178 ;
               RECT 33.894 50.382 33.946 50.418 ;
               RECT 33.894 54.702 33.946 54.738 ;
               RECT 33.894 54.942 33.946 54.978 ;
               RECT 33.894 57.478 33.946 57.514 ;
               RECT 33.894 58.678 33.946 58.714 ;
               RECT 33.894 59.878 33.946 59.914 ;
               RECT 33.894 61.078 33.946 61.114 ;
               RECT 33.894 62.278 33.946 62.314 ;
               RECT 33.894 63.478 33.946 63.514 ;
               RECT 33.894 64.678 33.946 64.714 ;
               RECT 33.894 65.878 33.946 65.914 ;
               RECT 33.894 67.078 33.946 67.114 ;
               RECT 33.894 68.278 33.946 68.314 ;
               RECT 33.894 69.478 33.946 69.514 ;
               RECT 33.894 70.678 33.946 70.714 ;
               RECT 33.894 71.878 33.946 71.914 ;
               RECT 33.894 73.078 33.946 73.114 ;
               RECT 33.894 74.278 33.946 74.314 ;
               RECT 33.894 75.478 33.946 75.514 ;
               RECT 33.894 76.678 33.946 76.714 ;
               RECT 33.894 77.878 33.946 77.914 ;
               RECT 33.894 79.078 33.946 79.114 ;
               RECT 33.894 80.278 33.946 80.314 ;
               RECT 33.894 81.478 33.946 81.514 ;
               RECT 33.894 82.678 33.946 82.714 ;
               RECT 33.894 83.878 33.946 83.914 ;
               RECT 33.894 85.078 33.946 85.114 ;
               RECT 33.894 86.278 33.946 86.314 ;
               RECT 33.894 87.478 33.946 87.514 ;
               RECT 33.894 88.678 33.946 88.714 ;
               RECT 33.894 89.878 33.946 89.914 ;
               RECT 33.894 91.078 33.946 91.114 ;
               RECT 33.894 92.278 33.946 92.314 ;
               RECT 33.894 93.478 33.946 93.514 ;
               RECT 33.894 94.678 33.946 94.714 ;
               RECT 33.894 95.878 33.946 95.914 ;
               RECT 33.894 97.078 33.946 97.114 ;
               RECT 33.894 98.278 33.946 98.314 ;
               RECT 33.894 99.478 33.946 99.514 ;
               RECT 33.894 100.678 33.946 100.714 ;
               RECT 33.894 101.878 33.946 101.914 ;
               RECT 33.894 103.078 33.946 103.114 ;
               RECT 33.894 104.278 33.946 104.314 ;
               RECT 33.974 0.281 34.026 0.317 ;
               RECT 33.974 104.803 34.026 104.839 ;
               RECT 34.054 0.806 34.106 0.842 ;
               RECT 34.054 2.006 34.106 2.042 ;
               RECT 34.054 3.206 34.106 3.242 ;
               RECT 34.054 4.406 34.106 4.442 ;
               RECT 34.054 5.606 34.106 5.642 ;
               RECT 34.054 6.806 34.106 6.842 ;
               RECT 34.054 8.006 34.106 8.042 ;
               RECT 34.054 9.206 34.106 9.242 ;
               RECT 34.054 10.406 34.106 10.442 ;
               RECT 34.054 11.606 34.106 11.642 ;
               RECT 34.054 12.806 34.106 12.842 ;
               RECT 34.054 14.006 34.106 14.042 ;
               RECT 34.054 15.206 34.106 15.242 ;
               RECT 34.054 16.406 34.106 16.442 ;
               RECT 34.054 17.606 34.106 17.642 ;
               RECT 34.054 18.806 34.106 18.842 ;
               RECT 34.054 20.006 34.106 20.042 ;
               RECT 34.054 21.206 34.106 21.242 ;
               RECT 34.054 22.406 34.106 22.442 ;
               RECT 34.054 23.606 34.106 23.642 ;
               RECT 34.054 24.806 34.106 24.842 ;
               RECT 34.054 26.006 34.106 26.042 ;
               RECT 34.054 27.206 34.106 27.242 ;
               RECT 34.054 28.406 34.106 28.442 ;
               RECT 34.054 29.606 34.106 29.642 ;
               RECT 34.054 30.806 34.106 30.842 ;
               RECT 34.054 32.006 34.106 32.042 ;
               RECT 34.054 33.206 34.106 33.242 ;
               RECT 34.054 34.406 34.106 34.442 ;
               RECT 34.054 35.606 34.106 35.642 ;
               RECT 34.054 36.806 34.106 36.842 ;
               RECT 34.054 38.006 34.106 38.042 ;
               RECT 34.054 39.206 34.106 39.242 ;
               RECT 34.054 40.406 34.106 40.442 ;
               RECT 34.054 41.606 34.106 41.642 ;
               RECT 34.054 42.806 34.106 42.842 ;
               RECT 34.054 44.006 34.106 44.042 ;
               RECT 34.054 45.206 34.106 45.242 ;
               RECT 34.054 46.406 34.106 46.442 ;
               RECT 34.054 47.606 34.106 47.642 ;
               RECT 34.054 49.422 34.106 49.458 ;
               RECT 34.054 49.662 34.106 49.698 ;
               RECT 34.054 55.422 34.106 55.458 ;
               RECT 34.054 55.662 34.106 55.698 ;
               RECT 34.054 56.726 34.106 56.762 ;
               RECT 34.054 57.926 34.106 57.962 ;
               RECT 34.054 59.126 34.106 59.162 ;
               RECT 34.054 60.326 34.106 60.362 ;
               RECT 34.054 61.526 34.106 61.562 ;
               RECT 34.054 62.726 34.106 62.762 ;
               RECT 34.054 63.926 34.106 63.962 ;
               RECT 34.054 65.126 34.106 65.162 ;
               RECT 34.054 66.326 34.106 66.362 ;
               RECT 34.054 67.526 34.106 67.562 ;
               RECT 34.054 68.726 34.106 68.762 ;
               RECT 34.054 69.926 34.106 69.962 ;
               RECT 34.054 71.126 34.106 71.162 ;
               RECT 34.054 72.326 34.106 72.362 ;
               RECT 34.054 73.526 34.106 73.562 ;
               RECT 34.054 74.726 34.106 74.762 ;
               RECT 34.054 75.926 34.106 75.962 ;
               RECT 34.054 77.126 34.106 77.162 ;
               RECT 34.054 78.326 34.106 78.362 ;
               RECT 34.054 79.526 34.106 79.562 ;
               RECT 34.054 80.726 34.106 80.762 ;
               RECT 34.054 81.926 34.106 81.962 ;
               RECT 34.054 83.126 34.106 83.162 ;
               RECT 34.054 84.326 34.106 84.362 ;
               RECT 34.054 85.526 34.106 85.562 ;
               RECT 34.054 86.726 34.106 86.762 ;
               RECT 34.054 87.926 34.106 87.962 ;
               RECT 34.054 89.126 34.106 89.162 ;
               RECT 34.054 90.326 34.106 90.362 ;
               RECT 34.054 91.526 34.106 91.562 ;
               RECT 34.054 92.726 34.106 92.762 ;
               RECT 34.054 93.926 34.106 93.962 ;
               RECT 34.054 95.126 34.106 95.162 ;
               RECT 34.054 96.326 34.106 96.362 ;
               RECT 34.054 97.526 34.106 97.562 ;
               RECT 34.054 98.726 34.106 98.762 ;
               RECT 34.054 99.926 34.106 99.962 ;
               RECT 34.054 101.126 34.106 101.162 ;
               RECT 34.054 102.326 34.106 102.362 ;
               RECT 34.054 103.526 34.106 103.562 ;
               RECT 34.134 1.558 34.186 1.594 ;
               RECT 34.134 2.758 34.186 2.794 ;
               RECT 34.134 3.958 34.186 3.994 ;
               RECT 34.134 5.158 34.186 5.194 ;
               RECT 34.134 6.358 34.186 6.394 ;
               RECT 34.134 7.558 34.186 7.594 ;
               RECT 34.134 8.758 34.186 8.794 ;
               RECT 34.134 9.958 34.186 9.994 ;
               RECT 34.134 11.158 34.186 11.194 ;
               RECT 34.134 12.358 34.186 12.394 ;
               RECT 34.134 13.558 34.186 13.594 ;
               RECT 34.134 14.758 34.186 14.794 ;
               RECT 34.134 15.958 34.186 15.994 ;
               RECT 34.134 17.158 34.186 17.194 ;
               RECT 34.134 18.358 34.186 18.394 ;
               RECT 34.134 19.558 34.186 19.594 ;
               RECT 34.134 20.758 34.186 20.794 ;
               RECT 34.134 21.958 34.186 21.994 ;
               RECT 34.134 23.158 34.186 23.194 ;
               RECT 34.134 24.358 34.186 24.394 ;
               RECT 34.134 25.558 34.186 25.594 ;
               RECT 34.134 26.758 34.186 26.794 ;
               RECT 34.134 27.958 34.186 27.994 ;
               RECT 34.134 29.158 34.186 29.194 ;
               RECT 34.134 30.358 34.186 30.394 ;
               RECT 34.134 31.558 34.186 31.594 ;
               RECT 34.134 32.758 34.186 32.794 ;
               RECT 34.134 33.958 34.186 33.994 ;
               RECT 34.134 35.158 34.186 35.194 ;
               RECT 34.134 36.358 34.186 36.394 ;
               RECT 34.134 37.558 34.186 37.594 ;
               RECT 34.134 38.758 34.186 38.794 ;
               RECT 34.134 39.958 34.186 39.994 ;
               RECT 34.134 41.158 34.186 41.194 ;
               RECT 34.134 42.358 34.186 42.394 ;
               RECT 34.134 43.558 34.186 43.594 ;
               RECT 34.134 44.758 34.186 44.794 ;
               RECT 34.134 45.958 34.186 45.994 ;
               RECT 34.134 47.158 34.186 47.194 ;
               RECT 34.134 48.358 34.186 48.394 ;
               RECT 34.134 50.142 34.186 50.178 ;
               RECT 34.134 50.382 34.186 50.418 ;
               RECT 34.134 54.702 34.186 54.738 ;
               RECT 34.134 54.942 34.186 54.978 ;
               RECT 34.134 57.478 34.186 57.514 ;
               RECT 34.134 58.678 34.186 58.714 ;
               RECT 34.134 59.878 34.186 59.914 ;
               RECT 34.134 61.078 34.186 61.114 ;
               RECT 34.134 62.278 34.186 62.314 ;
               RECT 34.134 63.478 34.186 63.514 ;
               RECT 34.134 64.678 34.186 64.714 ;
               RECT 34.134 65.878 34.186 65.914 ;
               RECT 34.134 67.078 34.186 67.114 ;
               RECT 34.134 68.278 34.186 68.314 ;
               RECT 34.134 69.478 34.186 69.514 ;
               RECT 34.134 70.678 34.186 70.714 ;
               RECT 34.134 71.878 34.186 71.914 ;
               RECT 34.134 73.078 34.186 73.114 ;
               RECT 34.134 74.278 34.186 74.314 ;
               RECT 34.134 75.478 34.186 75.514 ;
               RECT 34.134 76.678 34.186 76.714 ;
               RECT 34.134 77.878 34.186 77.914 ;
               RECT 34.134 79.078 34.186 79.114 ;
               RECT 34.134 80.278 34.186 80.314 ;
               RECT 34.134 81.478 34.186 81.514 ;
               RECT 34.134 82.678 34.186 82.714 ;
               RECT 34.134 83.878 34.186 83.914 ;
               RECT 34.134 85.078 34.186 85.114 ;
               RECT 34.134 86.278 34.186 86.314 ;
               RECT 34.134 87.478 34.186 87.514 ;
               RECT 34.134 88.678 34.186 88.714 ;
               RECT 34.134 89.878 34.186 89.914 ;
               RECT 34.134 91.078 34.186 91.114 ;
               RECT 34.134 92.278 34.186 92.314 ;
               RECT 34.134 93.478 34.186 93.514 ;
               RECT 34.134 94.678 34.186 94.714 ;
               RECT 34.134 95.878 34.186 95.914 ;
               RECT 34.134 97.078 34.186 97.114 ;
               RECT 34.134 98.278 34.186 98.314 ;
               RECT 34.134 99.478 34.186 99.514 ;
               RECT 34.134 100.678 34.186 100.714 ;
               RECT 34.134 101.878 34.186 101.914 ;
               RECT 34.134 103.078 34.186 103.114 ;
               RECT 34.134 104.278 34.186 104.314 ;
               RECT 34.214 0.806 34.266 0.842 ;
               RECT 34.214 2.006 34.266 2.042 ;
               RECT 34.214 3.206 34.266 3.242 ;
               RECT 34.214 4.406 34.266 4.442 ;
               RECT 34.214 5.606 34.266 5.642 ;
               RECT 34.214 6.806 34.266 6.842 ;
               RECT 34.214 8.006 34.266 8.042 ;
               RECT 34.214 9.206 34.266 9.242 ;
               RECT 34.214 10.406 34.266 10.442 ;
               RECT 34.214 11.606 34.266 11.642 ;
               RECT 34.214 12.806 34.266 12.842 ;
               RECT 34.214 14.006 34.266 14.042 ;
               RECT 34.214 15.206 34.266 15.242 ;
               RECT 34.214 16.406 34.266 16.442 ;
               RECT 34.214 17.606 34.266 17.642 ;
               RECT 34.214 18.806 34.266 18.842 ;
               RECT 34.214 20.006 34.266 20.042 ;
               RECT 34.214 21.206 34.266 21.242 ;
               RECT 34.214 22.406 34.266 22.442 ;
               RECT 34.214 23.606 34.266 23.642 ;
               RECT 34.214 24.806 34.266 24.842 ;
               RECT 34.214 26.006 34.266 26.042 ;
               RECT 34.214 27.206 34.266 27.242 ;
               RECT 34.214 28.406 34.266 28.442 ;
               RECT 34.214 29.606 34.266 29.642 ;
               RECT 34.214 30.806 34.266 30.842 ;
               RECT 34.214 32.006 34.266 32.042 ;
               RECT 34.214 33.206 34.266 33.242 ;
               RECT 34.214 34.406 34.266 34.442 ;
               RECT 34.214 35.606 34.266 35.642 ;
               RECT 34.214 36.806 34.266 36.842 ;
               RECT 34.214 38.006 34.266 38.042 ;
               RECT 34.214 39.206 34.266 39.242 ;
               RECT 34.214 40.406 34.266 40.442 ;
               RECT 34.214 41.606 34.266 41.642 ;
               RECT 34.214 42.806 34.266 42.842 ;
               RECT 34.214 44.006 34.266 44.042 ;
               RECT 34.214 45.206 34.266 45.242 ;
               RECT 34.214 46.406 34.266 46.442 ;
               RECT 34.214 47.606 34.266 47.642 ;
               RECT 34.214 49.422 34.266 49.458 ;
               RECT 34.214 49.662 34.266 49.698 ;
               RECT 34.214 55.422 34.266 55.458 ;
               RECT 34.214 55.662 34.266 55.698 ;
               RECT 34.214 56.726 34.266 56.762 ;
               RECT 34.214 57.926 34.266 57.962 ;
               RECT 34.214 59.126 34.266 59.162 ;
               RECT 34.214 60.326 34.266 60.362 ;
               RECT 34.214 61.526 34.266 61.562 ;
               RECT 34.214 62.726 34.266 62.762 ;
               RECT 34.214 63.926 34.266 63.962 ;
               RECT 34.214 65.126 34.266 65.162 ;
               RECT 34.214 66.326 34.266 66.362 ;
               RECT 34.214 67.526 34.266 67.562 ;
               RECT 34.214 68.726 34.266 68.762 ;
               RECT 34.214 69.926 34.266 69.962 ;
               RECT 34.214 71.126 34.266 71.162 ;
               RECT 34.214 72.326 34.266 72.362 ;
               RECT 34.214 73.526 34.266 73.562 ;
               RECT 34.214 74.726 34.266 74.762 ;
               RECT 34.214 75.926 34.266 75.962 ;
               RECT 34.214 77.126 34.266 77.162 ;
               RECT 34.214 78.326 34.266 78.362 ;
               RECT 34.214 79.526 34.266 79.562 ;
               RECT 34.214 80.726 34.266 80.762 ;
               RECT 34.214 81.926 34.266 81.962 ;
               RECT 34.214 83.126 34.266 83.162 ;
               RECT 34.214 84.326 34.266 84.362 ;
               RECT 34.214 85.526 34.266 85.562 ;
               RECT 34.214 86.726 34.266 86.762 ;
               RECT 34.214 87.926 34.266 87.962 ;
               RECT 34.214 89.126 34.266 89.162 ;
               RECT 34.214 90.326 34.266 90.362 ;
               RECT 34.214 91.526 34.266 91.562 ;
               RECT 34.214 92.726 34.266 92.762 ;
               RECT 34.214 93.926 34.266 93.962 ;
               RECT 34.214 95.126 34.266 95.162 ;
               RECT 34.214 96.326 34.266 96.362 ;
               RECT 34.214 97.526 34.266 97.562 ;
               RECT 34.214 98.726 34.266 98.762 ;
               RECT 34.214 99.926 34.266 99.962 ;
               RECT 34.214 101.126 34.266 101.162 ;
               RECT 34.214 102.326 34.266 102.362 ;
               RECT 34.214 103.526 34.266 103.562 ;
               RECT 34.294 1.558 34.346 1.594 ;
               RECT 34.294 2.758 34.346 2.794 ;
               RECT 34.294 3.958 34.346 3.994 ;
               RECT 34.294 5.158 34.346 5.194 ;
               RECT 34.294 6.358 34.346 6.394 ;
               RECT 34.294 7.558 34.346 7.594 ;
               RECT 34.294 8.758 34.346 8.794 ;
               RECT 34.294 9.958 34.346 9.994 ;
               RECT 34.294 11.158 34.346 11.194 ;
               RECT 34.294 12.358 34.346 12.394 ;
               RECT 34.294 13.558 34.346 13.594 ;
               RECT 34.294 14.758 34.346 14.794 ;
               RECT 34.294 15.958 34.346 15.994 ;
               RECT 34.294 17.158 34.346 17.194 ;
               RECT 34.294 18.358 34.346 18.394 ;
               RECT 34.294 19.558 34.346 19.594 ;
               RECT 34.294 20.758 34.346 20.794 ;
               RECT 34.294 21.958 34.346 21.994 ;
               RECT 34.294 23.158 34.346 23.194 ;
               RECT 34.294 24.358 34.346 24.394 ;
               RECT 34.294 25.558 34.346 25.594 ;
               RECT 34.294 26.758 34.346 26.794 ;
               RECT 34.294 27.958 34.346 27.994 ;
               RECT 34.294 29.158 34.346 29.194 ;
               RECT 34.294 30.358 34.346 30.394 ;
               RECT 34.294 31.558 34.346 31.594 ;
               RECT 34.294 32.758 34.346 32.794 ;
               RECT 34.294 33.958 34.346 33.994 ;
               RECT 34.294 35.158 34.346 35.194 ;
               RECT 34.294 36.358 34.346 36.394 ;
               RECT 34.294 37.558 34.346 37.594 ;
               RECT 34.294 38.758 34.346 38.794 ;
               RECT 34.294 39.958 34.346 39.994 ;
               RECT 34.294 41.158 34.346 41.194 ;
               RECT 34.294 42.358 34.346 42.394 ;
               RECT 34.294 43.558 34.346 43.594 ;
               RECT 34.294 44.758 34.346 44.794 ;
               RECT 34.294 45.958 34.346 45.994 ;
               RECT 34.294 47.158 34.346 47.194 ;
               RECT 34.294 48.358 34.346 48.394 ;
               RECT 34.294 50.142 34.346 50.178 ;
               RECT 34.294 50.382 34.346 50.418 ;
               RECT 34.294 54.702 34.346 54.738 ;
               RECT 34.294 54.942 34.346 54.978 ;
               RECT 34.294 57.478 34.346 57.514 ;
               RECT 34.294 58.678 34.346 58.714 ;
               RECT 34.294 59.878 34.346 59.914 ;
               RECT 34.294 61.078 34.346 61.114 ;
               RECT 34.294 62.278 34.346 62.314 ;
               RECT 34.294 63.478 34.346 63.514 ;
               RECT 34.294 64.678 34.346 64.714 ;
               RECT 34.294 65.878 34.346 65.914 ;
               RECT 34.294 67.078 34.346 67.114 ;
               RECT 34.294 68.278 34.346 68.314 ;
               RECT 34.294 69.478 34.346 69.514 ;
               RECT 34.294 70.678 34.346 70.714 ;
               RECT 34.294 71.878 34.346 71.914 ;
               RECT 34.294 73.078 34.346 73.114 ;
               RECT 34.294 74.278 34.346 74.314 ;
               RECT 34.294 75.478 34.346 75.514 ;
               RECT 34.294 76.678 34.346 76.714 ;
               RECT 34.294 77.878 34.346 77.914 ;
               RECT 34.294 79.078 34.346 79.114 ;
               RECT 34.294 80.278 34.346 80.314 ;
               RECT 34.294 81.478 34.346 81.514 ;
               RECT 34.294 82.678 34.346 82.714 ;
               RECT 34.294 83.878 34.346 83.914 ;
               RECT 34.294 85.078 34.346 85.114 ;
               RECT 34.294 86.278 34.346 86.314 ;
               RECT 34.294 87.478 34.346 87.514 ;
               RECT 34.294 88.678 34.346 88.714 ;
               RECT 34.294 89.878 34.346 89.914 ;
               RECT 34.294 91.078 34.346 91.114 ;
               RECT 34.294 92.278 34.346 92.314 ;
               RECT 34.294 93.478 34.346 93.514 ;
               RECT 34.294 94.678 34.346 94.714 ;
               RECT 34.294 95.878 34.346 95.914 ;
               RECT 34.294 97.078 34.346 97.114 ;
               RECT 34.294 98.278 34.346 98.314 ;
               RECT 34.294 99.478 34.346 99.514 ;
               RECT 34.294 100.678 34.346 100.714 ;
               RECT 34.294 101.878 34.346 101.914 ;
               RECT 34.294 103.078 34.346 103.114 ;
               RECT 34.294 104.278 34.346 104.314 ;
               RECT 34.374 0.281 34.426 0.317 ;
               RECT 34.374 104.803 34.426 104.839 ;
               RECT 34.454 0.806 34.506 0.842 ;
               RECT 34.454 2.006 34.506 2.042 ;
               RECT 34.454 3.206 34.506 3.242 ;
               RECT 34.454 4.406 34.506 4.442 ;
               RECT 34.454 5.606 34.506 5.642 ;
               RECT 34.454 6.806 34.506 6.842 ;
               RECT 34.454 8.006 34.506 8.042 ;
               RECT 34.454 9.206 34.506 9.242 ;
               RECT 34.454 10.406 34.506 10.442 ;
               RECT 34.454 11.606 34.506 11.642 ;
               RECT 34.454 12.806 34.506 12.842 ;
               RECT 34.454 14.006 34.506 14.042 ;
               RECT 34.454 15.206 34.506 15.242 ;
               RECT 34.454 16.406 34.506 16.442 ;
               RECT 34.454 17.606 34.506 17.642 ;
               RECT 34.454 18.806 34.506 18.842 ;
               RECT 34.454 20.006 34.506 20.042 ;
               RECT 34.454 21.206 34.506 21.242 ;
               RECT 34.454 22.406 34.506 22.442 ;
               RECT 34.454 23.606 34.506 23.642 ;
               RECT 34.454 24.806 34.506 24.842 ;
               RECT 34.454 26.006 34.506 26.042 ;
               RECT 34.454 27.206 34.506 27.242 ;
               RECT 34.454 28.406 34.506 28.442 ;
               RECT 34.454 29.606 34.506 29.642 ;
               RECT 34.454 30.806 34.506 30.842 ;
               RECT 34.454 32.006 34.506 32.042 ;
               RECT 34.454 33.206 34.506 33.242 ;
               RECT 34.454 34.406 34.506 34.442 ;
               RECT 34.454 35.606 34.506 35.642 ;
               RECT 34.454 36.806 34.506 36.842 ;
               RECT 34.454 38.006 34.506 38.042 ;
               RECT 34.454 39.206 34.506 39.242 ;
               RECT 34.454 40.406 34.506 40.442 ;
               RECT 34.454 41.606 34.506 41.642 ;
               RECT 34.454 42.806 34.506 42.842 ;
               RECT 34.454 44.006 34.506 44.042 ;
               RECT 34.454 45.206 34.506 45.242 ;
               RECT 34.454 46.406 34.506 46.442 ;
               RECT 34.454 47.606 34.506 47.642 ;
               RECT 34.454 49.422 34.506 49.458 ;
               RECT 34.454 49.662 34.506 49.698 ;
               RECT 34.454 51.102 34.506 51.138 ;
               RECT 34.454 51.582 34.506 51.618 ;
               RECT 34.454 53.502 34.506 53.538 ;
               RECT 34.454 53.982 34.506 54.018 ;
               RECT 34.454 55.422 34.506 55.458 ;
               RECT 34.454 55.662 34.506 55.698 ;
               RECT 34.454 56.726 34.506 56.762 ;
               RECT 34.454 57.926 34.506 57.962 ;
               RECT 34.454 59.126 34.506 59.162 ;
               RECT 34.454 60.326 34.506 60.362 ;
               RECT 34.454 61.526 34.506 61.562 ;
               RECT 34.454 62.726 34.506 62.762 ;
               RECT 34.454 63.926 34.506 63.962 ;
               RECT 34.454 65.126 34.506 65.162 ;
               RECT 34.454 66.326 34.506 66.362 ;
               RECT 34.454 67.526 34.506 67.562 ;
               RECT 34.454 68.726 34.506 68.762 ;
               RECT 34.454 69.926 34.506 69.962 ;
               RECT 34.454 71.126 34.506 71.162 ;
               RECT 34.454 72.326 34.506 72.362 ;
               RECT 34.454 73.526 34.506 73.562 ;
               RECT 34.454 74.726 34.506 74.762 ;
               RECT 34.454 75.926 34.506 75.962 ;
               RECT 34.454 77.126 34.506 77.162 ;
               RECT 34.454 78.326 34.506 78.362 ;
               RECT 34.454 79.526 34.506 79.562 ;
               RECT 34.454 80.726 34.506 80.762 ;
               RECT 34.454 81.926 34.506 81.962 ;
               RECT 34.454 83.126 34.506 83.162 ;
               RECT 34.454 84.326 34.506 84.362 ;
               RECT 34.454 85.526 34.506 85.562 ;
               RECT 34.454 86.726 34.506 86.762 ;
               RECT 34.454 87.926 34.506 87.962 ;
               RECT 34.454 89.126 34.506 89.162 ;
               RECT 34.454 90.326 34.506 90.362 ;
               RECT 34.454 91.526 34.506 91.562 ;
               RECT 34.454 92.726 34.506 92.762 ;
               RECT 34.454 93.926 34.506 93.962 ;
               RECT 34.454 95.126 34.506 95.162 ;
               RECT 34.454 96.326 34.506 96.362 ;
               RECT 34.454 97.526 34.506 97.562 ;
               RECT 34.454 98.726 34.506 98.762 ;
               RECT 34.454 99.926 34.506 99.962 ;
               RECT 34.454 101.126 34.506 101.162 ;
               RECT 34.454 102.326 34.506 102.362 ;
               RECT 34.454 103.526 34.506 103.562 ;
               RECT 34.534 1.558 34.586 1.594 ;
               RECT 34.534 2.758 34.586 2.794 ;
               RECT 34.534 3.958 34.586 3.994 ;
               RECT 34.534 5.158 34.586 5.194 ;
               RECT 34.534 6.358 34.586 6.394 ;
               RECT 34.534 7.558 34.586 7.594 ;
               RECT 34.534 8.758 34.586 8.794 ;
               RECT 34.534 9.958 34.586 9.994 ;
               RECT 34.534 11.158 34.586 11.194 ;
               RECT 34.534 12.358 34.586 12.394 ;
               RECT 34.534 13.558 34.586 13.594 ;
               RECT 34.534 14.758 34.586 14.794 ;
               RECT 34.534 15.958 34.586 15.994 ;
               RECT 34.534 17.158 34.586 17.194 ;
               RECT 34.534 18.358 34.586 18.394 ;
               RECT 34.534 19.558 34.586 19.594 ;
               RECT 34.534 20.758 34.586 20.794 ;
               RECT 34.534 21.958 34.586 21.994 ;
               RECT 34.534 23.158 34.586 23.194 ;
               RECT 34.534 24.358 34.586 24.394 ;
               RECT 34.534 25.558 34.586 25.594 ;
               RECT 34.534 26.758 34.586 26.794 ;
               RECT 34.534 27.958 34.586 27.994 ;
               RECT 34.534 29.158 34.586 29.194 ;
               RECT 34.534 30.358 34.586 30.394 ;
               RECT 34.534 31.558 34.586 31.594 ;
               RECT 34.534 32.758 34.586 32.794 ;
               RECT 34.534 33.958 34.586 33.994 ;
               RECT 34.534 35.158 34.586 35.194 ;
               RECT 34.534 36.358 34.586 36.394 ;
               RECT 34.534 37.558 34.586 37.594 ;
               RECT 34.534 38.758 34.586 38.794 ;
               RECT 34.534 39.958 34.586 39.994 ;
               RECT 34.534 41.158 34.586 41.194 ;
               RECT 34.534 42.358 34.586 42.394 ;
               RECT 34.534 43.558 34.586 43.594 ;
               RECT 34.534 44.758 34.586 44.794 ;
               RECT 34.534 45.958 34.586 45.994 ;
               RECT 34.534 47.158 34.586 47.194 ;
               RECT 34.534 48.358 34.586 48.394 ;
               RECT 34.534 50.142 34.586 50.178 ;
               RECT 34.534 50.382 34.586 50.418 ;
               RECT 34.534 54.702 34.586 54.738 ;
               RECT 34.534 54.942 34.586 54.978 ;
               RECT 34.534 57.478 34.586 57.514 ;
               RECT 34.534 58.678 34.586 58.714 ;
               RECT 34.534 59.878 34.586 59.914 ;
               RECT 34.534 61.078 34.586 61.114 ;
               RECT 34.534 62.278 34.586 62.314 ;
               RECT 34.534 63.478 34.586 63.514 ;
               RECT 34.534 64.678 34.586 64.714 ;
               RECT 34.534 65.878 34.586 65.914 ;
               RECT 34.534 67.078 34.586 67.114 ;
               RECT 34.534 68.278 34.586 68.314 ;
               RECT 34.534 69.478 34.586 69.514 ;
               RECT 34.534 70.678 34.586 70.714 ;
               RECT 34.534 71.878 34.586 71.914 ;
               RECT 34.534 73.078 34.586 73.114 ;
               RECT 34.534 74.278 34.586 74.314 ;
               RECT 34.534 75.478 34.586 75.514 ;
               RECT 34.534 76.678 34.586 76.714 ;
               RECT 34.534 77.878 34.586 77.914 ;
               RECT 34.534 79.078 34.586 79.114 ;
               RECT 34.534 80.278 34.586 80.314 ;
               RECT 34.534 81.478 34.586 81.514 ;
               RECT 34.534 82.678 34.586 82.714 ;
               RECT 34.534 83.878 34.586 83.914 ;
               RECT 34.534 85.078 34.586 85.114 ;
               RECT 34.534 86.278 34.586 86.314 ;
               RECT 34.534 87.478 34.586 87.514 ;
               RECT 34.534 88.678 34.586 88.714 ;
               RECT 34.534 89.878 34.586 89.914 ;
               RECT 34.534 91.078 34.586 91.114 ;
               RECT 34.534 92.278 34.586 92.314 ;
               RECT 34.534 93.478 34.586 93.514 ;
               RECT 34.534 94.678 34.586 94.714 ;
               RECT 34.534 95.878 34.586 95.914 ;
               RECT 34.534 97.078 34.586 97.114 ;
               RECT 34.534 98.278 34.586 98.314 ;
               RECT 34.534 99.478 34.586 99.514 ;
               RECT 34.534 100.678 34.586 100.714 ;
               RECT 34.534 101.878 34.586 101.914 ;
               RECT 34.534 103.078 34.586 103.114 ;
               RECT 34.534 104.278 34.586 104.314 ;
               RECT 34.614 0.806 34.666 0.842 ;
               RECT 34.614 2.006 34.666 2.042 ;
               RECT 34.614 3.206 34.666 3.242 ;
               RECT 34.614 4.406 34.666 4.442 ;
               RECT 34.614 5.606 34.666 5.642 ;
               RECT 34.614 6.806 34.666 6.842 ;
               RECT 34.614 8.006 34.666 8.042 ;
               RECT 34.614 9.206 34.666 9.242 ;
               RECT 34.614 10.406 34.666 10.442 ;
               RECT 34.614 11.606 34.666 11.642 ;
               RECT 34.614 12.806 34.666 12.842 ;
               RECT 34.614 14.006 34.666 14.042 ;
               RECT 34.614 15.206 34.666 15.242 ;
               RECT 34.614 16.406 34.666 16.442 ;
               RECT 34.614 17.606 34.666 17.642 ;
               RECT 34.614 18.806 34.666 18.842 ;
               RECT 34.614 20.006 34.666 20.042 ;
               RECT 34.614 21.206 34.666 21.242 ;
               RECT 34.614 22.406 34.666 22.442 ;
               RECT 34.614 23.606 34.666 23.642 ;
               RECT 34.614 24.806 34.666 24.842 ;
               RECT 34.614 26.006 34.666 26.042 ;
               RECT 34.614 27.206 34.666 27.242 ;
               RECT 34.614 28.406 34.666 28.442 ;
               RECT 34.614 29.606 34.666 29.642 ;
               RECT 34.614 30.806 34.666 30.842 ;
               RECT 34.614 32.006 34.666 32.042 ;
               RECT 34.614 33.206 34.666 33.242 ;
               RECT 34.614 34.406 34.666 34.442 ;
               RECT 34.614 35.606 34.666 35.642 ;
               RECT 34.614 36.806 34.666 36.842 ;
               RECT 34.614 38.006 34.666 38.042 ;
               RECT 34.614 39.206 34.666 39.242 ;
               RECT 34.614 40.406 34.666 40.442 ;
               RECT 34.614 41.606 34.666 41.642 ;
               RECT 34.614 42.806 34.666 42.842 ;
               RECT 34.614 44.006 34.666 44.042 ;
               RECT 34.614 45.206 34.666 45.242 ;
               RECT 34.614 46.406 34.666 46.442 ;
               RECT 34.614 47.606 34.666 47.642 ;
               RECT 34.614 49.422 34.666 49.458 ;
               RECT 34.614 49.662 34.666 49.698 ;
               RECT 34.614 55.422 34.666 55.458 ;
               RECT 34.614 55.662 34.666 55.698 ;
               RECT 34.614 56.726 34.666 56.762 ;
               RECT 34.614 57.926 34.666 57.962 ;
               RECT 34.614 59.126 34.666 59.162 ;
               RECT 34.614 60.326 34.666 60.362 ;
               RECT 34.614 61.526 34.666 61.562 ;
               RECT 34.614 62.726 34.666 62.762 ;
               RECT 34.614 63.926 34.666 63.962 ;
               RECT 34.614 65.126 34.666 65.162 ;
               RECT 34.614 66.326 34.666 66.362 ;
               RECT 34.614 67.526 34.666 67.562 ;
               RECT 34.614 68.726 34.666 68.762 ;
               RECT 34.614 69.926 34.666 69.962 ;
               RECT 34.614 71.126 34.666 71.162 ;
               RECT 34.614 72.326 34.666 72.362 ;
               RECT 34.614 73.526 34.666 73.562 ;
               RECT 34.614 74.726 34.666 74.762 ;
               RECT 34.614 75.926 34.666 75.962 ;
               RECT 34.614 77.126 34.666 77.162 ;
               RECT 34.614 78.326 34.666 78.362 ;
               RECT 34.614 79.526 34.666 79.562 ;
               RECT 34.614 80.726 34.666 80.762 ;
               RECT 34.614 81.926 34.666 81.962 ;
               RECT 34.614 83.126 34.666 83.162 ;
               RECT 34.614 84.326 34.666 84.362 ;
               RECT 34.614 85.526 34.666 85.562 ;
               RECT 34.614 86.726 34.666 86.762 ;
               RECT 34.614 87.926 34.666 87.962 ;
               RECT 34.614 89.126 34.666 89.162 ;
               RECT 34.614 90.326 34.666 90.362 ;
               RECT 34.614 91.526 34.666 91.562 ;
               RECT 34.614 92.726 34.666 92.762 ;
               RECT 34.614 93.926 34.666 93.962 ;
               RECT 34.614 95.126 34.666 95.162 ;
               RECT 34.614 96.326 34.666 96.362 ;
               RECT 34.614 97.526 34.666 97.562 ;
               RECT 34.614 98.726 34.666 98.762 ;
               RECT 34.614 99.926 34.666 99.962 ;
               RECT 34.614 101.126 34.666 101.162 ;
               RECT 34.614 102.326 34.666 102.362 ;
               RECT 34.614 103.526 34.666 103.562 ;
               RECT 34.694 1.558 34.746 1.594 ;
               RECT 34.694 2.758 34.746 2.794 ;
               RECT 34.694 3.958 34.746 3.994 ;
               RECT 34.694 5.158 34.746 5.194 ;
               RECT 34.694 6.358 34.746 6.394 ;
               RECT 34.694 7.558 34.746 7.594 ;
               RECT 34.694 8.758 34.746 8.794 ;
               RECT 34.694 9.958 34.746 9.994 ;
               RECT 34.694 11.158 34.746 11.194 ;
               RECT 34.694 12.358 34.746 12.394 ;
               RECT 34.694 13.558 34.746 13.594 ;
               RECT 34.694 14.758 34.746 14.794 ;
               RECT 34.694 15.958 34.746 15.994 ;
               RECT 34.694 17.158 34.746 17.194 ;
               RECT 34.694 18.358 34.746 18.394 ;
               RECT 34.694 19.558 34.746 19.594 ;
               RECT 34.694 20.758 34.746 20.794 ;
               RECT 34.694 21.958 34.746 21.994 ;
               RECT 34.694 23.158 34.746 23.194 ;
               RECT 34.694 24.358 34.746 24.394 ;
               RECT 34.694 25.558 34.746 25.594 ;
               RECT 34.694 26.758 34.746 26.794 ;
               RECT 34.694 27.958 34.746 27.994 ;
               RECT 34.694 29.158 34.746 29.194 ;
               RECT 34.694 30.358 34.746 30.394 ;
               RECT 34.694 31.558 34.746 31.594 ;
               RECT 34.694 32.758 34.746 32.794 ;
               RECT 34.694 33.958 34.746 33.994 ;
               RECT 34.694 35.158 34.746 35.194 ;
               RECT 34.694 36.358 34.746 36.394 ;
               RECT 34.694 37.558 34.746 37.594 ;
               RECT 34.694 38.758 34.746 38.794 ;
               RECT 34.694 39.958 34.746 39.994 ;
               RECT 34.694 41.158 34.746 41.194 ;
               RECT 34.694 42.358 34.746 42.394 ;
               RECT 34.694 43.558 34.746 43.594 ;
               RECT 34.694 44.758 34.746 44.794 ;
               RECT 34.694 45.958 34.746 45.994 ;
               RECT 34.694 47.158 34.746 47.194 ;
               RECT 34.694 48.358 34.746 48.394 ;
               RECT 34.694 50.142 34.746 50.178 ;
               RECT 34.694 50.382 34.746 50.418 ;
               RECT 34.694 54.702 34.746 54.738 ;
               RECT 34.694 54.942 34.746 54.978 ;
               RECT 34.694 57.478 34.746 57.514 ;
               RECT 34.694 58.678 34.746 58.714 ;
               RECT 34.694 59.878 34.746 59.914 ;
               RECT 34.694 61.078 34.746 61.114 ;
               RECT 34.694 62.278 34.746 62.314 ;
               RECT 34.694 63.478 34.746 63.514 ;
               RECT 34.694 64.678 34.746 64.714 ;
               RECT 34.694 65.878 34.746 65.914 ;
               RECT 34.694 67.078 34.746 67.114 ;
               RECT 34.694 68.278 34.746 68.314 ;
               RECT 34.694 69.478 34.746 69.514 ;
               RECT 34.694 70.678 34.746 70.714 ;
               RECT 34.694 71.878 34.746 71.914 ;
               RECT 34.694 73.078 34.746 73.114 ;
               RECT 34.694 74.278 34.746 74.314 ;
               RECT 34.694 75.478 34.746 75.514 ;
               RECT 34.694 76.678 34.746 76.714 ;
               RECT 34.694 77.878 34.746 77.914 ;
               RECT 34.694 79.078 34.746 79.114 ;
               RECT 34.694 80.278 34.746 80.314 ;
               RECT 34.694 81.478 34.746 81.514 ;
               RECT 34.694 82.678 34.746 82.714 ;
               RECT 34.694 83.878 34.746 83.914 ;
               RECT 34.694 85.078 34.746 85.114 ;
               RECT 34.694 86.278 34.746 86.314 ;
               RECT 34.694 87.478 34.746 87.514 ;
               RECT 34.694 88.678 34.746 88.714 ;
               RECT 34.694 89.878 34.746 89.914 ;
               RECT 34.694 91.078 34.746 91.114 ;
               RECT 34.694 92.278 34.746 92.314 ;
               RECT 34.694 93.478 34.746 93.514 ;
               RECT 34.694 94.678 34.746 94.714 ;
               RECT 34.694 95.878 34.746 95.914 ;
               RECT 34.694 97.078 34.746 97.114 ;
               RECT 34.694 98.278 34.746 98.314 ;
               RECT 34.694 99.478 34.746 99.514 ;
               RECT 34.694 100.678 34.746 100.714 ;
               RECT 34.694 101.878 34.746 101.914 ;
               RECT 34.694 103.078 34.746 103.114 ;
               RECT 34.694 104.278 34.746 104.314 ;
               RECT 34.774 0.281 34.826 0.317 ;
               RECT 34.774 104.803 34.826 104.839 ;
               RECT 34.854 0.806 34.906 0.842 ;
               RECT 34.854 2.006 34.906 2.042 ;
               RECT 34.854 3.206 34.906 3.242 ;
               RECT 34.854 4.406 34.906 4.442 ;
               RECT 34.854 5.606 34.906 5.642 ;
               RECT 34.854 6.806 34.906 6.842 ;
               RECT 34.854 8.006 34.906 8.042 ;
               RECT 34.854 9.206 34.906 9.242 ;
               RECT 34.854 10.406 34.906 10.442 ;
               RECT 34.854 11.606 34.906 11.642 ;
               RECT 34.854 12.806 34.906 12.842 ;
               RECT 34.854 14.006 34.906 14.042 ;
               RECT 34.854 15.206 34.906 15.242 ;
               RECT 34.854 16.406 34.906 16.442 ;
               RECT 34.854 17.606 34.906 17.642 ;
               RECT 34.854 18.806 34.906 18.842 ;
               RECT 34.854 20.006 34.906 20.042 ;
               RECT 34.854 21.206 34.906 21.242 ;
               RECT 34.854 22.406 34.906 22.442 ;
               RECT 34.854 23.606 34.906 23.642 ;
               RECT 34.854 24.806 34.906 24.842 ;
               RECT 34.854 26.006 34.906 26.042 ;
               RECT 34.854 27.206 34.906 27.242 ;
               RECT 34.854 28.406 34.906 28.442 ;
               RECT 34.854 29.606 34.906 29.642 ;
               RECT 34.854 30.806 34.906 30.842 ;
               RECT 34.854 32.006 34.906 32.042 ;
               RECT 34.854 33.206 34.906 33.242 ;
               RECT 34.854 34.406 34.906 34.442 ;
               RECT 34.854 35.606 34.906 35.642 ;
               RECT 34.854 36.806 34.906 36.842 ;
               RECT 34.854 38.006 34.906 38.042 ;
               RECT 34.854 39.206 34.906 39.242 ;
               RECT 34.854 40.406 34.906 40.442 ;
               RECT 34.854 41.606 34.906 41.642 ;
               RECT 34.854 42.806 34.906 42.842 ;
               RECT 34.854 44.006 34.906 44.042 ;
               RECT 34.854 45.206 34.906 45.242 ;
               RECT 34.854 46.406 34.906 46.442 ;
               RECT 34.854 47.606 34.906 47.642 ;
               RECT 34.854 49.422 34.906 49.458 ;
               RECT 34.854 49.662 34.906 49.698 ;
               RECT 34.854 55.422 34.906 55.458 ;
               RECT 34.854 55.662 34.906 55.698 ;
               RECT 34.854 56.726 34.906 56.762 ;
               RECT 34.854 57.926 34.906 57.962 ;
               RECT 34.854 59.126 34.906 59.162 ;
               RECT 34.854 60.326 34.906 60.362 ;
               RECT 34.854 61.526 34.906 61.562 ;
               RECT 34.854 62.726 34.906 62.762 ;
               RECT 34.854 63.926 34.906 63.962 ;
               RECT 34.854 65.126 34.906 65.162 ;
               RECT 34.854 66.326 34.906 66.362 ;
               RECT 34.854 67.526 34.906 67.562 ;
               RECT 34.854 68.726 34.906 68.762 ;
               RECT 34.854 69.926 34.906 69.962 ;
               RECT 34.854 71.126 34.906 71.162 ;
               RECT 34.854 72.326 34.906 72.362 ;
               RECT 34.854 73.526 34.906 73.562 ;
               RECT 34.854 74.726 34.906 74.762 ;
               RECT 34.854 75.926 34.906 75.962 ;
               RECT 34.854 77.126 34.906 77.162 ;
               RECT 34.854 78.326 34.906 78.362 ;
               RECT 34.854 79.526 34.906 79.562 ;
               RECT 34.854 80.726 34.906 80.762 ;
               RECT 34.854 81.926 34.906 81.962 ;
               RECT 34.854 83.126 34.906 83.162 ;
               RECT 34.854 84.326 34.906 84.362 ;
               RECT 34.854 85.526 34.906 85.562 ;
               RECT 34.854 86.726 34.906 86.762 ;
               RECT 34.854 87.926 34.906 87.962 ;
               RECT 34.854 89.126 34.906 89.162 ;
               RECT 34.854 90.326 34.906 90.362 ;
               RECT 34.854 91.526 34.906 91.562 ;
               RECT 34.854 92.726 34.906 92.762 ;
               RECT 34.854 93.926 34.906 93.962 ;
               RECT 34.854 95.126 34.906 95.162 ;
               RECT 34.854 96.326 34.906 96.362 ;
               RECT 34.854 97.526 34.906 97.562 ;
               RECT 34.854 98.726 34.906 98.762 ;
               RECT 34.854 99.926 34.906 99.962 ;
               RECT 34.854 101.126 34.906 101.162 ;
               RECT 34.854 102.326 34.906 102.362 ;
               RECT 34.854 103.526 34.906 103.562 ;
               RECT 34.934 1.558 34.986 1.594 ;
               RECT 34.934 2.758 34.986 2.794 ;
               RECT 34.934 3.958 34.986 3.994 ;
               RECT 34.934 5.158 34.986 5.194 ;
               RECT 34.934 6.358 34.986 6.394 ;
               RECT 34.934 7.558 34.986 7.594 ;
               RECT 34.934 8.758 34.986 8.794 ;
               RECT 34.934 9.958 34.986 9.994 ;
               RECT 34.934 11.158 34.986 11.194 ;
               RECT 34.934 12.358 34.986 12.394 ;
               RECT 34.934 13.558 34.986 13.594 ;
               RECT 34.934 14.758 34.986 14.794 ;
               RECT 34.934 15.958 34.986 15.994 ;
               RECT 34.934 17.158 34.986 17.194 ;
               RECT 34.934 18.358 34.986 18.394 ;
               RECT 34.934 19.558 34.986 19.594 ;
               RECT 34.934 20.758 34.986 20.794 ;
               RECT 34.934 21.958 34.986 21.994 ;
               RECT 34.934 23.158 34.986 23.194 ;
               RECT 34.934 24.358 34.986 24.394 ;
               RECT 34.934 25.558 34.986 25.594 ;
               RECT 34.934 26.758 34.986 26.794 ;
               RECT 34.934 27.958 34.986 27.994 ;
               RECT 34.934 29.158 34.986 29.194 ;
               RECT 34.934 30.358 34.986 30.394 ;
               RECT 34.934 31.558 34.986 31.594 ;
               RECT 34.934 32.758 34.986 32.794 ;
               RECT 34.934 33.958 34.986 33.994 ;
               RECT 34.934 35.158 34.986 35.194 ;
               RECT 34.934 36.358 34.986 36.394 ;
               RECT 34.934 37.558 34.986 37.594 ;
               RECT 34.934 38.758 34.986 38.794 ;
               RECT 34.934 39.958 34.986 39.994 ;
               RECT 34.934 41.158 34.986 41.194 ;
               RECT 34.934 42.358 34.986 42.394 ;
               RECT 34.934 43.558 34.986 43.594 ;
               RECT 34.934 44.758 34.986 44.794 ;
               RECT 34.934 45.958 34.986 45.994 ;
               RECT 34.934 47.158 34.986 47.194 ;
               RECT 34.934 48.358 34.986 48.394 ;
               RECT 34.934 50.142 34.986 50.178 ;
               RECT 34.934 50.382 34.986 50.418 ;
               RECT 34.934 54.702 34.986 54.738 ;
               RECT 34.934 54.942 34.986 54.978 ;
               RECT 34.934 57.478 34.986 57.514 ;
               RECT 34.934 58.678 34.986 58.714 ;
               RECT 34.934 59.878 34.986 59.914 ;
               RECT 34.934 61.078 34.986 61.114 ;
               RECT 34.934 62.278 34.986 62.314 ;
               RECT 34.934 63.478 34.986 63.514 ;
               RECT 34.934 64.678 34.986 64.714 ;
               RECT 34.934 65.878 34.986 65.914 ;
               RECT 34.934 67.078 34.986 67.114 ;
               RECT 34.934 68.278 34.986 68.314 ;
               RECT 34.934 69.478 34.986 69.514 ;
               RECT 34.934 70.678 34.986 70.714 ;
               RECT 34.934 71.878 34.986 71.914 ;
               RECT 34.934 73.078 34.986 73.114 ;
               RECT 34.934 74.278 34.986 74.314 ;
               RECT 34.934 75.478 34.986 75.514 ;
               RECT 34.934 76.678 34.986 76.714 ;
               RECT 34.934 77.878 34.986 77.914 ;
               RECT 34.934 79.078 34.986 79.114 ;
               RECT 34.934 80.278 34.986 80.314 ;
               RECT 34.934 81.478 34.986 81.514 ;
               RECT 34.934 82.678 34.986 82.714 ;
               RECT 34.934 83.878 34.986 83.914 ;
               RECT 34.934 85.078 34.986 85.114 ;
               RECT 34.934 86.278 34.986 86.314 ;
               RECT 34.934 87.478 34.986 87.514 ;
               RECT 34.934 88.678 34.986 88.714 ;
               RECT 34.934 89.878 34.986 89.914 ;
               RECT 34.934 91.078 34.986 91.114 ;
               RECT 34.934 92.278 34.986 92.314 ;
               RECT 34.934 93.478 34.986 93.514 ;
               RECT 34.934 94.678 34.986 94.714 ;
               RECT 34.934 95.878 34.986 95.914 ;
               RECT 34.934 97.078 34.986 97.114 ;
               RECT 34.934 98.278 34.986 98.314 ;
               RECT 34.934 99.478 34.986 99.514 ;
               RECT 34.934 100.678 34.986 100.714 ;
               RECT 34.934 101.878 34.986 101.914 ;
               RECT 34.934 103.078 34.986 103.114 ;
               RECT 34.934 104.278 34.986 104.314 ;
               RECT 35.014 0.806 35.066 0.842 ;
               RECT 35.014 2.006 35.066 2.042 ;
               RECT 35.014 3.206 35.066 3.242 ;
               RECT 35.014 4.406 35.066 4.442 ;
               RECT 35.014 5.606 35.066 5.642 ;
               RECT 35.014 6.806 35.066 6.842 ;
               RECT 35.014 8.006 35.066 8.042 ;
               RECT 35.014 9.206 35.066 9.242 ;
               RECT 35.014 10.406 35.066 10.442 ;
               RECT 35.014 11.606 35.066 11.642 ;
               RECT 35.014 12.806 35.066 12.842 ;
               RECT 35.014 14.006 35.066 14.042 ;
               RECT 35.014 15.206 35.066 15.242 ;
               RECT 35.014 16.406 35.066 16.442 ;
               RECT 35.014 17.606 35.066 17.642 ;
               RECT 35.014 18.806 35.066 18.842 ;
               RECT 35.014 20.006 35.066 20.042 ;
               RECT 35.014 21.206 35.066 21.242 ;
               RECT 35.014 22.406 35.066 22.442 ;
               RECT 35.014 23.606 35.066 23.642 ;
               RECT 35.014 24.806 35.066 24.842 ;
               RECT 35.014 26.006 35.066 26.042 ;
               RECT 35.014 27.206 35.066 27.242 ;
               RECT 35.014 28.406 35.066 28.442 ;
               RECT 35.014 29.606 35.066 29.642 ;
               RECT 35.014 30.806 35.066 30.842 ;
               RECT 35.014 32.006 35.066 32.042 ;
               RECT 35.014 33.206 35.066 33.242 ;
               RECT 35.014 34.406 35.066 34.442 ;
               RECT 35.014 35.606 35.066 35.642 ;
               RECT 35.014 36.806 35.066 36.842 ;
               RECT 35.014 38.006 35.066 38.042 ;
               RECT 35.014 39.206 35.066 39.242 ;
               RECT 35.014 40.406 35.066 40.442 ;
               RECT 35.014 41.606 35.066 41.642 ;
               RECT 35.014 42.806 35.066 42.842 ;
               RECT 35.014 44.006 35.066 44.042 ;
               RECT 35.014 45.206 35.066 45.242 ;
               RECT 35.014 46.406 35.066 46.442 ;
               RECT 35.014 47.606 35.066 47.642 ;
               RECT 35.014 49.422 35.066 49.458 ;
               RECT 35.014 49.662 35.066 49.698 ;
               RECT 35.014 55.422 35.066 55.458 ;
               RECT 35.014 55.662 35.066 55.698 ;
               RECT 35.014 56.726 35.066 56.762 ;
               RECT 35.014 57.926 35.066 57.962 ;
               RECT 35.014 59.126 35.066 59.162 ;
               RECT 35.014 60.326 35.066 60.362 ;
               RECT 35.014 61.526 35.066 61.562 ;
               RECT 35.014 62.726 35.066 62.762 ;
               RECT 35.014 63.926 35.066 63.962 ;
               RECT 35.014 65.126 35.066 65.162 ;
               RECT 35.014 66.326 35.066 66.362 ;
               RECT 35.014 67.526 35.066 67.562 ;
               RECT 35.014 68.726 35.066 68.762 ;
               RECT 35.014 69.926 35.066 69.962 ;
               RECT 35.014 71.126 35.066 71.162 ;
               RECT 35.014 72.326 35.066 72.362 ;
               RECT 35.014 73.526 35.066 73.562 ;
               RECT 35.014 74.726 35.066 74.762 ;
               RECT 35.014 75.926 35.066 75.962 ;
               RECT 35.014 77.126 35.066 77.162 ;
               RECT 35.014 78.326 35.066 78.362 ;
               RECT 35.014 79.526 35.066 79.562 ;
               RECT 35.014 80.726 35.066 80.762 ;
               RECT 35.014 81.926 35.066 81.962 ;
               RECT 35.014 83.126 35.066 83.162 ;
               RECT 35.014 84.326 35.066 84.362 ;
               RECT 35.014 85.526 35.066 85.562 ;
               RECT 35.014 86.726 35.066 86.762 ;
               RECT 35.014 87.926 35.066 87.962 ;
               RECT 35.014 89.126 35.066 89.162 ;
               RECT 35.014 90.326 35.066 90.362 ;
               RECT 35.014 91.526 35.066 91.562 ;
               RECT 35.014 92.726 35.066 92.762 ;
               RECT 35.014 93.926 35.066 93.962 ;
               RECT 35.014 95.126 35.066 95.162 ;
               RECT 35.014 96.326 35.066 96.362 ;
               RECT 35.014 97.526 35.066 97.562 ;
               RECT 35.014 98.726 35.066 98.762 ;
               RECT 35.014 99.926 35.066 99.962 ;
               RECT 35.014 101.126 35.066 101.162 ;
               RECT 35.014 102.326 35.066 102.362 ;
               RECT 35.014 103.526 35.066 103.562 ;
               RECT 35.094 1.558 35.146 1.594 ;
               RECT 35.094 2.758 35.146 2.794 ;
               RECT 35.094 3.958 35.146 3.994 ;
               RECT 35.094 5.158 35.146 5.194 ;
               RECT 35.094 6.358 35.146 6.394 ;
               RECT 35.094 7.558 35.146 7.594 ;
               RECT 35.094 8.758 35.146 8.794 ;
               RECT 35.094 9.958 35.146 9.994 ;
               RECT 35.094 11.158 35.146 11.194 ;
               RECT 35.094 12.358 35.146 12.394 ;
               RECT 35.094 13.558 35.146 13.594 ;
               RECT 35.094 14.758 35.146 14.794 ;
               RECT 35.094 15.958 35.146 15.994 ;
               RECT 35.094 17.158 35.146 17.194 ;
               RECT 35.094 18.358 35.146 18.394 ;
               RECT 35.094 19.558 35.146 19.594 ;
               RECT 35.094 20.758 35.146 20.794 ;
               RECT 35.094 21.958 35.146 21.994 ;
               RECT 35.094 23.158 35.146 23.194 ;
               RECT 35.094 24.358 35.146 24.394 ;
               RECT 35.094 25.558 35.146 25.594 ;
               RECT 35.094 26.758 35.146 26.794 ;
               RECT 35.094 27.958 35.146 27.994 ;
               RECT 35.094 29.158 35.146 29.194 ;
               RECT 35.094 30.358 35.146 30.394 ;
               RECT 35.094 31.558 35.146 31.594 ;
               RECT 35.094 32.758 35.146 32.794 ;
               RECT 35.094 33.958 35.146 33.994 ;
               RECT 35.094 35.158 35.146 35.194 ;
               RECT 35.094 36.358 35.146 36.394 ;
               RECT 35.094 37.558 35.146 37.594 ;
               RECT 35.094 38.758 35.146 38.794 ;
               RECT 35.094 39.958 35.146 39.994 ;
               RECT 35.094 41.158 35.146 41.194 ;
               RECT 35.094 42.358 35.146 42.394 ;
               RECT 35.094 43.558 35.146 43.594 ;
               RECT 35.094 44.758 35.146 44.794 ;
               RECT 35.094 45.958 35.146 45.994 ;
               RECT 35.094 47.158 35.146 47.194 ;
               RECT 35.094 48.358 35.146 48.394 ;
               RECT 35.094 50.142 35.146 50.178 ;
               RECT 35.094 50.382 35.146 50.418 ;
               RECT 35.094 54.702 35.146 54.738 ;
               RECT 35.094 54.942 35.146 54.978 ;
               RECT 35.094 57.478 35.146 57.514 ;
               RECT 35.094 58.678 35.146 58.714 ;
               RECT 35.094 59.878 35.146 59.914 ;
               RECT 35.094 61.078 35.146 61.114 ;
               RECT 35.094 62.278 35.146 62.314 ;
               RECT 35.094 63.478 35.146 63.514 ;
               RECT 35.094 64.678 35.146 64.714 ;
               RECT 35.094 65.878 35.146 65.914 ;
               RECT 35.094 67.078 35.146 67.114 ;
               RECT 35.094 68.278 35.146 68.314 ;
               RECT 35.094 69.478 35.146 69.514 ;
               RECT 35.094 70.678 35.146 70.714 ;
               RECT 35.094 71.878 35.146 71.914 ;
               RECT 35.094 73.078 35.146 73.114 ;
               RECT 35.094 74.278 35.146 74.314 ;
               RECT 35.094 75.478 35.146 75.514 ;
               RECT 35.094 76.678 35.146 76.714 ;
               RECT 35.094 77.878 35.146 77.914 ;
               RECT 35.094 79.078 35.146 79.114 ;
               RECT 35.094 80.278 35.146 80.314 ;
               RECT 35.094 81.478 35.146 81.514 ;
               RECT 35.094 82.678 35.146 82.714 ;
               RECT 35.094 83.878 35.146 83.914 ;
               RECT 35.094 85.078 35.146 85.114 ;
               RECT 35.094 86.278 35.146 86.314 ;
               RECT 35.094 87.478 35.146 87.514 ;
               RECT 35.094 88.678 35.146 88.714 ;
               RECT 35.094 89.878 35.146 89.914 ;
               RECT 35.094 91.078 35.146 91.114 ;
               RECT 35.094 92.278 35.146 92.314 ;
               RECT 35.094 93.478 35.146 93.514 ;
               RECT 35.094 94.678 35.146 94.714 ;
               RECT 35.094 95.878 35.146 95.914 ;
               RECT 35.094 97.078 35.146 97.114 ;
               RECT 35.094 98.278 35.146 98.314 ;
               RECT 35.094 99.478 35.146 99.514 ;
               RECT 35.094 100.678 35.146 100.714 ;
               RECT 35.094 101.878 35.146 101.914 ;
               RECT 35.094 103.078 35.146 103.114 ;
               RECT 35.094 104.278 35.146 104.314 ;
               RECT 35.174 0.281 35.226 0.317 ;
               RECT 35.174 104.803 35.226 104.839 ;
               RECT 35.254 0.806 35.306 0.842 ;
               RECT 35.254 2.006 35.306 2.042 ;
               RECT 35.254 3.206 35.306 3.242 ;
               RECT 35.254 4.406 35.306 4.442 ;
               RECT 35.254 5.606 35.306 5.642 ;
               RECT 35.254 6.806 35.306 6.842 ;
               RECT 35.254 8.006 35.306 8.042 ;
               RECT 35.254 9.206 35.306 9.242 ;
               RECT 35.254 10.406 35.306 10.442 ;
               RECT 35.254 11.606 35.306 11.642 ;
               RECT 35.254 12.806 35.306 12.842 ;
               RECT 35.254 14.006 35.306 14.042 ;
               RECT 35.254 15.206 35.306 15.242 ;
               RECT 35.254 16.406 35.306 16.442 ;
               RECT 35.254 17.606 35.306 17.642 ;
               RECT 35.254 18.806 35.306 18.842 ;
               RECT 35.254 20.006 35.306 20.042 ;
               RECT 35.254 21.206 35.306 21.242 ;
               RECT 35.254 22.406 35.306 22.442 ;
               RECT 35.254 23.606 35.306 23.642 ;
               RECT 35.254 24.806 35.306 24.842 ;
               RECT 35.254 26.006 35.306 26.042 ;
               RECT 35.254 27.206 35.306 27.242 ;
               RECT 35.254 28.406 35.306 28.442 ;
               RECT 35.254 29.606 35.306 29.642 ;
               RECT 35.254 30.806 35.306 30.842 ;
               RECT 35.254 32.006 35.306 32.042 ;
               RECT 35.254 33.206 35.306 33.242 ;
               RECT 35.254 34.406 35.306 34.442 ;
               RECT 35.254 35.606 35.306 35.642 ;
               RECT 35.254 36.806 35.306 36.842 ;
               RECT 35.254 38.006 35.306 38.042 ;
               RECT 35.254 39.206 35.306 39.242 ;
               RECT 35.254 40.406 35.306 40.442 ;
               RECT 35.254 41.606 35.306 41.642 ;
               RECT 35.254 42.806 35.306 42.842 ;
               RECT 35.254 44.006 35.306 44.042 ;
               RECT 35.254 45.206 35.306 45.242 ;
               RECT 35.254 46.406 35.306 46.442 ;
               RECT 35.254 47.606 35.306 47.642 ;
               RECT 35.254 49.422 35.306 49.458 ;
               RECT 35.254 49.662 35.306 49.698 ;
               RECT 35.254 51.102 35.306 51.138 ;
               RECT 35.254 51.582 35.306 51.618 ;
               RECT 35.254 53.502 35.306 53.538 ;
               RECT 35.254 53.982 35.306 54.018 ;
               RECT 35.254 55.422 35.306 55.458 ;
               RECT 35.254 55.662 35.306 55.698 ;
               RECT 35.254 56.726 35.306 56.762 ;
               RECT 35.254 57.926 35.306 57.962 ;
               RECT 35.254 59.126 35.306 59.162 ;
               RECT 35.254 60.326 35.306 60.362 ;
               RECT 35.254 61.526 35.306 61.562 ;
               RECT 35.254 62.726 35.306 62.762 ;
               RECT 35.254 63.926 35.306 63.962 ;
               RECT 35.254 65.126 35.306 65.162 ;
               RECT 35.254 66.326 35.306 66.362 ;
               RECT 35.254 67.526 35.306 67.562 ;
               RECT 35.254 68.726 35.306 68.762 ;
               RECT 35.254 69.926 35.306 69.962 ;
               RECT 35.254 71.126 35.306 71.162 ;
               RECT 35.254 72.326 35.306 72.362 ;
               RECT 35.254 73.526 35.306 73.562 ;
               RECT 35.254 74.726 35.306 74.762 ;
               RECT 35.254 75.926 35.306 75.962 ;
               RECT 35.254 77.126 35.306 77.162 ;
               RECT 35.254 78.326 35.306 78.362 ;
               RECT 35.254 79.526 35.306 79.562 ;
               RECT 35.254 80.726 35.306 80.762 ;
               RECT 35.254 81.926 35.306 81.962 ;
               RECT 35.254 83.126 35.306 83.162 ;
               RECT 35.254 84.326 35.306 84.362 ;
               RECT 35.254 85.526 35.306 85.562 ;
               RECT 35.254 86.726 35.306 86.762 ;
               RECT 35.254 87.926 35.306 87.962 ;
               RECT 35.254 89.126 35.306 89.162 ;
               RECT 35.254 90.326 35.306 90.362 ;
               RECT 35.254 91.526 35.306 91.562 ;
               RECT 35.254 92.726 35.306 92.762 ;
               RECT 35.254 93.926 35.306 93.962 ;
               RECT 35.254 95.126 35.306 95.162 ;
               RECT 35.254 96.326 35.306 96.362 ;
               RECT 35.254 97.526 35.306 97.562 ;
               RECT 35.254 98.726 35.306 98.762 ;
               RECT 35.254 99.926 35.306 99.962 ;
               RECT 35.254 101.126 35.306 101.162 ;
               RECT 35.254 102.326 35.306 102.362 ;
               RECT 35.254 103.526 35.306 103.562 ;
               RECT 35.334 1.558 35.386 1.594 ;
               RECT 35.334 2.758 35.386 2.794 ;
               RECT 35.334 3.958 35.386 3.994 ;
               RECT 35.334 5.158 35.386 5.194 ;
               RECT 35.334 6.358 35.386 6.394 ;
               RECT 35.334 7.558 35.386 7.594 ;
               RECT 35.334 8.758 35.386 8.794 ;
               RECT 35.334 9.958 35.386 9.994 ;
               RECT 35.334 11.158 35.386 11.194 ;
               RECT 35.334 12.358 35.386 12.394 ;
               RECT 35.334 13.558 35.386 13.594 ;
               RECT 35.334 14.758 35.386 14.794 ;
               RECT 35.334 15.958 35.386 15.994 ;
               RECT 35.334 17.158 35.386 17.194 ;
               RECT 35.334 18.358 35.386 18.394 ;
               RECT 35.334 19.558 35.386 19.594 ;
               RECT 35.334 20.758 35.386 20.794 ;
               RECT 35.334 21.958 35.386 21.994 ;
               RECT 35.334 23.158 35.386 23.194 ;
               RECT 35.334 24.358 35.386 24.394 ;
               RECT 35.334 25.558 35.386 25.594 ;
               RECT 35.334 26.758 35.386 26.794 ;
               RECT 35.334 27.958 35.386 27.994 ;
               RECT 35.334 29.158 35.386 29.194 ;
               RECT 35.334 30.358 35.386 30.394 ;
               RECT 35.334 31.558 35.386 31.594 ;
               RECT 35.334 32.758 35.386 32.794 ;
               RECT 35.334 33.958 35.386 33.994 ;
               RECT 35.334 35.158 35.386 35.194 ;
               RECT 35.334 36.358 35.386 36.394 ;
               RECT 35.334 37.558 35.386 37.594 ;
               RECT 35.334 38.758 35.386 38.794 ;
               RECT 35.334 39.958 35.386 39.994 ;
               RECT 35.334 41.158 35.386 41.194 ;
               RECT 35.334 42.358 35.386 42.394 ;
               RECT 35.334 43.558 35.386 43.594 ;
               RECT 35.334 44.758 35.386 44.794 ;
               RECT 35.334 45.958 35.386 45.994 ;
               RECT 35.334 47.158 35.386 47.194 ;
               RECT 35.334 48.358 35.386 48.394 ;
               RECT 35.334 50.142 35.386 50.178 ;
               RECT 35.334 50.382 35.386 50.418 ;
               RECT 35.334 54.702 35.386 54.738 ;
               RECT 35.334 54.942 35.386 54.978 ;
               RECT 35.334 57.478 35.386 57.514 ;
               RECT 35.334 58.678 35.386 58.714 ;
               RECT 35.334 59.878 35.386 59.914 ;
               RECT 35.334 61.078 35.386 61.114 ;
               RECT 35.334 62.278 35.386 62.314 ;
               RECT 35.334 63.478 35.386 63.514 ;
               RECT 35.334 64.678 35.386 64.714 ;
               RECT 35.334 65.878 35.386 65.914 ;
               RECT 35.334 67.078 35.386 67.114 ;
               RECT 35.334 68.278 35.386 68.314 ;
               RECT 35.334 69.478 35.386 69.514 ;
               RECT 35.334 70.678 35.386 70.714 ;
               RECT 35.334 71.878 35.386 71.914 ;
               RECT 35.334 73.078 35.386 73.114 ;
               RECT 35.334 74.278 35.386 74.314 ;
               RECT 35.334 75.478 35.386 75.514 ;
               RECT 35.334 76.678 35.386 76.714 ;
               RECT 35.334 77.878 35.386 77.914 ;
               RECT 35.334 79.078 35.386 79.114 ;
               RECT 35.334 80.278 35.386 80.314 ;
               RECT 35.334 81.478 35.386 81.514 ;
               RECT 35.334 82.678 35.386 82.714 ;
               RECT 35.334 83.878 35.386 83.914 ;
               RECT 35.334 85.078 35.386 85.114 ;
               RECT 35.334 86.278 35.386 86.314 ;
               RECT 35.334 87.478 35.386 87.514 ;
               RECT 35.334 88.678 35.386 88.714 ;
               RECT 35.334 89.878 35.386 89.914 ;
               RECT 35.334 91.078 35.386 91.114 ;
               RECT 35.334 92.278 35.386 92.314 ;
               RECT 35.334 93.478 35.386 93.514 ;
               RECT 35.334 94.678 35.386 94.714 ;
               RECT 35.334 95.878 35.386 95.914 ;
               RECT 35.334 97.078 35.386 97.114 ;
               RECT 35.334 98.278 35.386 98.314 ;
               RECT 35.334 99.478 35.386 99.514 ;
               RECT 35.334 100.678 35.386 100.714 ;
               RECT 35.334 101.878 35.386 101.914 ;
               RECT 35.334 103.078 35.386 103.114 ;
               RECT 35.334 104.278 35.386 104.314 ;
               RECT 35.414 0.806 35.466 0.842 ;
               RECT 35.414 2.006 35.466 2.042 ;
               RECT 35.414 3.206 35.466 3.242 ;
               RECT 35.414 4.406 35.466 4.442 ;
               RECT 35.414 5.606 35.466 5.642 ;
               RECT 35.414 6.806 35.466 6.842 ;
               RECT 35.414 8.006 35.466 8.042 ;
               RECT 35.414 9.206 35.466 9.242 ;
               RECT 35.414 10.406 35.466 10.442 ;
               RECT 35.414 11.606 35.466 11.642 ;
               RECT 35.414 12.806 35.466 12.842 ;
               RECT 35.414 14.006 35.466 14.042 ;
               RECT 35.414 15.206 35.466 15.242 ;
               RECT 35.414 16.406 35.466 16.442 ;
               RECT 35.414 17.606 35.466 17.642 ;
               RECT 35.414 18.806 35.466 18.842 ;
               RECT 35.414 20.006 35.466 20.042 ;
               RECT 35.414 21.206 35.466 21.242 ;
               RECT 35.414 22.406 35.466 22.442 ;
               RECT 35.414 23.606 35.466 23.642 ;
               RECT 35.414 24.806 35.466 24.842 ;
               RECT 35.414 26.006 35.466 26.042 ;
               RECT 35.414 27.206 35.466 27.242 ;
               RECT 35.414 28.406 35.466 28.442 ;
               RECT 35.414 29.606 35.466 29.642 ;
               RECT 35.414 30.806 35.466 30.842 ;
               RECT 35.414 32.006 35.466 32.042 ;
               RECT 35.414 33.206 35.466 33.242 ;
               RECT 35.414 34.406 35.466 34.442 ;
               RECT 35.414 35.606 35.466 35.642 ;
               RECT 35.414 36.806 35.466 36.842 ;
               RECT 35.414 38.006 35.466 38.042 ;
               RECT 35.414 39.206 35.466 39.242 ;
               RECT 35.414 40.406 35.466 40.442 ;
               RECT 35.414 41.606 35.466 41.642 ;
               RECT 35.414 42.806 35.466 42.842 ;
               RECT 35.414 44.006 35.466 44.042 ;
               RECT 35.414 45.206 35.466 45.242 ;
               RECT 35.414 46.406 35.466 46.442 ;
               RECT 35.414 47.606 35.466 47.642 ;
               RECT 35.414 49.422 35.466 49.458 ;
               RECT 35.414 49.662 35.466 49.698 ;
               RECT 35.414 55.422 35.466 55.458 ;
               RECT 35.414 55.662 35.466 55.698 ;
               RECT 35.414 56.726 35.466 56.762 ;
               RECT 35.414 57.926 35.466 57.962 ;
               RECT 35.414 59.126 35.466 59.162 ;
               RECT 35.414 60.326 35.466 60.362 ;
               RECT 35.414 61.526 35.466 61.562 ;
               RECT 35.414 62.726 35.466 62.762 ;
               RECT 35.414 63.926 35.466 63.962 ;
               RECT 35.414 65.126 35.466 65.162 ;
               RECT 35.414 66.326 35.466 66.362 ;
               RECT 35.414 67.526 35.466 67.562 ;
               RECT 35.414 68.726 35.466 68.762 ;
               RECT 35.414 69.926 35.466 69.962 ;
               RECT 35.414 71.126 35.466 71.162 ;
               RECT 35.414 72.326 35.466 72.362 ;
               RECT 35.414 73.526 35.466 73.562 ;
               RECT 35.414 74.726 35.466 74.762 ;
               RECT 35.414 75.926 35.466 75.962 ;
               RECT 35.414 77.126 35.466 77.162 ;
               RECT 35.414 78.326 35.466 78.362 ;
               RECT 35.414 79.526 35.466 79.562 ;
               RECT 35.414 80.726 35.466 80.762 ;
               RECT 35.414 81.926 35.466 81.962 ;
               RECT 35.414 83.126 35.466 83.162 ;
               RECT 35.414 84.326 35.466 84.362 ;
               RECT 35.414 85.526 35.466 85.562 ;
               RECT 35.414 86.726 35.466 86.762 ;
               RECT 35.414 87.926 35.466 87.962 ;
               RECT 35.414 89.126 35.466 89.162 ;
               RECT 35.414 90.326 35.466 90.362 ;
               RECT 35.414 91.526 35.466 91.562 ;
               RECT 35.414 92.726 35.466 92.762 ;
               RECT 35.414 93.926 35.466 93.962 ;
               RECT 35.414 95.126 35.466 95.162 ;
               RECT 35.414 96.326 35.466 96.362 ;
               RECT 35.414 97.526 35.466 97.562 ;
               RECT 35.414 98.726 35.466 98.762 ;
               RECT 35.414 99.926 35.466 99.962 ;
               RECT 35.414 101.126 35.466 101.162 ;
               RECT 35.414 102.326 35.466 102.362 ;
               RECT 35.414 103.526 35.466 103.562 ;
               RECT 35.494 1.558 35.546 1.594 ;
               RECT 35.494 2.758 35.546 2.794 ;
               RECT 35.494 3.958 35.546 3.994 ;
               RECT 35.494 5.158 35.546 5.194 ;
               RECT 35.494 6.358 35.546 6.394 ;
               RECT 35.494 7.558 35.546 7.594 ;
               RECT 35.494 8.758 35.546 8.794 ;
               RECT 35.494 9.958 35.546 9.994 ;
               RECT 35.494 11.158 35.546 11.194 ;
               RECT 35.494 12.358 35.546 12.394 ;
               RECT 35.494 13.558 35.546 13.594 ;
               RECT 35.494 14.758 35.546 14.794 ;
               RECT 35.494 15.958 35.546 15.994 ;
               RECT 35.494 17.158 35.546 17.194 ;
               RECT 35.494 18.358 35.546 18.394 ;
               RECT 35.494 19.558 35.546 19.594 ;
               RECT 35.494 20.758 35.546 20.794 ;
               RECT 35.494 21.958 35.546 21.994 ;
               RECT 35.494 23.158 35.546 23.194 ;
               RECT 35.494 24.358 35.546 24.394 ;
               RECT 35.494 25.558 35.546 25.594 ;
               RECT 35.494 26.758 35.546 26.794 ;
               RECT 35.494 27.958 35.546 27.994 ;
               RECT 35.494 29.158 35.546 29.194 ;
               RECT 35.494 30.358 35.546 30.394 ;
               RECT 35.494 31.558 35.546 31.594 ;
               RECT 35.494 32.758 35.546 32.794 ;
               RECT 35.494 33.958 35.546 33.994 ;
               RECT 35.494 35.158 35.546 35.194 ;
               RECT 35.494 36.358 35.546 36.394 ;
               RECT 35.494 37.558 35.546 37.594 ;
               RECT 35.494 38.758 35.546 38.794 ;
               RECT 35.494 39.958 35.546 39.994 ;
               RECT 35.494 41.158 35.546 41.194 ;
               RECT 35.494 42.358 35.546 42.394 ;
               RECT 35.494 43.558 35.546 43.594 ;
               RECT 35.494 44.758 35.546 44.794 ;
               RECT 35.494 45.958 35.546 45.994 ;
               RECT 35.494 47.158 35.546 47.194 ;
               RECT 35.494 48.358 35.546 48.394 ;
               RECT 35.494 50.142 35.546 50.178 ;
               RECT 35.494 50.382 35.546 50.418 ;
               RECT 35.494 54.702 35.546 54.738 ;
               RECT 35.494 54.942 35.546 54.978 ;
               RECT 35.494 57.478 35.546 57.514 ;
               RECT 35.494 58.678 35.546 58.714 ;
               RECT 35.494 59.878 35.546 59.914 ;
               RECT 35.494 61.078 35.546 61.114 ;
               RECT 35.494 62.278 35.546 62.314 ;
               RECT 35.494 63.478 35.546 63.514 ;
               RECT 35.494 64.678 35.546 64.714 ;
               RECT 35.494 65.878 35.546 65.914 ;
               RECT 35.494 67.078 35.546 67.114 ;
               RECT 35.494 68.278 35.546 68.314 ;
               RECT 35.494 69.478 35.546 69.514 ;
               RECT 35.494 70.678 35.546 70.714 ;
               RECT 35.494 71.878 35.546 71.914 ;
               RECT 35.494 73.078 35.546 73.114 ;
               RECT 35.494 74.278 35.546 74.314 ;
               RECT 35.494 75.478 35.546 75.514 ;
               RECT 35.494 76.678 35.546 76.714 ;
               RECT 35.494 77.878 35.546 77.914 ;
               RECT 35.494 79.078 35.546 79.114 ;
               RECT 35.494 80.278 35.546 80.314 ;
               RECT 35.494 81.478 35.546 81.514 ;
               RECT 35.494 82.678 35.546 82.714 ;
               RECT 35.494 83.878 35.546 83.914 ;
               RECT 35.494 85.078 35.546 85.114 ;
               RECT 35.494 86.278 35.546 86.314 ;
               RECT 35.494 87.478 35.546 87.514 ;
               RECT 35.494 88.678 35.546 88.714 ;
               RECT 35.494 89.878 35.546 89.914 ;
               RECT 35.494 91.078 35.546 91.114 ;
               RECT 35.494 92.278 35.546 92.314 ;
               RECT 35.494 93.478 35.546 93.514 ;
               RECT 35.494 94.678 35.546 94.714 ;
               RECT 35.494 95.878 35.546 95.914 ;
               RECT 35.494 97.078 35.546 97.114 ;
               RECT 35.494 98.278 35.546 98.314 ;
               RECT 35.494 99.478 35.546 99.514 ;
               RECT 35.494 100.678 35.546 100.714 ;
               RECT 35.494 101.878 35.546 101.914 ;
               RECT 35.494 103.078 35.546 103.114 ;
               RECT 35.494 104.278 35.546 104.314 ;
               RECT 35.574 0.281 35.626 0.317 ;
               RECT 35.574 104.803 35.626 104.839 ;
               RECT 35.946 0.582 35.994 0.618 ;
               RECT 35.946 0.882 35.994 0.918 ;
               RECT 35.946 1.182 35.994 1.218 ;
               RECT 35.946 1.482 35.994 1.518 ;
               RECT 35.946 1.782 35.994 1.818 ;
               RECT 35.946 2.082 35.994 2.118 ;
               RECT 35.946 2.382 35.994 2.418 ;
               RECT 35.946 2.682 35.994 2.718 ;
               RECT 35.946 2.982 35.994 3.018 ;
               RECT 35.946 3.282 35.994 3.318 ;
               RECT 35.946 3.582 35.994 3.618 ;
               RECT 35.946 3.882 35.994 3.918 ;
               RECT 35.946 4.182 35.994 4.218 ;
               RECT 35.946 4.482 35.994 4.518 ;
               RECT 35.946 4.782 35.994 4.818 ;
               RECT 35.946 5.082 35.994 5.118 ;
               RECT 35.946 5.382 35.994 5.418 ;
               RECT 35.946 5.682 35.994 5.718 ;
               RECT 35.946 5.982 35.994 6.018 ;
               RECT 35.946 6.282 35.994 6.318 ;
               RECT 35.946 6.582 35.994 6.618 ;
               RECT 35.946 6.882 35.994 6.918 ;
               RECT 35.946 7.182 35.994 7.218 ;
               RECT 35.946 7.482 35.994 7.518 ;
               RECT 35.946 7.782 35.994 7.818 ;
               RECT 35.946 8.082 35.994 8.118 ;
               RECT 35.946 8.382 35.994 8.418 ;
               RECT 35.946 8.682 35.994 8.718 ;
               RECT 35.946 8.982 35.994 9.018 ;
               RECT 35.946 9.282 35.994 9.318 ;
               RECT 35.946 9.582 35.994 9.618 ;
               RECT 35.946 9.882 35.994 9.918 ;
               RECT 35.946 10.182 35.994 10.218 ;
               RECT 35.946 10.482 35.994 10.518 ;
               RECT 35.946 10.782 35.994 10.818 ;
               RECT 35.946 11.082 35.994 11.118 ;
               RECT 35.946 11.382 35.994 11.418 ;
               RECT 35.946 11.682 35.994 11.718 ;
               RECT 35.946 11.982 35.994 12.018 ;
               RECT 35.946 12.282 35.994 12.318 ;
               RECT 35.946 12.582 35.994 12.618 ;
               RECT 35.946 12.882 35.994 12.918 ;
               RECT 35.946 13.182 35.994 13.218 ;
               RECT 35.946 13.482 35.994 13.518 ;
               RECT 35.946 13.782 35.994 13.818 ;
               RECT 35.946 14.082 35.994 14.118 ;
               RECT 35.946 14.382 35.994 14.418 ;
               RECT 35.946 14.682 35.994 14.718 ;
               RECT 35.946 14.982 35.994 15.018 ;
               RECT 35.946 15.282 35.994 15.318 ;
               RECT 35.946 15.582 35.994 15.618 ;
               RECT 35.946 15.882 35.994 15.918 ;
               RECT 35.946 16.182 35.994 16.218 ;
               RECT 35.946 16.482 35.994 16.518 ;
               RECT 35.946 16.782 35.994 16.818 ;
               RECT 35.946 17.082 35.994 17.118 ;
               RECT 35.946 17.382 35.994 17.418 ;
               RECT 35.946 17.682 35.994 17.718 ;
               RECT 35.946 17.982 35.994 18.018 ;
               RECT 35.946 18.282 35.994 18.318 ;
               RECT 35.946 18.582 35.994 18.618 ;
               RECT 35.946 18.882 35.994 18.918 ;
               RECT 35.946 19.182 35.994 19.218 ;
               RECT 35.946 19.482 35.994 19.518 ;
               RECT 35.946 19.782 35.994 19.818 ;
               RECT 35.946 20.082 35.994 20.118 ;
               RECT 35.946 20.382 35.994 20.418 ;
               RECT 35.946 20.682 35.994 20.718 ;
               RECT 35.946 20.982 35.994 21.018 ;
               RECT 35.946 21.282 35.994 21.318 ;
               RECT 35.946 21.582 35.994 21.618 ;
               RECT 35.946 21.882 35.994 21.918 ;
               RECT 35.946 22.182 35.994 22.218 ;
               RECT 35.946 22.482 35.994 22.518 ;
               RECT 35.946 22.782 35.994 22.818 ;
               RECT 35.946 23.082 35.994 23.118 ;
               RECT 35.946 23.382 35.994 23.418 ;
               RECT 35.946 23.682 35.994 23.718 ;
               RECT 35.946 23.982 35.994 24.018 ;
               RECT 35.946 24.282 35.994 24.318 ;
               RECT 35.946 24.582 35.994 24.618 ;
               RECT 35.946 24.882 35.994 24.918 ;
               RECT 35.946 25.182 35.994 25.218 ;
               RECT 35.946 25.482 35.994 25.518 ;
               RECT 35.946 25.782 35.994 25.818 ;
               RECT 35.946 26.082 35.994 26.118 ;
               RECT 35.946 26.382 35.994 26.418 ;
               RECT 35.946 26.682 35.994 26.718 ;
               RECT 35.946 26.982 35.994 27.018 ;
               RECT 35.946 27.282 35.994 27.318 ;
               RECT 35.946 27.582 35.994 27.618 ;
               RECT 35.946 27.882 35.994 27.918 ;
               RECT 35.946 28.182 35.994 28.218 ;
               RECT 35.946 28.482 35.994 28.518 ;
               RECT 35.946 28.782 35.994 28.818 ;
               RECT 35.946 29.082 35.994 29.118 ;
               RECT 35.946 29.382 35.994 29.418 ;
               RECT 35.946 29.682 35.994 29.718 ;
               RECT 35.946 29.982 35.994 30.018 ;
               RECT 35.946 30.282 35.994 30.318 ;
               RECT 35.946 30.582 35.994 30.618 ;
               RECT 35.946 30.882 35.994 30.918 ;
               RECT 35.946 31.182 35.994 31.218 ;
               RECT 35.946 31.482 35.994 31.518 ;
               RECT 35.946 31.782 35.994 31.818 ;
               RECT 35.946 32.082 35.994 32.118 ;
               RECT 35.946 32.382 35.994 32.418 ;
               RECT 35.946 32.682 35.994 32.718 ;
               RECT 35.946 32.982 35.994 33.018 ;
               RECT 35.946 33.282 35.994 33.318 ;
               RECT 35.946 33.582 35.994 33.618 ;
               RECT 35.946 33.882 35.994 33.918 ;
               RECT 35.946 34.182 35.994 34.218 ;
               RECT 35.946 34.482 35.994 34.518 ;
               RECT 35.946 34.782 35.994 34.818 ;
               RECT 35.946 35.082 35.994 35.118 ;
               RECT 35.946 35.382 35.994 35.418 ;
               RECT 35.946 35.682 35.994 35.718 ;
               RECT 35.946 35.982 35.994 36.018 ;
               RECT 35.946 36.282 35.994 36.318 ;
               RECT 35.946 36.582 35.994 36.618 ;
               RECT 35.946 36.882 35.994 36.918 ;
               RECT 35.946 37.182 35.994 37.218 ;
               RECT 35.946 37.482 35.994 37.518 ;
               RECT 35.946 37.782 35.994 37.818 ;
               RECT 35.946 38.082 35.994 38.118 ;
               RECT 35.946 38.382 35.994 38.418 ;
               RECT 35.946 38.682 35.994 38.718 ;
               RECT 35.946 38.982 35.994 39.018 ;
               RECT 35.946 39.282 35.994 39.318 ;
               RECT 35.946 39.582 35.994 39.618 ;
               RECT 35.946 39.882 35.994 39.918 ;
               RECT 35.946 40.182 35.994 40.218 ;
               RECT 35.946 40.482 35.994 40.518 ;
               RECT 35.946 40.782 35.994 40.818 ;
               RECT 35.946 41.082 35.994 41.118 ;
               RECT 35.946 41.382 35.994 41.418 ;
               RECT 35.946 41.682 35.994 41.718 ;
               RECT 35.946 41.982 35.994 42.018 ;
               RECT 35.946 42.282 35.994 42.318 ;
               RECT 35.946 42.582 35.994 42.618 ;
               RECT 35.946 42.882 35.994 42.918 ;
               RECT 35.946 43.182 35.994 43.218 ;
               RECT 35.946 43.482 35.994 43.518 ;
               RECT 35.946 43.782 35.994 43.818 ;
               RECT 35.946 44.082 35.994 44.118 ;
               RECT 35.946 44.382 35.994 44.418 ;
               RECT 35.946 44.682 35.994 44.718 ;
               RECT 35.946 44.982 35.994 45.018 ;
               RECT 35.946 45.282 35.994 45.318 ;
               RECT 35.946 45.582 35.994 45.618 ;
               RECT 35.946 45.882 35.994 45.918 ;
               RECT 35.946 46.182 35.994 46.218 ;
               RECT 35.946 46.482 35.994 46.518 ;
               RECT 35.946 46.782 35.994 46.818 ;
               RECT 35.946 47.082 35.994 47.118 ;
               RECT 35.946 47.382 35.994 47.418 ;
               RECT 35.946 47.682 35.994 47.718 ;
               RECT 35.946 47.982 35.994 48.018 ;
               RECT 35.946 48.282 35.994 48.318 ;
               RECT 35.946 48.582 35.994 48.618 ;
               RECT 35.946 49.1235 35.994 49.1595 ;
               RECT 35.946 49.422 35.994 49.458 ;
               RECT 35.946 49.7205 35.994 49.7565 ;
               RECT 35.946 50.022 35.994 50.058 ;
               RECT 35.946 50.3235 35.994 50.3595 ;
               RECT 35.946 50.622 35.994 50.658 ;
               RECT 35.946 50.9205 35.994 50.9565 ;
               RECT 35.946 51.222 35.994 51.258 ;
               RECT 35.946 51.5235 35.994 51.5595 ;
               RECT 35.946 52.062 35.994 52.098 ;
               RECT 35.946 52.662 35.994 52.698 ;
               RECT 35.946 52.9635 35.994 52.9995 ;
               RECT 35.946 53.262 35.994 53.298 ;
               RECT 35.946 53.5605 35.994 53.5965 ;
               RECT 35.946 53.862 35.994 53.898 ;
               RECT 35.946 54.1635 35.994 54.1995 ;
               RECT 35.946 54.462 35.994 54.498 ;
               RECT 35.946 54.7605 35.994 54.7965 ;
               RECT 35.946 55.062 35.994 55.098 ;
               RECT 35.946 55.3635 35.994 55.3995 ;
               RECT 35.946 55.662 35.994 55.698 ;
               RECT 35.946 55.9605 35.994 55.9965 ;
               RECT 35.946 56.502 35.994 56.538 ;
               RECT 35.946 56.802 35.994 56.838 ;
               RECT 35.946 57.102 35.994 57.138 ;
               RECT 35.946 57.402 35.994 57.438 ;
               RECT 35.946 57.702 35.994 57.738 ;
               RECT 35.946 58.002 35.994 58.038 ;
               RECT 35.946 58.302 35.994 58.338 ;
               RECT 35.946 58.602 35.994 58.638 ;
               RECT 35.946 58.902 35.994 58.938 ;
               RECT 35.946 59.202 35.994 59.238 ;
               RECT 35.946 59.502 35.994 59.538 ;
               RECT 35.946 59.802 35.994 59.838 ;
               RECT 35.946 60.102 35.994 60.138 ;
               RECT 35.946 60.402 35.994 60.438 ;
               RECT 35.946 60.702 35.994 60.738 ;
               RECT 35.946 61.002 35.994 61.038 ;
               RECT 35.946 61.302 35.994 61.338 ;
               RECT 35.946 61.602 35.994 61.638 ;
               RECT 35.946 61.902 35.994 61.938 ;
               RECT 35.946 62.202 35.994 62.238 ;
               RECT 35.946 62.502 35.994 62.538 ;
               RECT 35.946 62.802 35.994 62.838 ;
               RECT 35.946 63.102 35.994 63.138 ;
               RECT 35.946 63.402 35.994 63.438 ;
               RECT 35.946 63.702 35.994 63.738 ;
               RECT 35.946 64.002 35.994 64.038 ;
               RECT 35.946 64.302 35.994 64.338 ;
               RECT 35.946 64.602 35.994 64.638 ;
               RECT 35.946 64.902 35.994 64.938 ;
               RECT 35.946 65.202 35.994 65.238 ;
               RECT 35.946 65.502 35.994 65.538 ;
               RECT 35.946 65.802 35.994 65.838 ;
               RECT 35.946 66.102 35.994 66.138 ;
               RECT 35.946 66.402 35.994 66.438 ;
               RECT 35.946 66.702 35.994 66.738 ;
               RECT 35.946 67.002 35.994 67.038 ;
               RECT 35.946 67.302 35.994 67.338 ;
               RECT 35.946 67.602 35.994 67.638 ;
               RECT 35.946 67.902 35.994 67.938 ;
               RECT 35.946 68.202 35.994 68.238 ;
               RECT 35.946 68.502 35.994 68.538 ;
               RECT 35.946 68.802 35.994 68.838 ;
               RECT 35.946 69.102 35.994 69.138 ;
               RECT 35.946 69.402 35.994 69.438 ;
               RECT 35.946 69.702 35.994 69.738 ;
               RECT 35.946 70.002 35.994 70.038 ;
               RECT 35.946 70.302 35.994 70.338 ;
               RECT 35.946 70.602 35.994 70.638 ;
               RECT 35.946 70.902 35.994 70.938 ;
               RECT 35.946 71.202 35.994 71.238 ;
               RECT 35.946 71.502 35.994 71.538 ;
               RECT 35.946 71.802 35.994 71.838 ;
               RECT 35.946 72.102 35.994 72.138 ;
               RECT 35.946 72.402 35.994 72.438 ;
               RECT 35.946 72.702 35.994 72.738 ;
               RECT 35.946 73.002 35.994 73.038 ;
               RECT 35.946 73.302 35.994 73.338 ;
               RECT 35.946 73.602 35.994 73.638 ;
               RECT 35.946 73.902 35.994 73.938 ;
               RECT 35.946 74.202 35.994 74.238 ;
               RECT 35.946 74.502 35.994 74.538 ;
               RECT 35.946 74.802 35.994 74.838 ;
               RECT 35.946 75.102 35.994 75.138 ;
               RECT 35.946 75.402 35.994 75.438 ;
               RECT 35.946 75.702 35.994 75.738 ;
               RECT 35.946 76.002 35.994 76.038 ;
               RECT 35.946 76.302 35.994 76.338 ;
               RECT 35.946 76.602 35.994 76.638 ;
               RECT 35.946 76.902 35.994 76.938 ;
               RECT 35.946 77.202 35.994 77.238 ;
               RECT 35.946 77.502 35.994 77.538 ;
               RECT 35.946 77.802 35.994 77.838 ;
               RECT 35.946 78.102 35.994 78.138 ;
               RECT 35.946 78.402 35.994 78.438 ;
               RECT 35.946 78.702 35.994 78.738 ;
               RECT 35.946 79.002 35.994 79.038 ;
               RECT 35.946 79.302 35.994 79.338 ;
               RECT 35.946 79.602 35.994 79.638 ;
               RECT 35.946 79.902 35.994 79.938 ;
               RECT 35.946 80.202 35.994 80.238 ;
               RECT 35.946 80.502 35.994 80.538 ;
               RECT 35.946 80.802 35.994 80.838 ;
               RECT 35.946 81.102 35.994 81.138 ;
               RECT 35.946 81.402 35.994 81.438 ;
               RECT 35.946 81.702 35.994 81.738 ;
               RECT 35.946 82.002 35.994 82.038 ;
               RECT 35.946 82.302 35.994 82.338 ;
               RECT 35.946 82.602 35.994 82.638 ;
               RECT 35.946 82.902 35.994 82.938 ;
               RECT 35.946 83.202 35.994 83.238 ;
               RECT 35.946 83.502 35.994 83.538 ;
               RECT 35.946 83.802 35.994 83.838 ;
               RECT 35.946 84.102 35.994 84.138 ;
               RECT 35.946 84.402 35.994 84.438 ;
               RECT 35.946 84.702 35.994 84.738 ;
               RECT 35.946 85.002 35.994 85.038 ;
               RECT 35.946 85.302 35.994 85.338 ;
               RECT 35.946 85.602 35.994 85.638 ;
               RECT 35.946 85.902 35.994 85.938 ;
               RECT 35.946 86.202 35.994 86.238 ;
               RECT 35.946 86.502 35.994 86.538 ;
               RECT 35.946 86.802 35.994 86.838 ;
               RECT 35.946 87.102 35.994 87.138 ;
               RECT 35.946 87.402 35.994 87.438 ;
               RECT 35.946 87.702 35.994 87.738 ;
               RECT 35.946 88.002 35.994 88.038 ;
               RECT 35.946 88.302 35.994 88.338 ;
               RECT 35.946 88.602 35.994 88.638 ;
               RECT 35.946 88.902 35.994 88.938 ;
               RECT 35.946 89.202 35.994 89.238 ;
               RECT 35.946 89.502 35.994 89.538 ;
               RECT 35.946 89.802 35.994 89.838 ;
               RECT 35.946 90.102 35.994 90.138 ;
               RECT 35.946 90.402 35.994 90.438 ;
               RECT 35.946 90.702 35.994 90.738 ;
               RECT 35.946 91.002 35.994 91.038 ;
               RECT 35.946 91.302 35.994 91.338 ;
               RECT 35.946 91.602 35.994 91.638 ;
               RECT 35.946 91.902 35.994 91.938 ;
               RECT 35.946 92.202 35.994 92.238 ;
               RECT 35.946 92.502 35.994 92.538 ;
               RECT 35.946 92.802 35.994 92.838 ;
               RECT 35.946 93.102 35.994 93.138 ;
               RECT 35.946 93.402 35.994 93.438 ;
               RECT 35.946 93.702 35.994 93.738 ;
               RECT 35.946 94.002 35.994 94.038 ;
               RECT 35.946 94.302 35.994 94.338 ;
               RECT 35.946 94.602 35.994 94.638 ;
               RECT 35.946 94.902 35.994 94.938 ;
               RECT 35.946 95.202 35.994 95.238 ;
               RECT 35.946 95.502 35.994 95.538 ;
               RECT 35.946 95.802 35.994 95.838 ;
               RECT 35.946 96.102 35.994 96.138 ;
               RECT 35.946 96.402 35.994 96.438 ;
               RECT 35.946 96.702 35.994 96.738 ;
               RECT 35.946 97.002 35.994 97.038 ;
               RECT 35.946 97.302 35.994 97.338 ;
               RECT 35.946 97.602 35.994 97.638 ;
               RECT 35.946 97.902 35.994 97.938 ;
               RECT 35.946 98.202 35.994 98.238 ;
               RECT 35.946 98.502 35.994 98.538 ;
               RECT 35.946 98.802 35.994 98.838 ;
               RECT 35.946 99.102 35.994 99.138 ;
               RECT 35.946 99.402 35.994 99.438 ;
               RECT 35.946 99.702 35.994 99.738 ;
               RECT 35.946 100.002 35.994 100.038 ;
               RECT 35.946 100.302 35.994 100.338 ;
               RECT 35.946 100.602 35.994 100.638 ;
               RECT 35.946 100.902 35.994 100.938 ;
               RECT 35.946 101.202 35.994 101.238 ;
               RECT 35.946 101.502 35.994 101.538 ;
               RECT 35.946 101.802 35.994 101.838 ;
               RECT 35.946 102.102 35.994 102.138 ;
               RECT 35.946 102.402 35.994 102.438 ;
               RECT 35.946 102.702 35.994 102.738 ;
               RECT 35.946 103.002 35.994 103.038 ;
               RECT 35.946 103.302 35.994 103.338 ;
               RECT 35.946 103.602 35.994 103.638 ;
               RECT 35.946 103.902 35.994 103.938 ;
               RECT 35.946 104.202 35.994 104.238 ;
               RECT 35.946 104.502 35.994 104.538 ;
     END
END ip764hduspsr2048x39m8b2s0r2p0d0
END LIBRARY
