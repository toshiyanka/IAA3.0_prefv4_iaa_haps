VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf132b256e1r1w0cbbehcaa4acw
  CLASS BLOCK ;
  FOREIGN arf132b256e1r1w0cbbehcaa4acw ;
  ORIGIN 0 0 ;
  SIZE 86.4 BY 29.76 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 16.68 42.772 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 14.76 42.128 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 16.68 43.672 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 16.68 42.128 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 16.68 42.216 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 16.68 42.428 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 16.68 42.516 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 18.6 42.772 19.8 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 18.6 43.028 19.8 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 18.6 43.116 19.8 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 16.68 43.028 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 16.68 43.116 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 16.68 43.328 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 16.68 43.416 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 14.76 43.116 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 14.76 43.328 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 14.76 43.416 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 14.76 43.672 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 12.84 42.128 14.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 12.84 42.216 14.04 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 12.84 42.428 14.04 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 12.84 42.516 14.04 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 14.76 42.216 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 14.76 42.428 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 22.56 20.828 23.76 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 22.56 20.916 23.76 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 22.56 64.372 23.76 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 22.56 64.628 23.76 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 23.28 22.328 24.48 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 23.28 22.416 24.48 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 23.28 65.828 24.48 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 23.28 65.916 24.48 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 24 18.816 25.2 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 24 19.028 25.2 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.572 1.68 65.616 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.784 24 62.828 25.2 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.872 24 62.916 25.2 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 24.72 20.916 25.92 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 24.72 21.172 25.92 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 24.72 64.628 25.92 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 24.72 64.716 25.92 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 25.44 22.416 26.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 25.44 22.628 26.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 25.44 65.916 26.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 25.44 61.328 26.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 1.68 65.828 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.16 19.028 27.36 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 26.16 19.116 27.36 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.084 26.16 63.128 27.36 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.172 26.16 63.216 27.36 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 26.88 21.172 28.08 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 26.88 21.428 28.08 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 26.88 64.716 28.08 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 26.88 64.928 28.08 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 27.6 22.628 28.8 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 27.6 22.716 28.8 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 2.4 18.728 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 27.6 61.416 28.8 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 27.6 61.672 28.8 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 28.32 19.628 29.52 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 28.32 19.716 29.52 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.684 28.32 63.728 29.52 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.772 28.32 63.816 29.52 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 2.4 18.816 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 2.4 62.316 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 2.4 62.572 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 3.12 20.828 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 3.12 20.916 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 3.12 64.372 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 3.12 64.628 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 3.84 22.328 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 3.84 22.416 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 3.84 65.828 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 3.84 65.916 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 4.56 18.816 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 4.56 19.028 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.784 4.56 62.828 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.872 4.56 62.916 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 5.28 20.916 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 5.28 21.172 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 0.24 62.016 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 5.28 64.628 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 5.28 64.716 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 6 22.416 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 6 22.628 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 6 65.916 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 6 61.328 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 6.72 19.028 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 6.72 19.116 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.084 6.72 63.128 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.172 6.72 63.216 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 0.24 62.228 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 7.44 21.172 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 7.44 21.428 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 7.44 64.716 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 7.44 64.928 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 8.16 22.628 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 8.16 22.716 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 8.16 61.416 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 8.16 61.672 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 8.88 19.628 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 8.88 19.716 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 0.96 20.616 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.684 8.88 63.728 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.772 8.88 63.816 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 9.6 21.516 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 9.6 21.728 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.972 9.6 65.016 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.228 9.6 65.272 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 10.32 22.972 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 10.32 18.472 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.884 10.32 61.928 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 10.32 62.016 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 0.96 20.828 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 11.04 20.272 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 11.04 20.528 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.984 11.04 64.028 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 11.04 64.116 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 11.76 21.816 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 11.76 22.072 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.484 11.76 65.528 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.572 11.76 65.616 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 12.48 18.472 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 12.48 18.728 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 0.96 64.116 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 12.48 62.016 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 12.48 62.228 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 13.2 20.616 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 13.2 20.828 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 13.2 64.116 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 13.2 64.372 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 18.24 19.716 19.44 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 18.24 19.928 19.44 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.172 18.24 63.216 19.44 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.428 18.24 63.472 19.44 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 0.96 64.372 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 18.96 21.816 20.16 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 18.96 22.072 20.16 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.484 18.96 65.528 20.16 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.572 18.96 65.616 20.16 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 19.68 18.472 20.88 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 19.68 18.728 20.88 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 19.68 62.016 20.88 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 19.68 62.228 20.88 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 20.4 20.616 21.6 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 20.4 20.828 21.6 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 1.68 22.072 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 20.4 64.116 21.6 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 20.4 64.372 21.6 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 21.12 22.072 22.32 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 21.12 22.328 22.32 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.572 21.12 65.616 22.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 21.12 65.828 22.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 21.84 18.728 23.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 21.84 18.816 23.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 21.84 62.316 23.04 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 21.84 62.572 23.04 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 1.68 22.328 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 14.76 42.772 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 14.76 43.028 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 14.76 42.516 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 22.56 21.172 23.76 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 22.56 21.428 23.76 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 22.56 64.716 23.76 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 22.56 64.928 23.76 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 23.28 22.628 24.48 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 23.28 22.716 24.48 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 23.28 61.328 24.48 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 23.28 61.416 24.48 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 24 19.116 25.2 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 24 19.372 25.2 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 1.68 65.916 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.084 24 63.128 25.2 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.172 24 63.216 25.2 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 24.72 21.428 25.92 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 24.72 21.516 25.92 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 24.72 64.928 25.92 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.972 24.72 65.016 25.92 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 25.44 22.716 26.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 25.44 22.972 26.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 25.44 61.416 26.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 25.44 61.672 26.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 1.68 61.328 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 26.16 19.372 27.36 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 26.16 19.628 27.36 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.428 26.16 63.472 27.36 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.684 26.16 63.728 27.36 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 26.88 21.516 28.08 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 26.88 21.728 28.08 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.972 26.88 65.016 28.08 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.228 26.88 65.272 28.08 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 27.6 22.972 28.8 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 27.6 18.472 28.8 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 2.4 19.028 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.884 27.6 61.928 28.8 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 27.6 62.016 28.8 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 28.32 19.928 29.52 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 28.32 20.016 29.52 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.984 28.32 64.028 29.52 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 28.32 64.116 29.52 ;
    END
  END rddatap0[135]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 2.4 19.116 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.784 2.4 62.828 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.872 2.4 62.916 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 3.12 21.172 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 3.12 21.428 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 3.12 64.716 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 3.12 64.928 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 3.84 22.628 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 3.84 22.716 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 3.84 61.328 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 3.84 61.416 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 4.56 19.116 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 4.56 19.372 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.084 4.56 63.128 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.172 4.56 63.216 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 5.28 21.428 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 5.28 21.516 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 0.24 62.316 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.884 5.28 64.928 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.972 5.28 65.016 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 6 22.716 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 6 22.972 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.372 6 61.416 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.628 6 61.672 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 6.72 19.372 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 6.72 19.628 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.428 6.72 63.472 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.684 6.72 63.728 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 0.24 62.572 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 7.44 21.516 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 7.44 21.728 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.972 7.44 65.016 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.228 7.44 65.272 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 8.16 22.972 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 8.16 18.472 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.884 8.16 61.928 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.972 8.16 62.016 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 8.88 19.928 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 8.88 20.016 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 0.96 20.916 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.984 8.88 64.028 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.072 8.88 64.116 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 9.6 21.816 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 9.6 22.072 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.484 9.6 65.528 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.572 9.6 65.616 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 10.32 18.728 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 10.32 18.816 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.184 10.32 62.228 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 10.32 62.316 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 0.96 21.172 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 11.04 20.616 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 11.04 20.828 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.328 11.04 64.372 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 11.04 64.628 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 11.76 22.328 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 11.76 22.416 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 11.76 65.828 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 11.76 65.916 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 12.48 18.816 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 12.48 19.028 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 0.96 64.628 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 12.48 62.316 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 12.48 62.572 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 13.2 20.916 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 13.2 21.172 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 13.2 64.628 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 13.2 64.716 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 18.24 20.016 19.44 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 18.24 20.272 19.44 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.684 18.24 63.728 19.44 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 63.772 18.24 63.816 19.44 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 0.96 64.716 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 18.96 22.328 20.16 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 18.96 22.416 20.16 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.784 18.96 65.828 20.16 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 18.96 65.916 20.16 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 19.68 18.816 20.88 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 19.68 19.028 20.88 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.272 19.68 62.316 20.88 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.528 19.68 62.572 20.88 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 20.4 20.916 21.6 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 20.4 21.172 21.6 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 1.68 22.416 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.584 20.4 64.628 21.6 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 64.672 20.4 64.716 21.6 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 21.12 22.416 22.32 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 21.12 22.628 22.32 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 65.872 21.12 65.916 22.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 61.284 21.12 61.328 22.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 21.84 19.028 23.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 21.84 19.116 23.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.784 21.84 62.828 23.04 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 62.872 21.84 62.916 23.04 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 1.68 22.628 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 29.7 ;
        RECT 2.662 0.06 2.738 29.7 ;
        RECT 4.462 0.06 4.538 29.7 ;
        RECT 6.262 0.06 6.338 29.7 ;
        RECT 8.062 0.06 8.138 29.7 ;
        RECT 9.862 0.06 9.938 29.7 ;
        RECT 11.662 0.06 11.738 29.7 ;
        RECT 13.462 0.06 13.538 29.7 ;
        RECT 15.262 0.06 15.338 29.7 ;
        RECT 17.062 0.06 17.138 29.7 ;
        RECT 18.862 0.06 18.938 29.7 ;
        RECT 20.662 0.06 20.738 29.7 ;
        RECT 22.462 0.06 22.538 29.7 ;
        RECT 24.262 0.06 24.338 29.7 ;
        RECT 26.062 0.06 26.138 29.7 ;
        RECT 27.862 0.06 27.938 29.7 ;
        RECT 29.662 0.06 29.738 29.7 ;
        RECT 31.462 0.06 31.538 29.7 ;
        RECT 33.262 0.06 33.338 29.7 ;
        RECT 35.062 0.06 35.138 29.7 ;
        RECT 36.862 0.06 36.938 29.7 ;
        RECT 38.662 0.06 38.738 29.7 ;
        RECT 40.462 0.06 40.538 29.7 ;
        RECT 42.262 0.06 42.338 29.7 ;
        RECT 44.062 0.06 44.138 29.7 ;
        RECT 45.862 0.06 45.938 29.7 ;
        RECT 47.662 0.06 47.738 29.7 ;
        RECT 49.462 0.06 49.538 29.7 ;
        RECT 51.262 0.06 51.338 29.7 ;
        RECT 53.062 0.06 53.138 29.7 ;
        RECT 54.862 0.06 54.938 29.7 ;
        RECT 56.662 0.06 56.738 29.7 ;
        RECT 58.462 0.06 58.538 29.7 ;
        RECT 60.262 0.06 60.338 29.7 ;
        RECT 62.062 0.06 62.138 29.7 ;
        RECT 63.862 0.06 63.938 29.7 ;
        RECT 65.662 0.06 65.738 29.7 ;
        RECT 67.462 0.06 67.538 29.7 ;
        RECT 69.262 0.06 69.338 29.7 ;
        RECT 71.062 0.06 71.138 29.7 ;
        RECT 72.862 0.06 72.938 29.7 ;
        RECT 74.662 0.06 74.738 29.7 ;
        RECT 76.462 0.06 76.538 29.7 ;
        RECT 78.262 0.06 78.338 29.7 ;
        RECT 80.062 0.06 80.138 29.7 ;
        RECT 81.862 0.06 81.938 29.7 ;
        RECT 83.662 0.06 83.738 29.7 ;
        RECT 85.462 0.06 85.538 29.7 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 29.7 ;
        RECT 3.562 0.06 3.638 29.7 ;
        RECT 5.362 0.06 5.438 29.7 ;
        RECT 7.162 0.06 7.238 29.7 ;
        RECT 8.962 0.06 9.038 29.7 ;
        RECT 10.762 0.06 10.838 29.7 ;
        RECT 12.562 0.06 12.638 29.7 ;
        RECT 14.362 0.06 14.438 29.7 ;
        RECT 16.162 0.06 16.238 29.7 ;
        RECT 17.962 0.06 18.038 29.7 ;
        RECT 19.762 0.06 19.838 29.7 ;
        RECT 21.562 0.06 21.638 29.7 ;
        RECT 23.362 0.06 23.438 29.7 ;
        RECT 25.162 0.06 25.238 29.7 ;
        RECT 26.962 0.06 27.038 29.7 ;
        RECT 28.762 0.06 28.838 29.7 ;
        RECT 30.562 0.06 30.638 29.7 ;
        RECT 32.362 0.06 32.438 29.7 ;
        RECT 34.162 0.06 34.238 29.7 ;
        RECT 35.962 0.06 36.038 29.7 ;
        RECT 37.762 0.06 37.838 29.7 ;
        RECT 39.562 0.06 39.638 29.7 ;
        RECT 41.362 0.06 41.438 29.7 ;
        RECT 43.162 0.06 43.238 29.7 ;
        RECT 44.962 0.06 45.038 29.7 ;
        RECT 46.762 0.06 46.838 29.7 ;
        RECT 48.562 0.06 48.638 29.7 ;
        RECT 50.362 0.06 50.438 29.7 ;
        RECT 52.162 0.06 52.238 29.7 ;
        RECT 53.962 0.06 54.038 29.7 ;
        RECT 55.762 0.06 55.838 29.7 ;
        RECT 57.562 0.06 57.638 29.7 ;
        RECT 59.362 0.06 59.438 29.7 ;
        RECT 61.162 0.06 61.238 29.7 ;
        RECT 62.962 0.06 63.038 29.7 ;
        RECT 64.762 0.06 64.838 29.7 ;
        RECT 66.562 0.06 66.638 29.7 ;
        RECT 68.362 0.06 68.438 29.7 ;
        RECT 70.162 0.06 70.238 29.7 ;
        RECT 71.962 0.06 72.038 29.7 ;
        RECT 73.762 0.06 73.838 29.7 ;
        RECT 75.562 0.06 75.638 29.7 ;
        RECT 77.362 0.06 77.438 29.7 ;
        RECT 79.162 0.06 79.238 29.7 ;
        RECT 80.962 0.06 81.038 29.7 ;
        RECT 82.762 0.06 82.838 29.7 ;
        RECT 84.562 0.06 84.638 29.7 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 86.416 29.774 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 86.42 29.78 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 86.4705 29.798 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 86.435 29.83 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 86.47 29.798 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 86.459 29.85 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 86.49 29.822 ;
    LAYER m7 SPACING 0 ;
      RECT 85.538 29.82 86.44 29.88 ;
      RECT 85.538 -0.06 86.492 29.82 ;
      RECT 85.538 -0.12 86.44 -0.06 ;
      RECT 84.638 -0.12 85.462 29.88 ;
      RECT 83.738 -0.12 84.562 29.88 ;
      RECT 82.838 -0.12 83.662 29.88 ;
      RECT 81.938 -0.12 82.762 29.88 ;
      RECT 81.038 -0.12 81.862 29.88 ;
      RECT 80.138 -0.12 80.962 29.88 ;
      RECT 79.238 -0.12 80.062 29.88 ;
      RECT 78.338 -0.12 79.162 29.88 ;
      RECT 77.438 -0.12 78.262 29.88 ;
      RECT 76.538 -0.12 77.362 29.88 ;
      RECT 75.638 -0.12 76.462 29.88 ;
      RECT 74.738 -0.12 75.562 29.88 ;
      RECT 73.838 -0.12 74.662 29.88 ;
      RECT 72.938 -0.12 73.762 29.88 ;
      RECT 72.038 -0.12 72.862 29.88 ;
      RECT 71.138 -0.12 71.962 29.88 ;
      RECT 70.238 -0.12 71.062 29.88 ;
      RECT 69.338 -0.12 70.162 29.88 ;
      RECT 68.438 -0.12 69.262 29.88 ;
      RECT 67.538 -0.12 68.362 29.88 ;
      RECT 66.638 -0.12 67.462 29.88 ;
      RECT 65.738 26.64 66.562 29.88 ;
      RECT 65.738 25.44 65.872 26.64 ;
      RECT 65.916 25.44 66.562 26.64 ;
      RECT 65.738 24.48 66.562 25.44 ;
      RECT 65.738 23.28 65.784 24.48 ;
      RECT 65.828 23.28 65.872 24.48 ;
      RECT 65.916 23.28 66.562 24.48 ;
      RECT 65.738 22.32 66.562 23.28 ;
      RECT 65.738 21.12 65.784 22.32 ;
      RECT 65.828 21.12 65.872 22.32 ;
      RECT 65.916 21.12 66.562 22.32 ;
      RECT 65.738 20.16 66.562 21.12 ;
      RECT 65.738 18.96 65.784 20.16 ;
      RECT 65.828 18.96 65.872 20.16 ;
      RECT 65.916 18.96 66.562 20.16 ;
      RECT 65.738 12.96 66.562 18.96 ;
      RECT 65.738 11.76 65.784 12.96 ;
      RECT 65.828 11.76 65.872 12.96 ;
      RECT 65.916 11.76 66.562 12.96 ;
      RECT 65.738 7.2 66.562 11.76 ;
      RECT 65.738 6 65.872 7.2 ;
      RECT 65.916 6 66.562 7.2 ;
      RECT 65.738 5.04 66.562 6 ;
      RECT 65.738 3.84 65.784 5.04 ;
      RECT 65.828 3.84 65.872 5.04 ;
      RECT 65.916 3.84 66.562 5.04 ;
      RECT 65.738 2.88 66.562 3.84 ;
      RECT 65.738 1.68 65.784 2.88 ;
      RECT 65.828 1.68 65.872 2.88 ;
      RECT 65.916 1.68 66.562 2.88 ;
      RECT 65.738 -0.12 66.562 1.68 ;
      RECT 64.838 28.08 65.662 29.88 ;
      RECT 64.838 26.88 64.884 28.08 ;
      RECT 64.928 26.88 64.972 28.08 ;
      RECT 65.016 26.88 65.228 28.08 ;
      RECT 65.272 26.88 65.662 28.08 ;
      RECT 64.838 25.92 65.662 26.88 ;
      RECT 64.838 24.72 64.884 25.92 ;
      RECT 64.928 24.72 64.972 25.92 ;
      RECT 65.016 24.72 65.662 25.92 ;
      RECT 64.838 23.76 65.662 24.72 ;
      RECT 64.838 22.56 64.884 23.76 ;
      RECT 64.928 22.56 65.662 23.76 ;
      RECT 64.838 22.32 65.662 22.56 ;
      RECT 64.838 21.12 65.572 22.32 ;
      RECT 65.616 21.12 65.662 22.32 ;
      RECT 64.838 20.16 65.662 21.12 ;
      RECT 64.838 18.96 65.484 20.16 ;
      RECT 65.528 18.96 65.572 20.16 ;
      RECT 65.616 18.96 65.662 20.16 ;
      RECT 64.838 12.96 65.662 18.96 ;
      RECT 64.838 11.76 65.484 12.96 ;
      RECT 65.528 11.76 65.572 12.96 ;
      RECT 65.616 11.76 65.662 12.96 ;
      RECT 64.838 10.8 65.662 11.76 ;
      RECT 64.838 9.6 64.972 10.8 ;
      RECT 65.016 9.6 65.228 10.8 ;
      RECT 65.272 9.6 65.484 10.8 ;
      RECT 65.528 9.6 65.572 10.8 ;
      RECT 65.616 9.6 65.662 10.8 ;
      RECT 64.838 8.64 65.662 9.6 ;
      RECT 64.838 7.44 64.884 8.64 ;
      RECT 64.928 7.44 64.972 8.64 ;
      RECT 65.016 7.44 65.228 8.64 ;
      RECT 65.272 7.44 65.662 8.64 ;
      RECT 64.838 6.48 65.662 7.44 ;
      RECT 64.838 5.28 64.884 6.48 ;
      RECT 64.928 5.28 64.972 6.48 ;
      RECT 65.016 5.28 65.662 6.48 ;
      RECT 64.838 4.32 65.662 5.28 ;
      RECT 64.838 3.12 64.884 4.32 ;
      RECT 64.928 3.12 65.662 4.32 ;
      RECT 64.838 2.88 65.662 3.12 ;
      RECT 64.838 1.68 65.572 2.88 ;
      RECT 65.616 1.68 65.662 2.88 ;
      RECT 64.838 -0.12 65.662 1.68 ;
      RECT 63.938 29.52 64.762 29.88 ;
      RECT 63.938 28.32 63.984 29.52 ;
      RECT 64.028 28.32 64.072 29.52 ;
      RECT 64.116 28.32 64.762 29.52 ;
      RECT 63.938 28.08 64.762 28.32 ;
      RECT 63.938 26.88 64.672 28.08 ;
      RECT 64.716 26.88 64.762 28.08 ;
      RECT 63.938 25.92 64.762 26.88 ;
      RECT 63.938 24.72 64.584 25.92 ;
      RECT 64.628 24.72 64.672 25.92 ;
      RECT 64.716 24.72 64.762 25.92 ;
      RECT 63.938 23.76 64.762 24.72 ;
      RECT 63.938 22.56 64.328 23.76 ;
      RECT 64.372 22.56 64.584 23.76 ;
      RECT 64.628 22.56 64.672 23.76 ;
      RECT 64.716 22.56 64.762 23.76 ;
      RECT 63.938 21.6 64.762 22.56 ;
      RECT 63.938 20.4 64.072 21.6 ;
      RECT 64.116 20.4 64.328 21.6 ;
      RECT 64.372 20.4 64.584 21.6 ;
      RECT 64.628 20.4 64.672 21.6 ;
      RECT 64.716 20.4 64.762 21.6 ;
      RECT 63.938 14.4 64.762 20.4 ;
      RECT 63.938 13.2 64.072 14.4 ;
      RECT 64.116 13.2 64.328 14.4 ;
      RECT 64.372 13.2 64.584 14.4 ;
      RECT 64.628 13.2 64.672 14.4 ;
      RECT 64.716 13.2 64.762 14.4 ;
      RECT 63.938 12.24 64.762 13.2 ;
      RECT 63.938 11.04 63.984 12.24 ;
      RECT 64.028 11.04 64.072 12.24 ;
      RECT 64.116 11.04 64.328 12.24 ;
      RECT 64.372 11.04 64.584 12.24 ;
      RECT 64.628 11.04 64.762 12.24 ;
      RECT 63.938 10.08 64.762 11.04 ;
      RECT 63.938 8.88 63.984 10.08 ;
      RECT 64.028 8.88 64.072 10.08 ;
      RECT 64.116 8.88 64.762 10.08 ;
      RECT 63.938 8.64 64.762 8.88 ;
      RECT 63.938 7.44 64.672 8.64 ;
      RECT 64.716 7.44 64.762 8.64 ;
      RECT 63.938 6.48 64.762 7.44 ;
      RECT 63.938 5.28 64.584 6.48 ;
      RECT 64.628 5.28 64.672 6.48 ;
      RECT 64.716 5.28 64.762 6.48 ;
      RECT 63.938 4.32 64.762 5.28 ;
      RECT 63.938 3.12 64.328 4.32 ;
      RECT 64.372 3.12 64.584 4.32 ;
      RECT 64.628 3.12 64.672 4.32 ;
      RECT 64.716 3.12 64.762 4.32 ;
      RECT 63.938 2.16 64.762 3.12 ;
      RECT 63.938 0.96 64.072 2.16 ;
      RECT 64.116 0.96 64.328 2.16 ;
      RECT 64.372 0.96 64.584 2.16 ;
      RECT 64.628 0.96 64.672 2.16 ;
      RECT 64.716 0.96 64.762 2.16 ;
      RECT 63.938 -0.12 64.762 0.96 ;
      RECT 63.038 29.52 63.862 29.88 ;
      RECT 63.038 28.32 63.684 29.52 ;
      RECT 63.728 28.32 63.772 29.52 ;
      RECT 63.816 28.32 63.862 29.52 ;
      RECT 63.038 27.36 63.862 28.32 ;
      RECT 63.038 26.16 63.084 27.36 ;
      RECT 63.128 26.16 63.172 27.36 ;
      RECT 63.216 26.16 63.428 27.36 ;
      RECT 63.472 26.16 63.684 27.36 ;
      RECT 63.728 26.16 63.862 27.36 ;
      RECT 63.038 25.2 63.862 26.16 ;
      RECT 63.038 24 63.084 25.2 ;
      RECT 63.128 24 63.172 25.2 ;
      RECT 63.216 24 63.862 25.2 ;
      RECT 63.038 19.44 63.862 24 ;
      RECT 63.038 18.24 63.172 19.44 ;
      RECT 63.216 18.24 63.428 19.44 ;
      RECT 63.472 18.24 63.684 19.44 ;
      RECT 63.728 18.24 63.772 19.44 ;
      RECT 63.816 18.24 63.862 19.44 ;
      RECT 63.038 10.08 63.862 18.24 ;
      RECT 63.038 8.88 63.684 10.08 ;
      RECT 63.728 8.88 63.772 10.08 ;
      RECT 63.816 8.88 63.862 10.08 ;
      RECT 63.038 7.92 63.862 8.88 ;
      RECT 63.038 6.72 63.084 7.92 ;
      RECT 63.128 6.72 63.172 7.92 ;
      RECT 63.216 6.72 63.428 7.92 ;
      RECT 63.472 6.72 63.684 7.92 ;
      RECT 63.728 6.72 63.862 7.92 ;
      RECT 63.038 5.76 63.862 6.72 ;
      RECT 63.038 4.56 63.084 5.76 ;
      RECT 63.128 4.56 63.172 5.76 ;
      RECT 63.216 4.56 63.862 5.76 ;
      RECT 63.038 -0.12 63.862 4.56 ;
      RECT 62.138 25.2 62.962 29.88 ;
      RECT 62.138 24 62.784 25.2 ;
      RECT 62.828 24 62.872 25.2 ;
      RECT 62.916 24 62.962 25.2 ;
      RECT 62.138 23.04 62.962 24 ;
      RECT 62.138 21.84 62.272 23.04 ;
      RECT 62.316 21.84 62.528 23.04 ;
      RECT 62.572 21.84 62.784 23.04 ;
      RECT 62.828 21.84 62.872 23.04 ;
      RECT 62.916 21.84 62.962 23.04 ;
      RECT 62.138 20.88 62.962 21.84 ;
      RECT 62.138 19.68 62.184 20.88 ;
      RECT 62.228 19.68 62.272 20.88 ;
      RECT 62.316 19.68 62.528 20.88 ;
      RECT 62.572 19.68 62.962 20.88 ;
      RECT 62.138 13.68 62.962 19.68 ;
      RECT 62.138 12.48 62.184 13.68 ;
      RECT 62.228 12.48 62.272 13.68 ;
      RECT 62.316 12.48 62.528 13.68 ;
      RECT 62.572 12.48 62.962 13.68 ;
      RECT 62.138 11.52 62.962 12.48 ;
      RECT 62.138 10.32 62.184 11.52 ;
      RECT 62.228 10.32 62.272 11.52 ;
      RECT 62.316 10.32 62.962 11.52 ;
      RECT 62.138 5.76 62.962 10.32 ;
      RECT 62.138 4.56 62.784 5.76 ;
      RECT 62.828 4.56 62.872 5.76 ;
      RECT 62.916 4.56 62.962 5.76 ;
      RECT 62.138 3.6 62.962 4.56 ;
      RECT 62.138 2.4 62.272 3.6 ;
      RECT 62.316 2.4 62.528 3.6 ;
      RECT 62.572 2.4 62.784 3.6 ;
      RECT 62.828 2.4 62.872 3.6 ;
      RECT 62.916 2.4 62.962 3.6 ;
      RECT 62.138 1.44 62.962 2.4 ;
      RECT 62.138 0.24 62.184 1.44 ;
      RECT 62.228 0.24 62.272 1.44 ;
      RECT 62.316 0.24 62.528 1.44 ;
      RECT 62.572 0.24 62.962 1.44 ;
      RECT 62.138 -0.12 62.962 0.24 ;
      RECT 61.238 28.8 62.062 29.88 ;
      RECT 61.238 27.6 61.372 28.8 ;
      RECT 61.416 27.6 61.628 28.8 ;
      RECT 61.672 27.6 61.884 28.8 ;
      RECT 61.928 27.6 61.972 28.8 ;
      RECT 62.016 27.6 62.062 28.8 ;
      RECT 61.238 26.64 62.062 27.6 ;
      RECT 61.238 25.44 61.284 26.64 ;
      RECT 61.328 25.44 61.372 26.64 ;
      RECT 61.416 25.44 61.628 26.64 ;
      RECT 61.672 25.44 62.062 26.64 ;
      RECT 61.238 24.48 62.062 25.44 ;
      RECT 61.238 23.28 61.284 24.48 ;
      RECT 61.328 23.28 61.372 24.48 ;
      RECT 61.416 23.28 62.062 24.48 ;
      RECT 61.238 22.32 62.062 23.28 ;
      RECT 61.238 21.12 61.284 22.32 ;
      RECT 61.328 21.12 62.062 22.32 ;
      RECT 61.238 20.88 62.062 21.12 ;
      RECT 61.238 19.68 61.972 20.88 ;
      RECT 62.016 19.68 62.062 20.88 ;
      RECT 61.238 13.68 62.062 19.68 ;
      RECT 61.238 12.48 61.972 13.68 ;
      RECT 62.016 12.48 62.062 13.68 ;
      RECT 61.238 11.52 62.062 12.48 ;
      RECT 61.238 10.32 61.884 11.52 ;
      RECT 61.928 10.32 61.972 11.52 ;
      RECT 62.016 10.32 62.062 11.52 ;
      RECT 61.238 9.36 62.062 10.32 ;
      RECT 61.238 8.16 61.372 9.36 ;
      RECT 61.416 8.16 61.628 9.36 ;
      RECT 61.672 8.16 61.884 9.36 ;
      RECT 61.928 8.16 61.972 9.36 ;
      RECT 62.016 8.16 62.062 9.36 ;
      RECT 61.238 7.2 62.062 8.16 ;
      RECT 61.238 6 61.284 7.2 ;
      RECT 61.328 6 61.372 7.2 ;
      RECT 61.416 6 61.628 7.2 ;
      RECT 61.672 6 62.062 7.2 ;
      RECT 61.238 5.04 62.062 6 ;
      RECT 61.238 3.84 61.284 5.04 ;
      RECT 61.328 3.84 61.372 5.04 ;
      RECT 61.416 3.84 62.062 5.04 ;
      RECT 61.238 2.88 62.062 3.84 ;
      RECT 61.238 1.68 61.284 2.88 ;
      RECT 61.328 1.68 62.062 2.88 ;
      RECT 61.238 1.44 62.062 1.68 ;
      RECT 61.238 0.24 61.972 1.44 ;
      RECT 62.016 0.24 62.062 1.44 ;
      RECT 61.238 -0.12 62.062 0.24 ;
      RECT 60.338 -0.12 61.162 29.88 ;
      RECT 59.438 -0.12 60.262 29.88 ;
      RECT 58.538 -0.12 59.362 29.88 ;
      RECT 57.638 -0.12 58.462 29.88 ;
      RECT 56.738 -0.12 57.562 29.88 ;
      RECT 55.838 -0.12 56.662 29.88 ;
      RECT 54.938 -0.12 55.762 29.88 ;
      RECT 54.038 -0.12 54.862 29.88 ;
      RECT 53.138 -0.12 53.962 29.88 ;
      RECT 52.238 -0.12 53.062 29.88 ;
      RECT 51.338 -0.12 52.162 29.88 ;
      RECT 50.438 -0.12 51.262 29.88 ;
      RECT 49.538 -0.12 50.362 29.88 ;
      RECT 48.638 -0.12 49.462 29.88 ;
      RECT 47.738 -0.12 48.562 29.88 ;
      RECT 46.838 -0.12 47.662 29.88 ;
      RECT 45.938 -0.12 46.762 29.88 ;
      RECT 45.038 -0.12 45.862 29.88 ;
      RECT 44.138 -0.12 44.962 29.88 ;
      RECT 43.238 17.88 44.062 29.88 ;
      RECT 43.238 16.68 43.284 17.88 ;
      RECT 43.328 16.68 43.372 17.88 ;
      RECT 43.416 16.68 43.628 17.88 ;
      RECT 43.672 16.68 44.062 17.88 ;
      RECT 43.238 15.96 44.062 16.68 ;
      RECT 43.238 14.76 43.284 15.96 ;
      RECT 43.328 14.76 43.372 15.96 ;
      RECT 43.416 14.76 43.628 15.96 ;
      RECT 43.672 14.76 44.062 15.96 ;
      RECT 43.238 -0.12 44.062 14.76 ;
      RECT 42.338 19.8 43.162 29.88 ;
      RECT 42.338 18.6 42.728 19.8 ;
      RECT 42.772 18.6 42.984 19.8 ;
      RECT 43.028 18.6 43.072 19.8 ;
      RECT 43.116 18.6 43.162 19.8 ;
      RECT 42.338 17.88 43.162 18.6 ;
      RECT 42.338 16.68 42.384 17.88 ;
      RECT 42.428 16.68 42.472 17.88 ;
      RECT 42.516 16.68 42.728 17.88 ;
      RECT 42.772 16.68 42.984 17.88 ;
      RECT 43.028 16.68 43.072 17.88 ;
      RECT 43.116 16.68 43.162 17.88 ;
      RECT 42.338 15.96 43.162 16.68 ;
      RECT 42.338 14.76 42.384 15.96 ;
      RECT 42.428 14.76 42.472 15.96 ;
      RECT 42.516 14.76 42.728 15.96 ;
      RECT 42.772 14.76 42.984 15.96 ;
      RECT 43.028 14.76 43.072 15.96 ;
      RECT 43.116 14.76 43.162 15.96 ;
      RECT 42.338 14.04 43.162 14.76 ;
      RECT 42.338 12.84 42.384 14.04 ;
      RECT 42.428 12.84 42.472 14.04 ;
      RECT 42.516 12.84 43.162 14.04 ;
      RECT 42.338 -0.12 43.162 12.84 ;
      RECT 41.438 17.88 42.262 29.88 ;
      RECT 41.438 16.68 42.084 17.88 ;
      RECT 42.128 16.68 42.172 17.88 ;
      RECT 42.216 16.68 42.262 17.88 ;
      RECT 41.438 15.96 42.262 16.68 ;
      RECT 41.438 14.76 42.084 15.96 ;
      RECT 42.128 14.76 42.172 15.96 ;
      RECT 42.216 14.76 42.262 15.96 ;
      RECT 41.438 14.04 42.262 14.76 ;
      RECT 41.438 12.84 42.084 14.04 ;
      RECT 42.128 12.84 42.172 14.04 ;
      RECT 42.216 12.84 42.262 14.04 ;
      RECT 41.438 -0.12 42.262 12.84 ;
      RECT 40.538 -0.12 41.362 29.88 ;
      RECT 39.638 -0.12 40.462 29.88 ;
      RECT 38.738 -0.12 39.562 29.88 ;
      RECT 37.838 -0.12 38.662 29.88 ;
      RECT 36.938 -0.12 37.762 29.88 ;
      RECT 36.038 -0.12 36.862 29.88 ;
      RECT 35.138 -0.12 35.962 29.88 ;
      RECT 34.238 -0.12 35.062 29.88 ;
      RECT 33.338 -0.12 34.162 29.88 ;
      RECT 32.438 -0.12 33.262 29.88 ;
      RECT 31.538 -0.12 32.362 29.88 ;
      RECT 30.638 -0.12 31.462 29.88 ;
      RECT 29.738 -0.12 30.562 29.88 ;
      RECT 28.838 -0.12 29.662 29.88 ;
      RECT 27.938 -0.12 28.762 29.88 ;
      RECT 27.038 -0.12 27.862 29.88 ;
      RECT 26.138 -0.12 26.962 29.88 ;
      RECT 25.238 -0.12 26.062 29.88 ;
      RECT 24.338 -0.12 25.162 29.88 ;
      RECT 23.438 -0.12 24.262 29.88 ;
      RECT 22.538 28.8 23.362 29.88 ;
      RECT 22.538 27.6 22.584 28.8 ;
      RECT 22.628 27.6 22.672 28.8 ;
      RECT 22.716 27.6 22.928 28.8 ;
      RECT 22.972 27.6 23.362 28.8 ;
      RECT 22.538 26.64 23.362 27.6 ;
      RECT 22.538 25.44 22.584 26.64 ;
      RECT 22.628 25.44 22.672 26.64 ;
      RECT 22.716 25.44 22.928 26.64 ;
      RECT 22.972 25.44 23.362 26.64 ;
      RECT 22.538 24.48 23.362 25.44 ;
      RECT 22.538 23.28 22.584 24.48 ;
      RECT 22.628 23.28 22.672 24.48 ;
      RECT 22.716 23.28 23.362 24.48 ;
      RECT 22.538 22.32 23.362 23.28 ;
      RECT 22.538 21.12 22.584 22.32 ;
      RECT 22.628 21.12 23.362 22.32 ;
      RECT 22.538 11.52 23.362 21.12 ;
      RECT 22.538 10.32 22.928 11.52 ;
      RECT 22.972 10.32 23.362 11.52 ;
      RECT 22.538 9.36 23.362 10.32 ;
      RECT 22.538 8.16 22.584 9.36 ;
      RECT 22.628 8.16 22.672 9.36 ;
      RECT 22.716 8.16 22.928 9.36 ;
      RECT 22.972 8.16 23.362 9.36 ;
      RECT 22.538 7.2 23.362 8.16 ;
      RECT 22.538 6 22.584 7.2 ;
      RECT 22.628 6 22.672 7.2 ;
      RECT 22.716 6 22.928 7.2 ;
      RECT 22.972 6 23.362 7.2 ;
      RECT 22.538 5.04 23.362 6 ;
      RECT 22.538 3.84 22.584 5.04 ;
      RECT 22.628 3.84 22.672 5.04 ;
      RECT 22.716 3.84 23.362 5.04 ;
      RECT 22.538 2.88 23.362 3.84 ;
      RECT 22.538 1.68 22.584 2.88 ;
      RECT 22.628 1.68 23.362 2.88 ;
      RECT 22.538 -0.12 23.362 1.68 ;
      RECT 21.638 28.08 22.462 29.88 ;
      RECT 21.638 26.88 21.684 28.08 ;
      RECT 21.728 26.88 22.462 28.08 ;
      RECT 21.638 26.64 22.462 26.88 ;
      RECT 21.638 25.44 22.372 26.64 ;
      RECT 22.416 25.44 22.462 26.64 ;
      RECT 21.638 24.48 22.462 25.44 ;
      RECT 21.638 23.28 22.284 24.48 ;
      RECT 22.328 23.28 22.372 24.48 ;
      RECT 22.416 23.28 22.462 24.48 ;
      RECT 21.638 22.32 22.462 23.28 ;
      RECT 21.638 21.12 22.028 22.32 ;
      RECT 22.072 21.12 22.284 22.32 ;
      RECT 22.328 21.12 22.372 22.32 ;
      RECT 22.416 21.12 22.462 22.32 ;
      RECT 21.638 20.16 22.462 21.12 ;
      RECT 21.638 18.96 21.772 20.16 ;
      RECT 21.816 18.96 22.028 20.16 ;
      RECT 22.072 18.96 22.284 20.16 ;
      RECT 22.328 18.96 22.372 20.16 ;
      RECT 22.416 18.96 22.462 20.16 ;
      RECT 21.638 12.96 22.462 18.96 ;
      RECT 21.638 11.76 21.772 12.96 ;
      RECT 21.816 11.76 22.028 12.96 ;
      RECT 22.072 11.76 22.284 12.96 ;
      RECT 22.328 11.76 22.372 12.96 ;
      RECT 22.416 11.76 22.462 12.96 ;
      RECT 21.638 10.8 22.462 11.76 ;
      RECT 21.638 9.6 21.684 10.8 ;
      RECT 21.728 9.6 21.772 10.8 ;
      RECT 21.816 9.6 22.028 10.8 ;
      RECT 22.072 9.6 22.462 10.8 ;
      RECT 21.638 8.64 22.462 9.6 ;
      RECT 21.638 7.44 21.684 8.64 ;
      RECT 21.728 7.44 22.462 8.64 ;
      RECT 21.638 7.2 22.462 7.44 ;
      RECT 21.638 6 22.372 7.2 ;
      RECT 22.416 6 22.462 7.2 ;
      RECT 21.638 5.04 22.462 6 ;
      RECT 21.638 3.84 22.284 5.04 ;
      RECT 22.328 3.84 22.372 5.04 ;
      RECT 22.416 3.84 22.462 5.04 ;
      RECT 21.638 2.88 22.462 3.84 ;
      RECT 21.638 1.68 22.028 2.88 ;
      RECT 22.072 1.68 22.284 2.88 ;
      RECT 22.328 1.68 22.372 2.88 ;
      RECT 22.416 1.68 22.462 2.88 ;
      RECT 21.638 -0.12 22.462 1.68 ;
      RECT 20.738 28.08 21.562 29.88 ;
      RECT 20.738 26.88 21.128 28.08 ;
      RECT 21.172 26.88 21.384 28.08 ;
      RECT 21.428 26.88 21.472 28.08 ;
      RECT 21.516 26.88 21.562 28.08 ;
      RECT 20.738 25.92 21.562 26.88 ;
      RECT 20.738 24.72 20.872 25.92 ;
      RECT 20.916 24.72 21.128 25.92 ;
      RECT 21.172 24.72 21.384 25.92 ;
      RECT 21.428 24.72 21.472 25.92 ;
      RECT 21.516 24.72 21.562 25.92 ;
      RECT 20.738 23.76 21.562 24.72 ;
      RECT 20.738 22.56 20.784 23.76 ;
      RECT 20.828 22.56 20.872 23.76 ;
      RECT 20.916 22.56 21.128 23.76 ;
      RECT 21.172 22.56 21.384 23.76 ;
      RECT 21.428 22.56 21.562 23.76 ;
      RECT 20.738 21.6 21.562 22.56 ;
      RECT 20.738 20.4 20.784 21.6 ;
      RECT 20.828 20.4 20.872 21.6 ;
      RECT 20.916 20.4 21.128 21.6 ;
      RECT 21.172 20.4 21.562 21.6 ;
      RECT 20.738 14.4 21.562 20.4 ;
      RECT 20.738 13.2 20.784 14.4 ;
      RECT 20.828 13.2 20.872 14.4 ;
      RECT 20.916 13.2 21.128 14.4 ;
      RECT 21.172 13.2 21.562 14.4 ;
      RECT 20.738 12.24 21.562 13.2 ;
      RECT 20.738 11.04 20.784 12.24 ;
      RECT 20.828 11.04 21.562 12.24 ;
      RECT 20.738 10.8 21.562 11.04 ;
      RECT 20.738 9.6 21.472 10.8 ;
      RECT 21.516 9.6 21.562 10.8 ;
      RECT 20.738 8.64 21.562 9.6 ;
      RECT 20.738 7.44 21.128 8.64 ;
      RECT 21.172 7.44 21.384 8.64 ;
      RECT 21.428 7.44 21.472 8.64 ;
      RECT 21.516 7.44 21.562 8.64 ;
      RECT 20.738 6.48 21.562 7.44 ;
      RECT 20.738 5.28 20.872 6.48 ;
      RECT 20.916 5.28 21.128 6.48 ;
      RECT 21.172 5.28 21.384 6.48 ;
      RECT 21.428 5.28 21.472 6.48 ;
      RECT 21.516 5.28 21.562 6.48 ;
      RECT 20.738 4.32 21.562 5.28 ;
      RECT 20.738 3.12 20.784 4.32 ;
      RECT 20.828 3.12 20.872 4.32 ;
      RECT 20.916 3.12 21.128 4.32 ;
      RECT 21.172 3.12 21.384 4.32 ;
      RECT 21.428 3.12 21.562 4.32 ;
      RECT 20.738 2.16 21.562 3.12 ;
      RECT 20.738 0.96 20.784 2.16 ;
      RECT 20.828 0.96 20.872 2.16 ;
      RECT 20.916 0.96 21.128 2.16 ;
      RECT 21.172 0.96 21.562 2.16 ;
      RECT 20.738 -0.12 21.562 0.96 ;
      RECT 19.838 29.52 20.662 29.88 ;
      RECT 19.838 28.32 19.884 29.52 ;
      RECT 19.928 28.32 19.972 29.52 ;
      RECT 20.016 28.32 20.662 29.52 ;
      RECT 19.838 21.6 20.662 28.32 ;
      RECT 19.838 20.4 20.572 21.6 ;
      RECT 20.616 20.4 20.662 21.6 ;
      RECT 19.838 19.44 20.662 20.4 ;
      RECT 19.838 18.24 19.884 19.44 ;
      RECT 19.928 18.24 19.972 19.44 ;
      RECT 20.016 18.24 20.228 19.44 ;
      RECT 20.272 18.24 20.662 19.44 ;
      RECT 19.838 14.4 20.662 18.24 ;
      RECT 19.838 13.2 20.572 14.4 ;
      RECT 20.616 13.2 20.662 14.4 ;
      RECT 19.838 12.24 20.662 13.2 ;
      RECT 19.838 11.04 20.228 12.24 ;
      RECT 20.272 11.04 20.484 12.24 ;
      RECT 20.528 11.04 20.572 12.24 ;
      RECT 20.616 11.04 20.662 12.24 ;
      RECT 19.838 10.08 20.662 11.04 ;
      RECT 19.838 8.88 19.884 10.08 ;
      RECT 19.928 8.88 19.972 10.08 ;
      RECT 20.016 8.88 20.662 10.08 ;
      RECT 19.838 2.16 20.662 8.88 ;
      RECT 19.838 0.96 20.572 2.16 ;
      RECT 20.616 0.96 20.662 2.16 ;
      RECT 19.838 -0.12 20.662 0.96 ;
      RECT 18.938 29.52 19.762 29.88 ;
      RECT 18.938 28.32 19.584 29.52 ;
      RECT 19.628 28.32 19.672 29.52 ;
      RECT 19.716 28.32 19.762 29.52 ;
      RECT 18.938 27.36 19.762 28.32 ;
      RECT 18.938 26.16 18.984 27.36 ;
      RECT 19.028 26.16 19.072 27.36 ;
      RECT 19.116 26.16 19.328 27.36 ;
      RECT 19.372 26.16 19.584 27.36 ;
      RECT 19.628 26.16 19.762 27.36 ;
      RECT 18.938 25.2 19.762 26.16 ;
      RECT 18.938 24 18.984 25.2 ;
      RECT 19.028 24 19.072 25.2 ;
      RECT 19.116 24 19.328 25.2 ;
      RECT 19.372 24 19.762 25.2 ;
      RECT 18.938 23.04 19.762 24 ;
      RECT 18.938 21.84 18.984 23.04 ;
      RECT 19.028 21.84 19.072 23.04 ;
      RECT 19.116 21.84 19.762 23.04 ;
      RECT 18.938 20.88 19.762 21.84 ;
      RECT 18.938 19.68 18.984 20.88 ;
      RECT 19.028 19.68 19.762 20.88 ;
      RECT 18.938 19.44 19.762 19.68 ;
      RECT 18.938 18.24 19.672 19.44 ;
      RECT 19.716 18.24 19.762 19.44 ;
      RECT 18.938 13.68 19.762 18.24 ;
      RECT 18.938 12.48 18.984 13.68 ;
      RECT 19.028 12.48 19.762 13.68 ;
      RECT 18.938 10.08 19.762 12.48 ;
      RECT 18.938 8.88 19.584 10.08 ;
      RECT 19.628 8.88 19.672 10.08 ;
      RECT 19.716 8.88 19.762 10.08 ;
      RECT 18.938 7.92 19.762 8.88 ;
      RECT 18.938 6.72 18.984 7.92 ;
      RECT 19.028 6.72 19.072 7.92 ;
      RECT 19.116 6.72 19.328 7.92 ;
      RECT 19.372 6.72 19.584 7.92 ;
      RECT 19.628 6.72 19.762 7.92 ;
      RECT 18.938 5.76 19.762 6.72 ;
      RECT 18.938 4.56 18.984 5.76 ;
      RECT 19.028 4.56 19.072 5.76 ;
      RECT 19.116 4.56 19.328 5.76 ;
      RECT 19.372 4.56 19.762 5.76 ;
      RECT 18.938 3.6 19.762 4.56 ;
      RECT 18.938 2.4 18.984 3.6 ;
      RECT 19.028 2.4 19.072 3.6 ;
      RECT 19.116 2.4 19.762 3.6 ;
      RECT 18.938 1.44 19.762 2.4 ;
      RECT 18.938 0.24 18.984 1.44 ;
      RECT 19.028 0.24 19.762 1.44 ;
      RECT 18.938 -0.12 19.762 0.24 ;
      RECT 18.038 28.8 18.862 29.88 ;
      RECT 18.038 27.6 18.428 28.8 ;
      RECT 18.472 27.6 18.862 28.8 ;
      RECT 18.038 25.2 18.862 27.6 ;
      RECT 18.038 24 18.772 25.2 ;
      RECT 18.816 24 18.862 25.2 ;
      RECT 18.038 23.04 18.862 24 ;
      RECT 18.038 21.84 18.684 23.04 ;
      RECT 18.728 21.84 18.772 23.04 ;
      RECT 18.816 21.84 18.862 23.04 ;
      RECT 18.038 20.88 18.862 21.84 ;
      RECT 18.038 19.68 18.428 20.88 ;
      RECT 18.472 19.68 18.684 20.88 ;
      RECT 18.728 19.68 18.772 20.88 ;
      RECT 18.816 19.68 18.862 20.88 ;
      RECT 18.038 13.68 18.862 19.68 ;
      RECT 18.038 12.48 18.428 13.68 ;
      RECT 18.472 12.48 18.684 13.68 ;
      RECT 18.728 12.48 18.772 13.68 ;
      RECT 18.816 12.48 18.862 13.68 ;
      RECT 18.038 11.52 18.862 12.48 ;
      RECT 18.038 10.32 18.428 11.52 ;
      RECT 18.472 10.32 18.684 11.52 ;
      RECT 18.728 10.32 18.772 11.52 ;
      RECT 18.816 10.32 18.862 11.52 ;
      RECT 18.038 9.36 18.862 10.32 ;
      RECT 18.038 8.16 18.428 9.36 ;
      RECT 18.472 8.16 18.862 9.36 ;
      RECT 18.038 5.76 18.862 8.16 ;
      RECT 18.038 4.56 18.772 5.76 ;
      RECT 18.816 4.56 18.862 5.76 ;
      RECT 18.038 3.6 18.862 4.56 ;
      RECT 18.038 2.4 18.684 3.6 ;
      RECT 18.728 2.4 18.772 3.6 ;
      RECT 18.816 2.4 18.862 3.6 ;
      RECT 18.038 1.44 18.862 2.4 ;
      RECT 18.038 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.772 1.44 ;
      RECT 18.816 0.24 18.862 1.44 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 29.88 ;
      RECT 16.238 -0.12 17.062 29.88 ;
      RECT 15.338 -0.12 16.162 29.88 ;
      RECT 14.438 -0.12 15.262 29.88 ;
      RECT 13.538 -0.12 14.362 29.88 ;
      RECT 12.638 -0.12 13.462 29.88 ;
      RECT 11.738 -0.12 12.562 29.88 ;
      RECT 10.838 -0.12 11.662 29.88 ;
      RECT 9.938 -0.12 10.762 29.88 ;
      RECT 9.038 -0.12 9.862 29.88 ;
      RECT 8.138 -0.12 8.962 29.88 ;
      RECT 7.238 -0.12 8.062 29.88 ;
      RECT 6.338 -0.12 7.162 29.88 ;
      RECT 5.438 -0.12 6.262 29.88 ;
      RECT 4.538 -0.12 5.362 29.88 ;
      RECT 3.638 -0.12 4.462 29.88 ;
      RECT 2.738 -0.12 3.562 29.88 ;
      RECT 1.838 -0.12 2.662 29.88 ;
      RECT 0.938 -0.12 1.762 29.88 ;
      RECT -0.04 29.82 0.862 29.88 ;
      RECT -0.092 -0.06 0.862 29.82 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 85.658 0 86.32 29.76 ;
      RECT 84.758 0 85.342 29.76 ;
      RECT 83.858 0 84.442 29.76 ;
      RECT 82.958 0 83.542 29.76 ;
      RECT 82.058 0 82.642 29.76 ;
      RECT 81.158 0 81.742 29.76 ;
      RECT 80.258 0 80.842 29.76 ;
      RECT 79.358 0 79.942 29.76 ;
      RECT 78.458 0 79.042 29.76 ;
      RECT 77.558 0 78.142 29.76 ;
      RECT 76.658 0 77.242 29.76 ;
      RECT 75.758 0 76.342 29.76 ;
      RECT 74.858 0 75.442 29.76 ;
      RECT 73.958 0 74.542 29.76 ;
      RECT 73.058 0 73.642 29.76 ;
      RECT 72.158 0 72.742 29.76 ;
      RECT 71.258 0 71.842 29.76 ;
      RECT 70.358 0 70.942 29.76 ;
      RECT 69.458 0 70.042 29.76 ;
      RECT 68.558 0 69.142 29.76 ;
      RECT 67.658 0 68.242 29.76 ;
      RECT 66.758 0 67.342 29.76 ;
      RECT 65.858 26.76 66.442 29.76 ;
      RECT 66.036 25.32 66.442 26.76 ;
      RECT 65.858 24.6 66.442 25.32 ;
      RECT 66.036 23.16 66.442 24.6 ;
      RECT 65.858 22.44 66.442 23.16 ;
      RECT 66.036 21 66.442 22.44 ;
      RECT 65.858 20.28 66.442 21 ;
      RECT 66.036 18.84 66.442 20.28 ;
      RECT 65.858 13.08 66.442 18.84 ;
      RECT 66.036 11.64 66.442 13.08 ;
      RECT 65.858 7.32 66.442 11.64 ;
      RECT 66.036 5.88 66.442 7.32 ;
      RECT 65.858 5.16 66.442 5.88 ;
      RECT 66.036 3.72 66.442 5.16 ;
      RECT 65.858 3 66.442 3.72 ;
      RECT 66.036 1.56 66.442 3 ;
      RECT 65.858 0 66.442 1.56 ;
      RECT 64.958 28.2 65.542 29.76 ;
      RECT 65.392 26.76 65.542 28.2 ;
      RECT 64.958 26.04 65.542 26.76 ;
      RECT 65.136 24.6 65.542 26.04 ;
      RECT 64.958 23.88 65.542 24.6 ;
      RECT 65.048 22.44 65.542 23.88 ;
      RECT 64.958 21 65.452 22.44 ;
      RECT 64.958 20.28 65.542 21 ;
      RECT 64.958 18.84 65.364 20.28 ;
      RECT 64.958 13.08 65.542 18.84 ;
      RECT 64.958 11.64 65.364 13.08 ;
      RECT 64.958 10.92 65.542 11.64 ;
      RECT 64.058 29.64 64.642 29.76 ;
      RECT 64.236 28.2 64.642 29.64 ;
      RECT 64.058 26.76 64.552 28.2 ;
      RECT 64.058 26.04 64.642 26.76 ;
      RECT 64.058 24.6 64.464 26.04 ;
      RECT 64.058 23.88 64.642 24.6 ;
      RECT 64.058 22.44 64.208 23.88 ;
      RECT 64.058 21.72 64.642 22.44 ;
      RECT 63.158 29.64 63.742 29.76 ;
      RECT 63.158 28.2 63.564 29.64 ;
      RECT 63.158 27.48 63.742 28.2 ;
      RECT 62.258 25.32 62.842 29.76 ;
      RECT 62.258 23.88 62.664 25.32 ;
      RECT 62.258 23.16 62.842 23.88 ;
      RECT 61.358 28.92 61.942 29.76 ;
      RECT 60.458 0 61.042 29.76 ;
      RECT 59.558 0 60.142 29.76 ;
      RECT 58.658 0 59.242 29.76 ;
      RECT 57.758 0 58.342 29.76 ;
      RECT 56.858 0 57.442 29.76 ;
      RECT 55.958 0 56.542 29.76 ;
      RECT 55.058 0 55.642 29.76 ;
      RECT 54.158 0 54.742 29.76 ;
      RECT 53.258 0 53.842 29.76 ;
      RECT 52.358 0 52.942 29.76 ;
      RECT 51.458 0 52.042 29.76 ;
      RECT 50.558 0 51.142 29.76 ;
      RECT 49.658 0 50.242 29.76 ;
      RECT 48.758 0 49.342 29.76 ;
      RECT 47.858 0 48.442 29.76 ;
      RECT 46.958 0 47.542 29.76 ;
      RECT 46.058 0 46.642 29.76 ;
      RECT 45.158 0 45.742 29.76 ;
      RECT 44.258 0 44.842 29.76 ;
      RECT 43.358 18 43.942 29.76 ;
      RECT 43.792 16.56 43.942 18 ;
      RECT 43.358 16.08 43.942 16.56 ;
      RECT 43.792 14.64 43.942 16.08 ;
      RECT 43.358 0 43.942 14.64 ;
      RECT 42.458 19.92 43.042 29.76 ;
      RECT 42.458 18.48 42.608 19.92 ;
      RECT 42.458 18 43.042 18.48 ;
      RECT 41.558 18 42.142 29.76 ;
      RECT 41.558 16.56 41.964 18 ;
      RECT 41.558 16.08 42.142 16.56 ;
      RECT 41.558 14.64 41.964 16.08 ;
      RECT 41.558 14.16 42.142 14.64 ;
      RECT 41.558 12.72 41.964 14.16 ;
      RECT 41.558 0 42.142 12.72 ;
      RECT 40.658 0 41.242 29.76 ;
      RECT 39.758 0 40.342 29.76 ;
      RECT 38.858 0 39.442 29.76 ;
      RECT 37.958 0 38.542 29.76 ;
      RECT 37.058 0 37.642 29.76 ;
      RECT 36.158 0 36.742 29.76 ;
      RECT 35.258 0 35.842 29.76 ;
      RECT 34.358 0 34.942 29.76 ;
      RECT 33.458 0 34.042 29.76 ;
      RECT 32.558 0 33.142 29.76 ;
      RECT 31.658 0 32.242 29.76 ;
      RECT 30.758 0 31.342 29.76 ;
      RECT 29.858 0 30.442 29.76 ;
      RECT 28.958 0 29.542 29.76 ;
      RECT 28.058 0 28.642 29.76 ;
      RECT 27.158 0 27.742 29.76 ;
      RECT 26.258 0 26.842 29.76 ;
      RECT 25.358 0 25.942 29.76 ;
      RECT 24.458 0 25.042 29.76 ;
      RECT 23.558 0 24.142 29.76 ;
      RECT 22.658 28.92 23.242 29.76 ;
      RECT 23.092 27.48 23.242 28.92 ;
      RECT 22.658 26.76 23.242 27.48 ;
      RECT 23.092 25.32 23.242 26.76 ;
      RECT 22.658 24.6 23.242 25.32 ;
      RECT 22.836 23.16 23.242 24.6 ;
      RECT 22.658 22.44 23.242 23.16 ;
      RECT 22.748 21 23.242 22.44 ;
      RECT 22.658 11.64 23.242 21 ;
      RECT 22.658 10.2 22.808 11.64 ;
      RECT 23.092 10.2 23.242 11.64 ;
      RECT 22.658 9.48 23.242 10.2 ;
      RECT 23.092 8.04 23.242 9.48 ;
      RECT 22.658 7.32 23.242 8.04 ;
      RECT 23.092 5.88 23.242 7.32 ;
      RECT 22.658 5.16 23.242 5.88 ;
      RECT 22.836 3.72 23.242 5.16 ;
      RECT 22.658 3 23.242 3.72 ;
      RECT 22.748 1.56 23.242 3 ;
      RECT 22.658 0 23.242 1.56 ;
      RECT 21.758 28.2 22.342 29.76 ;
      RECT 21.848 26.76 22.342 28.2 ;
      RECT 21.758 25.32 22.252 26.76 ;
      RECT 21.758 24.6 22.342 25.32 ;
      RECT 21.758 23.16 22.164 24.6 ;
      RECT 21.758 22.44 22.342 23.16 ;
      RECT 21.758 21 21.908 22.44 ;
      RECT 21.758 20.28 22.342 21 ;
      RECT 20.858 28.2 21.442 29.76 ;
      RECT 20.858 26.76 21.008 28.2 ;
      RECT 20.858 26.04 21.442 26.76 ;
      RECT 19.958 29.64 20.542 29.76 ;
      RECT 20.136 28.2 20.542 29.64 ;
      RECT 19.958 21.72 20.542 28.2 ;
      RECT 19.958 20.28 20.452 21.72 ;
      RECT 19.958 19.56 20.542 20.28 ;
      RECT 20.392 18.12 20.542 19.56 ;
      RECT 19.958 14.52 20.542 18.12 ;
      RECT 19.958 13.08 20.452 14.52 ;
      RECT 19.958 12.36 20.542 13.08 ;
      RECT 19.958 10.92 20.108 12.36 ;
      RECT 19.958 10.2 20.542 10.92 ;
      RECT 20.136 8.76 20.542 10.2 ;
      RECT 19.958 2.28 20.542 8.76 ;
      RECT 19.958 0.84 20.452 2.28 ;
      RECT 19.958 0 20.542 0.84 ;
      RECT 19.058 29.64 19.642 29.76 ;
      RECT 19.058 28.2 19.464 29.64 ;
      RECT 19.058 27.48 19.642 28.2 ;
      RECT 18.158 28.92 18.742 29.76 ;
      RECT 18.158 27.48 18.308 28.92 ;
      RECT 18.592 27.48 18.742 28.92 ;
      RECT 18.158 25.32 18.742 27.48 ;
      RECT 18.158 23.88 18.652 25.32 ;
      RECT 18.158 23.16 18.742 23.88 ;
      RECT 18.158 21.72 18.564 23.16 ;
      RECT 18.158 21 18.742 21.72 ;
      RECT 18.158 19.56 18.308 21 ;
      RECT 18.158 13.8 18.742 19.56 ;
      RECT 18.158 12.36 18.308 13.8 ;
      RECT 18.158 11.64 18.742 12.36 ;
      RECT 18.158 10.2 18.308 11.64 ;
      RECT 18.158 9.48 18.742 10.2 ;
      RECT 18.158 8.04 18.308 9.48 ;
      RECT 18.592 8.04 18.742 9.48 ;
      RECT 18.158 5.88 18.742 8.04 ;
      RECT 18.158 4.44 18.652 5.88 ;
      RECT 18.158 3.72 18.742 4.44 ;
      RECT 18.158 2.28 18.564 3.72 ;
      RECT 18.158 1.56 18.742 2.28 ;
      RECT 18.158 0.12 18.308 1.56 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 29.76 ;
      RECT 16.358 0 16.942 29.76 ;
      RECT 15.458 0 16.042 29.76 ;
      RECT 14.558 0 15.142 29.76 ;
      RECT 13.658 0 14.242 29.76 ;
      RECT 12.758 0 13.342 29.76 ;
      RECT 11.858 0 12.442 29.76 ;
      RECT 10.958 0 11.542 29.76 ;
      RECT 10.058 0 10.642 29.76 ;
      RECT 9.158 0 9.742 29.76 ;
      RECT 8.258 0 8.842 29.76 ;
      RECT 7.358 0 7.942 29.76 ;
      RECT 6.458 0 7.042 29.76 ;
      RECT 5.558 0 6.142 29.76 ;
      RECT 4.658 0 5.242 29.76 ;
      RECT 3.758 0 4.342 29.76 ;
      RECT 2.858 0 3.442 29.76 ;
      RECT 1.958 0 2.542 29.76 ;
      RECT 1.058 0 1.642 29.76 ;
      RECT 0.08 0 0.742 29.76 ;
      RECT 61.358 26.76 61.942 27.48 ;
      RECT 61.792 25.32 61.942 26.76 ;
      RECT 61.358 24.6 61.942 25.32 ;
      RECT 61.536 23.16 61.942 24.6 ;
      RECT 61.358 22.44 61.942 23.16 ;
      RECT 61.448 21 61.942 22.44 ;
      RECT 61.358 19.56 61.852 21 ;
      RECT 61.358 13.8 61.942 19.56 ;
      RECT 61.358 12.36 61.852 13.8 ;
      RECT 61.358 11.64 61.942 12.36 ;
      RECT 61.358 10.2 61.764 11.64 ;
      RECT 61.358 9.48 61.942 10.2 ;
      RECT 63.158 25.32 63.742 26.04 ;
      RECT 63.336 23.88 63.742 25.32 ;
      RECT 63.158 19.56 63.742 23.88 ;
      RECT 19.058 25.32 19.642 26.04 ;
      RECT 19.492 23.88 19.642 25.32 ;
      RECT 19.058 23.16 19.642 23.88 ;
      RECT 19.236 21.72 19.642 23.16 ;
      RECT 19.058 21 19.642 21.72 ;
      RECT 19.148 19.56 19.642 21 ;
      RECT 19.058 18.12 19.552 19.56 ;
      RECT 19.058 13.8 19.642 18.12 ;
      RECT 19.148 12.36 19.642 13.8 ;
      RECT 19.058 10.2 19.642 12.36 ;
      RECT 19.058 8.76 19.464 10.2 ;
      RECT 19.058 8.04 19.642 8.76 ;
      RECT 20.858 23.88 21.442 24.6 ;
      RECT 20.858 21.72 21.442 22.44 ;
      RECT 21.292 20.28 21.442 21.72 ;
      RECT 20.858 14.52 21.442 20.28 ;
      RECT 21.292 13.08 21.442 14.52 ;
      RECT 20.858 12.36 21.442 13.08 ;
      RECT 20.948 10.92 21.442 12.36 ;
      RECT 20.858 9.48 21.352 10.92 ;
      RECT 20.858 8.76 21.442 9.48 ;
      RECT 20.858 7.32 21.008 8.76 ;
      RECT 20.858 6.6 21.442 7.32 ;
      RECT 62.258 21 62.842 21.72 ;
      RECT 62.692 19.56 62.842 21 ;
      RECT 62.258 13.8 62.842 19.56 ;
      RECT 62.692 12.36 62.842 13.8 ;
      RECT 62.258 11.64 62.842 12.36 ;
      RECT 62.436 10.2 62.842 11.64 ;
      RECT 62.258 5.88 62.842 10.2 ;
      RECT 62.258 4.44 62.664 5.88 ;
      RECT 62.258 3.72 62.842 4.44 ;
      RECT 64.058 14.52 64.642 20.28 ;
      RECT 21.758 13.08 22.342 18.84 ;
      RECT 63.158 10.2 63.742 18.12 ;
      RECT 63.158 8.76 63.564 10.2 ;
      RECT 63.158 8.04 63.742 8.76 ;
      RECT 42.458 16.08 43.042 16.56 ;
      RECT 42.458 14.16 43.042 14.64 ;
      RECT 42.636 12.72 43.042 14.16 ;
      RECT 42.458 0 43.042 12.72 ;
      RECT 64.058 12.36 64.642 13.08 ;
      RECT 21.758 10.92 22.342 11.64 ;
      RECT 22.192 9.48 22.342 10.92 ;
      RECT 21.758 8.76 22.342 9.48 ;
      RECT 21.848 7.32 22.342 8.76 ;
      RECT 21.758 5.88 22.252 7.32 ;
      RECT 21.758 5.16 22.342 5.88 ;
      RECT 21.758 3.72 22.164 5.16 ;
      RECT 21.758 3 22.342 3.72 ;
      RECT 21.758 1.56 21.908 3 ;
      RECT 21.758 0 22.342 1.56 ;
      RECT 64.058 10.2 64.642 10.92 ;
      RECT 64.236 8.76 64.642 10.2 ;
      RECT 64.058 7.32 64.552 8.76 ;
      RECT 64.058 6.6 64.642 7.32 ;
      RECT 64.058 5.16 64.464 6.6 ;
      RECT 64.058 4.44 64.642 5.16 ;
      RECT 64.058 3 64.208 4.44 ;
      RECT 64.058 2.28 64.642 3 ;
      RECT 64.958 8.76 65.542 9.48 ;
      RECT 65.392 7.32 65.542 8.76 ;
      RECT 64.958 6.6 65.542 7.32 ;
      RECT 65.136 5.16 65.542 6.6 ;
      RECT 64.958 4.44 65.542 5.16 ;
      RECT 65.048 3 65.542 4.44 ;
      RECT 64.958 1.56 65.452 3 ;
      RECT 64.958 0 65.542 1.56 ;
      RECT 61.358 7.32 61.942 8.04 ;
      RECT 61.792 5.88 61.942 7.32 ;
      RECT 61.358 5.16 61.942 5.88 ;
      RECT 61.536 3.72 61.942 5.16 ;
      RECT 61.358 3 61.942 3.72 ;
      RECT 61.448 1.56 61.942 3 ;
      RECT 61.358 0.12 61.852 1.56 ;
      RECT 61.358 0 61.942 0.12 ;
      RECT 63.158 5.88 63.742 6.6 ;
      RECT 63.336 4.44 63.742 5.88 ;
      RECT 63.158 0 63.742 4.44 ;
      RECT 19.058 5.88 19.642 6.6 ;
      RECT 19.492 4.44 19.642 5.88 ;
      RECT 19.058 3.72 19.642 4.44 ;
      RECT 19.236 2.28 19.642 3.72 ;
      RECT 19.058 1.56 19.642 2.28 ;
      RECT 19.148 0.12 19.642 1.56 ;
      RECT 19.058 0 19.642 0.12 ;
      RECT 20.858 4.44 21.442 5.16 ;
      RECT 20.858 2.28 21.442 3 ;
      RECT 21.292 0.84 21.442 2.28 ;
      RECT 20.858 0 21.442 0.84 ;
      RECT 62.258 1.56 62.842 2.28 ;
      RECT 62.692 0.12 62.842 1.56 ;
      RECT 62.258 0 62.842 0.12 ;
      RECT 64.058 0 64.642 0.84 ;
    LAYER m0 ;
      RECT 0 0.002 86.4 29.758 ;
    LAYER m1 ;
      RECT 0 0 86.4 29.76 ;
    LAYER m2 ;
      RECT 0 0.015 86.4 29.745 ;
    LAYER m3 ;
      RECT 0.015 0 86.385 29.76 ;
    LAYER m4 ;
      RECT 0 0.02 86.4 29.74 ;
    LAYER m5 ;
      RECT 0.012 0 86.388 29.76 ;
    LAYER m6 ;
      RECT 0 0.012 86.4 29.748 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf132b256e1r1w0cbbehcaa4acw

END LIBRARY
