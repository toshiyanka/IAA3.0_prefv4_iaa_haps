        //packets used 
      `include_typ("cfg_packet.sv")
      `include_typ("cfg_errcheck_packet.sv")
      `include_typ("mem_packet.sv")
      `include_typ("msg_packet.sv")
      `include_typ("mix_packet.sv")
      `include_typ("mem_badtxn_packet.sv")
      `include_typ("mem_errcheck_packet.sv")

                
      //generic sequence
      `include_typ("hqm_iosf_prim_memory_rd_seq.sv")
      `include_typ("hqm_iosf_config_rd_seq.sv")
      `include_typ("hqm_iosf_config_wr_seq.sv")
      `include_typ("hqm_iosf_config_rd_UR_seq.sv")
      `include_typ("hqm_iosf_config_wr_UR_seq.sv")
      `include_typ("hqm_iosf_config_wr_rqid_seq.sv")
      `include_typ("hqm_iosf_config_rd_rqid_seq.sv")
      `include_typ("hqm_iosf_prim_mem_rd_rqid_seq.sv")
      `include_typ("hqm_iosf_prim_mem_wr_rqid_seq.sv")
      `include_typ("hqm_iosf_config_seq11.sv")
      `include_typ("mix_generic_seq.sv")
      `include_typ("mix_generic_seq1.sv")
      `include_typ("cfg_genric_seq11.sv")
      //`include_typ("back2back_cfgrdwr_seq1.sv")
      `include_typ("cfg_common_seq.sv")
      `include_typ("error_common_seq.sv")



      //back2back sequence
      `include_typ("back2back_posted_wrd_rqid_seq.sv")
      `include_typ("back2back_cfgwr_rd_seq.sv")

       //stress sequences
      `include_typ("np_p_seq.sv")
      `include_typ("np_p_seq1.sv")
      `include_typ("np_np_seq1.sv")

      //badparity and badtxn sequences
      `include_typ("hqm_iosf_prim_cfg_rd_badparity_seq.sv")
      `include_typ("hqm_iosf_prim_cfg_wr_badparity_seq.sv")
      `include_typ("hqm_iosf_prim_mem_wr_badparity_seq.sv")
      `include_typ("hqm_iosf_prim_mem_rd_badparity_seq.sv")
      `include_typ("hqm_iosf_prim_cfg_wr_badLength_seq.sv")
      `include_typ("hqm_iosf_prim_cfg_wr_badtxn_seq.sv")

      //`include_typ("back2back_cfgwr_badDataparity_seq1.sv")
      //`include_typ("back2back_cfgrd_badCmdparity_seq.sv")
      `include_typ("back2back_posted_badDataparity_seq2.sv")

      //back2back memrd
      //`include_typ("back2back_memrdwr_seq2.sv")
      `include_typ("back2back_cfgrd_param_seq.sv")

      //poison sequence
      `include_typ("hqm_iosf_prim_cfg_wr_poisoned_seq.sv")
      `include_typ("back2back_cfgwr_poison_seq.sv")
      `include_typ("hqm_iosf_prim_mem_wr_poison_seq.sv")
      `include_typ("back2back_posted_poison_seq.sv")
      `include_typ("back2back_posted_poison_seq1.sv")
      `include_typ("back2back_posted_poison_seq2.sv")



      //ecrc sequence
      `include_typ("hqm_iosf_prim_cfg_rd_badecrc_seq.sv") 
      `include_typ("back2back_cfgrd_ecrc_seq.sv")
      `include_typ("hqm_iosf_prim_cfg_wr_badecrc_seq.sv") 
      `include_typ("back2back_cfgwr_ecrc_seq.sv")
      `include_typ("hqm_iosf_tb_file_seq.sv")
      `include_typ("back2back_cfgrd_badCmdparity_seq1.sv")

      //unsupported sequence
      `include_typ("back2back_posted_unsupported_seq.sv")
      `include_typ("back2back_memrd_unsupported_seq.sv")
      `include_typ("back2back_cfgrd_unsupported_seq.sv")
      `include_typ("back2back_cfgwr_unsupported_seq.sv")
      `include_typ("back2back_unaligned_seq.sv")

      //badlength sequence
      //`include_typ("back2back_cfgwr_badtxn_seq.sv")
      `include_typ("back2back_cfgwr_badlength_seq.sv")
      `include_typ("hqm_iosf_prim_mem_wr_badtxn_seq.sv")
      `include_typ("back2back_cfgwr_badlength_seq11.sv")
      `include_typ("back2back_cfgwr_badlength_seq22.sv")
 
      //LBE check
      `include_typ("hqm_iosf_config_wr_URlbe_seq.sv")
      `include_typ("hqm_iosf_config_rd_URlbe_seq.sv")
      `include_typ("hqm_iosf_prim_memory_rd_lbe_seq.sv")
      `include_typ("hqm_iosf_prim_mem_wr_badlbe_seq.sv")
      `include_typ("back2back_cfgwr_badlbe_seq1.sv")
      `include_typ("back2back_memwr_badtxn_seq.sv")


      //SAI sequences
      `include_typ("hqm_sai_config_rd_seq.sv")
      `include_typ("hqm_sai_config_wr_seq.sv")
      `include_typ("hqm_sai_memory_rd_seq.sv")
      `include_typ("hqm_sai_memory_wr_seq.sv")
      `include_typ("sai_packet.sv")
      `include_typ("SAI_seq.sv")
      `include_typ("SAI_invalid_seq.sv")
      `include_typ("SAI_invalid_all_seq.sv")
      `include_typ("SAI_valid_seq.sv")

     // `include_typ("SAI_meminvalid_seq.sv")
      `include_typ("SAI_invalid_seq1.sv")
      `include_typ("SAI_memrdinvalid_seq.sv")
      `include_typ("SAI_memrdinvalid_feature_seq.sv")
      `include_typ("SAI_memrdinvalid_dbg_seq.sv")
      `include_typ("SAI_memwrinvalid_feature_seq.sv")
      `include_typ("SAI_memwrinvalid_dbg_seq.sv")
      `include_typ("SAI_memwrinvalid_csr_seq.sv")
      `include_typ("SAI_UR_seq.sv")
 
      //unsupported commands seq
      `include_typ("hqm_iosf_prim_msg_seq.sv")
      `include_typ("hqm_iosf_config1_rd_seq.sv")
      `include_typ("hqm_iosf_config1_wr_seq.sv")
      `include_typ("hqm_iosf_unsupport_transaction_seq.sv")
      `include_typ("hqm_iosf_unsupport_memory_seq.sv")
      `include_typ("hqm_iosf_unsupport_memwr_seq.sv")
      `include_typ("hqm_iosf_unsupport_atomic_seq.sv")
      `include_typ("back2back_posted_msg_seq.sv")
      `include_typ("back2back_unsupport_memrd_seq.sv")
      `include_typ("back2back_unsupport_memwr_seq.sv")
      `include_typ("back2back_cfg1_seq.sv")

      //unexpected completion 
       `include_typ( "hqm_iosf_cplLk_seq.sv")

     
   //sideband sequences
   `include_typ("iosf_sb_file_seq.sv")
   `include_typ("cfg_sb_packet.sv") 
   `include_typ("mem_sb_packet.sv")
   `include_typ("hqm_iosf_sb_cfgrd_seq.sv")
   `include_typ("hqm_iosf_sb_cfgwr_seq.sv")
   `include_typ("hqm_iosf_sb_memwr_seq.sv")
   `include_typ("hqm_iosf_sb_memwr_np_seq1.sv")
   `include_typ("hqm_iosf_sb_memwr32_seq.sv")
   `include_typ("hqm_iosf_sb_memrd32_seq.sv")
   `include_typ("hqm_iosf_sb_unsupport_cfgrd_seq.sv")
   `include_typ("hqm_iosf_sb_unsupport_cfgwr_seq.sv")
   //`include_typ("hqm_iosf_sb_cfgrd_loopback_seq.sv")
   `include_typ("hqm_iosf_sb_forcewake_seq.sv")  // `include_mid
   `include_typ("hqm_iosf_sb_resetPrep_seq.sv")  // `include_mid
   `include_typ("hqm_iosf_sb_fuse_download_seq.sv")
   `include_typ("back2back_sb_fw_seq.sv")
   `include_typ("back2back_sb_nak_seq.sv")
   `include_typ("back2back_sb_memwr32_seq.sv")
   `include_typ("hqm_iosf_memrd_bar_seq.sv")
   `include_typ("hqm_iosf_sb_memwr_bar_seq.sv")
  // `include_typ("hqm_iosf_sb_memwr_brdcast_seq.sv")

   //broadcast sequence
   `include_typ("hqm_iosf_sb_cfgrd_brdcast_seq.sv")
   `include_typ("hqm_iosf_sb_cfgrd_brdcast1_seq.sv")
   `include_typ("hqm_iosf_sb_cfgrd_brdcast2_seq.sv")

   `include_typ("hqm_iosf_sb_cfgwr_brdcast_seq.sv")
   `include_typ("hqm_iosf_sb_cfgwr_brdcast1_seq.sv")
   `include_typ("hqm_iosf_sb_cfgwr_brdcast2_seq.sv")
   `include_typ("hqm_iosf_sb_cfgwr_brdcast3_seq.sv")

   `include_typ("hqm_iosf_sb_memwr_brdcast_seq.sv")
   `include_typ("hqm_iosf_sb_memrd_brdcast1_seq.sv")
   `include_typ("hqm_iosf_sb_memrd_brdcast2_seq.sv")

   `include_typ("hqm_iosf_sb_memrd_brdcast_seq.sv")
   `include_typ("hqm_iosf_sb_memwr_mcast_seq.sv")
   `include_typ("back2back_sb_cfgrd_brdcast_seq.sv")
   `include_typ("back2back_sb_mem_brdcast_seq.sv")

   


  //sideband SAI sequeces
  `include_typ("sai_sb_packet.sv")
  `include_typ("hqm_iosf_sb_cfgrd_sai_seq.sv")
  `include_typ("hqm_iosf_sb_cfgwr_sai_seq.sv")
  `include_typ("hqm_iosf_sb_memrd_sai_seq.sv")
  `include_typ("hqm_iosf_sb_memwr_sai_seq.sv")
  `include_typ("hqm_iosf_sb_npmemwr_sai_seq.sv")
  `include_typ("back2back_sb_cfgrd_sai_seq.sv")
  `include_typ("back2back_sb_cfgwr_sai_seq.sv")
  `include_typ("SAI_sb_cfgrd_csr_seq.sv")
  `include_typ("SAI_sb_cfgwr_csr_seq.sv")
  `include_typ("back2back_sb_memrd_sai_seq.sv")
  `include_typ("back2back_sb_memrd_dbg_seq.sv")
  `include_typ("back2back_sb_memrd_feature_seq.sv")
  `include_typ("back2back_sb_memwr_sai_csr_seq.sv")
  `include_typ("back2back_sb_memwr_sai_dbg_seq.sv")
  `include_typ("back2back_sb_memwr_sai_feature_seq.sv")
   

    //mixed_sequences
      `include_typ("mix_cfg_mem_seq.sv")
      `include_typ("mix_mem_cfg_seq.sv")

    //unsupported transaction with invalid_sai
       `include_typ("hqm_iosf_prim_msg_sai_seq.sv")
       `include_typ("back2back_posted_msg_sai_seq.sv")  
       `include_typ("back2back_cfg1_sai_seq.sv")
       `include_typ("back2back_unsupport_memwr_sai_seq.sv")
       `include_typ("back2back_unsupport_memrd_sai_seq.sv")

    // setid_sequence
  `include_typ("hqm_iosf_sb_setid_seq.sv")  
