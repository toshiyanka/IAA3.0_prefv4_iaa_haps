// File output was printed on: Saturday, January 19, 2013 2:59:29 PM
// Chassis TAP Tool version: 0.6.0.0
//----------------------------------------------------------------------
parameter NUMBER_OF_HIER  = 0;
parameter NUMBER_OF_STAPS = 0;
parameter NUMBER_OF_TERTIARY_PORTS = 0;
