//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// AW_pipe_rate_limit
//
// This module is responsible for gating the input valid to a pipeline based on the status of the
// pipeline's valid bits to limit the rate things are input to the pipeline.  Setting a CFG input bit
// requires that the associated pipeline valid be off before the input valid will be passed to the
// output valid.  Setting the CFG input to all ones ensures the pipeline must be completely empty before
// the input valid is propagated to the output.
//
// The following parameters are supported:
//
//  WIDTH       Width of the valid signal to gate
//  DEPTH       Depth of the pipeline to rate limit
//
//-----------------------------------------------------------------------------------------------------

module hqm_AW_pipe_rate_limit

     import hqm_AW_pkg::*;
#(
     parameter WIDTH = 1
    ,parameter DEPTH = 1
) (
     input  logic   [DEPTH-1:0] cfg
    ,input  logic   [DEPTH-1:0] pipe_v

    ,input  logic   [WIDTH-1:0] v_in

    ,output logic   [WIDTH-1:0] v_out
);

//-----------------------------------------------------------------------------------------------------

logic   allow_valid;

assign allow_valid = &{1'b1, ~(cfg & pipe_v)};

assign v_out = v_in & {WIDTH{allow_valid}};

endmodule // AW_pipe_rate_limit

