// File output was printed on: Thursday, March 21, 2013 4:21:02 PM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
// ENUM DECLARATIONS
//------------------------------------------------------------------------
typedef enum int {
   IPLEVEL_STAP   =  'd0,
   NOTAP          =  'hFFFF_FFFF
} Tap_t;


