`define I_HQM_CONTROL_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_CONTROL `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general
`define I_HQM_CONTROL_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_CONTROL `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general
`define I_HQM_CONTROL_MASTER_CORE_CONTROL_TARGET_CFG_MASTER_CORE_CONTROL_CSR_CONTROL `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general
`define I_HQM_CONTROL_CREDIT_HIST_00_TARGET_CFG_CREDIT_HIST_00_CSR_CONTROL `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00
`define I_HQM_CONTROL_CREDIT_HIST_01_TARGET_CFG_CREDIT_HIST_01_CSR_CONTROL `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_01
`define I_HQM_CONTROL_CREDIT_HIST_02_TARGET_CFG_CREDIT_HIST_02_CSR_CONTROL `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02
`define I_HQM_CONTROL_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_CONTROL `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_control_general
`define I_HQM_CONTROL_LIST_SEL_0_TARGET_CFG_LIST_SEL_0_CSR_CONTROL `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0
`define I_HQM_CONTROL_LIST_SEL_1_TARGET_CFG_LIST_SEL_1_CSR_CONTROL `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1
`define I_HQM_CONTROL_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_CONTROL `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_control_general
`define I_HQM_CONTROL_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_CONTROL `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_control_general
`define I_HQM_CONTROL_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_CONTROL `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_control_general_0
`define I_HQM_STATUS_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_STATUS `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status
`define I_HQM_STATUS_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_STATUS `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status
`define I_HQM_STATUS_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_STATUS `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status
`define I_HQM_STATUS_LIST_SEL_INTERFACE_TARGET_CFG_LIST_SEL_INTERFACE_CSR_STATUS `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status
`define I_HQM_STATUS_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_STATUS `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status
`define I_HQM_STATUS_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_STATUS `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status
`define I_HQM_STATUS_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_STATUS `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status
`define I_HQM_STATUS_MASTER_CORE_DIAGNOSTIC_1_TARGET_CFG_MASTER_CORE_DIAGNOSTIC_1_CSR_STATUS `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1
`define I_HQM_STATUS_LIST_SEL_DIAGNOSTIC_0_TARGET_CFG_LIST_SEL_DIAGNOSTIC_0_CSR_STATUS `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0
`define INT_CONTROL_AQED_PIPE_CHICKEN_SIM `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[0:0]
`define INT_CONTROL_AQED_PIPE_CHICKEN_50 `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[1:1]
`define INT_CONTROL_AQED_PIPE_FID_DECREMENT `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[4:4]
`define INT_CONTROL_AQED_PIPE_FID_SIM `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[5:5]
`define INT_CONTROL_AQED_PIPE_AQED_LSP_STOP_ATQATM `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[21:8]
`define INT_CONTROL_AQED_PIPE_AQED_CHICKEN_ONEPRI `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_control_general.internal_f[30:30]
`define INT_CONTROL_ATM_PIPE_CHICKEN_SIM `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[0:0]
`define INT_CONTROL_ATM_PIPE_CHICKEN_50 `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[1:1]
`define INT_CONTROL_ATM_PIPE_CHICKEN_33 `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[2:2]
`define INT_CONTROL_ATM_PIPE_CHICKEN_25 `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[3:3]
`define INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQSTALL `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[7:7]
`define INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQ_AFULL_HP_MODE `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[8:8]
`define INT_CONTROL_ATM_PIPE_CHICKEN_EN_ALWAYSBLAST `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[9:9]
`define INT_CONTROL_ATM_PIPE_CHICKEN_EN_ENQBLOCKRLST `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[10:10]
`define INT_CONTROL_ATM_PIPE_CHICKEN_MAX_ENQSTALL `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_control_general.internal_f[14:12]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_IDLE_DLY `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[15:0]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_PSLVERR_TIMEOUT `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[23:23]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_RDATA `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[24:24]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_ADDR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[25:25]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_WDATA `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[26:26]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_RING_PAR_CK `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[27:27]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_ALARMS `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[28:28]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_PM_ALLOW_ING_DROP `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[29:29]
`define INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_UNIT_IDLE `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[30:30]
`define INT_CONTROL_MASTER_CORE_CONTROL_IGNORE_PIPE_BUSY `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_control_general.internal_f[31:31]
`define INT_CONTROL_CREDIT_HIST_00_OUTBOUND_HCW_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[4:0]
`define INT_CONTROL_CREDIT_HIST_00_LSP_AP_CMP_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[9:5]
`define INT_CONTROL_CREDIT_HIST_00_LSP_TOK_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[14:10]
`define INT_CONTROL_CREDIT_HIST_00_ROP_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[19:15]
`define INT_CONTROL_CREDIT_HIST_00_EGRESS_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[23:20]
`define INT_CONTROL_CREDIT_HIST_00_QED_TO_CQ_PIPE_CREDIT_HWM `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[27:24]
`define INT_CONTROL_CREDIT_HIST_00_EGRESS_LSP_TOKEN_PIPE_CREDIT `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_00.internal_f[30:28]
`define INT_CONTROL_CREDIT_HIST_01_CHP_BLK_DUAL_ISSUE `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_01.internal_f[0:0]
`define INT_CONTROL_CREDIT_HIST_01_INCLUDE_CWDI_TIMER_IDLE_EN `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_01.internal_f[1:1]
`define INT_CONTROL_CREDIT_HIST_01_CIAL_CLOCK_GATE_CONTROL `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_01.internal_f[3:3]
`define INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[0:0]
`define INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[1:1]
`define INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[2:2]
`define INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[3:3]
`define INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[4:4]
`define INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[5:5]
`define INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[6:6]
`define INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[7:7]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[8:8]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[9:9]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[10:10]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[11:11]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[12:12]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[13:13]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[14:14]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[15:15]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[16:16]
`define INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[17:17]
`define INT_CONTROL_CREDIT_HIST_02_ENGPIPE_FLID_PARITY_ERROR_INJECTION `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[18:18]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_0 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[19:19]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_1 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[20:20]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_2 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[21:21]
`define INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_3 `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[22:22]
`define INT_CONTROL_CREDIT_HIST_02_CONTROL `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_credit_hist_pipe_register_pfcsr.i_hqm_chp_target_cfg_control_general_02.internal_f[31:23]
`define INT_CONTROL_DIR_PIPE_CHICKEN_SIM `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_control_general.internal_f[0:0]
`define INT_CONTROL_DIR_PIPE_CHICKEN_50 `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_control_general.internal_f[1:1]
`define INT_CONTROL_LIST_SEL_0_DISAB_ATQ_EMPTY_ARB `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[0:0]
`define INT_CONTROL_LIST_SEL_0_INC_TOK_UNIT_IDLE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[1:1]
`define INT_CONTROL_LIST_SEL_0_DISAB_RLIST_PRI `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[2:2]
`define INT_CONTROL_LIST_SEL_0_INC_CMP_UNIT_IDLE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[3:3]
`define INT_CONTROL_LIST_SEL_0_ENAB_IF_THRESH `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[4:4]
`define INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[6:6]
`define INT_CONTROL_LIST_SEL_0_DIR_HALF_BW `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[7:7]
`define INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OUT `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[8:8]
`define INT_CONTROL_LIST_SEL_0_DIR_DISAB_MULTI `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[9:9]
`define INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[10:10]
`define INT_CONTROL_LIST_SEL_0_ATQ_HALF_BW `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[11:11]
`define INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OUT `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[12:12]
`define INT_CONTROL_LIST_SEL_0_ATQ_DISAB_MULTI `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[13:13]
`define INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[14:14]
`define INT_CONTROL_LIST_SEL_0_DIRRPL_HALF_BW `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[15:15]
`define INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OUT `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[16:16]
`define INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[17:17]
`define INT_CONTROL_LIST_SEL_0_LBRPL_HALF_BW `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[18:18]
`define INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OUT `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[19:19]
`define INT_CONTROL_LIST_SEL_0_LDB_SINGLE_OP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[20:20]
`define INT_CONTROL_LIST_SEL_0_LDB_HALF_BW `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[21:21]
`define INT_CONTROL_LIST_SEL_0_LDB_DISAB_MULTI `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[22:22]
`define INT_CONTROL_LIST_SEL_0_ATM_SINGLE_SCH `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[23:23]
`define INT_CONTROL_LIST_SEL_0_ATM_SINGLE_CMP `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[24:24]
`define INT_CONTROL_LIST_SEL_0_LDB_CE_TOG_ARB `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[25:25]
`define INT_CONTROL_LIST_SEL_0_SMON0_VALID_SEL `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[28:27]
`define INT_CONTROL_LIST_SEL_0_SMON0_VALUE_SEL `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[29:29]
`define INT_CONTROL_LIST_SEL_0_SMON0_COMPARE_SEL `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_0.internal_f[31:30]
`define INT_CONTROL_LIST_SEL_1_QE_WT_FRC `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[1:0]
`define INT_CONTROL_LIST_SEL_1_QE_WT_FRCV `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[2:2]
`define INT_CONTROL_LIST_SEL_1_QE_WT_BLK `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[3:3]
`define INT_CONTROL_LIST_SEL_1_QED_DEQ_HIPRI_WM `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[8:4]
`define INT_CONTROL_LIST_SEL_1_DIS_WU_RES_CHK `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[9:9]
`define INT_CONTROL_LIST_SEL_1_AQED_DEQ_HIPRI_WM `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_control_general_1.internal_f[16:12]
`define INT_CONTROL_NALB_PIPE_CHICKEN_SIM `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_control_general.internal_f[0:0]
`define INT_CONTROL_NALB_PIPE_CHICKEN_50 `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_control_general.internal_f[1:1]
`define INT_CONTROL_QED_PIPE_REG_CHICKEN_SIM `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_control_general.internal_f[0:0]
`define INT_CONTROL_QED_PIPE_REG_CHICKEN_STRICT `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_control_general.internal_f[1:1]
`define INT_CONTROL_REORDER_PIPE_UNIT_SINGLE_STEP_MODE `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_control_general_0.internal_f[0:0]
`define INT_CONTROL_REORDER_PIPE_RR_EN `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_control_general_0.internal_f[1:1]
`define INT_CONTROL_REORDER_PIPE_RSZV0 `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_control_general_0.internal_f[31:2]
`define INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[1:0]
`define INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[5:4]
`define INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[9:8]
`define INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[13:12]
`define INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[17:16]
`define INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_DEPTH `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[21:20]
`define INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_READY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[22:22]
`define INT_STATUS_AQED_PIPE_FIFO_LSP_AQED_CMP_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[24:24]
`define INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_FID_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[25:25]
`define INT_STATUS_AQED_PIPE_FIFO_AQED_CHP_SCH_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[26:26]
`define INT_STATUS_AQED_PIPE_FIFO_AP_AQED_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[27:27]
`define INT_STATUS_AQED_PIPE_FIFO_AQED_AP_ENQ_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[28:28]
`define INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[29:29]
`define INT_STATUS_AQED_PIPE_FIFO_FREELIST_RETURN_EMPTY `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[30:30]
`define INT_STATUS_AQED_PIPE_AQED_CLK_IDLE `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_aqed_pipe_register_pfcsr.i_hqm_aqed_target_cfg_interface_status.internal_f[31:31]
`define INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[1:0]
`define INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_READY_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[5:4]
`define INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_READY `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[9:8]
`define INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_READY `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[13:12]
`define INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_READY `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_DEPTH `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[17:16]
`define INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_READY `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_ATM_PIPE_ATM_CLK_IDLE `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_ap_pipe_register_pfcsr.i_hqm_ap_target_cfg_interface_status.internal_f[31:31]
`define INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[1:0]
`define INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_DIR_PIPE_DP_DQED_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[5:4]
`define INT_STATUS_DIR_PIPE_DP_DQED_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[9:8]
`define INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[13:12]
`define INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[17:16]
`define INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[21:20]
`define INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[22:22]
`define INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_DEPTH `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[25:24]
`define INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_READY `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[26:26]
`define INT_STATUS_DIR_PIPE_INT_IDLE_B `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.i_hqm_dp_pipe_register_pfcsr.i_hqm_dp_target_cfg_interface_status.internal_f[31:31]
`define INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[0:0]
`define INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[1:1]
`define INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[3:3]
`define INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[4:4]
`define INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[5:5]
`define INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[7:7]
`define INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[8:8]
`define INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[9:9]
`define INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[11:11]
`define INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[12:12]
`define INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[13:13]
`define INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[15:15]
`define INT_STATUS_LIST_SEL_INTERFACE_INT_SER_CLOCK_NOT_IDLE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[16:16]
`define INT_STATUS_LIST_SEL_INTERFACE_AQED_CLOCK_NOT_IDLE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[17:17]
`define INT_STATUS_LIST_SEL_INTERFACE_AP_CLOCK_NOT_IDLE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[20:20]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[21:21]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[22:22]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[23:23]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[24:24]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[25:25]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[26:26]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[27:27]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[28:28]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[29:29]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[30:30]
`define INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_NOT_RDY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_interface_status.internal_f[31:31]
`define INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[1:0]
`define INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[5:4]
`define INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[9:8]
`define INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[13:12]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[17:16]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[21:20]
`define INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[22:22]
`define INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_DEPTH `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[25:24]
`define INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_READY `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[26:26]
`define INT_STATUS_NALB_PIPE_INT_IDLE_B `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.i_hqm_nalb_pipe_register_pfcsr.i_hqm_nalb_target_cfg_interface_status.internal_f[31:31]
`define INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[0:0]
`define INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[1:1]
`define INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[2:2]
`define INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[3:3]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[4:4]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[5:5]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[6:6]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[7:7]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[8:8]
`define INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[9:9]
`define INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[10:10]
`define INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[11:11]
`define INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[12:12]
`define INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[13:13]
`define INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[14:14]
`define INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[15:15]
`define INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[16:16]
`define INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[17:17]
`define INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[18:18]
`define INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[19:19]
`define INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[20:20]
`define INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[21:21]
`define INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[22:22]
`define INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[23:23]
`define INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[24:24]
`define INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[25:25]
`define INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[26:26]
`define INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[27:27]
`define INT_STATUS_QED_PIPE_REG_ROP_QED_ENQ_READY `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[28:28]
`define INT_STATUS_QED_PIPE_REG_ROP_QED_DQED_ENQ_V `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[29:29]
`define INT_STATUS_QED_PIPE_REG_INT_IDLE `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_qed_pipe_register_pfcsr.i_hqm_qed_target_cfg_interface_status.internal_f[30:30]
`define INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[0:0]
`define INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[1:1]
`define INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[2:2]
`define INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[3:3]
`define INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[4:4]
`define INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[5:5]
`define INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[6:6]
`define INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[7:7]
`define INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[8:8]
`define INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[9:9]
`define INT_STATUS_REORDER_PIPE_ROP_QED_ENQ_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[10:10]
`define INT_STATUS_REORDER_PIPE_ROP_QED_DQED_ENQ_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[11:11]
`define INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_READY `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[12:12]
`define INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_V `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[13:13]
`define INT_STATUS_REORDER_PIPE_INT_IDLE_B `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_register_pfcsr.i_hqm_rop_target_cfg_interface_status.status[31:31]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_TIMEOUT_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[0:0]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQRSP_UNSOL_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[1:1]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_PROTOCOL_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[2:2]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLV_PAR_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[3:3]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_PAR_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[4:4]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_DROP_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[16:16]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_UP_MISS_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[17:17]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[18:18]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_ACCESS_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[19:19]
`define INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_TIMEOUT_ERR `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_register_prim.i_hqm_mstr_target_cfg_diagnostic_status_1.internal_f[20:20]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[0:0]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_BLAST `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[1:1]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[2:2]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_BLAST `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[3:3]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[4:4]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_BLAST `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[5:5]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST_CHKV `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[6:6]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[7:7]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_QID_DIS `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[8:8]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_BUSY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[9:9]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_NO_SPACE `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[10:10]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_DIR_TOK_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[11:11]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_ACT `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[12:12]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AP_LSP_ATM_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[13:13]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_TOK_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[14:14]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CMP_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[15:15]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS0 `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[16:16]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS1 `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[17:17]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS2 `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[18:18]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS3 `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[19:19]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_STOP_ATQATM `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[23:23]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_SN_FCERR_RPTD `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[24:24]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_EMPTY `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[25:25]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATM_IF_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[26:26]
`define INT_STATUS_LIST_SEL_DIAGNOSTIC_0_TOT_IF_V `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_pipe_register_pfcsr.i_hqm_lsp_target_cfg_diagnostic_status_0.status[27:27]
