# Text_Tag % Vendor Intel % Product c73p4rfshdxrom % Techno P1273.1 % Tag_Spec 1.0 % ECCN US_3E002 % Signature 7d6e731266319034db308e638d9f2e55b99d318d % Version r1.0.0_m1.18 % _View_Id lef % Date_Time 20160303_050306 
################################################################################
# Intel Confidential                                                           #
################################################################################
# Copyright 2014 Intel Corporation.                                            #
# The information contained herein is the proprietary and confidential         #
# information of Intel or its licensors, and is supplied subject to, and       #
# may be used only in accordance with, previously executed agreements          #
# with Intel ,                                                                 #
# EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING:                                #
# (1) ALL MATERIALS FURNISHED BY INTEL HEREUNDER ARE PROVIDED "AS IS"          #
#      WITHOUT WARRANTY OF ANY KIND;                                           #
# (2) INTEL SPECIFICALLY DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS    #
#      FOR A PARTICULAR PURPOSE OR MERCHANTABILITY; AND                        #
# (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF SUBSTITUTES,    #
#      LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR                           #
#      FOR ANY OTHER SPECIAL, CONSEQUENTIAL OR INCIDENTAL DAMAGES,             #
#      HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY, CONTRACT,               #
#      TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                        #
################################################################################
################################################################################
#                                                                              #
# Vendor: Intel                                                                #
# Product: c73p4rfshdxrom                                                      #
# Version: r1.0.0_m1.18                                                        #
# Technology: p1273.1                                                          #
# Celltype: IP                                                                 #
# IP_Owner: Intel DTS CMO                                                      #
# Date_Time: YYYYMMDD_HHMMSS                                                   #
#                                                                              #
################################################################################
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

SITE c73p1rfshdxrom2048x16hb4img100
  SIZE 75.432 by 29.526 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END c73p1rfshdxrom2048x16hb4img100


MACRO c73p1rfshdxrom2048x16hb4img100
     FOREIGN c73p1rfshdxrom2048x16hb4img100 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 75.432 by 29.526 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE c73p1rfshdxrom2048x16hb4img100 ;
     PIN iar[10]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 10.932 0.308 10.964 ;
          END
     END iar[10]
     PIN iar[0]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 11.674 0.308 11.706 ;
          END
     END iar[0]
     PIN iar[1]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 12.472 0.308 12.504 ;
          END
     END iar[1]
     PIN iar[2]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 13.088 0.308 13.12 ;
          END
     END iar[2]
     PIN iar[4]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 13.774 0.308 13.806 ;
          END
     END iar[4]
     PIN iar[3]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 14.404 0.308 14.436 ;
          END
     END iar[3]
     PIN iar[7]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 15.72 0.308 15.752 ;
          END
     END iar[7]
     PIN iar[6]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 16.406 0.308 16.438 ;
          END
     END iar[6]
     PIN iar[5]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 16.966 0.308 16.998 ;
          END
     END iar[5]
     PIN iar[9]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 17.764 0.308 17.796 ;
          END
     END iar[9]
     PIN iar[8]
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 18.282 0.308 18.314 ;
          END
     END iar[8]
     PIN iren
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 15.146 0.308 15.178 ;
          END
     END iren
     PIN ickr
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 14.922 0.308 14.954 ;
          END
     END ickr
     PIN ipwreninb
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 28.544 0.308 28.576 ;
          END
     END ipwreninb
     PIN opwrenoutb
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 0.726 0.308 0.758 ;
          END
     END opwrenoutb
     PIN odout[0]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 0.95 0.308 0.982 ;
          END
     END odout[0]
     PIN odout[1]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 2.21 0.308 2.242 ;
          END
     END odout[1]
     PIN odout[2]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 3.456 0.308 3.488 ;
          END
     END odout[2]
     PIN odout[3]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 4.716 0.308 4.748 ;
          END
     END odout[3]
     PIN odout[4]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 5.85 0.308 5.882 ;
          END
     END odout[4]
     PIN odout[5]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 7.222 0.308 7.254 ;
          END
     END odout[5]
     PIN odout[6]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 8.482 0.308 8.514 ;
          END
     END odout[6]
     PIN odout[7]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 9.728 0.308 9.76 ;
          END
     END odout[7]
     PIN odout[8]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 19.08 0.308 19.112 ;
          END
     END odout[8]
     PIN odout[9]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 20.452 0.308 20.484 ;
          END
     END odout[9]
     PIN odout[10]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 21.698 0.308 21.73 ;
          END
     END odout[10]
     PIN odout[11]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 22.846 0.308 22.878 ;
          END
     END odout[11]
     PIN odout[12]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 24.092 0.308 24.124 ;
          END
     END odout[12]
     PIN odout[13]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 25.352 0.308 25.384 ;
          END
     END odout[13]
     PIN odout[14]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 26.836 0.308 26.868 ;
          END
     END odout[14]
     PIN odout[15]
     DIRECTION output ;
          PORT
               LAYER m4 ;
               RECT 0 28.194 0.308 28.226 ;
          END
     END odout[15]
     PIN vccd_1p0
     SHAPE ABUTMENT ;
     USE   POWER ;
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0.42 0.654 74.894 0.7 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.852 14.274 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.064 2.832 1.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.34 13.678 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.474 13.354 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.722 14 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.914 74.894 1.96 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.16 13.678 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.294 13.354 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.542 14 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.664 74.894 10.71 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.884 74.894 10.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.088 74.894 11.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.292 74.894 11.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.49 6.19 11.536 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.56 74.894 11.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.688 74.894 11.734 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.322 74.894 12.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.59 74.894 12.644 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.006 74.894 13.046 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.75 74.894 13.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.246 74.894 14.286 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.114 74.894 15.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.486 74.894 15.526 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.982 74.894 16.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.478 74.894 16.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.85 74.894 16.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.098 74.894 17.138 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.462 74.894 17.518 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.606 74.894 17.652 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.746 74.894 17.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.896 74.894 17.942 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.036 74.894 18.092 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.196 74.894 18.242 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.33 74.894 18.384 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.478 74.894 18.524 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.612 74.894 18.652 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.798 74.894 18.844 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.996 14.274 19.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.208 2.832 19.292 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.484 13.678 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.618 13.354 19.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.866 14 19.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.112 14.274 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.324 2.832 2.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.6 13.678 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.734 13.354 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.982 14 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.058 74.894 20.104 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.256 14.274 20.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.468 2.832 20.552 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.744 13.678 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.878 13.354 20.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.126 14 21.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.318 74.894 21.364 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.516 14.274 21.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.728 2.832 21.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.004 13.678 22.05 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.138 13.354 22.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.386 14 22.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.578 74.894 22.624 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.776 14.274 22.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.988 2.832 23.072 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.264 13.678 23.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.398 13.354 23.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.646 14 23.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.838 74.894 23.884 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.036 14.274 24.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.248 2.832 24.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.524 13.678 24.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.658 13.354 24.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.906 14 24.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.098 74.894 25.144 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.296 14.274 25.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.508 2.832 25.592 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.784 13.678 25.83 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.918 13.354 25.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.166 14 26.212 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.358 74.894 26.404 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.556 14.274 26.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.768 2.832 26.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.044 13.678 27.09 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.178 13.354 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.426 14 27.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.618 74.894 27.664 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.816 14.274 27.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.028 2.832 28.112 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.304 13.678 28.35 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.438 13.354 28.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.686 14 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.174 74.894 3.22 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.372 14.274 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.584 2.832 3.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.86 13.678 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.994 13.354 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.242 14 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.434 74.894 4.48 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.632 14.274 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.844 2.832 4.928 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.12 13.678 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.254 13.354 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.502 14 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.694 74.894 5.74 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.892 14.274 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.104 2.832 6.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.38 13.678 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.514 13.354 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.762 14 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.954 74.894 7 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.152 14.274 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.364 2.832 7.448 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.64 13.678 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.774 13.354 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.022 14 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.214 74.894 8.26 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.412 14.274 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.624 2.832 8.708 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.9 13.678 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.034 13.354 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.282 14 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.474 74.894 9.52 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.672 14.274 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.884 2.832 9.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 1.722 31.052 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 10.542 31.052 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 19.866 31.052 19.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 2.982 31.052 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 21.126 31.052 21.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 22.386 31.052 22.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 23.646 31.052 23.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 24.906 31.052 24.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 26.166 31.052 26.212 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 27.426 31.052 27.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 28.686 31.052 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 4.242 31.052 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 5.502 31.052 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 6.762 31.052 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 8.022 31.052 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 14.32 9.282 31.052 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 0.852 31.326 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 18.996 31.326 19.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 2.112 31.326 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 20.256 31.326 20.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 21.516 31.326 21.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 22.776 31.326 22.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 24.036 31.326 24.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 25.296 31.326 25.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 26.556 31.326 26.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 27.816 31.326 27.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 3.372 31.326 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 4.632 31.326 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 5.892 31.326 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 7.152 31.326 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 8.412 31.326 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 15.73 9.672 31.326 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 1.474 30.406 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 10.294 30.406 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 19.618 30.406 19.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 2.734 30.406 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 20.878 30.406 20.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 22.138 30.406 22.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 23.398 30.406 23.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 24.658 30.406 24.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 25.918 30.406 25.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 27.178 30.406 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 28.438 30.406 28.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 3.994 30.406 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 5.254 30.406 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 6.514 30.406 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 7.774 30.406 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.219 9.034 30.406 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 1.34 30.73 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 10.16 30.73 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 19.484 30.73 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 2.6 30.73 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 20.744 30.73 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 22.004 30.73 22.05 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 23.264 30.73 23.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 24.524 30.73 24.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 25.784 30.73 25.83 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 27.044 30.73 27.09 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 28.304 30.73 28.35 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 3.86 30.73 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 5.12 30.73 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 6.38 30.73 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 7.64 30.73 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.638 8.9 30.73 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 1.722 48.104 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 10.542 48.104 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 19.866 48.104 19.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 2.982 48.104 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 21.126 48.104 21.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 22.386 48.104 22.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 23.646 48.104 23.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 24.906 48.104 24.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 26.166 48.104 26.212 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 27.426 48.104 27.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 28.686 48.104 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 4.242 48.104 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 5.502 48.104 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 6.762 48.104 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 8.022 48.104 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 31.372 9.282 48.104 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 0.852 48.378 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 18.996 48.378 19.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 2.112 48.378 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 20.256 48.378 20.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 21.516 48.378 21.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 22.776 48.378 22.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 24.036 48.378 24.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 25.296 48.378 25.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 26.556 48.378 26.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 27.816 48.378 27.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 3.372 48.378 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 4.632 48.378 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 5.892 48.378 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 7.152 48.378 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 8.412 48.378 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.782 9.672 48.378 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 1.474 47.458 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 10.294 47.458 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 19.618 47.458 19.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 2.734 47.458 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 20.878 47.458 20.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 22.138 47.458 22.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 23.398 47.458 23.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 24.658 47.458 24.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 25.918 47.458 25.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 27.178 47.458 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 28.438 47.458 28.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 3.994 47.458 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 5.254 47.458 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 6.514 47.458 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 7.774 47.458 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.271 9.034 47.458 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 1.34 47.782 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 10.16 47.782 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 19.484 47.782 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 2.6 47.782 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 20.744 47.782 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 22.004 47.782 22.05 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 23.264 47.782 23.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 24.524 47.782 24.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 25.784 47.782 25.83 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 27.044 47.782 27.09 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 28.304 47.782 28.35 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 3.86 47.782 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 5.12 47.782 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 6.38 47.782 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 7.64 47.782 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.69 8.9 47.782 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 1.722 65.156 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 10.542 65.156 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 19.866 65.156 19.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 2.982 65.156 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 21.126 65.156 21.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 22.386 65.156 22.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 23.646 65.156 23.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 24.906 65.156 24.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 26.166 65.156 26.212 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 27.426 65.156 27.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 28.686 65.156 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 4.242 65.156 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 5.502 65.156 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 6.762 65.156 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 8.022 65.156 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.424 9.282 65.156 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 0.852 65.43 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 18.996 65.43 19.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 2.112 65.43 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 20.256 65.43 20.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 21.516 65.43 21.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 22.776 65.43 22.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 24.036 65.43 24.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 25.296 65.43 25.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 26.556 65.43 26.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 27.816 65.43 27.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 3.372 65.43 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 4.632 65.43 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 5.892 65.43 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 7.152 65.43 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 8.412 65.43 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.834 9.672 65.43 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 1.474 64.51 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 10.294 64.51 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 19.618 64.51 19.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 2.734 64.51 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 20.878 64.51 20.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 22.138 64.51 22.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 23.398 64.51 23.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 24.658 64.51 24.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 25.918 64.51 25.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 27.178 64.51 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 28.438 64.51 28.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 3.994 64.51 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 5.254 64.51 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 6.514 64.51 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 7.774 64.51 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.323 9.034 64.51 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 1.34 64.834 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 10.16 64.834 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 19.484 64.834 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 2.6 64.834 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 20.744 64.834 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 22.004 64.834 22.05 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 23.264 64.834 23.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 24.524 64.834 24.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 25.784 64.834 25.83 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 27.044 64.834 27.09 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 28.304 64.834 28.35 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 3.86 64.834 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 5.12 64.834 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 6.38 64.834 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 7.64 64.834 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.742 8.9 64.834 8.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 1.722 74.894 1.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 10.542 74.894 10.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 19.866 74.894 19.912 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 2.982 74.894 3.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 21.126 74.894 21.172 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 22.386 74.894 22.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 23.646 74.894 23.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 24.906 74.894 24.952 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 26.166 74.894 26.212 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 27.426 74.894 27.472 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 28.686 74.894 28.732 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 4.242 74.894 4.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 5.502 74.894 5.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 6.762 74.894 6.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 8.022 74.894 8.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 65.476 9.282 74.894 9.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 0.852 74.894 0.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 18.996 74.894 19.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 2.112 74.894 2.152 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 20.256 74.894 20.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 21.516 74.894 21.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 22.776 74.894 22.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 24.036 74.894 24.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 25.296 74.894 25.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 26.556 74.894 26.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 27.816 74.894 27.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 3.372 74.894 3.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 4.632 74.894 4.672 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 5.892 74.894 5.932 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 7.152 74.894 7.192 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 8.412 74.894 8.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 66.886 9.672 74.894 9.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 1.474 74.894 1.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 10.294 74.894 10.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 19.618 74.894 19.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 2.734 74.894 2.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 20.878 74.894 20.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 22.138 74.894 22.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 23.398 74.894 23.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 24.658 74.894 24.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 25.918 74.894 25.958 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 27.178 74.894 27.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 28.438 74.894 28.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 3.994 74.894 4.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 5.254 74.894 5.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 6.514 74.894 6.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 7.774 74.894 7.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.375 9.034 74.894 9.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 1.34 74.894 1.386 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 10.16 74.894 10.206 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 19.484 74.894 19.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 2.6 74.894 2.646 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 20.744 74.894 20.79 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 22.004 74.894 22.05 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 23.264 74.894 23.31 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 24.524 74.894 24.57 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 25.784 74.894 25.83 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 27.044 74.894 27.09 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 28.304 74.894 28.35 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 3.86 74.894 3.906 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 5.12 74.894 5.166 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 6.38 74.894 6.426 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 7.64 74.894 7.686 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.794 8.9 74.894 8.946 ;
          END
     END vccd_1p0
     PIN vss
     SHAPE ABUTMENT ;
     USE   GROUND ;
     DIRECTION input ;
          PORT
               LAYER m4 ;
               RECT 0 0.67 0.308 0.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 1.006 0.308 1.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 10.876 0.308 10.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 11.618 0.308 11.65 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 12.528 0.308 12.56 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 13.032 0.302 13.064 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 13.83 0.308 13.862 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 14.348 0.308 14.38 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 14.978 0.308 15.01 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 15.202 0.308 15.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 15.776 0.308 15.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 16.462 0.308 16.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 17.022 0.308 17.054 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 17.82 0.308 17.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 18.338 0.308 18.37 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 19.136 0.308 19.168 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 2.154 0.308 2.186 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 20.508 0.308 20.54 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 21.754 0.308 21.786 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 22.902 0.308 22.934 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 24.148 0.308 24.18 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 25.408 0.308 25.44 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 26.892 0.222 26.924 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 28.25 0.222 28.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 28.488 0.308 28.52 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 3.4 0.308 3.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 4.66 0.308 4.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 5.794 0.308 5.826 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 7.166 0.308 7.198 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 8.426 0.308 8.458 ;
          END
          PORT
               LAYER m4 ;
               RECT 0 9.672 0.308 9.704 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.584 14.184 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.788 74.894 0.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 0.986 74.894 1.04 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.262 74.894 1.316 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.538 74.894 1.578 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 1.844 14.184 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.082 74.894 10.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.358 74.894 10.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.814 74.894 10.86 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 10.954 74.894 11 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.426 74.894 11.466 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 11.818 74.894 11.864 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.068 74.894 12.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.446 74.894 12.486 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 12.668 74.894 12.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.13 74.894 13.17 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.378 74.894 13.418 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.626 74.894 13.666 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 13.998 74.894 14.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.494 74.894 14.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.742 74.894 14.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 14.99 74.894 15.03 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.362 74.894 15.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 15.858 74.894 15.898 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.106 74.894 16.146 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.354 74.894 16.394 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 16.602 74.894 16.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.372 74.894 17.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 17.676 74.894 17.722 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.408 74.894 18.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.728 14.184 18.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 18.932 74.894 18.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.13 74.894 19.184 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.406 74.894 19.46 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.682 74.894 19.722 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 19.988 14.184 20.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.048 74.894 2.088 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.246 74.894 2.3 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.522 74.894 2.576 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 2.798 74.894 2.838 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.192 74.894 20.232 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.39 74.894 20.444 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.666 74.894 20.72 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 20.942 74.894 20.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.248 14.184 21.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.452 74.894 21.492 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.65 74.894 21.704 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 21.926 74.894 21.98 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.202 74.894 22.242 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.508 14.184 22.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.712 74.894 22.752 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 22.91 74.894 22.964 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.186 74.894 23.24 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.462 74.894 23.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.768 14.184 23.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 23.972 74.894 24.012 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.17 74.894 24.224 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.446 74.894 24.5 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 24.722 74.894 24.762 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.028 14.184 25.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.232 74.894 25.272 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.43 74.894 25.484 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.706 74.894 25.76 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 25.982 74.894 26.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.288 14.184 26.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.492 74.894 26.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.69 74.894 26.744 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 26.966 74.894 27.02 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.242 74.894 27.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.548 14.184 27.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.752 74.894 27.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 27.95 74.894 28.004 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.226 74.894 28.28 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 28.502 74.894 28.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.104 14.184 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.308 74.894 3.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.506 74.894 3.56 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 3.782 74.894 3.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.058 74.894 4.098 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.364 14.184 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.568 74.894 4.608 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 4.766 74.894 4.82 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.042 74.894 5.096 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.318 74.894 5.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.624 14.184 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 5.828 74.894 5.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.026 74.894 6.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.302 74.894 6.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.578 74.894 6.618 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 6.884 14.184 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.088 74.894 7.128 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.286 74.894 7.34 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.562 74.894 7.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 7.838 74.894 7.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.144 14.184 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.348 74.894 8.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.546 74.894 8.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 8.822 74.894 8.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.098 74.894 9.138 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.404 14.184 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.608 74.894 9.648 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.42 9.806 74.894 9.86 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 0.584 31.236 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 1.844 31.236 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 18.728 31.236 18.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 19.988 31.236 20.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 21.248 31.236 21.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 22.508 31.236 22.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 23.768 31.236 23.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 25.028 31.236 25.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 26.288 31.236 26.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 27.548 31.236 27.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 3.104 31.236 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 4.364 31.236 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 5.624 31.236 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 6.884 31.236 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 8.144 31.236 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 16.718 9.404 31.236 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 0.584 48.288 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 1.844 48.288 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 18.728 48.288 18.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 19.988 48.288 20.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 21.248 48.288 21.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 22.508 48.288 22.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 23.768 48.288 23.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 25.028 48.288 25.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 26.288 48.288 26.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 27.548 48.288 27.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 3.104 48.288 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 4.364 48.288 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 5.624 48.288 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 6.884 48.288 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 8.144 48.288 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 33.77 9.404 48.288 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 0.584 65.34 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 1.844 65.34 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 18.728 65.34 18.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 19.988 65.34 20.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 21.248 65.34 21.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 22.508 65.34 22.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 23.768 65.34 23.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 25.028 65.34 25.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 26.288 65.34 26.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 27.548 65.34 27.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 3.104 65.34 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 4.364 65.34 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 5.624 65.34 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 6.884 65.34 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 8.144 65.34 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.822 9.404 65.34 9.45 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 0.584 74.894 0.63 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 1.844 74.894 1.89 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 18.728 74.894 18.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 19.988 74.894 20.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 21.248 74.894 21.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 22.508 74.894 22.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 23.768 74.894 23.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 25.028 74.894 25.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 26.288 74.894 26.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 27.548 74.894 27.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 3.104 74.894 3.15 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 4.364 74.894 4.41 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 5.624 74.894 5.67 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 6.884 74.894 6.93 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 8.144 74.894 8.19 ;
          END
          PORT
               LAYER m4 ;
               RECT 67.874 9.404 74.894 9.45 ;
          END
     END vss
     OBS
          LAYER m0 ;
               POLYGON
                    75.432 29.526 0 29.526 0 0 75.432 0 75.432 29.526 ;
          LAYER m1 ;
               POLYGON
                    75.432 29.526 0 29.526 0 0 75.432 0 75.432 29.526 ;
          LAYER m2 ;
               POLYGON
                    75.432 29.526 0 29.526 0 0 75.432 0 75.432 29.526 ;
          LAYER m3 ;
               POLYGON
                    75.432 29.526 0 29.526 0 0 75.432 0 75.432 29.526 ;
          LAYER m4 ;
               POLYGON
                    75.432 29.526 0 29.526 0 0 75.432 0 75.432 29.526 ;
     END
END c73p1rfshdxrom2048x16hb4img100
END LIBRARY
