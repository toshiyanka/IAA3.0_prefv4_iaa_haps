module hqm_reg_func_cov_groups import hqm_AW_pkg::*, hqm_pkg::*, hqm_core_pkg::*; ();


   
`ifdef HQM_COVER_ON

 covergroup CONTROL_AQED_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_AQED_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_AQED_PIPE_CHICKEN_SIM : coverpoint `INT_CONTROL_AQED_PIPE_CHICKEN_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_AQED_PIPE_CHICKEN_50 : coverpoint `INT_CONTROL_AQED_PIPE_CHICKEN_50   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_AQED_PIPE_FID_DECREMENT : coverpoint `INT_CONTROL_AQED_PIPE_FID_DECREMENT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_AQED_PIPE_FID_SIM : coverpoint `INT_CONTROL_AQED_PIPE_FID_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_AQED_PIPE_AQED_LSP_STOP_ATQATM : coverpoint `INT_CONTROL_AQED_PIPE_AQED_LSP_STOP_ATQATM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_AQED_PIPE_AQED_CHICKEN_ONEPRI : coverpoint `INT_CONTROL_AQED_PIPE_AQED_CHICKEN_ONEPRI   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_ATM_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_ATM_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_SIM : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_50 : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_50   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_33 : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_33   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_25 : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_25   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQSTALL : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQSTALL   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQ_AFULL_HP_MODE : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_DIS_ENQ_AFULL_HP_MODE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_EN_ALWAYSBLAST : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_EN_ALWAYSBLAST   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_EN_ENQBLOCKRLST : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_EN_ENQBLOCKRLST   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_ATM_PIPE_CHICKEN_MAX_ENQSTALL : coverpoint `INT_CONTROL_ATM_PIPE_CHICKEN_MAX_ENQSTALL   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_MASTER_CORE_CONTROL_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_MASTER_CORE_CONTROL_TARGET_CFG_MASTER_CORE_CONTROL_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_MASTER_CORE_CONTROL HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_IDLE_DLY : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_IDLE_DLY   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_PSLVERR_TIMEOUT : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_PSLVERR_TIMEOUT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_RDATA : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_RDATA   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_ADDR : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_ADDR   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_WDATA : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_INJ_PAR_ERR_WDATA   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_RING_PAR_CK : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_DISABLE_RING_PAR_CK   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_ALARMS : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_ALARMS   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_PM_ALLOW_ING_DROP : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_PM_ALLOW_ING_DROP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_UNIT_IDLE : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_CFG_ENABLE_UNIT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_MASTER_CORE_CONTROL_IGNORE_PIPE_BUSY : coverpoint `INT_CONTROL_MASTER_CORE_CONTROL_IGNORE_PIPE_BUSY   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_CREDIT_HIST_00_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_CREDIT_HIST_00_TARGET_CFG_CREDIT_HIST_00_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_CREDIT_HIST_00 HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_CREDIT_HIST_00_OUTBOUND_HCW_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_OUTBOUND_HCW_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_LSP_AP_CMP_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_LSP_AP_CMP_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_LSP_TOK_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_LSP_TOK_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_ROP_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_ROP_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_EGRESS_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_EGRESS_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_QED_TO_CQ_PIPE_CREDIT_HWM : coverpoint `INT_CONTROL_CREDIT_HIST_00_QED_TO_CQ_PIPE_CREDIT_HWM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_00_EGRESS_LSP_TOKEN_PIPE_CREDIT : coverpoint `INT_CONTROL_CREDIT_HIST_00_EGRESS_LSP_TOKEN_PIPE_CREDIT   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_CREDIT_HIST_01_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_CREDIT_HIST_01_TARGET_CFG_CREDIT_HIST_01_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_CREDIT_HIST_01 HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_CREDIT_HIST_01_CHP_BLK_DUAL_ISSUE : coverpoint `INT_CONTROL_CREDIT_HIST_01_CHP_BLK_DUAL_ISSUE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_01_INCLUDE_CWDI_TIMER_IDLE_EN : coverpoint `INT_CONTROL_CREDIT_HIST_01_INCLUDE_CWDI_TIMER_IDLE_EN   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_01_CIAL_CLOCK_GATE_CONTROL : coverpoint `INT_CONTROL_CREDIT_HIST_01_CIAL_CLOCK_GATE_CONTROL   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_CREDIT_HIST_02_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_CREDIT_HIST_02_TARGET_CFG_CREDIT_HIST_02_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_CREDIT_HIST_02 HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_L1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_ENQPIPE_ERROR_INJECTION_H1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_L1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_SCHPIPE_ERROR_INJECTION_H1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_L1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_ERROR_INJECTION_H1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_L1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_ERROR_INJECTION_H1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_INGRESS_FLID_PARITY_ERROR_INJECTION_1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_ENGPIPE_FLID_PARITY_ERROR_INJECTION : coverpoint `INT_CONTROL_CREDIT_HIST_02_ENGPIPE_FLID_PARITY_ERROR_INJECTION   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_0 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_0   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_1 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_1   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_2 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_2   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_3 : coverpoint `INT_CONTROL_CREDIT_HIST_02_EGRESS_WBO_ERROR_INJECTION_3   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_CREDIT_HIST_02_CONTROL : coverpoint `INT_CONTROL_CREDIT_HIST_02_CONTROL   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_DIR_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_DIR_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_DIR_PIPE_CHICKEN_SIM : coverpoint `INT_CONTROL_DIR_PIPE_CHICKEN_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_DIR_PIPE_CHICKEN_50 : coverpoint `INT_CONTROL_DIR_PIPE_CHICKEN_50   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_LIST_SEL_0_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_LIST_SEL_0_TARGET_CFG_LIST_SEL_0_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_LIST_SEL_0 HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_LIST_SEL_0_DISAB_ATQ_EMPTY_ARB : coverpoint `INT_CONTROL_LIST_SEL_0_DISAB_ATQ_EMPTY_ARB   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_INC_TOK_UNIT_IDLE : coverpoint `INT_CONTROL_LIST_SEL_0_INC_TOK_UNIT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DISAB_RLIST_PRI : coverpoint `INT_CONTROL_LIST_SEL_0_DISAB_RLIST_PRI   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_INC_CMP_UNIT_IDLE : coverpoint `INT_CONTROL_LIST_SEL_0_INC_CMP_UNIT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ENAB_IF_THRESH : coverpoint `INT_CONTROL_LIST_SEL_0_ENAB_IF_THRESH   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OP : coverpoint `INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIR_HALF_BW : coverpoint `INT_CONTROL_LIST_SEL_0_DIR_HALF_BW   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OUT : coverpoint `INT_CONTROL_LIST_SEL_0_DIR_SINGLE_OUT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIR_DISAB_MULTI : coverpoint `INT_CONTROL_LIST_SEL_0_DIR_DISAB_MULTI   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OP : coverpoint `INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATQ_HALF_BW : coverpoint `INT_CONTROL_LIST_SEL_0_ATQ_HALF_BW   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OUT : coverpoint `INT_CONTROL_LIST_SEL_0_ATQ_SINGLE_OUT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATQ_DISAB_MULTI : coverpoint `INT_CONTROL_LIST_SEL_0_ATQ_DISAB_MULTI   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OP : coverpoint `INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIRRPL_HALF_BW : coverpoint `INT_CONTROL_LIST_SEL_0_DIRRPL_HALF_BW   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OUT : coverpoint `INT_CONTROL_LIST_SEL_0_DIRRPL_SINGLE_OUT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OP : coverpoint `INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LBRPL_HALF_BW : coverpoint `INT_CONTROL_LIST_SEL_0_LBRPL_HALF_BW   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OUT : coverpoint `INT_CONTROL_LIST_SEL_0_LBRPL_SINGLE_OUT   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LDB_SINGLE_OP : coverpoint `INT_CONTROL_LIST_SEL_0_LDB_SINGLE_OP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LDB_HALF_BW : coverpoint `INT_CONTROL_LIST_SEL_0_LDB_HALF_BW   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LDB_DISAB_MULTI : coverpoint `INT_CONTROL_LIST_SEL_0_LDB_DISAB_MULTI   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATM_SINGLE_SCH : coverpoint `INT_CONTROL_LIST_SEL_0_ATM_SINGLE_SCH   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_ATM_SINGLE_CMP : coverpoint `INT_CONTROL_LIST_SEL_0_ATM_SINGLE_CMP   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_LDB_CE_TOG_ARB : coverpoint `INT_CONTROL_LIST_SEL_0_LDB_CE_TOG_ARB   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_SMON0_VALID_SEL : coverpoint `INT_CONTROL_LIST_SEL_0_SMON0_VALID_SEL   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_SMON0_VALUE_SEL : coverpoint `INT_CONTROL_LIST_SEL_0_SMON0_VALUE_SEL   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_0_SMON0_COMPARE_SEL : coverpoint `INT_CONTROL_LIST_SEL_0_SMON0_COMPARE_SEL   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_LIST_SEL_1_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_LIST_SEL_1_TARGET_CFG_LIST_SEL_1_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_LIST_SEL_1 HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_LIST_SEL_1_QE_WT_FRC : coverpoint `INT_CONTROL_LIST_SEL_1_QE_WT_FRC   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_1_QE_WT_FRCV : coverpoint `INT_CONTROL_LIST_SEL_1_QE_WT_FRCV   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_1_QE_WT_BLK : coverpoint `INT_CONTROL_LIST_SEL_1_QE_WT_BLK   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_1_QED_DEQ_HIPRI_WM : coverpoint `INT_CONTROL_LIST_SEL_1_QED_DEQ_HIPRI_WM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_1_DIS_WU_RES_CHK : coverpoint `INT_CONTROL_LIST_SEL_1_DIS_WU_RES_CHK   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_LIST_SEL_1_AQED_DEQ_HIPRI_WM : coverpoint `INT_CONTROL_LIST_SEL_1_AQED_DEQ_HIPRI_WM   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_NALB_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_NALB_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_NALB_PIPE_CHICKEN_SIM : coverpoint `INT_CONTROL_NALB_PIPE_CHICKEN_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_NALB_PIPE_CHICKEN_50 : coverpoint `INT_CONTROL_NALB_PIPE_CHICKEN_50   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_QED_PIPE_REG_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_QED_PIPE_REG HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_QED_PIPE_REG_CHICKEN_SIM : coverpoint `INT_CONTROL_QED_PIPE_REG_CHICKEN_SIM   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_QED_PIPE_REG_CHICKEN_STRICT : coverpoint `INT_CONTROL_QED_PIPE_REG_CHICKEN_STRICT   iff (rst_n & cfg_write) ;
endgroup 

covergroup CONTROL_REORDER_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_CONTROL_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_CONTROL.clk ) ;

 option.comment = "CONTROL_REORDER_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_CONTROL_REORDER_PIPE_UNIT_SINGLE_STEP_MODE : coverpoint `INT_CONTROL_REORDER_PIPE_UNIT_SINGLE_STEP_MODE   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_REORDER_PIPE_RR_EN : coverpoint `INT_CONTROL_REORDER_PIPE_RR_EN   iff (rst_n & cfg_write) ;
CP_REG_INT_CONTROL_REORDER_PIPE_RSZV0 : coverpoint `INT_CONTROL_REORDER_PIPE_RSZV0   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_AQED_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_AQED_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_LSP_SCH_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_CHP_SCH_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_AQED_AP_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_QED_AQED_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_AP_AQED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_DEPTH : coverpoint `INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_READY : coverpoint `INT_STATUS_AQED_PIPE_DB_LSP_AQED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_LSP_AQED_CMP_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_LSP_AQED_CMP_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_FID_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_FID_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_AQED_CHP_SCH_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_AQED_CHP_SCH_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_AP_AQED_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_AP_AQED_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_AQED_AP_ENQ_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_AQED_AP_ENQ_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_QED_AQED_ENQ_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_FIFO_FREELIST_RETURN_EMPTY : coverpoint `INT_STATUS_AQED_PIPE_FIFO_FREELIST_RETURN_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_AQED_PIPE_AQED_CLK_IDLE : coverpoint `INT_STATUS_AQED_PIPE_AQED_CLK_IDLE   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_ATM_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_ATM_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_READY_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_LSP_AP_SCH_ATM_STATUS_READY_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_READY : coverpoint `INT_STATUS_ATM_PIPE_DB_AP_LSP_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_READY : coverpoint `INT_STATUS_ATM_PIPE_DB_AQED_AP_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_READY : coverpoint `INT_STATUS_ATM_PIPE_DB_AP_AQED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_DEPTH : coverpoint `INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_READY : coverpoint `INT_STATUS_ATM_PIPE_DB_LSP_AQED_CMP_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_ATM_PIPE_ATM_CLK_IDLE : coverpoint `INT_STATUS_ATM_PIPE_ATM_CLK_IDLE   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_DIR_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_DIR_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_DQED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DP_DQED_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DP_DQED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DP_DQED_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DP_DQED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_RORPLY_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_DP_LSP_ENQ_DIR_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_RORPLY_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_LSP_DP_SCH_DIR_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_READY : coverpoint `INT_STATUS_DIR_PIPE_DB_ROP_DP_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_DIR_PIPE_INT_IDLE_B : coverpoint `INT_STATUS_DIR_PIPE_INT_IDLE_B   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_LIST_SEL_INTERFACE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_LIST_SEL_INTERFACE_TARGET_CFG_LIST_SEL_INTERFACE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_LIST_SEL_INTERFACE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_AQED_LSP_SENT_TO_CQ_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_RORPLY_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_DP_LSP_ENQ_DIR_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_RORPLY_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_NALB_LSP_ENQ_LDB_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_ROP_LSP_REORDCMP_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_CMP_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_CHP_LSP_TOK_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_INT_SER_CLOCK_NOT_IDLE : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_INT_SER_CLOCK_NOT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_AQED_CLOCK_NOT_IDLE : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_AQED_CLOCK_NOT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_AP_CLOCK_NOT_IDLE : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_AP_CLOCK_NOT_IDLE   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_RORPLY_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_RORPLY_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_DP_SCH_DIR_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_ATQ_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_NALB_SCH_UO_NOT_RDY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_V : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_NOT_RDY : coverpoint `INT_STATUS_LIST_SEL_INTERFACE_LSP_AP_ATM_NOT_RDY   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_NALB_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_NALB_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_QED_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_RORPLY_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_NALB_LSP_ENQ_LB_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_ATQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_RORPLY_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_LSP_NALB_SCH_UNOORD_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_DEPTH : coverpoint `INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_DEPTH   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_READY : coverpoint `INT_STATUS_NALB_PIPE_DB_ROP_NALB_ENQ_STATUS_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_NALB_PIPE_INT_IDLE_B : coverpoint `INT_STATUS_NALB_PIPE_INT_IDLE_B   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_QED_PIPE_REG_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_STATUS.clk ) ;

 option.comment = "STATUS_QED_PIPE_REG HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_READY : coverpoint `INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_V : coverpoint `INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_READY : coverpoint `INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_V : coverpoint `INT_STATUS_QED_PIPE_REG_NALB_LSP_ENQ_LB_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_READY : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_V : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_ATQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_READY : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_V : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_READY : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_V : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_NALB_SCH_UNOORD_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_READY : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_V : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_NALB_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_READY : coverpoint `INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_V : coverpoint `INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_READY : coverpoint `INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_V : coverpoint `INT_STATUS_QED_PIPE_REG_DP_LSP_ENQ_DIR_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_READY : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_V : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_RORPLY_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_READY : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_V : coverpoint `INT_STATUS_QED_PIPE_REG_LSP_DP_SCH_DIR_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_READY : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_V : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_DP_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_READY : coverpoint `INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_V : coverpoint `INT_STATUS_QED_PIPE_REG_DQED_CHP_SCH_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_READY : coverpoint `INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_V : coverpoint `INT_STATUS_QED_PIPE_REG_QED_AQED_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_READY : coverpoint `INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_V : coverpoint `INT_STATUS_QED_PIPE_REG_QED_CHP_SCH_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_QED_ENQ_READY : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_QED_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_ROP_QED_DQED_ENQ_V : coverpoint `INT_STATUS_QED_PIPE_REG_ROP_QED_DQED_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_QED_PIPE_REG_INT_IDLE : coverpoint `INT_STATUS_QED_PIPE_REG_INT_IDLE   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_REORDER_PIPE_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_STATUS.clk ) ;

 option.comment = "STATUS_REORDER_PIPE HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_ALARM_UP_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_ALARM_DOWN_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_READY : coverpoint `INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_V : coverpoint `INT_STATUS_REORDER_PIPE_CHP_ROP_HCW_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_DP_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_NALB_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_QED_ENQ_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_QED_ENQ_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_QED_DQED_ENQ_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_QED_DQED_ENQ_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_READY : coverpoint `INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_READY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_V : coverpoint `INT_STATUS_REORDER_PIPE_ROP_LSP_REORDERCMP_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_REORDER_PIPE_INT_IDLE_B : coverpoint `INT_STATUS_REORDER_PIPE_INT_IDLE_B   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_MASTER_CORE_DIAGNOSTIC_1_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_MASTER_CORE_DIAGNOSTIC_1_TARGET_CFG_MASTER_CORE_DIAGNOSTIC_1_CSR_STATUS.clk ) ;

 option.comment = "STATUS_MASTER_CORE_DIAGNOSTIC_1 HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_TIMEOUT_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_TIMEOUT_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQRSP_UNSOL_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQRSP_UNSOL_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_PROTOCOL_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_PROTOCOL_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLV_PAR_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLV_PAR_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_PAR_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_PAR_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_DROP_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_DROP_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_UP_MISS_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_REQ_UP_MISS_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_DECODE_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_ACCESS_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_ACCESS_ERR   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_TIMEOUT_ERR : coverpoint `INT_STATUS_MASTER_CORE_DIAGNOSTIC_1_CFG_SLAVE_TIMEOUT_ERR   iff (rst_n & cfg_write) ;
endgroup 

covergroup STATUS_LIST_SEL_DIAGNOSTIC_0_functional_reg_CG (ref logic rst_n, ref logic cfg_write ) @ (posedge ` I_HQM_STATUS_LIST_SEL_DIAGNOSTIC_0_TARGET_CFG_LIST_SEL_DIAGNOSTIC_0_CSR_STATUS.clk ) ;

 option.comment = "STATUS_LIST_SEL_DIAGNOSTIC_0 HQM Functional Register Coverage ";

 CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_BLAST : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_SLIST_BLAST   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_BLAST : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_RLIST_BLAST   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_BLAST : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_BLAST   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST_CHKV : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST_CHKV   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_CMPBLAST   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_QID_DIS : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_QID_DIS   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_BUSY : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_BUSY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_NO_SPACE : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_NO_SPACE   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_DIR_TOK_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_DIR_TOK_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_ACT : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_ACT   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AP_LSP_ATM_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AP_LSP_ATM_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_TOK_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_TOK_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CMP_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CMP_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS0 : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS0   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS1 : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS1   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS2 : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS2   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS3 : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_LDB_CQ_ARB_REQV_COS3   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_STOP_ATQATM : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATQ_STOP_ATQATM   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_SN_FCERR_RPTD : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_NALB_SN_FCERR_RPTD   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_EMPTY : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_AQED_EMPTY   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATM_IF_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_ATM_IF_V   iff (rst_n & cfg_write) ;
CP_REG_INT_STATUS_LIST_SEL_DIAGNOSTIC_0_TOT_IF_V : coverpoint `INT_STATUS_LIST_SEL_DIAGNOSTIC_0_TOT_IF_V   iff (rst_n & cfg_write) ;
endgroup 

initial begin

 CONTROL_AQED_PIPE_functional_reg_CG CONTROL_AQED_PIPE_functional_reg_CG_inst = new(` I_HQM_CONTROL_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_CONTROL.cfg_write);

 CONTROL_ATM_PIPE_functional_reg_CG CONTROL_ATM_PIPE_functional_reg_CG_inst = new(` I_HQM_CONTROL_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_CONTROL.cfg_write);

 CONTROL_MASTER_CORE_CONTROL_functional_reg_CG CONTROL_MASTER_CORE_CONTROL_functional_reg_CG_inst = new(` I_HQM_CONTROL_MASTER_CORE_CONTROL_TARGET_CFG_MASTER_CORE_CONTROL_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_MASTER_CORE_CONTROL_TARGET_CFG_MASTER_CORE_CONTROL_CSR_CONTROL.cfg_write);

 CONTROL_CREDIT_HIST_00_functional_reg_CG CONTROL_CREDIT_HIST_00_functional_reg_CG_inst = new(` I_HQM_CONTROL_CREDIT_HIST_00_TARGET_CFG_CREDIT_HIST_00_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_CREDIT_HIST_00_TARGET_CFG_CREDIT_HIST_00_CSR_CONTROL.cfg_write);

 CONTROL_CREDIT_HIST_01_functional_reg_CG CONTROL_CREDIT_HIST_01_functional_reg_CG_inst = new(` I_HQM_CONTROL_CREDIT_HIST_01_TARGET_CFG_CREDIT_HIST_01_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_CREDIT_HIST_01_TARGET_CFG_CREDIT_HIST_01_CSR_CONTROL.cfg_write);

 CONTROL_CREDIT_HIST_02_functional_reg_CG CONTROL_CREDIT_HIST_02_functional_reg_CG_inst = new(` I_HQM_CONTROL_CREDIT_HIST_02_TARGET_CFG_CREDIT_HIST_02_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_CREDIT_HIST_02_TARGET_CFG_CREDIT_HIST_02_CSR_CONTROL.cfg_write);

 CONTROL_DIR_PIPE_functional_reg_CG CONTROL_DIR_PIPE_functional_reg_CG_inst = new(` I_HQM_CONTROL_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_CONTROL.cfg_write);

 CONTROL_LIST_SEL_0_functional_reg_CG CONTROL_LIST_SEL_0_functional_reg_CG_inst = new(` I_HQM_CONTROL_LIST_SEL_0_TARGET_CFG_LIST_SEL_0_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_LIST_SEL_0_TARGET_CFG_LIST_SEL_0_CSR_CONTROL.cfg_write);

 CONTROL_LIST_SEL_1_functional_reg_CG CONTROL_LIST_SEL_1_functional_reg_CG_inst = new(` I_HQM_CONTROL_LIST_SEL_1_TARGET_CFG_LIST_SEL_1_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_LIST_SEL_1_TARGET_CFG_LIST_SEL_1_CSR_CONTROL.cfg_write);

 CONTROL_NALB_PIPE_functional_reg_CG CONTROL_NALB_PIPE_functional_reg_CG_inst = new(` I_HQM_CONTROL_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_CONTROL.cfg_write);

 CONTROL_QED_PIPE_REG_functional_reg_CG CONTROL_QED_PIPE_REG_functional_reg_CG_inst = new(` I_HQM_CONTROL_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_CONTROL.cfg_write);

 CONTROL_REORDER_PIPE_functional_reg_CG CONTROL_REORDER_PIPE_functional_reg_CG_inst = new(` I_HQM_CONTROL_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_CONTROL.rst_n, ` I_HQM_CONTROL_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_CONTROL.cfg_write);

 STATUS_AQED_PIPE_functional_reg_CG STATUS_AQED_PIPE_functional_reg_CG_inst = new(` I_HQM_STATUS_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_STATUS.rst_n, ` I_HQM_STATUS_AQED_PIPE_TARGET_CFG_AQED_PIPE_CSR_STATUS.cfg_write);

 STATUS_ATM_PIPE_functional_reg_CG STATUS_ATM_PIPE_functional_reg_CG_inst = new(` I_HQM_STATUS_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_STATUS.rst_n, ` I_HQM_STATUS_ATM_PIPE_TARGET_CFG_ATM_PIPE_CSR_STATUS.cfg_write);

 STATUS_DIR_PIPE_functional_reg_CG STATUS_DIR_PIPE_functional_reg_CG_inst = new(` I_HQM_STATUS_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_STATUS.rst_n, ` I_HQM_STATUS_DIR_PIPE_TARGET_CFG_DIR_PIPE_CSR_STATUS.cfg_write);

 STATUS_LIST_SEL_INTERFACE_functional_reg_CG STATUS_LIST_SEL_INTERFACE_functional_reg_CG_inst = new(` I_HQM_STATUS_LIST_SEL_INTERFACE_TARGET_CFG_LIST_SEL_INTERFACE_CSR_STATUS.rst_n, ` I_HQM_STATUS_LIST_SEL_INTERFACE_TARGET_CFG_LIST_SEL_INTERFACE_CSR_STATUS.cfg_write);

 STATUS_NALB_PIPE_functional_reg_CG STATUS_NALB_PIPE_functional_reg_CG_inst = new(` I_HQM_STATUS_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_STATUS.rst_n, ` I_HQM_STATUS_NALB_PIPE_TARGET_CFG_NALB_PIPE_CSR_STATUS.cfg_write);

 STATUS_QED_PIPE_REG_functional_reg_CG STATUS_QED_PIPE_REG_functional_reg_CG_inst = new(` I_HQM_STATUS_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_STATUS.rst_n, ` I_HQM_STATUS_QED_PIPE_REG_TARGET_CFG_QED_PIPE_REG_CSR_STATUS.cfg_write);

 STATUS_REORDER_PIPE_functional_reg_CG STATUS_REORDER_PIPE_functional_reg_CG_inst = new(` I_HQM_STATUS_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_STATUS.rst_n, ` I_HQM_STATUS_REORDER_PIPE_TARGET_CFG_REORDER_PIPE_CSR_STATUS.cfg_write);

 STATUS_MASTER_CORE_DIAGNOSTIC_1_functional_reg_CG STATUS_MASTER_CORE_DIAGNOSTIC_1_functional_reg_CG_inst = new(` I_HQM_STATUS_MASTER_CORE_DIAGNOSTIC_1_TARGET_CFG_MASTER_CORE_DIAGNOSTIC_1_CSR_STATUS.rst_n, ` I_HQM_STATUS_MASTER_CORE_DIAGNOSTIC_1_TARGET_CFG_MASTER_CORE_DIAGNOSTIC_1_CSR_STATUS.cfg_write);

 STATUS_LIST_SEL_DIAGNOSTIC_0_functional_reg_CG STATUS_LIST_SEL_DIAGNOSTIC_0_functional_reg_CG_inst = new(` I_HQM_STATUS_LIST_SEL_DIAGNOSTIC_0_TARGET_CFG_LIST_SEL_DIAGNOSTIC_0_CSR_STATUS.rst_n, ` I_HQM_STATUS_LIST_SEL_DIAGNOSTIC_0_TARGET_CFG_LIST_SEL_DIAGNOSTIC_0_CSR_STATUS.cfg_write);

end

 `endif

 endmodule

 
