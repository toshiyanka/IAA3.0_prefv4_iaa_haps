VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf198b128e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf198b128e1r1w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 43.2 BY 41.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 22.44 22.416 23.64 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 20.52 19.116 21.72 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 22.44 23.616 23.64 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 22.44 23.872 23.64 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 22.44 18.472 23.64 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 22.44 18.728 23.64 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 22.44 19.028 23.64 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 22.44 19.116 23.64 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 22.44 19.372 23.64 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 22.44 22.628 23.64 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 22.44 22.972 23.64 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 22.44 23.228 23.64 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.484 22.44 23.528 23.64 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 20.52 20.828 21.72 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 20.52 20.916 21.72 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 20.52 21.172 21.72 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 20.52 21.428 21.72 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 20.52 21.516 21.72 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 20.52 21.816 21.72 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 20.52 22.072 21.72 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 20.52 19.372 21.72 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 20.52 19.716 21.72 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 0.24 20.616 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 18.24 20.916 19.44 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 18.24 21.172 19.44 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 18.24 21.428 19.44 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 18.24 21.516 19.44 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 18.96 20.528 20.16 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 18.96 20.616 20.16 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 18.96 22.328 20.16 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 18.96 21.728 20.16 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 24 20.616 25.2 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 24 20.828 25.2 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 1.68 22.328 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 24 22.072 25.2 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 24 22.328 25.2 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 24.72 20.272 25.92 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 24.72 20.528 25.92 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 24.72 21.728 25.92 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 24.72 21.816 25.92 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 25.44 20.916 26.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 25.44 21.172 26.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 25.44 21.428 26.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 25.44 21.516 26.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 1.68 21.728 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 26.16 20.528 27.36 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 26.16 20.616 27.36 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 26.16 22.328 27.36 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 26.16 21.728 27.36 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 26.88 20.272 28.08 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 26.88 20.828 28.08 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 26.88 21.816 28.08 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 26.88 22.072 28.08 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 27.6 20.916 28.8 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 27.6 21.172 28.8 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 2.4 20.272 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 27.6 21.428 28.8 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 27.6 21.516 28.8 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 28.32 20.528 29.52 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 28.32 20.616 29.52 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 28.32 22.328 29.52 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 28.32 21.728 29.52 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 29.04 20.272 30.24 ;
    END
  END wrdatap0[136]
  PIN wrdatap0[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 29.04 20.828 30.24 ;
    END
  END wrdatap0[137]
  PIN wrdatap0[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 29.04 21.816 30.24 ;
    END
  END wrdatap0[138]
  PIN wrdatap0[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 29.04 22.072 30.24 ;
    END
  END wrdatap0[139]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 2.4 20.828 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 29.76 20.916 30.96 ;
    END
  END wrdatap0[140]
  PIN wrdatap0[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 29.76 21.172 30.96 ;
    END
  END wrdatap0[141]
  PIN wrdatap0[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 29.76 21.428 30.96 ;
    END
  END wrdatap0[142]
  PIN wrdatap0[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 29.76 21.516 30.96 ;
    END
  END wrdatap0[143]
  PIN wrdatap0[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 30.48 20.528 31.68 ;
    END
  END wrdatap0[144]
  PIN wrdatap0[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 30.48 20.616 31.68 ;
    END
  END wrdatap0[145]
  PIN wrdatap0[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 30.48 22.328 31.68 ;
    END
  END wrdatap0[146]
  PIN wrdatap0[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 30.48 21.728 31.68 ;
    END
  END wrdatap0[147]
  PIN wrdatap0[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 31.2 20.272 32.4 ;
    END
  END wrdatap0[148]
  PIN wrdatap0[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 31.2 20.828 32.4 ;
    END
  END wrdatap0[149]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.4 21.816 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 31.2 21.816 32.4 ;
    END
  END wrdatap0[150]
  PIN wrdatap0[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 31.2 22.072 32.4 ;
    END
  END wrdatap0[151]
  PIN wrdatap0[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 31.92 20.916 33.12 ;
    END
  END wrdatap0[152]
  PIN wrdatap0[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 31.92 21.172 33.12 ;
    END
  END wrdatap0[153]
  PIN wrdatap0[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 31.92 21.428 33.12 ;
    END
  END wrdatap0[154]
  PIN wrdatap0[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 31.92 21.516 33.12 ;
    END
  END wrdatap0[155]
  PIN wrdatap0[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 32.64 20.528 33.84 ;
    END
  END wrdatap0[156]
  PIN wrdatap0[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 32.64 20.616 33.84 ;
    END
  END wrdatap0[157]
  PIN wrdatap0[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 32.64 22.328 33.84 ;
    END
  END wrdatap0[158]
  PIN wrdatap0[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 32.64 21.728 33.84 ;
    END
  END wrdatap0[159]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 2.4 22.072 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 33.36 20.272 34.56 ;
    END
  END wrdatap0[160]
  PIN wrdatap0[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 33.36 20.828 34.56 ;
    END
  END wrdatap0[161]
  PIN wrdatap0[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 33.36 21.816 34.56 ;
    END
  END wrdatap0[162]
  PIN wrdatap0[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 33.36 22.072 34.56 ;
    END
  END wrdatap0[163]
  PIN wrdatap0[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 34.08 20.916 35.28 ;
    END
  END wrdatap0[164]
  PIN wrdatap0[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 34.08 21.172 35.28 ;
    END
  END wrdatap0[165]
  PIN wrdatap0[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 34.08 21.428 35.28 ;
    END
  END wrdatap0[166]
  PIN wrdatap0[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 34.08 21.516 35.28 ;
    END
  END wrdatap0[167]
  PIN wrdatap0[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 34.8 20.528 36 ;
    END
  END wrdatap0[168]
  PIN wrdatap0[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 34.8 20.616 36 ;
    END
  END wrdatap0[169]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 3.12 20.916 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 34.8 22.328 36 ;
    END
  END wrdatap0[170]
  PIN wrdatap0[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 34.8 21.728 36 ;
    END
  END wrdatap0[171]
  PIN wrdatap0[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 35.52 20.272 36.72 ;
    END
  END wrdatap0[172]
  PIN wrdatap0[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 35.52 20.828 36.72 ;
    END
  END wrdatap0[173]
  PIN wrdatap0[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 35.52 21.816 36.72 ;
    END
  END wrdatap0[174]
  PIN wrdatap0[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 35.52 22.072 36.72 ;
    END
  END wrdatap0[175]
  PIN wrdatap0[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 36.24 20.916 37.44 ;
    END
  END wrdatap0[176]
  PIN wrdatap0[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 36.24 21.172 37.44 ;
    END
  END wrdatap0[177]
  PIN wrdatap0[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 36.24 21.428 37.44 ;
    END
  END wrdatap0[178]
  PIN wrdatap0[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 36.24 21.516 37.44 ;
    END
  END wrdatap0[179]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 3.12 21.172 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 36.96 20.528 38.16 ;
    END
  END wrdatap0[180]
  PIN wrdatap0[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 36.96 20.616 38.16 ;
    END
  END wrdatap0[181]
  PIN wrdatap0[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 36.96 22.328 38.16 ;
    END
  END wrdatap0[182]
  PIN wrdatap0[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 36.96 21.728 38.16 ;
    END
  END wrdatap0[183]
  PIN wrdatap0[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 37.68 20.272 38.88 ;
    END
  END wrdatap0[184]
  PIN wrdatap0[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 37.68 20.828 38.88 ;
    END
  END wrdatap0[185]
  PIN wrdatap0[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 37.68 21.816 38.88 ;
    END
  END wrdatap0[186]
  PIN wrdatap0[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 37.68 22.072 38.88 ;
    END
  END wrdatap0[187]
  PIN wrdatap0[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 38.4 20.916 39.6 ;
    END
  END wrdatap0[188]
  PIN wrdatap0[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 38.4 21.172 39.6 ;
    END
  END wrdatap0[189]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 3.12 21.428 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 38.4 21.428 39.6 ;
    END
  END wrdatap0[190]
  PIN wrdatap0[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 38.4 21.516 39.6 ;
    END
  END wrdatap0[191]
  PIN wrdatap0[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 39.12 20.528 40.32 ;
    END
  END wrdatap0[192]
  PIN wrdatap0[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 39.12 20.616 40.32 ;
    END
  END wrdatap0[193]
  PIN wrdatap0[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 39.12 22.328 40.32 ;
    END
  END wrdatap0[194]
  PIN wrdatap0[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 39.12 21.728 40.32 ;
    END
  END wrdatap0[195]
  PIN wrdatap0[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 39.84 20.272 41.04 ;
    END
  END wrdatap0[196]
  PIN wrdatap0[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 39.84 20.828 41.04 ;
    END
  END wrdatap0[197]
  PIN wrdatap0[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 39.84 21.816 41.04 ;
    END
  END wrdatap0[198]
  PIN wrdatap0[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 39.84 22.072 41.04 ;
    END
  END wrdatap0[199]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 3.12 21.516 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 0.24 20.828 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 3.84 20.528 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 3.84 20.616 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 3.84 22.328 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 3.84 21.728 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 4.56 20.272 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 4.56 20.828 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 4.56 21.816 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 4.56 22.072 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 5.28 20.916 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 5.28 21.172 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 0.24 22.072 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 5.28 21.428 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 5.28 21.516 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 6 20.528 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 6 20.616 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 6 22.328 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 6 21.728 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 6.72 20.272 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 6.72 20.828 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 6.72 21.816 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 6.72 22.072 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 0.24 22.328 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 7.44 20.916 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 7.44 21.172 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 7.44 21.428 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 7.44 21.516 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 8.16 20.528 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 8.16 20.616 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 8.16 22.328 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 8.16 21.728 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 8.88 20.272 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 8.88 20.828 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 0.96 20.916 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 8.88 21.816 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 8.88 22.072 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 9.6 20.916 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 9.6 21.172 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 9.6 21.428 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 9.6 21.516 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 10.32 20.528 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 10.32 20.616 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 10.32 22.328 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 10.32 21.728 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 0.96 21.172 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 11.04 20.272 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 11.04 20.828 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 11.04 21.816 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 11.04 22.072 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 11.76 20.916 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 11.76 21.172 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 11.76 21.428 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 11.76 21.516 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 12.48 20.528 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 12.48 20.616 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 0.96 21.428 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 12.48 22.328 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 12.48 21.728 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 13.2 20.272 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 13.2 20.828 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 13.2 21.816 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 13.2 22.072 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 13.92 20.916 15.12 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 13.92 21.172 15.12 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 13.92 21.428 15.12 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 13.92 21.516 15.12 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 0.96 21.516 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 14.64 20.528 15.84 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 14.64 20.616 15.84 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 14.64 22.328 15.84 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 14.64 21.728 15.84 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 15.36 20.272 16.56 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 15.36 20.828 16.56 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 15.36 21.816 16.56 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 15.36 22.072 16.56 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 16.08 20.916 17.28 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 16.08 21.172 17.28 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 1.68 20.528 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 16.08 21.428 17.28 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 16.08 21.516 17.28 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 16.8 20.528 18 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 16.8 20.616 18 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 16.8 22.328 18 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 16.8 21.728 18 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 17.52 20.272 18.72 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 17.52 20.828 18.72 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 17.52 21.816 18.72 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 17.52 22.072 18.72 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.68 20.616 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 20.52 20.016 21.72 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 20.52 20.272 21.72 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 20.52 19.928 21.72 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 18.24 18.472 19.44 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 18.24 18.728 19.44 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 18.24 22.972 19.44 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 18.24 23.228 19.44 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 18.96 19.628 20.16 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 18.96 18.816 20.16 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 18.96 22.716 20.16 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 18.96 23.316 20.16 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 24 18.816 25.2 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 24 19.628 25.2 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 1.68 22.716 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 24 22.716 25.2 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 24 23.316 25.2 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 24.72 19.028 25.92 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 24.72 19.116 25.92 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 24.72 23.616 25.92 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 24.72 23.872 25.92 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 25.44 18.472 26.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 25.44 18.728 26.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 25.44 22.972 26.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 25.44 23.228 26.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 1.68 23.316 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 26.16 19.628 27.36 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.16 18.816 27.36 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 26.16 22.716 27.36 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 26.16 23.316 27.36 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 26.88 19.116 28.08 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 26.88 19.372 28.08 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 26.88 23.616 28.08 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 26.88 23.872 28.08 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 27.6 18.472 28.8 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 27.6 18.728 28.8 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 2.4 19.116 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 27.6 22.972 28.8 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 27.6 23.228 28.8 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 28.32 19.628 29.52 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 28.32 18.816 29.52 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 28.32 22.716 29.52 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 28.32 23.316 29.52 ;
    END
  END rddatap0[135]
  PIN rddatap0[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 29.04 19.116 30.24 ;
    END
  END rddatap0[136]
  PIN rddatap0[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 29.04 19.372 30.24 ;
    END
  END rddatap0[137]
  PIN rddatap0[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 29.04 23.616 30.24 ;
    END
  END rddatap0[138]
  PIN rddatap0[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 29.04 23.872 30.24 ;
    END
  END rddatap0[139]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 2.4 19.372 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 29.76 18.472 30.96 ;
    END
  END rddatap0[140]
  PIN rddatap0[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 29.76 18.728 30.96 ;
    END
  END rddatap0[141]
  PIN rddatap0[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 29.76 22.972 30.96 ;
    END
  END rddatap0[142]
  PIN rddatap0[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 29.76 23.228 30.96 ;
    END
  END rddatap0[143]
  PIN rddatap0[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 30.48 19.628 31.68 ;
    END
  END rddatap0[144]
  PIN rddatap0[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 30.48 18.816 31.68 ;
    END
  END rddatap0[145]
  PIN rddatap0[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 30.48 22.716 31.68 ;
    END
  END rddatap0[146]
  PIN rddatap0[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 30.48 23.316 31.68 ;
    END
  END rddatap0[147]
  PIN rddatap0[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 31.2 19.116 32.4 ;
    END
  END rddatap0[148]
  PIN rddatap0[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 31.2 19.372 32.4 ;
    END
  END rddatap0[149]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 2.4 23.616 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 31.2 23.616 32.4 ;
    END
  END rddatap0[150]
  PIN rddatap0[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 31.2 23.872 32.4 ;
    END
  END rddatap0[151]
  PIN rddatap0[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 31.92 18.472 33.12 ;
    END
  END rddatap0[152]
  PIN rddatap0[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 31.92 18.728 33.12 ;
    END
  END rddatap0[153]
  PIN rddatap0[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 31.92 22.972 33.12 ;
    END
  END rddatap0[154]
  PIN rddatap0[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 31.92 23.228 33.12 ;
    END
  END rddatap0[155]
  PIN rddatap0[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 32.64 19.628 33.84 ;
    END
  END rddatap0[156]
  PIN rddatap0[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 32.64 18.816 33.84 ;
    END
  END rddatap0[157]
  PIN rddatap0[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 32.64 22.716 33.84 ;
    END
  END rddatap0[158]
  PIN rddatap0[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 32.64 23.316 33.84 ;
    END
  END rddatap0[159]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 2.4 23.872 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 33.36 19.116 34.56 ;
    END
  END rddatap0[160]
  PIN rddatap0[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 33.36 19.372 34.56 ;
    END
  END rddatap0[161]
  PIN rddatap0[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 33.36 23.616 34.56 ;
    END
  END rddatap0[162]
  PIN rddatap0[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 33.36 23.872 34.56 ;
    END
  END rddatap0[163]
  PIN rddatap0[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 34.08 18.472 35.28 ;
    END
  END rddatap0[164]
  PIN rddatap0[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 34.08 18.728 35.28 ;
    END
  END rddatap0[165]
  PIN rddatap0[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 34.08 22.972 35.28 ;
    END
  END rddatap0[166]
  PIN rddatap0[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 34.08 23.228 35.28 ;
    END
  END rddatap0[167]
  PIN rddatap0[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 34.8 19.628 36 ;
    END
  END rddatap0[168]
  PIN rddatap0[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 34.8 18.816 36 ;
    END
  END rddatap0[169]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 3.12 18.472 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 34.8 22.716 36 ;
    END
  END rddatap0[170]
  PIN rddatap0[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 34.8 23.316 36 ;
    END
  END rddatap0[171]
  PIN rddatap0[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 35.52 19.116 36.72 ;
    END
  END rddatap0[172]
  PIN rddatap0[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 35.52 19.372 36.72 ;
    END
  END rddatap0[173]
  PIN rddatap0[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 35.52 23.616 36.72 ;
    END
  END rddatap0[174]
  PIN rddatap0[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 35.52 23.872 36.72 ;
    END
  END rddatap0[175]
  PIN rddatap0[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 36.24 18.472 37.44 ;
    END
  END rddatap0[176]
  PIN rddatap0[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 36.24 18.728 37.44 ;
    END
  END rddatap0[177]
  PIN rddatap0[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 36.24 22.972 37.44 ;
    END
  END rddatap0[178]
  PIN rddatap0[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 36.24 23.228 37.44 ;
    END
  END rddatap0[179]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 3.12 18.728 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 36.96 19.628 38.16 ;
    END
  END rddatap0[180]
  PIN rddatap0[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 36.96 18.816 38.16 ;
    END
  END rddatap0[181]
  PIN rddatap0[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 36.96 22.716 38.16 ;
    END
  END rddatap0[182]
  PIN rddatap0[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 36.96 23.316 38.16 ;
    END
  END rddatap0[183]
  PIN rddatap0[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 37.68 19.116 38.88 ;
    END
  END rddatap0[184]
  PIN rddatap0[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 37.68 19.372 38.88 ;
    END
  END rddatap0[185]
  PIN rddatap0[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 37.68 23.616 38.88 ;
    END
  END rddatap0[186]
  PIN rddatap0[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 37.68 23.872 38.88 ;
    END
  END rddatap0[187]
  PIN rddatap0[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 38.4 18.472 39.6 ;
    END
  END rddatap0[188]
  PIN rddatap0[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 38.4 18.728 39.6 ;
    END
  END rddatap0[189]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 3.12 22.972 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 38.4 22.972 39.6 ;
    END
  END rddatap0[190]
  PIN rddatap0[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 38.4 23.228 39.6 ;
    END
  END rddatap0[191]
  PIN rddatap0[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 39.12 19.628 40.32 ;
    END
  END rddatap0[192]
  PIN rddatap0[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 39.12 18.816 40.32 ;
    END
  END rddatap0[193]
  PIN rddatap0[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 39.12 22.716 40.32 ;
    END
  END rddatap0[194]
  PIN rddatap0[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 39.12 23.316 40.32 ;
    END
  END rddatap0[195]
  PIN rddatap0[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 39.84 19.116 41.04 ;
    END
  END rddatap0[196]
  PIN rddatap0[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 39.84 19.372 41.04 ;
    END
  END rddatap0[197]
  PIN rddatap0[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 39.84 23.616 41.04 ;
    END
  END rddatap0[198]
  PIN rddatap0[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 39.84 23.872 41.04 ;
    END
  END rddatap0[199]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 3.12 23.228 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 3.84 19.628 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 3.84 18.816 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 3.84 22.716 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 3.84 23.316 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 4.56 19.116 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 4.56 19.372 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 4.56 23.616 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 4.56 23.872 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 5.28 18.472 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 5.28 18.728 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 0.24 23.616 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 5.28 22.972 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 5.28 23.228 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 6 19.628 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 6 18.816 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 6 22.716 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 6 23.316 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 6.72 19.116 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 6.72 19.372 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 6.72 23.616 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 6.72 23.872 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 0.24 23.872 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 7.44 18.472 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 7.44 18.728 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 7.44 22.972 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 7.44 23.228 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 8.16 19.628 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.16 18.816 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 8.16 22.716 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 8.16 23.316 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 8.88 19.116 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 8.88 19.372 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.96 18.816 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 8.88 23.616 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 8.88 23.872 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 9.6 18.472 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 9.6 18.728 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 9.6 22.972 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 9.6 23.228 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 10.32 19.628 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 10.32 18.816 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 10.32 22.716 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 10.32 23.316 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.96 19.028 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 11.04 19.116 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 11.04 19.372 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 11.04 23.616 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 11.04 23.872 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 11.76 18.472 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.76 18.728 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 11.76 22.972 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 11.76 23.228 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 12.48 19.628 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 12.48 18.816 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 0.96 22.972 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 12.48 22.716 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 12.48 23.316 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 13.2 19.116 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 13.2 19.372 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 13.2 23.616 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 13.2 23.872 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 13.92 18.472 15.12 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 13.92 18.728 15.12 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 13.92 22.972 15.12 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 13.92 23.228 15.12 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 0.96 23.228 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 14.64 19.628 15.84 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 14.64 18.816 15.84 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 14.64 22.716 15.84 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 14.64 23.316 15.84 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 15.36 19.116 16.56 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 15.36 19.372 16.56 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 15.36 23.616 16.56 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 15.36 23.872 16.56 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 16.08 18.472 17.28 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 16.08 18.728 17.28 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 1.68 19.628 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 16.08 22.972 17.28 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 16.08 23.228 17.28 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 16.8 19.628 18 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 16.8 18.816 18 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 16.8 22.716 18 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 16.8 23.316 18 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 17.52 19.116 18.72 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 17.52 19.372 18.72 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 17.52 23.616 18.72 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 17.52 23.872 18.72 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 1.68 18.472 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 41.22 ;
        RECT 2.662 0.06 2.738 41.22 ;
        RECT 4.462 0.06 4.538 41.22 ;
        RECT 6.262 0.06 6.338 41.22 ;
        RECT 8.062 0.06 8.138 41.22 ;
        RECT 9.862 0.06 9.938 41.22 ;
        RECT 11.662 0.06 11.738 41.22 ;
        RECT 13.462 0.06 13.538 41.22 ;
        RECT 15.262 0.06 15.338 41.22 ;
        RECT 17.062 0.06 17.138 41.22 ;
        RECT 18.862 0.06 18.938 41.22 ;
        RECT 20.662 0.06 20.738 41.22 ;
        RECT 22.462 0.06 22.538 41.22 ;
        RECT 24.262 0.06 24.338 41.22 ;
        RECT 26.062 0.06 26.138 41.22 ;
        RECT 27.862 0.06 27.938 41.22 ;
        RECT 29.662 0.06 29.738 41.22 ;
        RECT 31.462 0.06 31.538 41.22 ;
        RECT 33.262 0.06 33.338 41.22 ;
        RECT 35.062 0.06 35.138 41.22 ;
        RECT 36.862 0.06 36.938 41.22 ;
        RECT 38.662 0.06 38.738 41.22 ;
        RECT 40.462 0.06 40.538 41.22 ;
        RECT 42.262 0.06 42.338 41.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 41.22 ;
        RECT 3.562 0.06 3.638 41.22 ;
        RECT 5.362 0.06 5.438 41.22 ;
        RECT 7.162 0.06 7.238 41.22 ;
        RECT 8.962 0.06 9.038 41.22 ;
        RECT 10.762 0.06 10.838 41.22 ;
        RECT 12.562 0.06 12.638 41.22 ;
        RECT 14.362 0.06 14.438 41.22 ;
        RECT 16.162 0.06 16.238 41.22 ;
        RECT 17.962 0.06 18.038 41.22 ;
        RECT 19.762 0.06 19.838 41.22 ;
        RECT 21.562 0.06 21.638 41.22 ;
        RECT 23.362 0.06 23.438 41.22 ;
        RECT 25.162 0.06 25.238 41.22 ;
        RECT 26.962 0.06 27.038 41.22 ;
        RECT 28.762 0.06 28.838 41.22 ;
        RECT 30.562 0.06 30.638 41.22 ;
        RECT 32.362 0.06 32.438 41.22 ;
        RECT 34.162 0.06 34.238 41.22 ;
        RECT 35.962 0.06 36.038 41.22 ;
        RECT 37.762 0.06 37.838 41.22 ;
        RECT 39.562 0.06 39.638 41.22 ;
        RECT 41.362 0.06 41.438 41.22 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 43.216 41.294 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 43.22 41.3 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 43.2705 41.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 43.235 41.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 43.27 41.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 43.259 41.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 43.29 41.342 ;
    LAYER m7 SPACING 0 ;
      RECT 42.338 41.34 43.24 41.4 ;
      RECT 42.338 -0.06 43.292 41.34 ;
      RECT 42.338 -0.12 43.24 -0.06 ;
      RECT 41.438 -0.12 42.262 41.4 ;
      RECT 40.538 -0.12 41.362 41.4 ;
      RECT 39.638 -0.12 40.462 41.4 ;
      RECT 38.738 -0.12 39.562 41.4 ;
      RECT 37.838 -0.12 38.662 41.4 ;
      RECT 36.938 -0.12 37.762 41.4 ;
      RECT 36.038 -0.12 36.862 41.4 ;
      RECT 35.138 -0.12 35.962 41.4 ;
      RECT 34.238 -0.12 35.062 41.4 ;
      RECT 33.338 -0.12 34.162 41.4 ;
      RECT 32.438 -0.12 33.262 41.4 ;
      RECT 31.538 -0.12 32.362 41.4 ;
      RECT 30.638 -0.12 31.462 41.4 ;
      RECT 29.738 -0.12 30.562 41.4 ;
      RECT 28.838 -0.12 29.662 41.4 ;
      RECT 27.938 -0.12 28.762 41.4 ;
      RECT 27.038 -0.12 27.862 41.4 ;
      RECT 26.138 -0.12 26.962 41.4 ;
      RECT 25.238 -0.12 26.062 41.4 ;
      RECT 24.338 -0.12 25.162 41.4 ;
      RECT 23.438 41.04 24.262 41.4 ;
      RECT 23.438 39.84 23.572 41.04 ;
      RECT 23.616 39.84 23.828 41.04 ;
      RECT 23.872 39.84 24.262 41.04 ;
      RECT 23.438 38.88 24.262 39.84 ;
      RECT 23.438 37.68 23.572 38.88 ;
      RECT 23.616 37.68 23.828 38.88 ;
      RECT 23.872 37.68 24.262 38.88 ;
      RECT 23.438 36.72 24.262 37.68 ;
      RECT 23.438 35.52 23.572 36.72 ;
      RECT 23.616 35.52 23.828 36.72 ;
      RECT 23.872 35.52 24.262 36.72 ;
      RECT 23.438 34.56 24.262 35.52 ;
      RECT 23.438 33.36 23.572 34.56 ;
      RECT 23.616 33.36 23.828 34.56 ;
      RECT 23.872 33.36 24.262 34.56 ;
      RECT 23.438 32.4 24.262 33.36 ;
      RECT 23.438 31.2 23.572 32.4 ;
      RECT 23.616 31.2 23.828 32.4 ;
      RECT 23.872 31.2 24.262 32.4 ;
      RECT 23.438 30.24 24.262 31.2 ;
      RECT 23.438 29.04 23.572 30.24 ;
      RECT 23.616 29.04 23.828 30.24 ;
      RECT 23.872 29.04 24.262 30.24 ;
      RECT 23.438 28.08 24.262 29.04 ;
      RECT 23.438 26.88 23.572 28.08 ;
      RECT 23.616 26.88 23.828 28.08 ;
      RECT 23.872 26.88 24.262 28.08 ;
      RECT 23.438 25.92 24.262 26.88 ;
      RECT 23.438 24.72 23.572 25.92 ;
      RECT 23.616 24.72 23.828 25.92 ;
      RECT 23.872 24.72 24.262 25.92 ;
      RECT 23.438 23.64 24.262 24.72 ;
      RECT 23.438 22.44 23.484 23.64 ;
      RECT 23.528 22.44 23.572 23.64 ;
      RECT 23.616 22.44 23.828 23.64 ;
      RECT 23.872 22.44 24.262 23.64 ;
      RECT 23.438 18.72 24.262 22.44 ;
      RECT 23.438 17.52 23.572 18.72 ;
      RECT 23.616 17.52 23.828 18.72 ;
      RECT 23.872 17.52 24.262 18.72 ;
      RECT 23.438 16.56 24.262 17.52 ;
      RECT 23.438 15.36 23.572 16.56 ;
      RECT 23.616 15.36 23.828 16.56 ;
      RECT 23.872 15.36 24.262 16.56 ;
      RECT 23.438 14.4 24.262 15.36 ;
      RECT 23.438 13.2 23.572 14.4 ;
      RECT 23.616 13.2 23.828 14.4 ;
      RECT 23.872 13.2 24.262 14.4 ;
      RECT 23.438 12.24 24.262 13.2 ;
      RECT 23.438 11.04 23.572 12.24 ;
      RECT 23.616 11.04 23.828 12.24 ;
      RECT 23.872 11.04 24.262 12.24 ;
      RECT 23.438 10.08 24.262 11.04 ;
      RECT 23.438 8.88 23.572 10.08 ;
      RECT 23.616 8.88 23.828 10.08 ;
      RECT 23.872 8.88 24.262 10.08 ;
      RECT 23.438 7.92 24.262 8.88 ;
      RECT 23.438 6.72 23.572 7.92 ;
      RECT 23.616 6.72 23.828 7.92 ;
      RECT 23.872 6.72 24.262 7.92 ;
      RECT 23.438 5.76 24.262 6.72 ;
      RECT 23.438 4.56 23.572 5.76 ;
      RECT 23.616 4.56 23.828 5.76 ;
      RECT 23.872 4.56 24.262 5.76 ;
      RECT 23.438 3.6 24.262 4.56 ;
      RECT 23.438 2.4 23.572 3.6 ;
      RECT 23.616 2.4 23.828 3.6 ;
      RECT 23.872 2.4 24.262 3.6 ;
      RECT 23.438 1.44 24.262 2.4 ;
      RECT 23.438 0.24 23.572 1.44 ;
      RECT 23.616 0.24 23.828 1.44 ;
      RECT 23.872 0.24 24.262 1.44 ;
      RECT 23.438 -0.12 24.262 0.24 ;
      RECT 22.538 40.32 23.362 41.4 ;
      RECT 22.716 39.6 23.272 40.32 ;
      RECT 22.538 39.12 22.672 40.32 ;
      RECT 23.316 39.12 23.362 40.32 ;
      RECT 22.716 39.12 22.928 39.6 ;
      RECT 23.228 39.12 23.272 39.6 ;
      RECT 22.972 38.4 23.184 39.6 ;
      RECT 22.538 38.4 22.928 39.12 ;
      RECT 23.228 38.4 23.362 39.12 ;
      RECT 22.538 38.16 23.362 38.4 ;
      RECT 22.716 37.44 23.272 38.16 ;
      RECT 22.538 36.96 22.672 38.16 ;
      RECT 23.316 36.96 23.362 38.16 ;
      RECT 22.716 36.96 22.928 37.44 ;
      RECT 23.228 36.96 23.272 37.44 ;
      RECT 22.972 36.24 23.184 37.44 ;
      RECT 22.538 36.24 22.928 36.96 ;
      RECT 23.228 36.24 23.362 36.96 ;
      RECT 22.538 36 23.362 36.24 ;
      RECT 22.716 35.28 23.272 36 ;
      RECT 22.538 34.8 22.672 36 ;
      RECT 23.316 34.8 23.362 36 ;
      RECT 22.716 34.8 22.928 35.28 ;
      RECT 23.228 34.8 23.272 35.28 ;
      RECT 22.972 34.08 23.184 35.28 ;
      RECT 22.538 34.08 22.928 34.8 ;
      RECT 23.228 34.08 23.362 34.8 ;
      RECT 22.538 33.84 23.362 34.08 ;
      RECT 22.716 33.12 23.272 33.84 ;
      RECT 22.538 32.64 22.672 33.84 ;
      RECT 23.316 32.64 23.362 33.84 ;
      RECT 22.716 32.64 22.928 33.12 ;
      RECT 23.228 32.64 23.272 33.12 ;
      RECT 22.972 31.92 23.184 33.12 ;
      RECT 22.538 31.92 22.928 32.64 ;
      RECT 23.228 31.92 23.362 32.64 ;
      RECT 22.538 31.68 23.362 31.92 ;
      RECT 22.716 30.96 23.272 31.68 ;
      RECT 22.538 30.48 22.672 31.68 ;
      RECT 23.316 30.48 23.362 31.68 ;
      RECT 22.716 30.48 22.928 30.96 ;
      RECT 23.228 30.48 23.272 30.96 ;
      RECT 22.972 29.76 23.184 30.96 ;
      RECT 22.538 29.76 22.928 30.48 ;
      RECT 23.228 29.76 23.362 30.48 ;
      RECT 22.538 29.52 23.362 29.76 ;
      RECT 22.716 28.8 23.272 29.52 ;
      RECT 22.538 28.32 22.672 29.52 ;
      RECT 23.316 28.32 23.362 29.52 ;
      RECT 22.716 28.32 22.928 28.8 ;
      RECT 23.228 28.32 23.272 28.8 ;
      RECT 22.972 27.6 23.184 28.8 ;
      RECT 22.538 27.6 22.928 28.32 ;
      RECT 23.228 27.6 23.362 28.32 ;
      RECT 22.538 27.36 23.362 27.6 ;
      RECT 22.716 26.64 23.272 27.36 ;
      RECT 22.538 26.16 22.672 27.36 ;
      RECT 23.316 26.16 23.362 27.36 ;
      RECT 22.716 26.16 22.928 26.64 ;
      RECT 23.228 26.16 23.272 26.64 ;
      RECT 22.972 25.44 23.184 26.64 ;
      RECT 22.538 25.44 22.928 26.16 ;
      RECT 23.228 25.44 23.362 26.16 ;
      RECT 22.538 25.2 23.362 25.44 ;
      RECT 22.538 24 22.672 25.2 ;
      RECT 22.716 24 23.272 25.2 ;
      RECT 23.316 24 23.362 25.2 ;
      RECT 22.538 23.64 23.362 24 ;
      RECT 22.538 22.44 22.584 23.64 ;
      RECT 22.628 22.44 22.928 23.64 ;
      RECT 22.972 22.44 23.184 23.64 ;
      RECT 23.228 22.44 23.362 23.64 ;
      RECT 22.538 20.16 23.362 22.44 ;
      RECT 22.716 19.44 23.272 20.16 ;
      RECT 22.538 18.96 22.672 20.16 ;
      RECT 23.316 18.96 23.362 20.16 ;
      RECT 22.716 18.96 22.928 19.44 ;
      RECT 23.228 18.96 23.272 19.44 ;
      RECT 22.972 18.24 23.184 19.44 ;
      RECT 22.538 18.24 22.928 18.96 ;
      RECT 23.228 18.24 23.362 18.96 ;
      RECT 22.538 18 23.362 18.24 ;
      RECT 22.716 17.28 23.272 18 ;
      RECT 22.538 16.8 22.672 18 ;
      RECT 23.316 16.8 23.362 18 ;
      RECT 22.716 16.8 22.928 17.28 ;
      RECT 23.228 16.8 23.272 17.28 ;
      RECT 22.972 16.08 23.184 17.28 ;
      RECT 22.538 16.08 22.928 16.8 ;
      RECT 23.228 16.08 23.362 16.8 ;
      RECT 22.538 15.84 23.362 16.08 ;
      RECT 22.716 15.12 23.272 15.84 ;
      RECT 22.538 14.64 22.672 15.84 ;
      RECT 23.316 14.64 23.362 15.84 ;
      RECT 22.716 14.64 22.928 15.12 ;
      RECT 23.228 14.64 23.272 15.12 ;
      RECT 22.972 13.92 23.184 15.12 ;
      RECT 22.538 13.92 22.928 14.64 ;
      RECT 23.228 13.92 23.362 14.64 ;
      RECT 22.538 13.68 23.362 13.92 ;
      RECT 22.716 12.96 23.272 13.68 ;
      RECT 22.538 12.48 22.672 13.68 ;
      RECT 23.316 12.48 23.362 13.68 ;
      RECT 22.716 12.48 22.928 12.96 ;
      RECT 23.228 12.48 23.272 12.96 ;
      RECT 22.972 11.76 23.184 12.96 ;
      RECT 22.538 11.76 22.928 12.48 ;
      RECT 23.228 11.76 23.362 12.48 ;
      RECT 22.538 11.52 23.362 11.76 ;
      RECT 22.716 10.8 23.272 11.52 ;
      RECT 22.538 10.32 22.672 11.52 ;
      RECT 23.316 10.32 23.362 11.52 ;
      RECT 22.716 10.32 22.928 10.8 ;
      RECT 23.228 10.32 23.272 10.8 ;
      RECT 22.972 9.6 23.184 10.8 ;
      RECT 22.538 9.6 22.928 10.32 ;
      RECT 23.228 9.6 23.362 10.32 ;
      RECT 22.538 9.36 23.362 9.6 ;
      RECT 22.716 8.64 23.272 9.36 ;
      RECT 22.538 8.16 22.672 9.36 ;
      RECT 23.316 8.16 23.362 9.36 ;
      RECT 22.716 8.16 22.928 8.64 ;
      RECT 23.228 8.16 23.272 8.64 ;
      RECT 22.972 7.44 23.184 8.64 ;
      RECT 22.538 7.44 22.928 8.16 ;
      RECT 23.228 7.44 23.362 8.16 ;
      RECT 22.538 7.2 23.362 7.44 ;
      RECT 22.716 6.48 23.272 7.2 ;
      RECT 22.538 6 22.672 7.2 ;
      RECT 23.316 6 23.362 7.2 ;
      RECT 22.716 6 22.928 6.48 ;
      RECT 23.228 6 23.272 6.48 ;
      RECT 22.972 5.28 23.184 6.48 ;
      RECT 22.538 5.28 22.928 6 ;
      RECT 23.228 5.28 23.362 6 ;
      RECT 22.538 5.04 23.362 5.28 ;
      RECT 22.716 4.32 23.272 5.04 ;
      RECT 22.538 3.84 22.672 5.04 ;
      RECT 23.316 3.84 23.362 5.04 ;
      RECT 22.716 3.84 22.928 4.32 ;
      RECT 23.228 3.84 23.272 4.32 ;
      RECT 22.972 3.12 23.184 4.32 ;
      RECT 22.538 3.12 22.928 3.84 ;
      RECT 23.228 3.12 23.362 3.84 ;
      RECT 22.538 2.88 23.362 3.12 ;
      RECT 22.716 2.16 23.272 2.88 ;
      RECT 22.538 1.68 22.672 2.88 ;
      RECT 23.316 1.68 23.362 2.88 ;
      RECT 22.716 1.68 22.928 2.16 ;
      RECT 23.228 1.68 23.272 2.16 ;
      RECT 22.972 0.96 23.184 2.16 ;
      RECT 22.538 0.96 22.928 1.68 ;
      RECT 23.228 0.96 23.362 1.68 ;
      RECT 22.538 -0.12 23.362 0.96 ;
      RECT 21.638 41.04 22.462 41.4 ;
      RECT 21.638 40.32 21.772 41.04 ;
      RECT 22.072 40.32 22.462 41.04 ;
      RECT 21.816 39.84 22.028 41.04 ;
      RECT 21.728 39.84 21.772 40.32 ;
      RECT 22.072 39.84 22.284 40.32 ;
      RECT 21.638 39.12 21.684 40.32 ;
      RECT 22.328 39.12 22.462 40.32 ;
      RECT 21.728 39.12 22.284 39.84 ;
      RECT 21.638 38.88 22.462 39.12 ;
      RECT 21.638 38.16 21.772 38.88 ;
      RECT 22.072 38.16 22.462 38.88 ;
      RECT 21.816 37.68 22.028 38.88 ;
      RECT 21.728 37.68 21.772 38.16 ;
      RECT 22.072 37.68 22.284 38.16 ;
      RECT 21.638 36.96 21.684 38.16 ;
      RECT 22.328 36.96 22.462 38.16 ;
      RECT 21.728 36.96 22.284 37.68 ;
      RECT 21.638 36.72 22.462 36.96 ;
      RECT 21.638 36 21.772 36.72 ;
      RECT 22.072 36 22.462 36.72 ;
      RECT 21.816 35.52 22.028 36.72 ;
      RECT 21.728 35.52 21.772 36 ;
      RECT 22.072 35.52 22.284 36 ;
      RECT 21.638 34.8 21.684 36 ;
      RECT 22.328 34.8 22.462 36 ;
      RECT 21.728 34.8 22.284 35.52 ;
      RECT 21.638 34.56 22.462 34.8 ;
      RECT 21.638 33.84 21.772 34.56 ;
      RECT 22.072 33.84 22.462 34.56 ;
      RECT 21.816 33.36 22.028 34.56 ;
      RECT 21.728 33.36 21.772 33.84 ;
      RECT 22.072 33.36 22.284 33.84 ;
      RECT 21.638 32.64 21.684 33.84 ;
      RECT 22.328 32.64 22.462 33.84 ;
      RECT 21.728 32.64 22.284 33.36 ;
      RECT 21.638 32.4 22.462 32.64 ;
      RECT 21.638 31.68 21.772 32.4 ;
      RECT 22.072 31.68 22.462 32.4 ;
      RECT 21.816 31.2 22.028 32.4 ;
      RECT 21.728 31.2 21.772 31.68 ;
      RECT 22.072 31.2 22.284 31.68 ;
      RECT 21.638 30.48 21.684 31.68 ;
      RECT 22.328 30.48 22.462 31.68 ;
      RECT 21.728 30.48 22.284 31.2 ;
      RECT 21.638 30.24 22.462 30.48 ;
      RECT 21.638 29.52 21.772 30.24 ;
      RECT 22.072 29.52 22.462 30.24 ;
      RECT 21.816 29.04 22.028 30.24 ;
      RECT 21.728 29.04 21.772 29.52 ;
      RECT 22.072 29.04 22.284 29.52 ;
      RECT 21.638 28.32 21.684 29.52 ;
      RECT 22.328 28.32 22.462 29.52 ;
      RECT 21.728 28.32 22.284 29.04 ;
      RECT 21.638 28.08 22.462 28.32 ;
      RECT 21.638 27.36 21.772 28.08 ;
      RECT 22.072 27.36 22.462 28.08 ;
      RECT 21.816 26.88 22.028 28.08 ;
      RECT 21.728 26.88 21.772 27.36 ;
      RECT 22.072 26.88 22.284 27.36 ;
      RECT 21.638 26.16 21.684 27.36 ;
      RECT 22.328 26.16 22.462 27.36 ;
      RECT 21.728 26.16 22.284 26.88 ;
      RECT 21.638 25.92 22.462 26.16 ;
      RECT 21.816 25.2 22.462 25.92 ;
      RECT 21.638 24.72 21.684 25.92 ;
      RECT 21.728 24.72 21.772 25.92 ;
      RECT 21.816 24.72 22.028 25.2 ;
      RECT 22.072 24 22.284 25.2 ;
      RECT 22.328 24 22.462 25.2 ;
      RECT 21.638 24 22.028 24.72 ;
      RECT 21.638 23.64 22.462 24 ;
      RECT 21.638 22.44 22.372 23.64 ;
      RECT 22.416 22.44 22.462 23.64 ;
      RECT 21.638 21.72 22.462 22.44 ;
      RECT 21.638 20.52 21.772 21.72 ;
      RECT 21.816 20.52 22.028 21.72 ;
      RECT 22.072 20.52 22.462 21.72 ;
      RECT 21.638 20.16 22.462 20.52 ;
      RECT 21.638 18.96 21.684 20.16 ;
      RECT 21.728 18.96 22.284 20.16 ;
      RECT 22.328 18.96 22.462 20.16 ;
      RECT 21.638 18.72 22.462 18.96 ;
      RECT 21.638 18 21.772 18.72 ;
      RECT 22.072 18 22.462 18.72 ;
      RECT 21.816 17.52 22.028 18.72 ;
      RECT 21.728 17.52 21.772 18 ;
      RECT 22.072 17.52 22.284 18 ;
      RECT 21.638 16.8 21.684 18 ;
      RECT 22.328 16.8 22.462 18 ;
      RECT 21.728 16.8 22.284 17.52 ;
      RECT 21.638 16.56 22.462 16.8 ;
      RECT 21.638 15.84 21.772 16.56 ;
      RECT 22.072 15.84 22.462 16.56 ;
      RECT 21.816 15.36 22.028 16.56 ;
      RECT 21.728 15.36 21.772 15.84 ;
      RECT 22.072 15.36 22.284 15.84 ;
      RECT 21.638 14.64 21.684 15.84 ;
      RECT 22.328 14.64 22.462 15.84 ;
      RECT 21.728 14.64 22.284 15.36 ;
      RECT 21.638 14.4 22.462 14.64 ;
      RECT 21.638 13.68 21.772 14.4 ;
      RECT 22.072 13.68 22.462 14.4 ;
      RECT 21.816 13.2 22.028 14.4 ;
      RECT 21.728 13.2 21.772 13.68 ;
      RECT 22.072 13.2 22.284 13.68 ;
      RECT 21.638 12.48 21.684 13.68 ;
      RECT 22.328 12.48 22.462 13.68 ;
      RECT 21.728 12.48 22.284 13.2 ;
      RECT 21.638 12.24 22.462 12.48 ;
      RECT 21.638 11.52 21.772 12.24 ;
      RECT 22.072 11.52 22.462 12.24 ;
      RECT 21.816 11.04 22.028 12.24 ;
      RECT 21.728 11.04 21.772 11.52 ;
      RECT 22.072 11.04 22.284 11.52 ;
      RECT 21.638 10.32 21.684 11.52 ;
      RECT 22.328 10.32 22.462 11.52 ;
      RECT 21.728 10.32 22.284 11.04 ;
      RECT 21.638 10.08 22.462 10.32 ;
      RECT 21.638 9.36 21.772 10.08 ;
      RECT 22.072 9.36 22.462 10.08 ;
      RECT 21.816 8.88 22.028 10.08 ;
      RECT 21.728 8.88 21.772 9.36 ;
      RECT 22.072 8.88 22.284 9.36 ;
      RECT 21.638 8.16 21.684 9.36 ;
      RECT 22.328 8.16 22.462 9.36 ;
      RECT 21.728 8.16 22.284 8.88 ;
      RECT 21.638 7.92 22.462 8.16 ;
      RECT 21.638 7.2 21.772 7.92 ;
      RECT 22.072 7.2 22.462 7.92 ;
      RECT 21.816 6.72 22.028 7.92 ;
      RECT 21.728 6.72 21.772 7.2 ;
      RECT 22.072 6.72 22.284 7.2 ;
      RECT 21.638 6 21.684 7.2 ;
      RECT 22.328 6 22.462 7.2 ;
      RECT 21.728 6 22.284 6.72 ;
      RECT 21.638 5.76 22.462 6 ;
      RECT 21.638 5.04 21.772 5.76 ;
      RECT 22.072 5.04 22.462 5.76 ;
      RECT 21.816 4.56 22.028 5.76 ;
      RECT 21.728 4.56 21.772 5.04 ;
      RECT 22.072 4.56 22.284 5.04 ;
      RECT 21.638 3.84 21.684 5.04 ;
      RECT 22.328 3.84 22.462 5.04 ;
      RECT 21.728 3.84 22.284 4.56 ;
      RECT 21.638 3.6 22.462 3.84 ;
      RECT 21.638 2.88 21.772 3.6 ;
      RECT 22.072 2.88 22.462 3.6 ;
      RECT 21.816 2.4 22.028 3.6 ;
      RECT 21.728 2.4 21.772 2.88 ;
      RECT 22.072 2.4 22.284 2.88 ;
      RECT 21.638 1.68 21.684 2.88 ;
      RECT 22.328 1.68 22.462 2.88 ;
      RECT 21.728 1.68 22.284 2.4 ;
      RECT 21.638 1.44 22.462 1.68 ;
      RECT 21.638 0.24 22.028 1.44 ;
      RECT 22.072 0.24 22.284 1.44 ;
      RECT 22.328 0.24 22.462 1.44 ;
      RECT 21.638 -0.12 22.462 0.24 ;
      RECT 20.738 41.04 21.562 41.4 ;
      RECT 20.738 39.84 20.784 41.04 ;
      RECT 20.828 39.84 21.562 41.04 ;
      RECT 20.738 39.6 21.562 39.84 ;
      RECT 20.738 38.88 20.872 39.6 ;
      RECT 20.916 38.4 21.128 39.6 ;
      RECT 21.172 38.4 21.384 39.6 ;
      RECT 21.428 38.4 21.472 39.6 ;
      RECT 21.516 38.4 21.562 39.6 ;
      RECT 20.828 38.4 20.872 38.88 ;
      RECT 20.738 37.68 20.784 38.88 ;
      RECT 20.828 37.68 21.562 38.4 ;
      RECT 20.738 37.44 21.562 37.68 ;
      RECT 20.738 36.72 20.872 37.44 ;
      RECT 20.916 36.24 21.128 37.44 ;
      RECT 21.172 36.24 21.384 37.44 ;
      RECT 21.428 36.24 21.472 37.44 ;
      RECT 21.516 36.24 21.562 37.44 ;
      RECT 20.828 36.24 20.872 36.72 ;
      RECT 20.738 35.52 20.784 36.72 ;
      RECT 20.828 35.52 21.562 36.24 ;
      RECT 20.738 35.28 21.562 35.52 ;
      RECT 20.738 34.56 20.872 35.28 ;
      RECT 20.916 34.08 21.128 35.28 ;
      RECT 21.172 34.08 21.384 35.28 ;
      RECT 21.428 34.08 21.472 35.28 ;
      RECT 21.516 34.08 21.562 35.28 ;
      RECT 20.828 34.08 20.872 34.56 ;
      RECT 20.738 33.36 20.784 34.56 ;
      RECT 20.828 33.36 21.562 34.08 ;
      RECT 20.738 33.12 21.562 33.36 ;
      RECT 20.738 32.4 20.872 33.12 ;
      RECT 20.916 31.92 21.128 33.12 ;
      RECT 21.172 31.92 21.384 33.12 ;
      RECT 21.428 31.92 21.472 33.12 ;
      RECT 21.516 31.92 21.562 33.12 ;
      RECT 20.828 31.92 20.872 32.4 ;
      RECT 20.738 31.2 20.784 32.4 ;
      RECT 20.828 31.2 21.562 31.92 ;
      RECT 20.738 30.96 21.562 31.2 ;
      RECT 20.738 30.24 20.872 30.96 ;
      RECT 20.916 29.76 21.128 30.96 ;
      RECT 21.172 29.76 21.384 30.96 ;
      RECT 21.428 29.76 21.472 30.96 ;
      RECT 21.516 29.76 21.562 30.96 ;
      RECT 20.828 29.76 20.872 30.24 ;
      RECT 20.738 29.04 20.784 30.24 ;
      RECT 20.828 29.04 21.562 29.76 ;
      RECT 20.738 28.8 21.562 29.04 ;
      RECT 20.738 28.08 20.872 28.8 ;
      RECT 20.916 27.6 21.128 28.8 ;
      RECT 21.172 27.6 21.384 28.8 ;
      RECT 21.428 27.6 21.472 28.8 ;
      RECT 21.516 27.6 21.562 28.8 ;
      RECT 20.828 27.6 20.872 28.08 ;
      RECT 20.738 26.88 20.784 28.08 ;
      RECT 20.828 26.88 21.562 27.6 ;
      RECT 20.738 26.64 21.562 26.88 ;
      RECT 20.738 25.44 20.872 26.64 ;
      RECT 20.916 25.44 21.128 26.64 ;
      RECT 21.172 25.44 21.384 26.64 ;
      RECT 21.428 25.44 21.472 26.64 ;
      RECT 21.516 25.44 21.562 26.64 ;
      RECT 20.738 25.2 21.562 25.44 ;
      RECT 20.738 24 20.784 25.2 ;
      RECT 20.828 24 21.562 25.2 ;
      RECT 20.738 21.72 21.562 24 ;
      RECT 20.738 20.52 20.784 21.72 ;
      RECT 20.828 20.52 20.872 21.72 ;
      RECT 20.916 20.52 21.128 21.72 ;
      RECT 21.172 20.52 21.384 21.72 ;
      RECT 21.428 20.52 21.472 21.72 ;
      RECT 21.516 20.52 21.562 21.72 ;
      RECT 20.738 19.44 21.562 20.52 ;
      RECT 20.738 18.72 20.872 19.44 ;
      RECT 20.916 18.24 21.128 19.44 ;
      RECT 21.172 18.24 21.384 19.44 ;
      RECT 21.428 18.24 21.472 19.44 ;
      RECT 21.516 18.24 21.562 19.44 ;
      RECT 20.828 18.24 20.872 18.72 ;
      RECT 20.738 17.52 20.784 18.72 ;
      RECT 20.828 17.52 21.562 18.24 ;
      RECT 20.738 17.28 21.562 17.52 ;
      RECT 20.738 16.56 20.872 17.28 ;
      RECT 20.916 16.08 21.128 17.28 ;
      RECT 21.172 16.08 21.384 17.28 ;
      RECT 21.428 16.08 21.472 17.28 ;
      RECT 21.516 16.08 21.562 17.28 ;
      RECT 20.828 16.08 20.872 16.56 ;
      RECT 20.738 15.36 20.784 16.56 ;
      RECT 20.828 15.36 21.562 16.08 ;
      RECT 20.738 15.12 21.562 15.36 ;
      RECT 20.738 14.4 20.872 15.12 ;
      RECT 20.916 13.92 21.128 15.12 ;
      RECT 21.172 13.92 21.384 15.12 ;
      RECT 21.428 13.92 21.472 15.12 ;
      RECT 21.516 13.92 21.562 15.12 ;
      RECT 20.828 13.92 20.872 14.4 ;
      RECT 20.738 13.2 20.784 14.4 ;
      RECT 20.828 13.2 21.562 13.92 ;
      RECT 20.738 12.96 21.562 13.2 ;
      RECT 20.738 12.24 20.872 12.96 ;
      RECT 20.916 11.76 21.128 12.96 ;
      RECT 21.172 11.76 21.384 12.96 ;
      RECT 21.428 11.76 21.472 12.96 ;
      RECT 21.516 11.76 21.562 12.96 ;
      RECT 20.828 11.76 20.872 12.24 ;
      RECT 20.738 11.04 20.784 12.24 ;
      RECT 20.828 11.04 21.562 11.76 ;
      RECT 20.738 10.8 21.562 11.04 ;
      RECT 20.738 10.08 20.872 10.8 ;
      RECT 20.916 9.6 21.128 10.8 ;
      RECT 21.172 9.6 21.384 10.8 ;
      RECT 21.428 9.6 21.472 10.8 ;
      RECT 21.516 9.6 21.562 10.8 ;
      RECT 20.828 9.6 20.872 10.08 ;
      RECT 20.738 8.88 20.784 10.08 ;
      RECT 20.828 8.88 21.562 9.6 ;
      RECT 20.738 8.64 21.562 8.88 ;
      RECT 20.738 7.92 20.872 8.64 ;
      RECT 20.916 7.44 21.128 8.64 ;
      RECT 21.172 7.44 21.384 8.64 ;
      RECT 21.428 7.44 21.472 8.64 ;
      RECT 21.516 7.44 21.562 8.64 ;
      RECT 20.828 7.44 20.872 7.92 ;
      RECT 20.738 6.72 20.784 7.92 ;
      RECT 20.828 6.72 21.562 7.44 ;
      RECT 20.738 6.48 21.562 6.72 ;
      RECT 20.738 5.76 20.872 6.48 ;
      RECT 20.916 5.28 21.128 6.48 ;
      RECT 21.172 5.28 21.384 6.48 ;
      RECT 21.428 5.28 21.472 6.48 ;
      RECT 21.516 5.28 21.562 6.48 ;
      RECT 20.828 5.28 20.872 5.76 ;
      RECT 20.738 4.56 20.784 5.76 ;
      RECT 20.828 4.56 21.562 5.28 ;
      RECT 20.738 4.32 21.562 4.56 ;
      RECT 20.738 3.6 20.872 4.32 ;
      RECT 20.916 3.12 21.128 4.32 ;
      RECT 21.172 3.12 21.384 4.32 ;
      RECT 21.428 3.12 21.472 4.32 ;
      RECT 21.516 3.12 21.562 4.32 ;
      RECT 20.828 3.12 20.872 3.6 ;
      RECT 20.738 2.4 20.784 3.6 ;
      RECT 20.828 2.4 21.562 3.12 ;
      RECT 20.738 2.16 21.562 2.4 ;
      RECT 20.738 1.44 20.872 2.16 ;
      RECT 20.916 0.96 21.128 2.16 ;
      RECT 21.172 0.96 21.384 2.16 ;
      RECT 21.428 0.96 21.472 2.16 ;
      RECT 21.516 0.96 21.562 2.16 ;
      RECT 20.828 0.96 20.872 1.44 ;
      RECT 20.738 0.24 20.784 1.44 ;
      RECT 20.828 0.24 21.562 0.96 ;
      RECT 20.738 -0.12 21.562 0.24 ;
      RECT 19.838 41.04 20.662 41.4 ;
      RECT 20.272 40.32 20.662 41.04 ;
      RECT 19.838 39.84 20.228 41.04 ;
      RECT 20.272 39.84 20.484 40.32 ;
      RECT 20.528 39.12 20.572 40.32 ;
      RECT 20.616 39.12 20.662 40.32 ;
      RECT 19.838 39.12 20.484 39.84 ;
      RECT 19.838 38.88 20.662 39.12 ;
      RECT 20.272 38.16 20.662 38.88 ;
      RECT 19.838 37.68 20.228 38.88 ;
      RECT 20.272 37.68 20.484 38.16 ;
      RECT 20.528 36.96 20.572 38.16 ;
      RECT 20.616 36.96 20.662 38.16 ;
      RECT 19.838 36.96 20.484 37.68 ;
      RECT 19.838 36.72 20.662 36.96 ;
      RECT 20.272 36 20.662 36.72 ;
      RECT 19.838 35.52 20.228 36.72 ;
      RECT 20.272 35.52 20.484 36 ;
      RECT 20.528 34.8 20.572 36 ;
      RECT 20.616 34.8 20.662 36 ;
      RECT 19.838 34.8 20.484 35.52 ;
      RECT 19.838 34.56 20.662 34.8 ;
      RECT 20.272 33.84 20.662 34.56 ;
      RECT 19.838 33.36 20.228 34.56 ;
      RECT 20.272 33.36 20.484 33.84 ;
      RECT 20.528 32.64 20.572 33.84 ;
      RECT 20.616 32.64 20.662 33.84 ;
      RECT 19.838 32.64 20.484 33.36 ;
      RECT 19.838 32.4 20.662 32.64 ;
      RECT 20.272 31.68 20.662 32.4 ;
      RECT 19.838 31.2 20.228 32.4 ;
      RECT 20.272 31.2 20.484 31.68 ;
      RECT 20.528 30.48 20.572 31.68 ;
      RECT 20.616 30.48 20.662 31.68 ;
      RECT 19.838 30.48 20.484 31.2 ;
      RECT 19.838 30.24 20.662 30.48 ;
      RECT 20.272 29.52 20.662 30.24 ;
      RECT 19.838 29.04 20.228 30.24 ;
      RECT 20.272 29.04 20.484 29.52 ;
      RECT 20.528 28.32 20.572 29.52 ;
      RECT 20.616 28.32 20.662 29.52 ;
      RECT 19.838 28.32 20.484 29.04 ;
      RECT 19.838 28.08 20.662 28.32 ;
      RECT 20.272 27.36 20.662 28.08 ;
      RECT 19.838 26.88 20.228 28.08 ;
      RECT 20.272 26.88 20.484 27.36 ;
      RECT 20.528 26.16 20.572 27.36 ;
      RECT 20.616 26.16 20.662 27.36 ;
      RECT 19.838 26.16 20.484 26.88 ;
      RECT 19.838 25.92 20.662 26.16 ;
      RECT 20.528 25.2 20.662 25.92 ;
      RECT 19.838 24.72 20.228 25.92 ;
      RECT 20.272 24.72 20.484 25.92 ;
      RECT 20.528 24.72 20.572 25.2 ;
      RECT 20.616 24 20.662 25.2 ;
      RECT 19.838 24 20.572 24.72 ;
      RECT 19.838 21.72 20.662 24 ;
      RECT 19.838 20.52 19.884 21.72 ;
      RECT 19.928 20.52 19.972 21.72 ;
      RECT 20.016 20.52 20.228 21.72 ;
      RECT 20.272 20.52 20.662 21.72 ;
      RECT 19.838 20.16 20.662 20.52 ;
      RECT 19.838 18.96 20.484 20.16 ;
      RECT 20.528 18.96 20.572 20.16 ;
      RECT 20.616 18.96 20.662 20.16 ;
      RECT 19.838 18.72 20.662 18.96 ;
      RECT 20.272 18 20.662 18.72 ;
      RECT 19.838 17.52 20.228 18.72 ;
      RECT 20.272 17.52 20.484 18 ;
      RECT 20.528 16.8 20.572 18 ;
      RECT 20.616 16.8 20.662 18 ;
      RECT 19.838 16.8 20.484 17.52 ;
      RECT 19.838 16.56 20.662 16.8 ;
      RECT 20.272 15.84 20.662 16.56 ;
      RECT 19.838 15.36 20.228 16.56 ;
      RECT 20.272 15.36 20.484 15.84 ;
      RECT 20.528 14.64 20.572 15.84 ;
      RECT 20.616 14.64 20.662 15.84 ;
      RECT 19.838 14.64 20.484 15.36 ;
      RECT 19.838 14.4 20.662 14.64 ;
      RECT 20.272 13.68 20.662 14.4 ;
      RECT 19.838 13.2 20.228 14.4 ;
      RECT 20.272 13.2 20.484 13.68 ;
      RECT 20.528 12.48 20.572 13.68 ;
      RECT 20.616 12.48 20.662 13.68 ;
      RECT 19.838 12.48 20.484 13.2 ;
      RECT 19.838 12.24 20.662 12.48 ;
      RECT 20.272 11.52 20.662 12.24 ;
      RECT 19.838 11.04 20.228 12.24 ;
      RECT 20.272 11.04 20.484 11.52 ;
      RECT 20.528 10.32 20.572 11.52 ;
      RECT 20.616 10.32 20.662 11.52 ;
      RECT 19.838 10.32 20.484 11.04 ;
      RECT 19.838 10.08 20.662 10.32 ;
      RECT 20.272 9.36 20.662 10.08 ;
      RECT 19.838 8.88 20.228 10.08 ;
      RECT 20.272 8.88 20.484 9.36 ;
      RECT 20.528 8.16 20.572 9.36 ;
      RECT 20.616 8.16 20.662 9.36 ;
      RECT 19.838 8.16 20.484 8.88 ;
      RECT 19.838 7.92 20.662 8.16 ;
      RECT 20.272 7.2 20.662 7.92 ;
      RECT 19.838 6.72 20.228 7.92 ;
      RECT 20.272 6.72 20.484 7.2 ;
      RECT 20.528 6 20.572 7.2 ;
      RECT 20.616 6 20.662 7.2 ;
      RECT 19.838 6 20.484 6.72 ;
      RECT 19.838 5.76 20.662 6 ;
      RECT 20.272 5.04 20.662 5.76 ;
      RECT 19.838 4.56 20.228 5.76 ;
      RECT 20.272 4.56 20.484 5.04 ;
      RECT 20.528 3.84 20.572 5.04 ;
      RECT 20.616 3.84 20.662 5.04 ;
      RECT 19.838 3.84 20.484 4.56 ;
      RECT 19.838 3.6 20.662 3.84 ;
      RECT 20.272 2.88 20.662 3.6 ;
      RECT 19.838 2.4 20.228 3.6 ;
      RECT 20.272 2.4 20.484 2.88 ;
      RECT 20.528 1.68 20.572 2.88 ;
      RECT 20.616 1.68 20.662 2.88 ;
      RECT 19.838 1.68 20.484 2.4 ;
      RECT 19.838 1.44 20.662 1.68 ;
      RECT 19.838 0.24 20.572 1.44 ;
      RECT 20.616 0.24 20.662 1.44 ;
      RECT 19.838 -0.12 20.662 0.24 ;
      RECT 18.938 41.04 19.762 41.4 ;
      RECT 19.372 40.32 19.762 41.04 ;
      RECT 18.938 39.84 19.072 41.04 ;
      RECT 19.116 39.84 19.328 41.04 ;
      RECT 19.372 39.84 19.584 40.32 ;
      RECT 19.628 39.12 19.762 40.32 ;
      RECT 18.938 39.12 19.584 39.84 ;
      RECT 18.938 38.88 19.762 39.12 ;
      RECT 19.372 38.16 19.762 38.88 ;
      RECT 18.938 37.68 19.072 38.88 ;
      RECT 19.116 37.68 19.328 38.88 ;
      RECT 19.372 37.68 19.584 38.16 ;
      RECT 19.628 36.96 19.762 38.16 ;
      RECT 18.938 36.96 19.584 37.68 ;
      RECT 18.938 36.72 19.762 36.96 ;
      RECT 19.372 36 19.762 36.72 ;
      RECT 18.938 35.52 19.072 36.72 ;
      RECT 19.116 35.52 19.328 36.72 ;
      RECT 19.372 35.52 19.584 36 ;
      RECT 19.628 34.8 19.762 36 ;
      RECT 18.938 34.8 19.584 35.52 ;
      RECT 18.938 34.56 19.762 34.8 ;
      RECT 19.372 33.84 19.762 34.56 ;
      RECT 18.938 33.36 19.072 34.56 ;
      RECT 19.116 33.36 19.328 34.56 ;
      RECT 19.372 33.36 19.584 33.84 ;
      RECT 19.628 32.64 19.762 33.84 ;
      RECT 18.938 32.64 19.584 33.36 ;
      RECT 18.938 32.4 19.762 32.64 ;
      RECT 19.372 31.68 19.762 32.4 ;
      RECT 18.938 31.2 19.072 32.4 ;
      RECT 19.116 31.2 19.328 32.4 ;
      RECT 19.372 31.2 19.584 31.68 ;
      RECT 19.628 30.48 19.762 31.68 ;
      RECT 18.938 30.48 19.584 31.2 ;
      RECT 18.938 30.24 19.762 30.48 ;
      RECT 19.372 29.52 19.762 30.24 ;
      RECT 18.938 29.04 19.072 30.24 ;
      RECT 19.116 29.04 19.328 30.24 ;
      RECT 19.372 29.04 19.584 29.52 ;
      RECT 19.628 28.32 19.762 29.52 ;
      RECT 18.938 28.32 19.584 29.04 ;
      RECT 18.938 28.08 19.762 28.32 ;
      RECT 19.372 27.36 19.762 28.08 ;
      RECT 18.938 26.88 19.072 28.08 ;
      RECT 19.116 26.88 19.328 28.08 ;
      RECT 19.372 26.88 19.584 27.36 ;
      RECT 19.628 26.16 19.762 27.36 ;
      RECT 18.938 26.16 19.584 26.88 ;
      RECT 18.938 25.92 19.762 26.16 ;
      RECT 19.116 25.2 19.762 25.92 ;
      RECT 18.938 24.72 18.984 25.92 ;
      RECT 19.028 24.72 19.072 25.92 ;
      RECT 19.116 24.72 19.584 25.2 ;
      RECT 19.628 24 19.762 25.2 ;
      RECT 18.938 24 19.584 24.72 ;
      RECT 18.938 23.64 19.762 24 ;
      RECT 18.938 22.44 18.984 23.64 ;
      RECT 19.028 22.44 19.072 23.64 ;
      RECT 19.116 22.44 19.328 23.64 ;
      RECT 19.372 22.44 19.762 23.64 ;
      RECT 18.938 21.72 19.762 22.44 ;
      RECT 18.938 20.52 19.072 21.72 ;
      RECT 19.116 20.52 19.328 21.72 ;
      RECT 19.372 20.52 19.672 21.72 ;
      RECT 19.716 20.52 19.762 21.72 ;
      RECT 18.938 20.16 19.762 20.52 ;
      RECT 18.938 18.96 19.584 20.16 ;
      RECT 19.628 18.96 19.762 20.16 ;
      RECT 18.938 18.72 19.762 18.96 ;
      RECT 19.372 18 19.762 18.72 ;
      RECT 18.938 17.52 19.072 18.72 ;
      RECT 19.116 17.52 19.328 18.72 ;
      RECT 19.372 17.52 19.584 18 ;
      RECT 19.628 16.8 19.762 18 ;
      RECT 18.938 16.8 19.584 17.52 ;
      RECT 18.938 16.56 19.762 16.8 ;
      RECT 19.372 15.84 19.762 16.56 ;
      RECT 18.938 15.36 19.072 16.56 ;
      RECT 19.116 15.36 19.328 16.56 ;
      RECT 19.372 15.36 19.584 15.84 ;
      RECT 19.628 14.64 19.762 15.84 ;
      RECT 18.938 14.64 19.584 15.36 ;
      RECT 18.938 14.4 19.762 14.64 ;
      RECT 19.372 13.68 19.762 14.4 ;
      RECT 18.938 13.2 19.072 14.4 ;
      RECT 19.116 13.2 19.328 14.4 ;
      RECT 19.372 13.2 19.584 13.68 ;
      RECT 19.628 12.48 19.762 13.68 ;
      RECT 18.938 12.48 19.584 13.2 ;
      RECT 18.938 12.24 19.762 12.48 ;
      RECT 19.372 11.52 19.762 12.24 ;
      RECT 18.938 11.04 19.072 12.24 ;
      RECT 19.116 11.04 19.328 12.24 ;
      RECT 19.372 11.04 19.584 11.52 ;
      RECT 19.628 10.32 19.762 11.52 ;
      RECT 18.938 10.32 19.584 11.04 ;
      RECT 18.938 10.08 19.762 10.32 ;
      RECT 19.372 9.36 19.762 10.08 ;
      RECT 18.938 8.88 19.072 10.08 ;
      RECT 19.116 8.88 19.328 10.08 ;
      RECT 19.372 8.88 19.584 9.36 ;
      RECT 19.628 8.16 19.762 9.36 ;
      RECT 18.938 8.16 19.584 8.88 ;
      RECT 18.938 7.92 19.762 8.16 ;
      RECT 19.372 7.2 19.762 7.92 ;
      RECT 18.938 6.72 19.072 7.92 ;
      RECT 19.116 6.72 19.328 7.92 ;
      RECT 19.372 6.72 19.584 7.2 ;
      RECT 19.628 6 19.762 7.2 ;
      RECT 18.938 6 19.584 6.72 ;
      RECT 18.938 5.76 19.762 6 ;
      RECT 19.372 5.04 19.762 5.76 ;
      RECT 18.938 4.56 19.072 5.76 ;
      RECT 19.116 4.56 19.328 5.76 ;
      RECT 19.372 4.56 19.584 5.04 ;
      RECT 19.628 3.84 19.762 5.04 ;
      RECT 18.938 3.84 19.584 4.56 ;
      RECT 18.938 3.6 19.762 3.84 ;
      RECT 19.372 2.88 19.762 3.6 ;
      RECT 18.938 2.4 19.072 3.6 ;
      RECT 19.116 2.4 19.328 3.6 ;
      RECT 19.372 2.4 19.584 2.88 ;
      RECT 18.938 2.16 19.584 2.4 ;
      RECT 19.628 1.68 19.762 2.88 ;
      RECT 19.028 1.68 19.584 2.16 ;
      RECT 18.938 0.96 18.984 2.16 ;
      RECT 19.028 0.96 19.762 1.68 ;
      RECT 18.938 -0.12 19.762 0.96 ;
      RECT 18.038 40.32 18.862 41.4 ;
      RECT 18.038 39.6 18.772 40.32 ;
      RECT 18.816 39.12 18.862 40.32 ;
      RECT 18.728 39.12 18.772 39.6 ;
      RECT 18.038 38.4 18.428 39.6 ;
      RECT 18.472 38.4 18.684 39.6 ;
      RECT 18.728 38.4 18.862 39.12 ;
      RECT 18.038 38.16 18.862 38.4 ;
      RECT 18.038 37.44 18.772 38.16 ;
      RECT 18.816 36.96 18.862 38.16 ;
      RECT 18.728 36.96 18.772 37.44 ;
      RECT 18.038 36.24 18.428 37.44 ;
      RECT 18.472 36.24 18.684 37.44 ;
      RECT 18.728 36.24 18.862 36.96 ;
      RECT 18.038 36 18.862 36.24 ;
      RECT 18.038 35.28 18.772 36 ;
      RECT 18.816 34.8 18.862 36 ;
      RECT 18.728 34.8 18.772 35.28 ;
      RECT 18.038 34.08 18.428 35.28 ;
      RECT 18.472 34.08 18.684 35.28 ;
      RECT 18.728 34.08 18.862 34.8 ;
      RECT 18.038 33.84 18.862 34.08 ;
      RECT 18.038 33.12 18.772 33.84 ;
      RECT 18.816 32.64 18.862 33.84 ;
      RECT 18.728 32.64 18.772 33.12 ;
      RECT 18.038 31.92 18.428 33.12 ;
      RECT 18.472 31.92 18.684 33.12 ;
      RECT 18.728 31.92 18.862 32.64 ;
      RECT 18.038 31.68 18.862 31.92 ;
      RECT 18.038 30.96 18.772 31.68 ;
      RECT 18.816 30.48 18.862 31.68 ;
      RECT 18.728 30.48 18.772 30.96 ;
      RECT 18.038 29.76 18.428 30.96 ;
      RECT 18.472 29.76 18.684 30.96 ;
      RECT 18.728 29.76 18.862 30.48 ;
      RECT 18.038 29.52 18.862 29.76 ;
      RECT 18.038 28.8 18.772 29.52 ;
      RECT 18.816 28.32 18.862 29.52 ;
      RECT 18.728 28.32 18.772 28.8 ;
      RECT 18.038 27.6 18.428 28.8 ;
      RECT 18.472 27.6 18.684 28.8 ;
      RECT 18.728 27.6 18.862 28.32 ;
      RECT 18.038 27.36 18.862 27.6 ;
      RECT 18.038 26.64 18.772 27.36 ;
      RECT 18.816 26.16 18.862 27.36 ;
      RECT 18.728 26.16 18.772 26.64 ;
      RECT 18.038 25.44 18.428 26.64 ;
      RECT 18.472 25.44 18.684 26.64 ;
      RECT 18.728 25.44 18.862 26.16 ;
      RECT 18.038 25.2 18.862 25.44 ;
      RECT 18.038 24 18.772 25.2 ;
      RECT 18.816 24 18.862 25.2 ;
      RECT 18.038 23.64 18.862 24 ;
      RECT 18.038 22.44 18.428 23.64 ;
      RECT 18.472 22.44 18.684 23.64 ;
      RECT 18.728 22.44 18.862 23.64 ;
      RECT 18.038 20.16 18.862 22.44 ;
      RECT 18.038 19.44 18.772 20.16 ;
      RECT 18.816 18.96 18.862 20.16 ;
      RECT 18.728 18.96 18.772 19.44 ;
      RECT 18.038 18.24 18.428 19.44 ;
      RECT 18.472 18.24 18.684 19.44 ;
      RECT 18.728 18.24 18.862 18.96 ;
      RECT 18.038 18 18.862 18.24 ;
      RECT 18.038 17.28 18.772 18 ;
      RECT 18.816 16.8 18.862 18 ;
      RECT 18.728 16.8 18.772 17.28 ;
      RECT 18.038 16.08 18.428 17.28 ;
      RECT 18.472 16.08 18.684 17.28 ;
      RECT 18.728 16.08 18.862 16.8 ;
      RECT 18.038 15.84 18.862 16.08 ;
      RECT 18.038 15.12 18.772 15.84 ;
      RECT 18.816 14.64 18.862 15.84 ;
      RECT 18.728 14.64 18.772 15.12 ;
      RECT 18.038 13.92 18.428 15.12 ;
      RECT 18.472 13.92 18.684 15.12 ;
      RECT 18.728 13.92 18.862 14.64 ;
      RECT 18.038 13.68 18.862 13.92 ;
      RECT 18.038 12.96 18.772 13.68 ;
      RECT 18.816 12.48 18.862 13.68 ;
      RECT 18.728 12.48 18.772 12.96 ;
      RECT 18.038 11.76 18.428 12.96 ;
      RECT 18.472 11.76 18.684 12.96 ;
      RECT 18.728 11.76 18.862 12.48 ;
      RECT 18.038 11.52 18.862 11.76 ;
      RECT 18.038 10.8 18.772 11.52 ;
      RECT 18.816 10.32 18.862 11.52 ;
      RECT 18.728 10.32 18.772 10.8 ;
      RECT 18.038 9.6 18.428 10.8 ;
      RECT 18.472 9.6 18.684 10.8 ;
      RECT 18.728 9.6 18.862 10.32 ;
      RECT 18.038 9.36 18.862 9.6 ;
      RECT 18.038 8.64 18.772 9.36 ;
      RECT 18.816 8.16 18.862 9.36 ;
      RECT 18.728 8.16 18.772 8.64 ;
      RECT 18.038 7.44 18.428 8.64 ;
      RECT 18.472 7.44 18.684 8.64 ;
      RECT 18.728 7.44 18.862 8.16 ;
      RECT 18.038 7.2 18.862 7.44 ;
      RECT 18.038 6.48 18.772 7.2 ;
      RECT 18.816 6 18.862 7.2 ;
      RECT 18.728 6 18.772 6.48 ;
      RECT 18.038 5.28 18.428 6.48 ;
      RECT 18.472 5.28 18.684 6.48 ;
      RECT 18.728 5.28 18.862 6 ;
      RECT 18.038 5.04 18.862 5.28 ;
      RECT 18.038 4.32 18.772 5.04 ;
      RECT 18.816 3.84 18.862 5.04 ;
      RECT 18.728 3.84 18.772 4.32 ;
      RECT 18.038 3.12 18.428 4.32 ;
      RECT 18.472 3.12 18.684 4.32 ;
      RECT 18.728 3.12 18.862 3.84 ;
      RECT 18.038 2.88 18.862 3.12 ;
      RECT 18.472 2.16 18.862 2.88 ;
      RECT 18.038 1.68 18.428 2.88 ;
      RECT 18.472 1.68 18.772 2.16 ;
      RECT 18.038 1.44 18.772 1.68 ;
      RECT 18.816 0.96 18.862 2.16 ;
      RECT 18.728 0.96 18.772 1.44 ;
      RECT 18.038 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.862 0.96 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 41.4 ;
      RECT 16.238 -0.12 17.062 41.4 ;
      RECT 15.338 -0.12 16.162 41.4 ;
      RECT 14.438 -0.12 15.262 41.4 ;
      RECT 13.538 -0.12 14.362 41.4 ;
      RECT 12.638 -0.12 13.462 41.4 ;
      RECT 11.738 -0.12 12.562 41.4 ;
      RECT 10.838 -0.12 11.662 41.4 ;
      RECT 9.938 -0.12 10.762 41.4 ;
      RECT 9.038 -0.12 9.862 41.4 ;
      RECT 8.138 -0.12 8.962 41.4 ;
      RECT 7.238 -0.12 8.062 41.4 ;
      RECT 6.338 -0.12 7.162 41.4 ;
      RECT 5.438 -0.12 6.262 41.4 ;
      RECT 4.538 -0.12 5.362 41.4 ;
      RECT 3.638 -0.12 4.462 41.4 ;
      RECT 2.738 -0.12 3.562 41.4 ;
      RECT 1.838 -0.12 2.662 41.4 ;
      RECT 0.938 -0.12 1.762 41.4 ;
      RECT -0.04 41.34 0.862 41.4 ;
      RECT -0.092 -0.06 0.862 41.34 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 42.458 0 43.12 41.28 ;
      RECT 41.558 0 42.142 41.28 ;
      RECT 40.658 0 41.242 41.28 ;
      RECT 39.758 0 40.342 41.28 ;
      RECT 38.858 0 39.442 41.28 ;
      RECT 37.958 0 38.542 41.28 ;
      RECT 37.058 0 37.642 41.28 ;
      RECT 36.158 0 36.742 41.28 ;
      RECT 35.258 0 35.842 41.28 ;
      RECT 34.358 0 34.942 41.28 ;
      RECT 33.458 0 34.042 41.28 ;
      RECT 32.558 0 33.142 41.28 ;
      RECT 31.658 0 32.242 41.28 ;
      RECT 30.758 0 31.342 41.28 ;
      RECT 29.858 0 30.442 41.28 ;
      RECT 28.958 0 29.542 41.28 ;
      RECT 28.058 0 28.642 41.28 ;
      RECT 27.158 0 27.742 41.28 ;
      RECT 26.258 0 26.842 41.28 ;
      RECT 25.358 0 25.942 41.28 ;
      RECT 24.458 0 25.042 41.28 ;
      RECT 23.558 41.16 24.142 41.28 ;
      RECT 23.992 39.72 24.142 41.16 ;
      RECT 23.558 39 24.142 39.72 ;
      RECT 23.992 37.56 24.142 39 ;
      RECT 23.558 36.84 24.142 37.56 ;
      RECT 23.992 35.4 24.142 36.84 ;
      RECT 23.558 34.68 24.142 35.4 ;
      RECT 23.992 33.24 24.142 34.68 ;
      RECT 23.558 32.52 24.142 33.24 ;
      RECT 23.992 31.08 24.142 32.52 ;
      RECT 23.558 30.36 24.142 31.08 ;
      RECT 23.992 28.92 24.142 30.36 ;
      RECT 23.558 28.2 24.142 28.92 ;
      RECT 23.992 26.76 24.142 28.2 ;
      RECT 23.558 26.04 24.142 26.76 ;
      RECT 23.992 24.6 24.142 26.04 ;
      RECT 23.558 23.76 24.142 24.6 ;
      RECT 23.992 22.32 24.142 23.76 ;
      RECT 23.558 18.84 24.142 22.32 ;
      RECT 23.992 17.4 24.142 18.84 ;
      RECT 23.558 16.68 24.142 17.4 ;
      RECT 23.992 15.24 24.142 16.68 ;
      RECT 23.558 14.52 24.142 15.24 ;
      RECT 23.992 13.08 24.142 14.52 ;
      RECT 23.558 12.36 24.142 13.08 ;
      RECT 23.992 10.92 24.142 12.36 ;
      RECT 23.558 10.2 24.142 10.92 ;
      RECT 23.992 8.76 24.142 10.2 ;
      RECT 23.558 8.04 24.142 8.76 ;
      RECT 23.992 6.6 24.142 8.04 ;
      RECT 23.558 5.88 24.142 6.6 ;
      RECT 23.992 4.44 24.142 5.88 ;
      RECT 23.558 3.72 24.142 4.44 ;
      RECT 23.992 2.28 24.142 3.72 ;
      RECT 23.558 1.56 24.142 2.28 ;
      RECT 23.992 0.12 24.142 1.56 ;
      RECT 23.558 0 24.142 0.12 ;
      RECT 22.658 40.44 23.242 41.28 ;
      RECT 22.836 39.72 23.152 40.44 ;
      RECT 21.758 41.16 22.342 41.28 ;
      RECT 22.192 40.44 22.342 41.16 ;
      RECT 20.858 41.16 21.442 41.28 ;
      RECT 20.948 39.72 21.442 41.16 ;
      RECT 19.958 41.16 20.542 41.28 ;
      RECT 20.392 40.44 20.542 41.16 ;
      RECT 19.958 39.72 20.108 41.16 ;
      RECT 19.958 39 20.364 39.72 ;
      RECT 19.958 37.56 20.108 39 ;
      RECT 19.958 36.84 20.364 37.56 ;
      RECT 19.958 35.4 20.108 36.84 ;
      RECT 19.958 34.68 20.364 35.4 ;
      RECT 19.958 33.24 20.108 34.68 ;
      RECT 19.958 32.52 20.364 33.24 ;
      RECT 19.958 31.08 20.108 32.52 ;
      RECT 19.958 30.36 20.364 31.08 ;
      RECT 19.958 28.92 20.108 30.36 ;
      RECT 19.958 28.2 20.364 28.92 ;
      RECT 19.958 26.76 20.108 28.2 ;
      RECT 19.958 26.04 20.364 26.76 ;
      RECT 19.958 24.6 20.108 26.04 ;
      RECT 19.958 23.88 20.452 24.6 ;
      RECT 19.958 21.84 20.542 23.88 ;
      RECT 20.392 20.4 20.542 21.84 ;
      RECT 19.958 20.28 20.542 20.4 ;
      RECT 19.958 18.84 20.364 20.28 ;
      RECT 19.958 17.4 20.108 18.84 ;
      RECT 19.958 16.68 20.364 17.4 ;
      RECT 19.958 15.24 20.108 16.68 ;
      RECT 19.958 14.52 20.364 15.24 ;
      RECT 19.958 13.08 20.108 14.52 ;
      RECT 19.958 12.36 20.364 13.08 ;
      RECT 19.958 10.92 20.108 12.36 ;
      RECT 19.958 10.2 20.364 10.92 ;
      RECT 19.958 8.76 20.108 10.2 ;
      RECT 19.958 8.04 20.364 8.76 ;
      RECT 19.958 6.6 20.108 8.04 ;
      RECT 19.958 5.88 20.364 6.6 ;
      RECT 19.958 4.44 20.108 5.88 ;
      RECT 19.958 3.72 20.364 4.44 ;
      RECT 19.958 2.28 20.108 3.72 ;
      RECT 19.958 1.56 20.364 2.28 ;
      RECT 19.958 0.12 20.452 1.56 ;
      RECT 19.958 0 20.542 0.12 ;
      RECT 19.058 41.16 19.642 41.28 ;
      RECT 19.492 40.44 19.642 41.16 ;
      RECT 18.158 40.44 18.742 41.28 ;
      RECT 18.158 39.72 18.652 40.44 ;
      RECT 18.158 38.28 18.308 39.72 ;
      RECT 18.158 37.56 18.652 38.28 ;
      RECT 18.158 36.12 18.308 37.56 ;
      RECT 18.158 35.4 18.652 36.12 ;
      RECT 18.158 33.96 18.308 35.4 ;
      RECT 18.158 33.24 18.652 33.96 ;
      RECT 18.158 31.8 18.308 33.24 ;
      RECT 18.158 31.08 18.652 31.8 ;
      RECT 18.158 29.64 18.308 31.08 ;
      RECT 18.158 28.92 18.652 29.64 ;
      RECT 18.158 27.48 18.308 28.92 ;
      RECT 18.158 26.76 18.652 27.48 ;
      RECT 18.158 25.32 18.308 26.76 ;
      RECT 18.158 23.88 18.652 25.32 ;
      RECT 18.158 23.76 18.742 23.88 ;
      RECT 18.158 22.32 18.308 23.76 ;
      RECT 18.158 20.28 18.742 22.32 ;
      RECT 18.158 19.56 18.652 20.28 ;
      RECT 18.158 18.12 18.308 19.56 ;
      RECT 18.158 17.4 18.652 18.12 ;
      RECT 18.158 15.96 18.308 17.4 ;
      RECT 18.158 15.24 18.652 15.96 ;
      RECT 18.158 13.8 18.308 15.24 ;
      RECT 18.158 13.08 18.652 13.8 ;
      RECT 18.158 11.64 18.308 13.08 ;
      RECT 18.158 10.92 18.652 11.64 ;
      RECT 18.158 9.48 18.308 10.92 ;
      RECT 18.158 8.76 18.652 9.48 ;
      RECT 18.158 7.32 18.308 8.76 ;
      RECT 18.158 6.6 18.652 7.32 ;
      RECT 18.158 5.16 18.308 6.6 ;
      RECT 18.158 4.44 18.652 5.16 ;
      RECT 18.158 0.12 18.308 4.44 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 41.28 ;
      RECT 16.358 0 16.942 41.28 ;
      RECT 15.458 0 16.042 41.28 ;
      RECT 14.558 0 15.142 41.28 ;
      RECT 13.658 0 14.242 41.28 ;
      RECT 12.758 0 13.342 41.28 ;
      RECT 11.858 0 12.442 41.28 ;
      RECT 10.958 0 11.542 41.28 ;
      RECT 10.058 0 10.642 41.28 ;
      RECT 9.158 0 9.742 41.28 ;
      RECT 8.258 0 8.842 41.28 ;
      RECT 7.358 0 7.942 41.28 ;
      RECT 6.458 0 7.042 41.28 ;
      RECT 5.558 0 6.142 41.28 ;
      RECT 4.658 0 5.242 41.28 ;
      RECT 3.758 0 4.342 41.28 ;
      RECT 2.858 0 3.442 41.28 ;
      RECT 1.958 0 2.542 41.28 ;
      RECT 1.058 0 1.642 41.28 ;
      RECT 0.08 0 0.742 41.28 ;
      RECT 21.848 39 22.164 39.72 ;
      RECT 19.058 39 19.464 39.72 ;
      RECT 22.658 38.28 22.808 39 ;
      RECT 22.192 38.28 22.342 39 ;
      RECT 20.392 38.28 20.542 39 ;
      RECT 19.492 38.28 19.642 39 ;
      RECT 22.836 37.56 23.152 38.28 ;
      RECT 20.948 37.56 21.442 38.28 ;
      RECT 21.848 36.84 22.164 37.56 ;
      RECT 19.058 36.84 19.464 37.56 ;
      RECT 22.658 36.12 22.808 36.84 ;
      RECT 22.192 36.12 22.342 36.84 ;
      RECT 20.392 36.12 20.542 36.84 ;
      RECT 19.492 36.12 19.642 36.84 ;
      RECT 22.836 35.4 23.152 36.12 ;
      RECT 20.948 35.4 21.442 36.12 ;
      RECT 21.848 34.68 22.164 35.4 ;
      RECT 19.058 34.68 19.464 35.4 ;
      RECT 22.658 33.96 22.808 34.68 ;
      RECT 22.192 33.96 22.342 34.68 ;
      RECT 20.392 33.96 20.542 34.68 ;
      RECT 19.492 33.96 19.642 34.68 ;
      RECT 22.836 33.24 23.152 33.96 ;
      RECT 20.948 33.24 21.442 33.96 ;
      RECT 21.848 32.52 22.164 33.24 ;
      RECT 19.058 32.52 19.464 33.24 ;
      RECT 22.658 31.8 22.808 32.52 ;
      RECT 22.192 31.8 22.342 32.52 ;
      RECT 20.392 31.8 20.542 32.52 ;
      RECT 19.492 31.8 19.642 32.52 ;
      RECT 22.836 31.08 23.152 31.8 ;
      RECT 20.948 31.08 21.442 31.8 ;
      RECT 21.848 30.36 22.164 31.08 ;
      RECT 19.058 30.36 19.464 31.08 ;
      RECT 22.658 29.64 22.808 30.36 ;
      RECT 22.192 29.64 22.342 30.36 ;
      RECT 20.392 29.64 20.542 30.36 ;
      RECT 19.492 29.64 19.642 30.36 ;
      RECT 22.836 28.92 23.152 29.64 ;
      RECT 20.948 28.92 21.442 29.64 ;
      RECT 21.848 28.2 22.164 28.92 ;
      RECT 19.058 28.2 19.464 28.92 ;
      RECT 22.658 27.48 22.808 28.2 ;
      RECT 22.192 27.48 22.342 28.2 ;
      RECT 20.392 27.48 20.542 28.2 ;
      RECT 19.492 27.48 19.642 28.2 ;
      RECT 22.836 26.76 23.152 27.48 ;
      RECT 20.948 26.76 21.442 27.48 ;
      RECT 21.848 26.04 22.164 26.76 ;
      RECT 21.936 25.32 22.342 26.04 ;
      RECT 19.058 26.04 19.464 26.76 ;
      RECT 19.236 25.32 19.642 26.04 ;
      RECT 19.236 24.6 19.464 25.32 ;
      RECT 19.058 23.88 19.464 24.6 ;
      RECT 19.058 23.76 19.642 23.88 ;
      RECT 19.492 22.32 19.642 23.76 ;
      RECT 19.058 21.84 19.642 22.32 ;
      RECT 19.492 20.4 19.552 21.84 ;
      RECT 19.058 20.28 19.642 20.4 ;
      RECT 19.058 18.84 19.464 20.28 ;
      RECT 22.658 25.32 22.808 26.04 ;
      RECT 22.836 23.88 23.152 25.32 ;
      RECT 22.658 23.76 23.242 23.88 ;
      RECT 22.748 22.32 22.808 23.76 ;
      RECT 22.658 20.28 23.242 22.32 ;
      RECT 22.836 19.56 23.152 20.28 ;
      RECT 20.948 23.88 21.442 25.32 ;
      RECT 20.858 21.84 21.442 23.88 ;
      RECT 21.758 23.88 21.908 24.6 ;
      RECT 21.758 23.76 22.342 23.88 ;
      RECT 21.758 22.32 22.252 23.76 ;
      RECT 21.758 21.84 22.342 22.32 ;
      RECT 22.192 20.4 22.342 21.84 ;
      RECT 21.758 20.28 22.342 20.4 ;
      RECT 21.848 18.84 22.164 20.28 ;
      RECT 20.858 19.56 21.442 20.4 ;
      RECT 22.658 18.12 22.808 18.84 ;
      RECT 22.192 18.12 22.342 18.84 ;
      RECT 20.392 18.12 20.542 18.84 ;
      RECT 19.492 18.12 19.642 18.84 ;
      RECT 22.836 17.4 23.152 18.12 ;
      RECT 20.948 17.4 21.442 18.12 ;
      RECT 21.848 16.68 22.164 17.4 ;
      RECT 19.058 16.68 19.464 17.4 ;
      RECT 22.658 15.96 22.808 16.68 ;
      RECT 22.192 15.96 22.342 16.68 ;
      RECT 20.392 15.96 20.542 16.68 ;
      RECT 19.492 15.96 19.642 16.68 ;
      RECT 22.836 15.24 23.152 15.96 ;
      RECT 20.948 15.24 21.442 15.96 ;
      RECT 21.848 14.52 22.164 15.24 ;
      RECT 19.058 14.52 19.464 15.24 ;
      RECT 22.658 13.8 22.808 14.52 ;
      RECT 22.192 13.8 22.342 14.52 ;
      RECT 20.392 13.8 20.542 14.52 ;
      RECT 19.492 13.8 19.642 14.52 ;
      RECT 22.836 13.08 23.152 13.8 ;
      RECT 20.948 13.08 21.442 13.8 ;
      RECT 21.848 12.36 22.164 13.08 ;
      RECT 19.058 12.36 19.464 13.08 ;
      RECT 22.658 11.64 22.808 12.36 ;
      RECT 22.192 11.64 22.342 12.36 ;
      RECT 20.392 11.64 20.542 12.36 ;
      RECT 19.492 11.64 19.642 12.36 ;
      RECT 22.836 10.92 23.152 11.64 ;
      RECT 20.948 10.92 21.442 11.64 ;
      RECT 21.848 10.2 22.164 10.92 ;
      RECT 19.058 10.2 19.464 10.92 ;
      RECT 22.658 9.48 22.808 10.2 ;
      RECT 22.192 9.48 22.342 10.2 ;
      RECT 20.392 9.48 20.542 10.2 ;
      RECT 19.492 9.48 19.642 10.2 ;
      RECT 22.836 8.76 23.152 9.48 ;
      RECT 20.948 8.76 21.442 9.48 ;
      RECT 21.848 8.04 22.164 8.76 ;
      RECT 19.058 8.04 19.464 8.76 ;
      RECT 22.658 7.32 22.808 8.04 ;
      RECT 22.192 7.32 22.342 8.04 ;
      RECT 20.392 7.32 20.542 8.04 ;
      RECT 19.492 7.32 19.642 8.04 ;
      RECT 22.836 6.6 23.152 7.32 ;
      RECT 20.948 6.6 21.442 7.32 ;
      RECT 21.848 5.88 22.164 6.6 ;
      RECT 19.058 5.88 19.464 6.6 ;
      RECT 22.658 5.16 22.808 5.88 ;
      RECT 22.192 5.16 22.342 5.88 ;
      RECT 20.392 5.16 20.542 5.88 ;
      RECT 19.492 5.16 19.642 5.88 ;
      RECT 22.836 4.44 23.152 5.16 ;
      RECT 20.948 4.44 21.442 5.16 ;
      RECT 21.848 3.72 22.164 4.44 ;
      RECT 19.058 3.72 19.464 4.44 ;
      RECT 22.658 3 22.808 3.72 ;
      RECT 22.192 3 22.342 3.72 ;
      RECT 20.392 3 20.542 3.72 ;
      RECT 19.492 3 19.642 3.72 ;
      RECT 22.836 2.28 23.152 3 ;
      RECT 20.948 2.28 21.442 3 ;
      RECT 18.592 2.28 18.742 3 ;
      RECT 18.592 1.56 18.652 2.28 ;
      RECT 21.848 1.56 22.164 2.28 ;
      RECT 21.758 0.12 21.908 1.56 ;
      RECT 21.758 0 22.342 0.12 ;
      RECT 19.148 1.56 19.464 2.28 ;
      RECT 19.148 0.84 19.642 1.56 ;
      RECT 19.058 0 19.642 0.84 ;
      RECT 22.658 0.84 22.808 1.56 ;
      RECT 22.658 0 23.242 0.84 ;
      RECT 20.948 0.12 21.442 0.84 ;
      RECT 20.858 0 21.442 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 43.2 41.278 ;
    LAYER m1 ;
      RECT 0 0 43.2 41.28 ;
    LAYER m2 ;
      RECT 0 0.015 43.2 41.265 ;
    LAYER m3 ;
      RECT 0.015 0 43.185 41.28 ;
    LAYER m4 ;
      RECT 0 0.02 43.2 41.26 ;
    LAYER m5 ;
      RECT 0.012 0 43.188 41.28 ;
    LAYER m6 ;
      RECT 0 0.012 43.2 41.268 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf198b128e1r1w0cbbehbaa4acw

END LIBRARY
