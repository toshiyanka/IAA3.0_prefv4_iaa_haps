localparam int MAX_NUM_SLICES=512;
