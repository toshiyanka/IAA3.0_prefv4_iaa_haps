module ctech_lib_latch_async_set (clk, d, psb, o);
   input clk, d, psb;
   output o;
   logic o;
   d04lyn0cld0b0 ctech_lib_dcszo (.clk(clk),.d(d),.psb(psb),.o(o));
endmodule
