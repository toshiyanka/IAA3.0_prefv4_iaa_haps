parameter MATCHED_INTERNAL_WIDTH=0;
parameter MASTERREG=1;
parameter MAXPCMSTR=0;
parameter MAXNPMSTR=0;
parameter MAXMSTRDATA=63;
parameter MAXMSTRADDR=31;
parameter TARGETREG=1;
parameter MAXPCTRGT=0;
parameter MAXTRGTDATA=63;
parameter MAXNPTRGT=0;
parameter MAXTRGTADDR=47;
parameter ASYNCENDPT=1;
parameter ASYNCIQDEPTH=4;
parameter ASYNCEQDEPTH=4;
parameter NPQUEUEDEPTH=7;
parameter PCQUEUEDEPTH=7;
parameter LATCHQUEUES=0;
parameter MAXPLDBIT=31;
parameter RX_EXT_HEADER_IDS=0;
parameter RSWIDTH=3;
parameter SAIWIDTH=7;
parameter PIPEINPS=1;
parameter PIPEISMS=1;
parameter USYNC_ENABLE=0;
parameter SIDE_USYNC_DELAY=2;
parameter AGENT_USYNC_DELAY=2;
parameter FAB_CLK_PERIOD=2500ps;//899ps;
parameter AGT_CLK_PERIOD=1111ps;//9330ps;
parameter DISABLE_COMPLETION_FENCING=0;
parameter ISM_COMPLETION_FENCING=1;
parameter EXPECTED_COMPLETIONS_COUNTER=1;
parameter SKIP_ACTIVEREQ=1;
parameter TX_EXT_HEADER_SUPPORT=1;
parameter RX_EXT_HEADER_SUPPORT=1;
parameter UNIQUE_EXT_HEADERS=1;
parameter NUM_RX_EXT_HEADERS=1+0;
parameter NUM_TX_EXT_HEADERS=1+0;
parameter FBRC_EXT_HEADER_SUPPORT=1;
parameter AGT_EXT_HEADER_SUPPORT=0;
parameter VALONLYMODEL=0;
parameter DUMMY_CLKBUF=0;
parameter IOSFSB_EP_SPEC_REV=11;
parameter IOSFSB_FBRC_SPEC_REV=11;
parameter CUP2PUT1CYC=0;
parameter NUMBER_OF_OUTPUT_LANES=1;
parameter NUMBER_OF_BITS_PER_LANE=8;
parameter SBE_VISA_ID_PARAM=11;
parameter NUMBER_OF_VISAMUX_MODULES=1;
parameter VARIABLE_CLAIM_DELAY = 0;
parameter SB_PARITY_REQUIRED = 0;
parameter DO_SERR_MASTER=0;
parameter NUM_REPEATER=0;
parameter NUM_CLAIM_REPEATER=0;
parameter RELATIVE_PLACEMENT_EN=0;
parameter CLKREQDEFAULT=0;
parameter GLOBAL_EP=0;
parameter GLOBAL_EP_IS_STRAP=0;
parameter BULKRDWR=0;
parameter DEASSERT_CLK_SIGS=0;
