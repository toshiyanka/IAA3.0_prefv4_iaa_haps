VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf046b032e1r1w0cbbehraa4acw
  CLASS BLOCK ;
  FOREIGN arf046b032e1r1w0cbbehraa4acw ;
  ORIGIN 0 0 ;
  SIZE 12.6 BY 22.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 2.52 0.728 3.72 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 0.6 0.472 1.8 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.52 2.528 3.72 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 2.52 2.828 3.72 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 2.52 3.172 3.72 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 2.52 3.516 3.72 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 2.52 3.816 3.72 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 2.52 1.028 3.72 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 2.52 1.372 3.72 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 2.52 1.716 3.72 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 2.52 2.016 3.72 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 0.6 2.616 1.8 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.6 2.916 1.8 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.6 3.428 1.8 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.6 3.728 1.8 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 0.6 4.072 1.8 ;
    END
  END wraddrp0[4]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 0.6 0.816 1.8 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 0.6 1.116 1.8 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 4.08 2.272 5.28 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 7.68 2.528 8.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 7.68 2.828 8.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 8.4 2.272 9.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 8.4 2.616 9.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 9.12 2.528 10.32 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 9.12 2.828 10.32 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 9.84 2.272 11.04 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 9.84 2.616 11.04 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 10.56 2.528 11.76 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 10.56 2.828 11.76 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 4.08 2.616 5.28 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 11.28 2.272 12.48 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 11.28 2.616 12.48 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 12 2.528 13.2 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12 2.828 13.2 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 12.72 2.272 13.92 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 12.72 2.616 13.92 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 13.44 2.528 14.64 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 13.44 2.828 14.64 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 14.16 2.272 15.36 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.16 2.616 15.36 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 4.8 2.528 6 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 14.88 2.528 16.08 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 14.88 2.828 16.08 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 15.6 2.272 16.8 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 15.6 2.616 16.8 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 16.32 2.528 17.52 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 16.32 2.828 17.52 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 17.04 2.272 18.24 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 17.04 2.616 18.24 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 17.76 2.528 18.96 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 17.76 2.828 18.96 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 4.8 2.828 6 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 18.48 2.272 19.68 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 18.48 2.616 19.68 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 19.2 2.528 20.4 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 19.2 2.828 20.4 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 19.92 2.272 21.12 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.92 2.616 21.12 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 20.64 2.528 21.84 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 20.64 2.828 21.84 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 5.52 2.272 6.72 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.52 2.616 6.72 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6.24 2.528 7.44 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 6.24 2.828 7.44 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 6.96 2.272 8.16 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 6.96 2.616 8.16 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.6 1.928 1.8 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.6 2.272 1.8 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 0.6 1.628 1.8 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 4.08 4.328 5.28 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 7.68 4.072 8.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 7.68 3.428 8.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 8.4 4.328 9.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.4 3.516 9.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 9.12 4.072 10.32 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9.12 3.428 10.32 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.84 4.328 11.04 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 9.84 3.516 11.04 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 10.56 4.072 11.76 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 10.56 3.428 11.76 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 4.08 3.728 5.28 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 11.28 4.328 12.48 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.28 3.516 12.48 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 12 4.072 13.2 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 12 3.428 13.2 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 12.72 4.328 13.92 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.72 3.516 13.92 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 13.44 4.072 14.64 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 13.44 3.428 14.64 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 14.16 4.328 15.36 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 14.16 3.516 15.36 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 4.8 4.072 6 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 14.88 4.072 16.08 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 14.88 3.428 16.08 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 15.6 4.328 16.8 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 15.6 3.516 16.8 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.32 4.072 17.52 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.32 3.428 17.52 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 17.04 4.328 18.24 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 17.04 3.516 18.24 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 17.76 4.072 18.96 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 17.76 3.428 18.96 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.8 3.428 6 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 18.48 4.328 19.68 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 18.48 3.516 19.68 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 19.2 4.072 20.4 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 19.2 3.428 20.4 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 19.92 4.328 21.12 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.92 3.516 21.12 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 20.64 4.072 21.84 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.64 3.428 21.84 ;
    END
  END rddatap0[47]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 5.52 4.328 6.72 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.52 3.516 6.72 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.24 4.072 7.44 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6.24 3.428 7.44 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6.96 4.328 8.16 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 6.96 3.516 8.16 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 22.02 ;
        RECT 2.662 0.06 2.738 22.02 ;
        RECT 4.462 0.06 4.538 22.02 ;
        RECT 6.262 0.06 6.338 22.02 ;
        RECT 8.062 0.06 8.138 22.02 ;
        RECT 9.862 0.06 9.938 22.02 ;
        RECT 11.662 0.06 11.738 22.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 22.02 ;
        RECT 3.562 0.06 3.638 22.02 ;
        RECT 5.362 0.06 5.438 22.02 ;
        RECT 7.162 0.06 7.238 22.02 ;
        RECT 8.962 0.06 9.038 22.02 ;
        RECT 10.762 0.06 10.838 22.02 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 12.616 22.094 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 12.62 22.1 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 12.6705 22.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 12.635 22.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 12.67 22.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 12.659 22.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 12.69 22.142 ;
    LAYER m7 SPACING 0 ;
      RECT 11.738 22.14 12.64 22.2 ;
      RECT 11.738 -0.06 12.692 22.14 ;
      RECT 11.738 -0.12 12.64 -0.06 ;
      RECT 10.838 -0.12 11.662 22.2 ;
      RECT 9.938 -0.12 10.762 22.2 ;
      RECT 9.038 -0.12 9.862 22.2 ;
      RECT 8.138 -0.12 8.962 22.2 ;
      RECT 7.238 -0.12 8.062 22.2 ;
      RECT 6.338 -0.12 7.162 22.2 ;
      RECT 5.438 -0.12 6.262 22.2 ;
      RECT 4.538 -0.12 5.362 22.2 ;
      RECT 3.638 21.84 4.462 22.2 ;
      RECT 4.072 21.12 4.462 21.84 ;
      RECT 3.638 20.64 4.028 21.84 ;
      RECT 4.072 20.64 4.284 21.12 ;
      RECT 3.638 20.4 4.284 20.64 ;
      RECT 4.328 19.92 4.462 21.12 ;
      RECT 4.072 19.92 4.284 20.4 ;
      RECT 4.072 19.68 4.462 19.92 ;
      RECT 3.638 19.2 4.028 20.4 ;
      RECT 4.072 19.2 4.284 19.68 ;
      RECT 3.638 18.96 4.284 19.2 ;
      RECT 4.328 18.48 4.462 19.68 ;
      RECT 4.072 18.48 4.284 18.96 ;
      RECT 4.072 18.24 4.462 18.48 ;
      RECT 3.638 17.76 4.028 18.96 ;
      RECT 4.072 17.76 4.284 18.24 ;
      RECT 3.638 17.52 4.284 17.76 ;
      RECT 4.328 17.04 4.462 18.24 ;
      RECT 4.072 17.04 4.284 17.52 ;
      RECT 4.072 16.8 4.462 17.04 ;
      RECT 3.638 16.32 4.028 17.52 ;
      RECT 4.072 16.32 4.284 16.8 ;
      RECT 3.638 16.08 4.284 16.32 ;
      RECT 4.328 15.6 4.462 16.8 ;
      RECT 4.072 15.6 4.284 16.08 ;
      RECT 4.072 15.36 4.462 15.6 ;
      RECT 3.638 14.88 4.028 16.08 ;
      RECT 4.072 14.88 4.284 15.36 ;
      RECT 3.638 14.64 4.284 14.88 ;
      RECT 4.328 14.16 4.462 15.36 ;
      RECT 4.072 14.16 4.284 14.64 ;
      RECT 4.072 13.92 4.462 14.16 ;
      RECT 3.638 13.44 4.028 14.64 ;
      RECT 4.072 13.44 4.284 13.92 ;
      RECT 3.638 13.2 4.284 13.44 ;
      RECT 4.328 12.72 4.462 13.92 ;
      RECT 4.072 12.72 4.284 13.2 ;
      RECT 4.072 12.48 4.462 12.72 ;
      RECT 3.638 12 4.028 13.2 ;
      RECT 4.072 12 4.284 12.48 ;
      RECT 3.638 11.76 4.284 12 ;
      RECT 4.328 11.28 4.462 12.48 ;
      RECT 4.072 11.28 4.284 11.76 ;
      RECT 4.072 11.04 4.462 11.28 ;
      RECT 3.638 10.56 4.028 11.76 ;
      RECT 4.072 10.56 4.284 11.04 ;
      RECT 3.638 10.32 4.284 10.56 ;
      RECT 4.328 9.84 4.462 11.04 ;
      RECT 4.072 9.84 4.284 10.32 ;
      RECT 4.072 9.6 4.462 9.84 ;
      RECT 3.638 9.12 4.028 10.32 ;
      RECT 4.072 9.12 4.284 9.6 ;
      RECT 3.638 8.88 4.284 9.12 ;
      RECT 4.328 8.4 4.462 9.6 ;
      RECT 4.072 8.4 4.284 8.88 ;
      RECT 4.072 8.16 4.462 8.4 ;
      RECT 3.638 7.68 4.028 8.88 ;
      RECT 4.072 7.68 4.284 8.16 ;
      RECT 3.638 7.44 4.284 7.68 ;
      RECT 4.328 6.96 4.462 8.16 ;
      RECT 4.072 6.96 4.284 7.44 ;
      RECT 4.072 6.72 4.462 6.96 ;
      RECT 3.638 6.24 4.028 7.44 ;
      RECT 4.072 6.24 4.284 6.72 ;
      RECT 3.638 6 4.284 6.24 ;
      RECT 4.328 5.52 4.462 6.72 ;
      RECT 4.072 5.52 4.284 6 ;
      RECT 3.638 5.28 4.028 6 ;
      RECT 4.072 5.28 4.462 5.52 ;
      RECT 3.728 4.8 4.028 5.28 ;
      RECT 4.072 4.8 4.284 5.28 ;
      RECT 3.638 4.08 3.684 5.28 ;
      RECT 4.328 4.08 4.462 5.28 ;
      RECT 3.728 4.08 4.284 4.8 ;
      RECT 3.638 3.72 4.462 4.08 ;
      RECT 3.638 2.52 3.772 3.72 ;
      RECT 3.816 2.52 4.462 3.72 ;
      RECT 3.638 1.8 4.462 2.52 ;
      RECT 3.638 0.6 3.684 1.8 ;
      RECT 3.728 0.6 4.028 1.8 ;
      RECT 4.072 0.6 4.462 1.8 ;
      RECT 3.638 -0.12 4.462 0.6 ;
      RECT 2.738 21.84 3.562 22.2 ;
      RECT 3.428 21.12 3.562 21.84 ;
      RECT 2.738 20.64 2.784 21.84 ;
      RECT 2.828 20.64 3.384 21.84 ;
      RECT 3.428 20.64 3.472 21.12 ;
      RECT 2.738 20.4 3.472 20.64 ;
      RECT 3.516 19.92 3.562 21.12 ;
      RECT 3.428 19.92 3.472 20.4 ;
      RECT 3.428 19.68 3.562 19.92 ;
      RECT 2.738 19.2 2.784 20.4 ;
      RECT 2.828 19.2 3.384 20.4 ;
      RECT 3.428 19.2 3.472 19.68 ;
      RECT 2.738 18.96 3.472 19.2 ;
      RECT 3.516 18.48 3.562 19.68 ;
      RECT 3.428 18.48 3.472 18.96 ;
      RECT 3.428 18.24 3.562 18.48 ;
      RECT 2.738 17.76 2.784 18.96 ;
      RECT 2.828 17.76 3.384 18.96 ;
      RECT 3.428 17.76 3.472 18.24 ;
      RECT 2.738 17.52 3.472 17.76 ;
      RECT 3.516 17.04 3.562 18.24 ;
      RECT 3.428 17.04 3.472 17.52 ;
      RECT 3.428 16.8 3.562 17.04 ;
      RECT 2.738 16.32 2.784 17.52 ;
      RECT 2.828 16.32 3.384 17.52 ;
      RECT 3.428 16.32 3.472 16.8 ;
      RECT 2.738 16.08 3.472 16.32 ;
      RECT 3.516 15.6 3.562 16.8 ;
      RECT 3.428 15.6 3.472 16.08 ;
      RECT 3.428 15.36 3.562 15.6 ;
      RECT 2.738 14.88 2.784 16.08 ;
      RECT 2.828 14.88 3.384 16.08 ;
      RECT 3.428 14.88 3.472 15.36 ;
      RECT 2.738 14.64 3.472 14.88 ;
      RECT 3.516 14.16 3.562 15.36 ;
      RECT 3.428 14.16 3.472 14.64 ;
      RECT 3.428 13.92 3.562 14.16 ;
      RECT 2.738 13.44 2.784 14.64 ;
      RECT 2.828 13.44 3.384 14.64 ;
      RECT 3.428 13.44 3.472 13.92 ;
      RECT 2.738 13.2 3.472 13.44 ;
      RECT 3.516 12.72 3.562 13.92 ;
      RECT 3.428 12.72 3.472 13.2 ;
      RECT 3.428 12.48 3.562 12.72 ;
      RECT 2.738 12 2.784 13.2 ;
      RECT 2.828 12 3.384 13.2 ;
      RECT 3.428 12 3.472 12.48 ;
      RECT 2.738 11.76 3.472 12 ;
      RECT 3.516 11.28 3.562 12.48 ;
      RECT 3.428 11.28 3.472 11.76 ;
      RECT 3.428 11.04 3.562 11.28 ;
      RECT 2.738 10.56 2.784 11.76 ;
      RECT 2.828 10.56 3.384 11.76 ;
      RECT 3.428 10.56 3.472 11.04 ;
      RECT 2.738 10.32 3.472 10.56 ;
      RECT 3.516 9.84 3.562 11.04 ;
      RECT 3.428 9.84 3.472 10.32 ;
      RECT 3.428 9.6 3.562 9.84 ;
      RECT 2.738 9.12 2.784 10.32 ;
      RECT 2.828 9.12 3.384 10.32 ;
      RECT 3.428 9.12 3.472 9.6 ;
      RECT 2.738 8.88 3.472 9.12 ;
      RECT 3.516 8.4 3.562 9.6 ;
      RECT 3.428 8.4 3.472 8.88 ;
      RECT 3.428 8.16 3.562 8.4 ;
      RECT 2.738 7.68 2.784 8.88 ;
      RECT 2.828 7.68 3.384 8.88 ;
      RECT 3.428 7.68 3.472 8.16 ;
      RECT 2.738 7.44 3.472 7.68 ;
      RECT 3.516 6.96 3.562 8.16 ;
      RECT 3.428 6.96 3.472 7.44 ;
      RECT 3.428 6.72 3.562 6.96 ;
      RECT 2.738 6.24 2.784 7.44 ;
      RECT 2.828 6.24 3.384 7.44 ;
      RECT 3.428 6.24 3.472 6.72 ;
      RECT 2.738 6 3.472 6.24 ;
      RECT 3.516 5.52 3.562 6.72 ;
      RECT 3.428 5.52 3.472 6 ;
      RECT 2.738 4.8 2.784 6 ;
      RECT 2.828 4.8 3.384 6 ;
      RECT 3.428 4.8 3.562 5.52 ;
      RECT 2.738 3.72 3.562 4.8 ;
      RECT 2.738 2.52 2.784 3.72 ;
      RECT 2.828 2.52 3.128 3.72 ;
      RECT 3.172 2.52 3.472 3.72 ;
      RECT 3.516 2.52 3.562 3.72 ;
      RECT 2.738 1.8 3.562 2.52 ;
      RECT 2.738 0.6 2.872 1.8 ;
      RECT 2.916 0.6 3.384 1.8 ;
      RECT 3.428 0.6 3.562 1.8 ;
      RECT 2.738 -0.12 3.562 0.6 ;
      RECT 1.838 21.84 2.662 22.2 ;
      RECT 1.838 21.12 2.484 21.84 ;
      RECT 2.528 21.12 2.662 21.84 ;
      RECT 2.272 20.64 2.484 21.12 ;
      RECT 2.528 20.64 2.572 21.12 ;
      RECT 2.272 20.4 2.572 20.64 ;
      RECT 1.838 19.92 2.228 21.12 ;
      RECT 2.616 19.92 2.662 21.12 ;
      RECT 2.272 19.92 2.484 20.4 ;
      RECT 2.528 19.92 2.572 20.4 ;
      RECT 1.838 19.68 2.484 19.92 ;
      RECT 2.528 19.68 2.662 19.92 ;
      RECT 2.272 19.2 2.484 19.68 ;
      RECT 2.528 19.2 2.572 19.68 ;
      RECT 2.272 18.96 2.572 19.2 ;
      RECT 1.838 18.48 2.228 19.68 ;
      RECT 2.616 18.48 2.662 19.68 ;
      RECT 2.272 18.48 2.484 18.96 ;
      RECT 2.528 18.48 2.572 18.96 ;
      RECT 1.838 18.24 2.484 18.48 ;
      RECT 2.528 18.24 2.662 18.48 ;
      RECT 2.272 17.76 2.484 18.24 ;
      RECT 2.528 17.76 2.572 18.24 ;
      RECT 2.272 17.52 2.572 17.76 ;
      RECT 1.838 17.04 2.228 18.24 ;
      RECT 2.616 17.04 2.662 18.24 ;
      RECT 2.272 17.04 2.484 17.52 ;
      RECT 2.528 17.04 2.572 17.52 ;
      RECT 1.838 16.8 2.484 17.04 ;
      RECT 2.528 16.8 2.662 17.04 ;
      RECT 2.272 16.32 2.484 16.8 ;
      RECT 2.528 16.32 2.572 16.8 ;
      RECT 2.272 16.08 2.572 16.32 ;
      RECT 1.838 15.6 2.228 16.8 ;
      RECT 2.616 15.6 2.662 16.8 ;
      RECT 2.272 15.6 2.484 16.08 ;
      RECT 2.528 15.6 2.572 16.08 ;
      RECT 1.838 15.36 2.484 15.6 ;
      RECT 2.528 15.36 2.662 15.6 ;
      RECT 2.272 14.88 2.484 15.36 ;
      RECT 2.528 14.88 2.572 15.36 ;
      RECT 2.272 14.64 2.572 14.88 ;
      RECT 1.838 14.16 2.228 15.36 ;
      RECT 2.616 14.16 2.662 15.36 ;
      RECT 2.272 14.16 2.484 14.64 ;
      RECT 2.528 14.16 2.572 14.64 ;
      RECT 1.838 13.92 2.484 14.16 ;
      RECT 2.528 13.92 2.662 14.16 ;
      RECT 2.272 13.44 2.484 13.92 ;
      RECT 2.528 13.44 2.572 13.92 ;
      RECT 2.272 13.2 2.572 13.44 ;
      RECT 1.838 12.72 2.228 13.92 ;
      RECT 2.616 12.72 2.662 13.92 ;
      RECT 2.272 12.72 2.484 13.2 ;
      RECT 2.528 12.72 2.572 13.2 ;
      RECT 1.838 12.48 2.484 12.72 ;
      RECT 2.528 12.48 2.662 12.72 ;
      RECT 2.272 12 2.484 12.48 ;
      RECT 2.528 12 2.572 12.48 ;
      RECT 2.272 11.76 2.572 12 ;
      RECT 1.838 11.28 2.228 12.48 ;
      RECT 2.616 11.28 2.662 12.48 ;
      RECT 2.272 11.28 2.484 11.76 ;
      RECT 2.528 11.28 2.572 11.76 ;
      RECT 1.838 11.04 2.484 11.28 ;
      RECT 2.528 11.04 2.662 11.28 ;
      RECT 2.272 10.56 2.484 11.04 ;
      RECT 2.528 10.56 2.572 11.04 ;
      RECT 2.272 10.32 2.572 10.56 ;
      RECT 1.838 9.84 2.228 11.04 ;
      RECT 2.616 9.84 2.662 11.04 ;
      RECT 2.272 9.84 2.484 10.32 ;
      RECT 2.528 9.84 2.572 10.32 ;
      RECT 1.838 9.6 2.484 9.84 ;
      RECT 2.528 9.6 2.662 9.84 ;
      RECT 2.272 9.12 2.484 9.6 ;
      RECT 2.528 9.12 2.572 9.6 ;
      RECT 2.272 8.88 2.572 9.12 ;
      RECT 1.838 8.4 2.228 9.6 ;
      RECT 2.616 8.4 2.662 9.6 ;
      RECT 2.272 8.4 2.484 8.88 ;
      RECT 2.528 8.4 2.572 8.88 ;
      RECT 1.838 8.16 2.484 8.4 ;
      RECT 2.528 8.16 2.662 8.4 ;
      RECT 2.272 7.68 2.484 8.16 ;
      RECT 2.528 7.68 2.572 8.16 ;
      RECT 2.272 7.44 2.572 7.68 ;
      RECT 1.838 6.96 2.228 8.16 ;
      RECT 2.616 6.96 2.662 8.16 ;
      RECT 2.272 6.96 2.484 7.44 ;
      RECT 2.528 6.96 2.572 7.44 ;
      RECT 1.838 6.72 2.484 6.96 ;
      RECT 2.528 6.72 2.662 6.96 ;
      RECT 2.272 6.24 2.484 6.72 ;
      RECT 2.528 6.24 2.572 6.72 ;
      RECT 2.272 6 2.572 6.24 ;
      RECT 1.838 5.52 2.228 6.72 ;
      RECT 2.616 5.52 2.662 6.72 ;
      RECT 2.272 5.52 2.484 6 ;
      RECT 2.528 5.52 2.572 6 ;
      RECT 1.838 5.28 2.484 5.52 ;
      RECT 2.528 5.28 2.662 5.52 ;
      RECT 2.272 4.8 2.484 5.28 ;
      RECT 2.528 4.8 2.572 5.28 ;
      RECT 1.838 4.08 2.228 5.28 ;
      RECT 2.616 4.08 2.662 5.28 ;
      RECT 2.272 4.08 2.572 4.8 ;
      RECT 1.838 3.72 2.662 4.08 ;
      RECT 1.838 2.52 1.972 3.72 ;
      RECT 2.016 2.52 2.484 3.72 ;
      RECT 2.528 2.52 2.662 3.72 ;
      RECT 1.838 1.8 2.662 2.52 ;
      RECT 1.838 0.6 1.884 1.8 ;
      RECT 1.928 0.6 2.228 1.8 ;
      RECT 2.272 0.6 2.572 1.8 ;
      RECT 2.616 0.6 2.662 1.8 ;
      RECT 1.838 -0.12 2.662 0.6 ;
      RECT 0.938 3.72 1.762 22.2 ;
      RECT 0.938 2.52 0.984 3.72 ;
      RECT 1.028 2.52 1.328 3.72 ;
      RECT 1.372 2.52 1.672 3.72 ;
      RECT 1.716 2.52 1.762 3.72 ;
      RECT 0.938 1.8 1.762 2.52 ;
      RECT 0.938 0.6 1.072 1.8 ;
      RECT 1.116 0.6 1.584 1.8 ;
      RECT 1.628 0.6 1.762 1.8 ;
      RECT 0.938 -0.12 1.762 0.6 ;
      RECT -0.04 22.14 0.862 22.2 ;
      RECT -0.092 3.72 0.862 22.14 ;
      RECT -0.092 2.52 0.684 3.72 ;
      RECT 0.728 2.52 0.862 3.72 ;
      RECT -0.092 1.8 0.862 2.52 ;
      RECT -0.092 0.6 0.428 1.8 ;
      RECT 0.472 0.6 0.772 1.8 ;
      RECT 0.816 0.6 0.862 1.8 ;
      RECT -0.092 -0.06 0.862 0.6 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 11.858 0 12.52 22.08 ;
      RECT 10.958 0 11.542 22.08 ;
      RECT 10.058 0 10.642 22.08 ;
      RECT 9.158 0 9.742 22.08 ;
      RECT 8.258 0 8.842 22.08 ;
      RECT 7.358 0 7.942 22.08 ;
      RECT 6.458 0 7.042 22.08 ;
      RECT 5.558 0 6.142 22.08 ;
      RECT 4.658 0 5.242 22.08 ;
      RECT 3.758 21.96 4.342 22.08 ;
      RECT 4.192 21.24 4.342 21.96 ;
      RECT 3.758 5.4 3.908 21.96 ;
      RECT 3.848 4.68 3.908 5.4 ;
      RECT 3.848 3.96 4.164 4.68 ;
      RECT 3.758 3.84 4.342 3.96 ;
      RECT 3.936 2.4 4.342 3.84 ;
      RECT 3.758 1.92 4.342 2.4 ;
      RECT 3.848 0.48 3.908 1.92 ;
      RECT 4.192 0.48 4.342 1.92 ;
      RECT 3.758 0 4.342 0.48 ;
      RECT 2.858 21.96 3.442 22.08 ;
      RECT 2.948 4.68 3.264 21.96 ;
      RECT 2.858 3.84 3.442 4.68 ;
      RECT 2.948 2.4 3.008 3.84 ;
      RECT 3.292 2.4 3.352 3.84 ;
      RECT 2.858 1.92 3.442 2.4 ;
      RECT 3.036 0.48 3.264 1.92 ;
      RECT 2.858 0 3.442 0.48 ;
      RECT 1.958 21.96 2.542 22.08 ;
      RECT 1.958 21.24 2.364 21.96 ;
      RECT 1.958 3.96 2.108 21.24 ;
      RECT 2.392 3.96 2.452 4.68 ;
      RECT 1.958 3.84 2.542 3.96 ;
      RECT 2.136 2.4 2.364 3.84 ;
      RECT 1.958 1.92 2.542 2.4 ;
      RECT 2.048 0.48 2.108 1.92 ;
      RECT 2.392 0.48 2.452 1.92 ;
      RECT 1.958 0 2.542 0.48 ;
      RECT 1.058 3.84 1.642 22.08 ;
      RECT 1.148 2.4 1.208 3.84 ;
      RECT 1.492 2.4 1.552 3.84 ;
      RECT 1.058 1.92 1.642 2.4 ;
      RECT 1.236 0.48 1.464 1.92 ;
      RECT 1.058 0 1.642 0.48 ;
      RECT 0.08 3.84 0.742 22.08 ;
      RECT 0.08 2.4 0.564 3.84 ;
      RECT 0.08 1.92 0.742 2.4 ;
      RECT 0.08 0.48 0.308 1.92 ;
      RECT 0.592 0.48 0.652 1.92 ;
      RECT 0.08 0 0.742 0.48 ;
    LAYER m0 ;
      RECT 0 0.002 12.6 22.078 ;
    LAYER m1 ;
      RECT 0 0 12.6 22.08 ;
    LAYER m2 ;
      RECT 0 0.015 12.6 22.065 ;
    LAYER m3 ;
      RECT 0.015 0 12.585 22.08 ;
    LAYER m4 ;
      RECT 0 0.02 12.6 22.06 ;
    LAYER m5 ;
      RECT 0.012 0 12.588 22.08 ;
    LAYER m6 ;
      RECT 0 0.012 12.6 22.068 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf046b032e1r1w0cbbehraa4acw

END LIBRARY
