VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf028b256e2r2w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf028b256e2r2w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 81 BY 22.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 12.12 35.828 13.32 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 12.12 40.156 13.32 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 9.24 35.828 10.44 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 9.24 40.416 10.44 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 12.12 38.188 13.32 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 12.12 38.356 13.32 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 12.12 38.616 13.32 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 12.12 38.916 13.32 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 12.12 39.172 13.32 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 12.12 39.428 13.32 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 12.12 39.728 13.32 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 12.12 39.988 13.32 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.072 12.12 37.116 13.32 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.328 12.12 37.372 13.32 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 12.12 41.528 13.32 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 12.12 41.788 13.32 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 12.12 41.956 13.32 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 12.12 42.216 13.32 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 12.12 42.516 13.32 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 12.12 42.772 13.32 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 12.12 43.028 13.32 ;
    END
  END rdaddrp1[6]
  PIN rdaddrp1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 12.12 43.328 13.32 ;
    END
  END rdaddrp1[7]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 12.12 40.416 13.32 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 12.12 40.716 13.32 ;
    END
  END rdaddrp1_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.584 12.12 37.628 13.32 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 12.12 40.972 13.32 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 12.12 37.928 13.32 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 12.12 41.228 13.32 ;
    END
  END sdl_initp1
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 9.24 38.356 10.44 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 9.24 38.616 10.44 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 9.24 38.916 10.44 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 9.24 39.172 10.44 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 9.24 39.428 10.44 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 9.24 39.728 10.44 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 9.24 39.988 10.44 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 9.24 40.156 10.44 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.072 9.24 37.116 10.44 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.328 9.24 37.372 10.44 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 9.24 41.956 10.44 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 9.24 42.216 10.44 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 9.24 42.516 10.44 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 9.24 42.772 10.44 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 9.24 43.028 10.44 ;
    END
  END wraddrp1[4]
  PIN wraddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 9.24 43.328 10.44 ;
    END
  END wraddrp1[5]
  PIN wraddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 9.24 43.588 10.44 ;
    END
  END wraddrp1[6]
  PIN wraddrp1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 9.24 43.756 10.44 ;
    END
  END wraddrp1[7]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 9.24 40.716 10.44 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 9.24 40.972 10.44 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 0.36 35.828 1.56 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 5.16 41.956 6.36 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 5.16 42.128 6.36 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 6.12 43.028 7.32 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 6.12 43.116 7.32 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 7.08 35.916 8.28 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 7.08 36.128 8.28 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 14.28 36.128 15.48 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 14.28 36.216 15.48 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.972 15.24 38.016 16.44 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 15.24 38.188 16.44 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 0.36 35.916 1.56 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 16.2 39.088 17.4 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 16.2 39.172 17.4 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.028 17.16 40.072 18.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 17.16 40.156 18.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.012 18.12 41.056 19.32 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 18.12 41.228 19.32 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 19.08 42.128 20.28 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 19.08 42.216 20.28 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 20.04 43.116 21.24 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 20.04 43.328 21.24 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 1.32 37.928 2.52 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.972 1.32 38.016 2.52 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 2.28 38.916 3.48 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 2.28 39.088 3.48 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 3.24 39.988 4.44 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.028 3.24 40.072 4.44 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 4.2 40.972 5.4 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.012 4.2 41.056 5.4 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 9.24 37.928 10.44 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 9.24 38.188 10.44 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 0.36 36.128 1.56 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 5.16 42.216 6.36 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 5.16 42.428 6.36 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 6.12 43.328 7.32 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 6.12 43.416 7.32 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 7.08 36.216 8.28 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 7.08 36.388 8.28 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 14.28 36.388 15.48 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 14.28 36.472 15.48 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.228 15.24 38.272 16.44 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 15.24 38.356 16.44 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 0.36 36.216 1.56 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 16.2 39.256 17.4 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 16.2 39.428 17.4 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 17.16 40.328 18.36 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 17.16 40.416 18.36 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.272 18.12 41.316 19.32 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 18.12 41.528 19.32 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 19.08 42.428 20.28 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 19.08 42.516 20.28 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 20.04 43.416 21.24 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 20.04 43.588 21.24 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 1.32 38.188 2.52 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.228 1.32 38.272 2.52 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 2.28 39.172 3.48 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 2.28 39.256 3.48 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 3.24 40.156 4.44 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 3.24 40.328 4.44 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 4.2 41.228 5.4 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.272 4.2 41.316 5.4 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 9.24 41.528 10.44 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 9.24 41.788 10.44 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.584 9.24 37.628 10.44 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 9.24 41.228 10.44 ;
    END
  END wrenp1
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 0.36 36.388 1.56 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 5.16 42.516 6.36 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.644 5.16 42.688 6.36 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 6.12 43.588 7.32 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 6.12 43.672 7.32 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 7.08 36.472 8.28 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 7.08 36.556 8.28 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 14.28 36.556 15.48 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 14.28 36.728 15.48 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.484 15.24 38.528 16.44 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 15.24 38.616 16.44 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 0.36 36.472 1.56 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 16.2 39.516 17.4 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 16.2 39.728 17.4 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.584 17.16 40.628 18.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 17.16 40.716 18.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.572 18.12 41.616 19.32 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 18.12 41.788 19.32 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.644 19.08 42.688 20.28 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 19.08 42.772 20.28 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 20.04 43.672 21.24 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 20.04 43.756 21.24 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 1.32 38.356 2.52 ;
    END
  END rddatap0[2]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.484 1.32 38.528 2.52 ;
    END
  END rddatap0[3]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 2.28 39.428 3.48 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 2.28 39.516 3.48 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 3.24 40.416 4.44 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.584 3.24 40.628 4.44 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 4.2 41.528 5.4 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.572 4.2 41.616 5.4 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 0.36 36.556 1.56 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 5.16 42.772 6.36 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.812 5.16 42.856 6.36 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 6.12 43.756 7.32 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.884 6.12 43.928 7.32 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 7.08 36.728 8.28 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.772 7.08 36.816 8.28 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.772 14.28 36.816 15.48 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.984 14.28 37.028 15.48 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 15.24 38.828 16.44 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 15.24 38.916 16.44 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 0.36 36.728 1.56 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 16.2 39.816 17.4 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 16.2 39.988 17.4 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.844 17.16 40.888 18.36 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 17.16 40.972 18.36 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.828 18.12 41.872 19.32 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 18.12 41.956 19.32 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.812 19.08 42.856 20.28 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 19.08 43.028 20.28 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.884 20.04 43.928 21.24 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 20.04 35.916 21.24 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 1.32 38.616 2.52 ;
    END
  END rddatap1[2]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 1.32 38.828 2.52 ;
    END
  END rddatap1[3]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 2.28 39.728 3.48 ;
    END
  END rddatap1[4]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 2.28 39.816 3.48 ;
    END
  END rddatap1[5]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 3.24 40.716 4.44 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.844 3.24 40.888 4.44 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 4.2 41.788 5.4 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.828 4.2 41.872 5.4 ;
    END
  END rddatap1[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 22.02 ;
        RECT 2.662 0.06 2.738 22.02 ;
        RECT 4.462 0.06 4.538 22.02 ;
        RECT 6.262 0.06 6.338 22.02 ;
        RECT 8.062 0.06 8.138 22.02 ;
        RECT 9.862 0.06 9.938 22.02 ;
        RECT 11.662 0.06 11.738 22.02 ;
        RECT 13.462 0.06 13.538 22.02 ;
        RECT 15.262 0.06 15.338 22.02 ;
        RECT 17.062 0.06 17.138 22.02 ;
        RECT 18.862 0.06 18.938 22.02 ;
        RECT 20.662 0.06 20.738 22.02 ;
        RECT 22.462 0.06 22.538 22.02 ;
        RECT 24.262 0.06 24.338 22.02 ;
        RECT 26.062 0.06 26.138 22.02 ;
        RECT 27.862 0.06 27.938 22.02 ;
        RECT 29.662 0.06 29.738 22.02 ;
        RECT 31.462 0.06 31.538 22.02 ;
        RECT 33.262 0.06 33.338 22.02 ;
        RECT 35.062 0.06 35.138 22.02 ;
        RECT 36.862 0.06 36.938 22.02 ;
        RECT 38.662 0.06 38.738 22.02 ;
        RECT 40.462 0.06 40.538 22.02 ;
        RECT 42.262 0.06 42.338 22.02 ;
        RECT 44.062 0.06 44.138 22.02 ;
        RECT 45.862 0.06 45.938 22.02 ;
        RECT 47.662 0.06 47.738 22.02 ;
        RECT 49.462 0.06 49.538 22.02 ;
        RECT 51.262 0.06 51.338 22.02 ;
        RECT 53.062 0.06 53.138 22.02 ;
        RECT 54.862 0.06 54.938 22.02 ;
        RECT 56.662 0.06 56.738 22.02 ;
        RECT 58.462 0.06 58.538 22.02 ;
        RECT 60.262 0.06 60.338 22.02 ;
        RECT 62.062 0.06 62.138 22.02 ;
        RECT 63.862 0.06 63.938 22.02 ;
        RECT 65.662 0.06 65.738 22.02 ;
        RECT 67.462 0.06 67.538 22.02 ;
        RECT 69.262 0.06 69.338 22.02 ;
        RECT 71.062 0.06 71.138 22.02 ;
        RECT 72.862 0.06 72.938 22.02 ;
        RECT 74.662 0.06 74.738 22.02 ;
        RECT 76.462 0.06 76.538 22.02 ;
        RECT 78.262 0.06 78.338 22.02 ;
        RECT 80.062 0.06 80.138 22.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 22.02 ;
        RECT 3.562 0.06 3.638 22.02 ;
        RECT 5.362 0.06 5.438 22.02 ;
        RECT 7.162 0.06 7.238 22.02 ;
        RECT 8.962 0.06 9.038 22.02 ;
        RECT 10.762 0.06 10.838 22.02 ;
        RECT 12.562 0.06 12.638 22.02 ;
        RECT 14.362 0.06 14.438 22.02 ;
        RECT 16.162 0.06 16.238 22.02 ;
        RECT 17.962 0.06 18.038 22.02 ;
        RECT 19.762 0.06 19.838 22.02 ;
        RECT 21.562 0.06 21.638 22.02 ;
        RECT 23.362 0.06 23.438 22.02 ;
        RECT 25.162 0.06 25.238 22.02 ;
        RECT 26.962 0.06 27.038 22.02 ;
        RECT 28.762 0.06 28.838 22.02 ;
        RECT 30.562 0.06 30.638 22.02 ;
        RECT 32.362 0.06 32.438 22.02 ;
        RECT 34.162 0.06 34.238 22.02 ;
        RECT 35.962 0.06 36.038 22.02 ;
        RECT 37.762 0.06 37.838 22.02 ;
        RECT 39.562 0.06 39.638 22.02 ;
        RECT 41.362 0.06 41.438 22.02 ;
        RECT 43.162 0.06 43.238 22.02 ;
        RECT 44.962 0.06 45.038 22.02 ;
        RECT 46.762 0.06 46.838 22.02 ;
        RECT 48.562 0.06 48.638 22.02 ;
        RECT 50.362 0.06 50.438 22.02 ;
        RECT 52.162 0.06 52.238 22.02 ;
        RECT 53.962 0.06 54.038 22.02 ;
        RECT 55.762 0.06 55.838 22.02 ;
        RECT 57.562 0.06 57.638 22.02 ;
        RECT 59.362 0.06 59.438 22.02 ;
        RECT 61.162 0.06 61.238 22.02 ;
        RECT 62.962 0.06 63.038 22.02 ;
        RECT 64.762 0.06 64.838 22.02 ;
        RECT 66.562 0.06 66.638 22.02 ;
        RECT 68.362 0.06 68.438 22.02 ;
        RECT 70.162 0.06 70.238 22.02 ;
        RECT 71.962 0.06 72.038 22.02 ;
        RECT 73.762 0.06 73.838 22.02 ;
        RECT 75.562 0.06 75.638 22.02 ;
        RECT 77.362 0.06 77.438 22.02 ;
        RECT 79.162 0.06 79.238 22.02 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 81.016 22.094 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 81.02 22.1 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 81.0705 22.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 81.035 22.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 81.07 22.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 81.059 22.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 81.09 22.142 ;
    LAYER m7 SPACING 0 ;
      RECT 80.138 22.14 81.04 22.2 ;
      RECT 80.138 -0.06 81.092 22.14 ;
      RECT 80.138 -0.12 81.04 -0.06 ;
      RECT 79.238 -0.12 80.062 22.2 ;
      RECT 78.338 -0.12 79.162 22.2 ;
      RECT 77.438 -0.12 78.262 22.2 ;
      RECT 76.538 -0.12 77.362 22.2 ;
      RECT 75.638 -0.12 76.462 22.2 ;
      RECT 74.738 -0.12 75.562 22.2 ;
      RECT 73.838 -0.12 74.662 22.2 ;
      RECT 72.938 -0.12 73.762 22.2 ;
      RECT 72.038 -0.12 72.862 22.2 ;
      RECT 71.138 -0.12 71.962 22.2 ;
      RECT 70.238 -0.12 71.062 22.2 ;
      RECT 69.338 -0.12 70.162 22.2 ;
      RECT 68.438 -0.12 69.262 22.2 ;
      RECT 67.538 -0.12 68.362 22.2 ;
      RECT 66.638 -0.12 67.462 22.2 ;
      RECT 65.738 -0.12 66.562 22.2 ;
      RECT 64.838 -0.12 65.662 22.2 ;
      RECT 63.938 -0.12 64.762 22.2 ;
      RECT 63.038 -0.12 63.862 22.2 ;
      RECT 62.138 -0.12 62.962 22.2 ;
      RECT 61.238 -0.12 62.062 22.2 ;
      RECT 60.338 -0.12 61.162 22.2 ;
      RECT 59.438 -0.12 60.262 22.2 ;
      RECT 58.538 -0.12 59.362 22.2 ;
      RECT 57.638 -0.12 58.462 22.2 ;
      RECT 56.738 -0.12 57.562 22.2 ;
      RECT 55.838 -0.12 56.662 22.2 ;
      RECT 54.938 -0.12 55.762 22.2 ;
      RECT 54.038 -0.12 54.862 22.2 ;
      RECT 53.138 -0.12 53.962 22.2 ;
      RECT 52.238 -0.12 53.062 22.2 ;
      RECT 51.338 -0.12 52.162 22.2 ;
      RECT 50.438 -0.12 51.262 22.2 ;
      RECT 49.538 -0.12 50.362 22.2 ;
      RECT 48.638 -0.12 49.462 22.2 ;
      RECT 47.738 -0.12 48.562 22.2 ;
      RECT 46.838 -0.12 47.662 22.2 ;
      RECT 45.938 -0.12 46.762 22.2 ;
      RECT 45.038 -0.12 45.862 22.2 ;
      RECT 44.138 -0.12 44.962 22.2 ;
      RECT 43.238 21.24 44.062 22.2 ;
      RECT 43.238 20.04 43.284 21.24 ;
      RECT 43.328 20.04 43.372 21.24 ;
      RECT 43.416 20.04 43.544 21.24 ;
      RECT 43.588 20.04 43.628 21.24 ;
      RECT 43.672 20.04 43.712 21.24 ;
      RECT 43.756 20.04 43.884 21.24 ;
      RECT 43.928 20.04 44.062 21.24 ;
      RECT 43.238 13.32 44.062 20.04 ;
      RECT 43.238 12.12 43.284 13.32 ;
      RECT 43.328 12.12 44.062 13.32 ;
      RECT 43.238 10.44 44.062 12.12 ;
      RECT 43.238 9.24 43.284 10.44 ;
      RECT 43.328 9.24 43.544 10.44 ;
      RECT 43.588 9.24 43.712 10.44 ;
      RECT 43.756 9.24 44.062 10.44 ;
      RECT 43.238 7.32 44.062 9.24 ;
      RECT 43.238 6.12 43.284 7.32 ;
      RECT 43.328 6.12 43.372 7.32 ;
      RECT 43.416 6.12 43.544 7.32 ;
      RECT 43.588 6.12 43.628 7.32 ;
      RECT 43.672 6.12 43.712 7.32 ;
      RECT 43.756 6.12 43.884 7.32 ;
      RECT 43.928 6.12 44.062 7.32 ;
      RECT 43.238 -0.12 44.062 6.12 ;
      RECT 42.338 21.24 43.162 22.2 ;
      RECT 42.338 20.28 43.072 21.24 ;
      RECT 43.116 20.04 43.162 21.24 ;
      RECT 43.028 20.04 43.072 20.28 ;
      RECT 42.338 19.08 42.384 20.28 ;
      RECT 42.428 19.08 42.472 20.28 ;
      RECT 42.516 19.08 42.644 20.28 ;
      RECT 42.688 19.08 42.728 20.28 ;
      RECT 42.772 19.08 42.812 20.28 ;
      RECT 42.856 19.08 42.984 20.28 ;
      RECT 43.028 19.08 43.162 20.04 ;
      RECT 42.338 13.32 43.162 19.08 ;
      RECT 42.338 12.12 42.472 13.32 ;
      RECT 42.516 12.12 42.728 13.32 ;
      RECT 42.772 12.12 42.984 13.32 ;
      RECT 43.028 12.12 43.162 13.32 ;
      RECT 42.338 10.44 43.162 12.12 ;
      RECT 42.338 9.24 42.472 10.44 ;
      RECT 42.516 9.24 42.728 10.44 ;
      RECT 42.772 9.24 42.984 10.44 ;
      RECT 43.028 9.24 43.162 10.44 ;
      RECT 42.338 7.32 43.162 9.24 ;
      RECT 42.338 6.36 42.984 7.32 ;
      RECT 43.028 6.12 43.072 7.32 ;
      RECT 43.116 6.12 43.162 7.32 ;
      RECT 42.856 6.12 42.984 6.36 ;
      RECT 42.338 5.16 42.384 6.36 ;
      RECT 42.428 5.16 42.472 6.36 ;
      RECT 42.516 5.16 42.644 6.36 ;
      RECT 42.688 5.16 42.728 6.36 ;
      RECT 42.772 5.16 42.812 6.36 ;
      RECT 42.856 5.16 43.162 6.12 ;
      RECT 42.338 -0.12 43.162 5.16 ;
      RECT 41.438 20.28 42.262 22.2 ;
      RECT 41.438 19.32 42.084 20.28 ;
      RECT 42.128 19.08 42.172 20.28 ;
      RECT 42.216 19.08 42.262 20.28 ;
      RECT 41.956 19.08 42.084 19.32 ;
      RECT 41.438 18.12 41.484 19.32 ;
      RECT 41.528 18.12 41.572 19.32 ;
      RECT 41.616 18.12 41.744 19.32 ;
      RECT 41.788 18.12 41.828 19.32 ;
      RECT 41.872 18.12 41.912 19.32 ;
      RECT 41.956 18.12 42.262 19.08 ;
      RECT 41.438 13.32 42.262 18.12 ;
      RECT 41.438 12.12 41.484 13.32 ;
      RECT 41.528 12.12 41.744 13.32 ;
      RECT 41.788 12.12 41.912 13.32 ;
      RECT 41.956 12.12 42.172 13.32 ;
      RECT 42.216 12.12 42.262 13.32 ;
      RECT 41.438 10.44 42.262 12.12 ;
      RECT 41.438 9.24 41.484 10.44 ;
      RECT 41.528 9.24 41.744 10.44 ;
      RECT 41.788 9.24 41.912 10.44 ;
      RECT 41.956 9.24 42.172 10.44 ;
      RECT 42.216 9.24 42.262 10.44 ;
      RECT 41.438 6.36 42.262 9.24 ;
      RECT 41.438 5.4 41.912 6.36 ;
      RECT 41.956 5.16 42.084 6.36 ;
      RECT 42.128 5.16 42.172 6.36 ;
      RECT 42.216 5.16 42.262 6.36 ;
      RECT 41.872 5.16 41.912 5.4 ;
      RECT 41.438 4.2 41.484 5.4 ;
      RECT 41.528 4.2 41.572 5.4 ;
      RECT 41.616 4.2 41.744 5.4 ;
      RECT 41.788 4.2 41.828 5.4 ;
      RECT 41.872 4.2 42.262 5.16 ;
      RECT 41.438 -0.12 42.262 4.2 ;
      RECT 40.538 19.32 41.362 22.2 ;
      RECT 40.538 18.36 41.012 19.32 ;
      RECT 41.056 18.12 41.184 19.32 ;
      RECT 41.228 18.12 41.272 19.32 ;
      RECT 41.316 18.12 41.362 19.32 ;
      RECT 40.972 18.12 41.012 18.36 ;
      RECT 40.538 17.16 40.584 18.36 ;
      RECT 40.628 17.16 40.672 18.36 ;
      RECT 40.716 17.16 40.844 18.36 ;
      RECT 40.888 17.16 40.928 18.36 ;
      RECT 40.972 17.16 41.362 18.12 ;
      RECT 40.538 13.32 41.362 17.16 ;
      RECT 40.538 12.12 40.672 13.32 ;
      RECT 40.716 12.12 40.928 13.32 ;
      RECT 40.972 12.12 41.184 13.32 ;
      RECT 41.228 12.12 41.362 13.32 ;
      RECT 40.538 10.44 41.362 12.12 ;
      RECT 40.538 9.24 40.672 10.44 ;
      RECT 40.716 9.24 40.928 10.44 ;
      RECT 40.972 9.24 41.184 10.44 ;
      RECT 41.228 9.24 41.362 10.44 ;
      RECT 40.538 5.4 41.362 9.24 ;
      RECT 40.538 4.44 40.928 5.4 ;
      RECT 40.972 4.2 41.012 5.4 ;
      RECT 41.056 4.2 41.184 5.4 ;
      RECT 41.228 4.2 41.272 5.4 ;
      RECT 41.316 4.2 41.362 5.4 ;
      RECT 40.888 4.2 40.928 4.44 ;
      RECT 40.538 3.24 40.584 4.44 ;
      RECT 40.628 3.24 40.672 4.44 ;
      RECT 40.716 3.24 40.844 4.44 ;
      RECT 40.888 3.24 41.362 4.2 ;
      RECT 40.538 -0.12 41.362 3.24 ;
      RECT 39.638 18.36 40.462 22.2 ;
      RECT 39.638 17.4 40.028 18.36 ;
      RECT 40.072 17.16 40.112 18.36 ;
      RECT 40.156 17.16 40.284 18.36 ;
      RECT 40.328 17.16 40.372 18.36 ;
      RECT 40.416 17.16 40.462 18.36 ;
      RECT 39.988 17.16 40.028 17.4 ;
      RECT 39.638 16.2 39.684 17.4 ;
      RECT 39.728 16.2 39.772 17.4 ;
      RECT 39.816 16.2 39.944 17.4 ;
      RECT 39.988 16.2 40.462 17.16 ;
      RECT 39.638 13.32 40.462 16.2 ;
      RECT 39.638 12.12 39.684 13.32 ;
      RECT 39.728 12.12 39.944 13.32 ;
      RECT 39.988 12.12 40.112 13.32 ;
      RECT 40.156 12.12 40.372 13.32 ;
      RECT 40.416 12.12 40.462 13.32 ;
      RECT 39.638 10.44 40.462 12.12 ;
      RECT 39.638 9.24 39.684 10.44 ;
      RECT 39.728 9.24 39.944 10.44 ;
      RECT 39.988 9.24 40.112 10.44 ;
      RECT 40.156 9.24 40.372 10.44 ;
      RECT 40.416 9.24 40.462 10.44 ;
      RECT 39.638 4.44 40.462 9.24 ;
      RECT 39.638 3.48 39.944 4.44 ;
      RECT 39.988 3.24 40.028 4.44 ;
      RECT 40.072 3.24 40.112 4.44 ;
      RECT 40.156 3.24 40.284 4.44 ;
      RECT 40.328 3.24 40.372 4.44 ;
      RECT 40.416 3.24 40.462 4.44 ;
      RECT 39.816 3.24 39.944 3.48 ;
      RECT 39.638 2.28 39.684 3.48 ;
      RECT 39.728 2.28 39.772 3.48 ;
      RECT 39.816 2.28 40.462 3.24 ;
      RECT 39.638 -0.12 40.462 2.28 ;
      RECT 38.738 17.4 39.562 22.2 ;
      RECT 38.738 16.44 39.044 17.4 ;
      RECT 39.088 16.2 39.128 17.4 ;
      RECT 39.172 16.2 39.212 17.4 ;
      RECT 39.256 16.2 39.384 17.4 ;
      RECT 39.428 16.2 39.472 17.4 ;
      RECT 39.516 16.2 39.562 17.4 ;
      RECT 38.916 16.2 39.044 16.44 ;
      RECT 38.738 15.24 38.784 16.44 ;
      RECT 38.828 15.24 38.872 16.44 ;
      RECT 38.916 15.24 39.562 16.2 ;
      RECT 38.738 13.32 39.562 15.24 ;
      RECT 38.738 12.12 38.872 13.32 ;
      RECT 38.916 12.12 39.128 13.32 ;
      RECT 39.172 12.12 39.384 13.32 ;
      RECT 39.428 12.12 39.562 13.32 ;
      RECT 38.738 10.44 39.562 12.12 ;
      RECT 38.738 9.24 38.872 10.44 ;
      RECT 38.916 9.24 39.128 10.44 ;
      RECT 39.172 9.24 39.384 10.44 ;
      RECT 39.428 9.24 39.562 10.44 ;
      RECT 38.738 3.48 39.562 9.24 ;
      RECT 38.738 2.52 38.872 3.48 ;
      RECT 38.916 2.28 39.044 3.48 ;
      RECT 39.088 2.28 39.128 3.48 ;
      RECT 39.172 2.28 39.212 3.48 ;
      RECT 39.256 2.28 39.384 3.48 ;
      RECT 39.428 2.28 39.472 3.48 ;
      RECT 39.516 2.28 39.562 3.48 ;
      RECT 38.828 2.28 38.872 2.52 ;
      RECT 38.738 1.32 38.784 2.52 ;
      RECT 38.828 1.32 39.562 2.28 ;
      RECT 38.738 -0.12 39.562 1.32 ;
      RECT 37.838 16.44 38.662 22.2 ;
      RECT 37.838 15.24 37.972 16.44 ;
      RECT 38.016 15.24 38.144 16.44 ;
      RECT 38.188 15.24 38.228 16.44 ;
      RECT 38.272 15.24 38.312 16.44 ;
      RECT 38.356 15.24 38.484 16.44 ;
      RECT 38.528 15.24 38.572 16.44 ;
      RECT 38.616 15.24 38.662 16.44 ;
      RECT 37.838 13.32 38.662 15.24 ;
      RECT 37.838 12.12 37.884 13.32 ;
      RECT 37.928 12.12 38.144 13.32 ;
      RECT 38.188 12.12 38.312 13.32 ;
      RECT 38.356 12.12 38.572 13.32 ;
      RECT 38.616 12.12 38.662 13.32 ;
      RECT 37.838 10.44 38.662 12.12 ;
      RECT 37.838 9.24 37.884 10.44 ;
      RECT 37.928 9.24 38.144 10.44 ;
      RECT 38.188 9.24 38.312 10.44 ;
      RECT 38.356 9.24 38.572 10.44 ;
      RECT 38.616 9.24 38.662 10.44 ;
      RECT 37.838 2.52 38.662 9.24 ;
      RECT 37.838 1.32 37.884 2.52 ;
      RECT 37.928 1.32 37.972 2.52 ;
      RECT 38.016 1.32 38.144 2.52 ;
      RECT 38.188 1.32 38.228 2.52 ;
      RECT 38.272 1.32 38.312 2.52 ;
      RECT 38.356 1.32 38.484 2.52 ;
      RECT 38.528 1.32 38.572 2.52 ;
      RECT 38.616 1.32 38.662 2.52 ;
      RECT 37.838 -0.12 38.662 1.32 ;
      RECT 36.938 15.48 37.762 22.2 ;
      RECT 36.938 14.28 36.984 15.48 ;
      RECT 37.028 14.28 37.762 15.48 ;
      RECT 36.938 13.32 37.762 14.28 ;
      RECT 36.938 12.12 37.072 13.32 ;
      RECT 37.116 12.12 37.328 13.32 ;
      RECT 37.372 12.12 37.584 13.32 ;
      RECT 37.628 12.12 37.762 13.32 ;
      RECT 36.938 10.44 37.762 12.12 ;
      RECT 36.938 9.24 37.072 10.44 ;
      RECT 37.116 9.24 37.328 10.44 ;
      RECT 37.372 9.24 37.584 10.44 ;
      RECT 37.628 9.24 37.762 10.44 ;
      RECT 36.938 -0.12 37.762 9.24 ;
      RECT 36.038 15.48 36.862 22.2 ;
      RECT 36.038 14.28 36.084 15.48 ;
      RECT 36.128 14.28 36.172 15.48 ;
      RECT 36.216 14.28 36.344 15.48 ;
      RECT 36.388 14.28 36.428 15.48 ;
      RECT 36.472 14.28 36.512 15.48 ;
      RECT 36.556 14.28 36.684 15.48 ;
      RECT 36.728 14.28 36.772 15.48 ;
      RECT 36.816 14.28 36.862 15.48 ;
      RECT 36.038 8.28 36.862 14.28 ;
      RECT 36.038 7.08 36.084 8.28 ;
      RECT 36.128 7.08 36.172 8.28 ;
      RECT 36.216 7.08 36.344 8.28 ;
      RECT 36.388 7.08 36.428 8.28 ;
      RECT 36.472 7.08 36.512 8.28 ;
      RECT 36.556 7.08 36.684 8.28 ;
      RECT 36.728 7.08 36.772 8.28 ;
      RECT 36.816 7.08 36.862 8.28 ;
      RECT 36.038 1.56 36.862 7.08 ;
      RECT 36.038 0.36 36.084 1.56 ;
      RECT 36.128 0.36 36.172 1.56 ;
      RECT 36.216 0.36 36.344 1.56 ;
      RECT 36.388 0.36 36.428 1.56 ;
      RECT 36.472 0.36 36.512 1.56 ;
      RECT 36.556 0.36 36.684 1.56 ;
      RECT 36.728 0.36 36.862 1.56 ;
      RECT 36.038 -0.12 36.862 0.36 ;
      RECT 35.138 21.24 35.962 22.2 ;
      RECT 35.138 20.04 35.872 21.24 ;
      RECT 35.916 20.04 35.962 21.24 ;
      RECT 35.138 13.32 35.962 20.04 ;
      RECT 35.138 12.12 35.784 13.32 ;
      RECT 35.828 12.12 35.962 13.32 ;
      RECT 35.138 10.44 35.962 12.12 ;
      RECT 35.138 9.24 35.784 10.44 ;
      RECT 35.828 9.24 35.962 10.44 ;
      RECT 35.138 8.28 35.962 9.24 ;
      RECT 35.138 7.08 35.872 8.28 ;
      RECT 35.916 7.08 35.962 8.28 ;
      RECT 35.138 1.56 35.962 7.08 ;
      RECT 35.138 0.36 35.784 1.56 ;
      RECT 35.828 0.36 35.872 1.56 ;
      RECT 35.916 0.36 35.962 1.56 ;
      RECT 35.138 -0.12 35.962 0.36 ;
      RECT 34.238 -0.12 35.062 22.2 ;
      RECT 33.338 -0.12 34.162 22.2 ;
      RECT 32.438 -0.12 33.262 22.2 ;
      RECT 31.538 -0.12 32.362 22.2 ;
      RECT 30.638 -0.12 31.462 22.2 ;
      RECT 29.738 -0.12 30.562 22.2 ;
      RECT 28.838 -0.12 29.662 22.2 ;
      RECT 27.938 -0.12 28.762 22.2 ;
      RECT 27.038 -0.12 27.862 22.2 ;
      RECT 26.138 -0.12 26.962 22.2 ;
      RECT 25.238 -0.12 26.062 22.2 ;
      RECT 24.338 -0.12 25.162 22.2 ;
      RECT 23.438 -0.12 24.262 22.2 ;
      RECT 22.538 -0.12 23.362 22.2 ;
      RECT 21.638 -0.12 22.462 22.2 ;
      RECT 20.738 -0.12 21.562 22.2 ;
      RECT 19.838 -0.12 20.662 22.2 ;
      RECT 18.938 -0.12 19.762 22.2 ;
      RECT 18.038 -0.12 18.862 22.2 ;
      RECT 17.138 -0.12 17.962 22.2 ;
      RECT 16.238 -0.12 17.062 22.2 ;
      RECT 15.338 -0.12 16.162 22.2 ;
      RECT 14.438 -0.12 15.262 22.2 ;
      RECT 13.538 -0.12 14.362 22.2 ;
      RECT 12.638 -0.12 13.462 22.2 ;
      RECT 11.738 -0.12 12.562 22.2 ;
      RECT 10.838 -0.12 11.662 22.2 ;
      RECT 9.938 -0.12 10.762 22.2 ;
      RECT 9.038 -0.12 9.862 22.2 ;
      RECT 8.138 -0.12 8.962 22.2 ;
      RECT 7.238 -0.12 8.062 22.2 ;
      RECT 6.338 -0.12 7.162 22.2 ;
      RECT 5.438 -0.12 6.262 22.2 ;
      RECT 4.538 -0.12 5.362 22.2 ;
      RECT 3.638 -0.12 4.462 22.2 ;
      RECT 2.738 -0.12 3.562 22.2 ;
      RECT 1.838 -0.12 2.662 22.2 ;
      RECT 0.938 -0.12 1.762 22.2 ;
      RECT -0.04 22.14 0.862 22.2 ;
      RECT -0.092 -0.06 0.862 22.14 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 80.258 0 80.92 22.08 ;
      RECT 79.358 0 79.942 22.08 ;
      RECT 78.458 0 79.042 22.08 ;
      RECT 77.558 0 78.142 22.08 ;
      RECT 76.658 0 77.242 22.08 ;
      RECT 75.758 0 76.342 22.08 ;
      RECT 74.858 0 75.442 22.08 ;
      RECT 73.958 0 74.542 22.08 ;
      RECT 73.058 0 73.642 22.08 ;
      RECT 72.158 0 72.742 22.08 ;
      RECT 71.258 0 71.842 22.08 ;
      RECT 70.358 0 70.942 22.08 ;
      RECT 69.458 0 70.042 22.08 ;
      RECT 68.558 0 69.142 22.08 ;
      RECT 67.658 0 68.242 22.08 ;
      RECT 66.758 0 67.342 22.08 ;
      RECT 65.858 0 66.442 22.08 ;
      RECT 64.958 0 65.542 22.08 ;
      RECT 64.058 0 64.642 22.08 ;
      RECT 63.158 0 63.742 22.08 ;
      RECT 62.258 0 62.842 22.08 ;
      RECT 61.358 0 61.942 22.08 ;
      RECT 60.458 0 61.042 22.08 ;
      RECT 59.558 0 60.142 22.08 ;
      RECT 58.658 0 59.242 22.08 ;
      RECT 57.758 0 58.342 22.08 ;
      RECT 56.858 0 57.442 22.08 ;
      RECT 55.958 0 56.542 22.08 ;
      RECT 55.058 0 55.642 22.08 ;
      RECT 54.158 0 54.742 22.08 ;
      RECT 53.258 0 53.842 22.08 ;
      RECT 52.358 0 52.942 22.08 ;
      RECT 51.458 0 52.042 22.08 ;
      RECT 50.558 0 51.142 22.08 ;
      RECT 49.658 0 50.242 22.08 ;
      RECT 48.758 0 49.342 22.08 ;
      RECT 47.858 0 48.442 22.08 ;
      RECT 46.958 0 47.542 22.08 ;
      RECT 46.058 0 46.642 22.08 ;
      RECT 45.158 0 45.742 22.08 ;
      RECT 44.258 0 44.842 22.08 ;
      RECT 43.358 21.36 43.942 22.08 ;
      RECT 42.458 21.36 43.042 22.08 ;
      RECT 42.458 20.4 42.952 21.36 ;
      RECT 41.558 20.4 42.142 22.08 ;
      RECT 41.558 19.44 41.964 20.4 ;
      RECT 40.658 19.44 41.242 22.08 ;
      RECT 40.658 18.48 40.892 19.44 ;
      RECT 39.758 18.48 40.342 22.08 ;
      RECT 39.758 17.52 39.908 18.48 ;
      RECT 38.858 17.52 39.442 22.08 ;
      RECT 38.858 16.56 38.924 17.52 ;
      RECT 37.958 16.56 38.542 22.08 ;
      RECT 37.058 15.6 37.642 22.08 ;
      RECT 37.148 14.16 37.642 15.6 ;
      RECT 37.058 13.44 37.642 14.16 ;
      RECT 36.158 15.6 36.742 22.08 ;
      RECT 35.258 21.36 35.842 22.08 ;
      RECT 35.258 19.92 35.752 21.36 ;
      RECT 35.258 13.44 35.842 19.92 ;
      RECT 35.258 12 35.664 13.44 ;
      RECT 35.258 10.56 35.842 12 ;
      RECT 35.258 9.12 35.664 10.56 ;
      RECT 35.258 8.4 35.842 9.12 ;
      RECT 35.258 6.96 35.752 8.4 ;
      RECT 35.258 1.68 35.842 6.96 ;
      RECT 35.258 0.24 35.664 1.68 ;
      RECT 35.258 0 35.842 0.24 ;
      RECT 34.358 0 34.942 22.08 ;
      RECT 33.458 0 34.042 22.08 ;
      RECT 32.558 0 33.142 22.08 ;
      RECT 31.658 0 32.242 22.08 ;
      RECT 30.758 0 31.342 22.08 ;
      RECT 29.858 0 30.442 22.08 ;
      RECT 28.958 0 29.542 22.08 ;
      RECT 28.058 0 28.642 22.08 ;
      RECT 27.158 0 27.742 22.08 ;
      RECT 26.258 0 26.842 22.08 ;
      RECT 25.358 0 25.942 22.08 ;
      RECT 24.458 0 25.042 22.08 ;
      RECT 23.558 0 24.142 22.08 ;
      RECT 22.658 0 23.242 22.08 ;
      RECT 21.758 0 22.342 22.08 ;
      RECT 20.858 0 21.442 22.08 ;
      RECT 19.958 0 20.542 22.08 ;
      RECT 19.058 0 19.642 22.08 ;
      RECT 18.158 0 18.742 22.08 ;
      RECT 17.258 0 17.842 22.08 ;
      RECT 16.358 0 16.942 22.08 ;
      RECT 15.458 0 16.042 22.08 ;
      RECT 14.558 0 15.142 22.08 ;
      RECT 13.658 0 14.242 22.08 ;
      RECT 12.758 0 13.342 22.08 ;
      RECT 11.858 0 12.442 22.08 ;
      RECT 10.958 0 11.542 22.08 ;
      RECT 10.058 0 10.642 22.08 ;
      RECT 9.158 0 9.742 22.08 ;
      RECT 8.258 0 8.842 22.08 ;
      RECT 7.358 0 7.942 22.08 ;
      RECT 6.458 0 7.042 22.08 ;
      RECT 5.558 0 6.142 22.08 ;
      RECT 4.658 0 5.242 22.08 ;
      RECT 3.758 0 4.342 22.08 ;
      RECT 2.858 0 3.442 22.08 ;
      RECT 1.958 0 2.542 22.08 ;
      RECT 1.058 0 1.642 22.08 ;
      RECT 0.08 0 0.742 22.08 ;
      RECT 43.358 13.44 43.942 19.92 ;
      RECT 43.448 12 43.942 13.44 ;
      RECT 43.358 10.56 43.942 12 ;
      RECT 43.876 9.12 43.942 10.56 ;
      RECT 43.358 7.44 43.942 9.12 ;
      RECT 42.458 13.44 43.042 18.96 ;
      RECT 42.076 18 42.142 18.96 ;
      RECT 41.558 13.44 42.142 18 ;
      RECT 41.092 17.04 41.242 18 ;
      RECT 40.658 13.44 41.242 17.04 ;
      RECT 40.108 16.08 40.342 17.04 ;
      RECT 39.758 13.44 40.342 16.08 ;
      RECT 39.036 15.12 39.442 16.08 ;
      RECT 38.858 13.44 39.442 15.12 ;
      RECT 37.958 13.44 38.542 15.12 ;
      RECT 36.158 8.4 36.742 14.16 ;
      RECT 42.458 10.56 43.042 12 ;
      RECT 41.558 10.56 42.142 12 ;
      RECT 40.658 10.56 41.242 12 ;
      RECT 39.758 10.56 40.342 12 ;
      RECT 38.858 10.56 39.442 12 ;
      RECT 37.958 10.56 38.542 12 ;
      RECT 37.058 10.56 37.642 12 ;
      RECT 42.458 7.44 43.042 9.12 ;
      RECT 42.458 6.48 42.864 7.44 ;
      RECT 41.558 6.48 42.142 9.12 ;
      RECT 41.558 5.52 41.792 6.48 ;
      RECT 40.658 5.52 41.242 9.12 ;
      RECT 40.658 4.56 40.808 5.52 ;
      RECT 39.758 4.56 40.342 9.12 ;
      RECT 39.758 3.6 39.824 4.56 ;
      RECT 38.858 3.6 39.442 9.12 ;
      RECT 37.958 2.64 38.542 9.12 ;
      RECT 37.058 0 37.642 9.12 ;
      RECT 36.158 1.68 36.742 6.96 ;
      RECT 43.358 0 43.942 6 ;
      RECT 42.976 5.04 43.042 6 ;
      RECT 42.458 0 43.042 5.04 ;
      RECT 41.992 4.08 42.142 5.04 ;
      RECT 41.558 0 42.142 4.08 ;
      RECT 41.008 3.12 41.242 4.08 ;
      RECT 40.658 0 41.242 3.12 ;
      RECT 39.936 2.16 40.342 3.12 ;
      RECT 39.758 0 40.342 2.16 ;
      RECT 38.948 1.2 39.442 2.16 ;
      RECT 38.858 0 39.442 1.2 ;
      RECT 37.958 0 38.542 1.2 ;
      RECT 36.158 0 36.742 0.24 ;
    LAYER m0 ;
      RECT 0 0.002 81 22.078 ;
    LAYER m1 ;
      RECT 0 0 81 22.08 ;
    LAYER m2 ;
      RECT 0 0.015 81 22.065 ;
    LAYER m3 ;
      RECT 0.015 0 80.985 22.08 ;
    LAYER m4 ;
      RECT 0 0.02 81 22.06 ;
    LAYER m5 ;
      RECT 0.012 0 80.988 22.08 ;
    LAYER m6 ;
      RECT 0 0.012 81 22.068 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf028b256e2r2w0cbbeheaa4acw

END LIBRARY
