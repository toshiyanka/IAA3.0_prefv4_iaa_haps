//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr_b : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr_b
(
  // Synchronous Clock/Reset
  clk_100,
  rst_b_100,

  // Asynchronous Clock/Reset(s)
  clk_200,

  // Power Well Isolation Input Signals
  island0_pok,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  p3_fab_init_idle_exit,
  p3_fab_init_idle_exit_ack,
  p4_fab_init_idle_exit,
  p4_fab_init_idle_exit_ack,
  p5_fab_init_idle_exit,
  p5_fab_init_idle_exit_ack,
  p6_fab_init_idle_exit,
  p6_fab_init_idle_exit_ack,
  p7_fab_init_idle_exit,
  p7_fab_init_idle_exit_ack,
  p8_fab_init_idle_exit,
  p8_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_clk_100,
  visa_vp_clk_100,
  visa_p0_tier1_clk_100,
  visa_p0_tier2_clk_100,
  visa_p1_tier1_clk_100,
  visa_p1_tier2_clk_100,
  visa_p2_tier1_clk_100,
  visa_p2_tier2_clk_100,
  visa_p3_tier1_clk_100,
  visa_p3_tier2_clk_100,
  visa_p4_tier1_clk_100,
  visa_p4_tier2_clk_100,
  visa_p5_tier1_clk_100,
  visa_p5_tier2_clk_100,
  visa_p6_tier1_clk_200,
  visa_p6_tier2_clk_200,
  visa_p6_ififo_tier1_clk_100,
  visa_p6_ififo_tier2_clk_100,
  visa_p6_efifo_tier1_clk_100,
  visa_p6_efifo_tier2_clk_100,
  visa_p7_tier1_clk_100,
  visa_p7_tier2_clk_100,
  visa_p8_tier1_clk_200,
  visa_p8_tier2_clk_200,
  visa_p8_ififo_tier1_clk_100,
  visa_p8_ififo_tier2_clk_100,
  visa_p8_efifo_tier1_clk_100,
  visa_p8_efifo_tier2_clk_100,


  // Register wires
  cfg_sbr_b_cgovrd,
  cfg_sbr_b_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  sbr_a_sbr_b_side_ism_agent,
  sbr_b_sbr_a_side_ism_fabric,
  sbr_a_sbr_b_pccup,
  sbr_a_sbr_b_npcup,
  sbr_b_sbr_a_pcput,
  sbr_b_sbr_a_npput,
  sbr_b_sbr_a_eom,
  sbr_b_sbr_a_payload,
  sbr_b_sbr_a_pccup,
  sbr_b_sbr_a_npcup,
  sbr_a_sbr_b_pcput,
  sbr_a_sbr_b_npput,
  sbr_a_sbr_b_eom,
  sbr_a_sbr_b_payload,

  // Port 1 declarations
  pcie_afe_sbr_b_side_ism_agent,
  sbr_b_pcie_afe_side_ism_fabric,
  pcie_afe_sbr_b_pccup,
  pcie_afe_sbr_b_npcup,
  sbr_b_pcie_afe_pcput,
  sbr_b_pcie_afe_npput,
  sbr_b_pcie_afe_eom,
  sbr_b_pcie_afe_payload,
  sbr_b_pcie_afe_pccup,
  sbr_b_pcie_afe_npcup,
  pcie_afe_sbr_b_pcput,
  pcie_afe_sbr_b_npput,
  pcie_afe_sbr_b_eom,
  pcie_afe_sbr_b_payload,

  // Port 2 declarations
  sata_afe_sbr_b_side_ism_agent,
  sbr_b_sata_afe_side_ism_fabric,
  sata_afe_sbr_b_pccup,
  sata_afe_sbr_b_npcup,
  sbr_b_sata_afe_pcput,
  sbr_b_sata_afe_npput,
  sbr_b_sata_afe_eom,
  sbr_b_sata_afe_payload,
  sbr_b_sata_afe_pccup,
  sbr_b_sata_afe_npcup,
  sata_afe_sbr_b_pcput,
  sata_afe_sbr_b_npput,
  sata_afe_sbr_b_eom,
  sata_afe_sbr_b_payload,

  // Port 3 declarations
  usb_afe_sbr_b_side_ism_agent,
  sbr_b_usb_afe_side_ism_fabric,
  usb_afe_sbr_b_pccup,
  usb_afe_sbr_b_npcup,
  sbr_b_usb_afe_pcput,
  sbr_b_usb_afe_npput,
  sbr_b_usb_afe_eom,
  sbr_b_usb_afe_payload,
  sbr_b_usb_afe_pccup,
  sbr_b_usb_afe_npcup,
  usb_afe_sbr_b_pcput,
  usb_afe_sbr_b_npput,
  usb_afe_sbr_b_eom,
  usb_afe_sbr_b_payload,

  // Port 4 declarations
  sata_ctrl_sbr_b_side_ism_agent,
  sbr_b_sata_ctrl_side_ism_fabric,
  sata_ctrl_sbr_b_pccup,
  sata_ctrl_sbr_b_npcup,
  sbr_b_sata_ctrl_pcput,
  sbr_b_sata_ctrl_npput,
  sbr_b_sata_ctrl_eom,
  sbr_b_sata_ctrl_payload,
  sbr_b_sata_ctrl_pccup,
  sbr_b_sata_ctrl_npcup,
  sata_ctrl_sbr_b_pcput,
  sata_ctrl_sbr_b_npput,
  sata_ctrl_sbr_b_eom,
  sata_ctrl_sbr_b_payload,

  // Port 5 declarations
  pcie_ctrl_sbr_b_side_ism_agent,
  sbr_b_pcie_ctrl_side_ism_fabric,
  pcie_ctrl_sbr_b_pccup,
  pcie_ctrl_sbr_b_npcup,
  sbr_b_pcie_ctrl_pcput,
  sbr_b_pcie_ctrl_npput,
  sbr_b_pcie_ctrl_eom,
  sbr_b_pcie_ctrl_payload,
  sbr_b_pcie_ctrl_pccup,
  sbr_b_pcie_ctrl_npcup,
  pcie_ctrl_sbr_b_pcput,
  pcie_ctrl_sbr_b_npput,
  pcie_ctrl_sbr_b_eom,
  pcie_ctrl_sbr_b_payload,

  // Port 6 declarations
  psf_1_sbr_b_side_ism_agent,
  sbr_b_psf_1_side_ism_fabric,
  psf_1_sbr_b_pccup,
  psf_1_sbr_b_npcup,
  sbr_b_psf_1_pcput,
  sbr_b_psf_1_npput,
  sbr_b_psf_1_eom,
  sbr_b_psf_1_payload,
  sbr_b_psf_1_pccup,
  sbr_b_psf_1_npcup,
  psf_1_sbr_b_pcput,
  psf_1_sbr_b_npput,
  psf_1_sbr_b_eom,
  psf_1_sbr_b_payload,

  // Port 7 declarations
  psf_0_south_sbr_b_side_ism_agent,
  sbr_b_psf_0_south_side_ism_fabric,
  psf_0_south_sbr_b_pccup,
  psf_0_south_sbr_b_npcup,
  sbr_b_psf_0_south_pcput,
  sbr_b_psf_0_south_npput,
  sbr_b_psf_0_south_eom,
  sbr_b_psf_0_south_payload,
  sbr_b_psf_0_south_pccup,
  sbr_b_psf_0_south_npcup,
  psf_0_south_sbr_b_pcput,
  psf_0_south_sbr_b_npput,
  psf_0_south_sbr_b_eom,
  psf_0_south_sbr_b_payload,

  // Port 8 declarations
  psf_0_north_sbr_b_side_ism_agent,
  sbr_b_psf_0_north_side_ism_fabric,
  psf_0_north_sbr_b_pccup,
  psf_0_north_sbr_b_npcup,
  sbr_b_psf_0_north_pcput,
  sbr_b_psf_0_north_npput,
  sbr_b_psf_0_north_eom,
  sbr_b_psf_0_north_payload,
  sbr_b_psf_0_north_pccup,
  sbr_b_psf_0_north_npcup,
  psf_0_north_sbr_b_pcput,
  psf_0_north_sbr_b_npput,
  psf_0_north_sbr_b_eom,
  psf_0_north_sbr_b_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic clk_100;
  input logic rst_b_100;

  // Asynchronous Clock/Reset(s)
  input logic clk_200;

  // Power Well Isolation Input Signals
  input logic island0_pok;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic p3_fab_init_idle_exit;
  input logic p3_fab_init_idle_exit_ack;
  output logic p4_fab_init_idle_exit;
  input logic p4_fab_init_idle_exit_ack;
  output logic p5_fab_init_idle_exit;
  input logic p5_fab_init_idle_exit_ack;
  output logic p6_fab_init_idle_exit;
  input logic p6_fab_init_idle_exit_ack;
  output logic p7_fab_init_idle_exit;
  input logic p7_fab_init_idle_exit_ack;
  output logic p8_fab_init_idle_exit;
  input logic p8_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_clk_100;
  output visa_vp  visa_vp_clk_100;
  output visa_port_tier1 visa_p0_tier1_clk_100;
  output visa_port_tier2 visa_p0_tier2_clk_100;
  output visa_port_tier1 visa_p1_tier1_clk_100;
  output visa_port_tier2 visa_p1_tier2_clk_100;
  output visa_port_tier1 visa_p2_tier1_clk_100;
  output visa_port_tier2 visa_p2_tier2_clk_100;
  output visa_port_tier1 visa_p3_tier1_clk_100;
  output visa_port_tier2 visa_p3_tier2_clk_100;
  output visa_port_tier1 visa_p4_tier1_clk_100;
  output visa_port_tier2 visa_p4_tier2_clk_100;
  output visa_port_tier1 visa_p5_tier1_clk_100;
  output visa_port_tier2 visa_p5_tier2_clk_100;
  output visa_port_tier1 visa_p6_tier1_clk_200;
  output visa_port_tier2 visa_p6_tier2_clk_200;
  output visa_ififo_tier1 visa_p6_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p6_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p6_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p6_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p7_tier1_clk_100;
  output visa_port_tier2 visa_p7_tier2_clk_100;
  output visa_port_tier1 visa_p8_tier1_clk_200;
  output visa_port_tier2 visa_p8_tier2_clk_200;
  output visa_ififo_tier1 visa_p8_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p8_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p8_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p8_efifo_tier2_clk_100;

  // Register wires
  input logic [4:0]  cfg_sbr_b_cgovrd;
  input logic [15:0] cfg_sbr_b_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic fscan_rstbypen;
  input logic fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] sbr_a_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_sbr_a_side_ism_fabric;
  input logic sbr_a_sbr_b_pccup;
  input logic sbr_a_sbr_b_npcup;
  output logic sbr_b_sbr_a_pcput;
  output logic sbr_b_sbr_a_npput;
  output logic sbr_b_sbr_a_eom;
  output logic [7:0] sbr_b_sbr_a_payload;
  output logic sbr_b_sbr_a_pccup;
  output logic sbr_b_sbr_a_npcup;
  input logic sbr_a_sbr_b_pcput;
  input logic sbr_a_sbr_b_npput;
  input logic sbr_a_sbr_b_eom;
  input logic [7:0] sbr_a_sbr_b_payload;

  // Port 1 declarations
  input logic [2:0] pcie_afe_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_pcie_afe_side_ism_fabric;
  input logic pcie_afe_sbr_b_pccup;
  input logic pcie_afe_sbr_b_npcup;
  output logic sbr_b_pcie_afe_pcput;
  output logic sbr_b_pcie_afe_npput;
  output logic sbr_b_pcie_afe_eom;
  output logic [7:0] sbr_b_pcie_afe_payload;
  output logic sbr_b_pcie_afe_pccup;
  output logic sbr_b_pcie_afe_npcup;
  input logic pcie_afe_sbr_b_pcput;
  input logic pcie_afe_sbr_b_npput;
  input logic pcie_afe_sbr_b_eom;
  input logic [7:0] pcie_afe_sbr_b_payload;

  // Port 2 declarations
  input logic [2:0] sata_afe_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_sata_afe_side_ism_fabric;
  input logic sata_afe_sbr_b_pccup;
  input logic sata_afe_sbr_b_npcup;
  output logic sbr_b_sata_afe_pcput;
  output logic sbr_b_sata_afe_npput;
  output logic sbr_b_sata_afe_eom;
  output logic [7:0] sbr_b_sata_afe_payload;
  output logic sbr_b_sata_afe_pccup;
  output logic sbr_b_sata_afe_npcup;
  input logic sata_afe_sbr_b_pcput;
  input logic sata_afe_sbr_b_npput;
  input logic sata_afe_sbr_b_eom;
  input logic [7:0] sata_afe_sbr_b_payload;

  // Port 3 declarations
  input logic [2:0] usb_afe_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_usb_afe_side_ism_fabric;
  input logic usb_afe_sbr_b_pccup;
  input logic usb_afe_sbr_b_npcup;
  output logic sbr_b_usb_afe_pcput;
  output logic sbr_b_usb_afe_npput;
  output logic sbr_b_usb_afe_eom;
  output logic [7:0] sbr_b_usb_afe_payload;
  output logic sbr_b_usb_afe_pccup;
  output logic sbr_b_usb_afe_npcup;
  input logic usb_afe_sbr_b_pcput;
  input logic usb_afe_sbr_b_npput;
  input logic usb_afe_sbr_b_eom;
  input logic [7:0] usb_afe_sbr_b_payload;

  // Port 4 declarations
  input logic [2:0] sata_ctrl_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_sata_ctrl_side_ism_fabric;
  input logic sata_ctrl_sbr_b_pccup;
  input logic sata_ctrl_sbr_b_npcup;
  output logic sbr_b_sata_ctrl_pcput;
  output logic sbr_b_sata_ctrl_npput;
  output logic sbr_b_sata_ctrl_eom;
  output logic [7:0] sbr_b_sata_ctrl_payload;
  output logic sbr_b_sata_ctrl_pccup;
  output logic sbr_b_sata_ctrl_npcup;
  input logic sata_ctrl_sbr_b_pcput;
  input logic sata_ctrl_sbr_b_npput;
  input logic sata_ctrl_sbr_b_eom;
  input logic [7:0] sata_ctrl_sbr_b_payload;

  // Port 5 declarations
  input logic [2:0] pcie_ctrl_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_pcie_ctrl_side_ism_fabric;
  input logic pcie_ctrl_sbr_b_pccup;
  input logic pcie_ctrl_sbr_b_npcup;
  output logic sbr_b_pcie_ctrl_pcput;
  output logic sbr_b_pcie_ctrl_npput;
  output logic sbr_b_pcie_ctrl_eom;
  output logic [7:0] sbr_b_pcie_ctrl_payload;
  output logic sbr_b_pcie_ctrl_pccup;
  output logic sbr_b_pcie_ctrl_npcup;
  input logic pcie_ctrl_sbr_b_pcput;
  input logic pcie_ctrl_sbr_b_npput;
  input logic pcie_ctrl_sbr_b_eom;
  input logic [7:0] pcie_ctrl_sbr_b_payload;

  // Port 6 declarations
  input logic [2:0] psf_1_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_psf_1_side_ism_fabric;
  input logic psf_1_sbr_b_pccup;
  input logic psf_1_sbr_b_npcup;
  output logic sbr_b_psf_1_pcput;
  output logic sbr_b_psf_1_npput;
  output logic sbr_b_psf_1_eom;
  output logic [7:0] sbr_b_psf_1_payload;
  output logic sbr_b_psf_1_pccup;
  output logic sbr_b_psf_1_npcup;
  input logic psf_1_sbr_b_pcput;
  input logic psf_1_sbr_b_npput;
  input logic psf_1_sbr_b_eom;
  input logic [7:0] psf_1_sbr_b_payload;

  // Port 7 declarations
  input logic [2:0] psf_0_south_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_psf_0_south_side_ism_fabric;
  input logic psf_0_south_sbr_b_pccup;
  input logic psf_0_south_sbr_b_npcup;
  output logic sbr_b_psf_0_south_pcput;
  output logic sbr_b_psf_0_south_npput;
  output logic sbr_b_psf_0_south_eom;
  output logic [7:0] sbr_b_psf_0_south_payload;
  output logic sbr_b_psf_0_south_pccup;
  output logic sbr_b_psf_0_south_npcup;
  input logic psf_0_south_sbr_b_pcput;
  input logic psf_0_south_sbr_b_npput;
  input logic psf_0_south_sbr_b_eom;
  input logic [7:0] psf_0_south_sbr_b_payload;

  // Port 8 declarations
  input logic [2:0] psf_0_north_sbr_b_side_ism_agent;
  output logic [2:0] sbr_b_psf_0_north_side_ism_fabric;
  input logic psf_0_north_sbr_b_pccup;
  input logic psf_0_north_sbr_b_npcup;
  output logic sbr_b_psf_0_north_pcput;
  output logic sbr_b_psf_0_north_npput;
  output logic sbr_b_psf_0_north_eom;
  output logic [7:0] sbr_b_psf_0_north_payload;
  output logic sbr_b_psf_0_north_pccup;
  output logic sbr_b_psf_0_north_npcup;
  input logic psf_0_north_sbr_b_pcput;
  input logic psf_0_north_sbr_b_npput;
  input logic psf_0_north_sbr_b_eom;
  input logic [7:0] psf_0_north_sbr_b_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_b_sbcportmap;
always_comb sbr_b_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr_b (sbr_b)                                 SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  107 { 17'b0_0000_0000_0000_0000 }},   //   254:148      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //   147          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   146          SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //   145          SBCPORTMAPTABLE
               17'b0_0000_0000_1000_0000,      //   144          SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   143:140      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   139:136      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   135:132      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   131:128      SBCPORTMAPTABLE
      {   31 { 17'b0_0000_0000_0000_0000 }},   //   127: 97      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //    96          SBCPORTMAPTABLE
      {    6 { 17'b0_0000_0000_0000_0000 }},   //    95: 90      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //    89          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //    88          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    87: 86      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    85: 84      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0000 }},   //    83: 81      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    80          SBCPORTMAPTABLE
      {   13 { 17'b0_0000_0000_0000_0000 }},   //    79: 67      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //    66: 64      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0000 }},   //    63: 59      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0001 }},   //    58: 54      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //    53          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    52          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //    51          SBCPORTMAPTABLE
               17'b0_0000_0001_0000_0000,      //    50          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    49: 48      SBCPORTMAPTABLE
      {    9 { 17'b0_0000_0000_0000_0000 }},   //    47: 39      SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_0000_0001 }},   //    38: 32      SBCPORTMAPTABLE
      {   14 { 17'b0_0000_0000_0000_0000 }},   //    31: 18      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //    17          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //    16          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    15: 14      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //    13: 10      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //     7          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     6:  5      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0001 }}    //     4:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  8;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;
logic                              p7_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic                              p7_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;
logic                              p7_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              p3_ism_idle;
logic                              p3_cg_inprogress;
logic                              p3_credit_reinit;
logic                              p4_ism_idle;
logic                              p4_cg_inprogress;
logic                              p4_credit_reinit;
logic                              p5_ism_idle;
logic                              p5_cg_inprogress;
logic                              p5_credit_reinit;
logic                              p6_ism_idle;
logic                              p6_cg_inprogress;
logic                              p6_credit_reinit;
logic                              p7_ism_idle;
logic                              p7_cg_inprogress;
logic                              p7_credit_reinit;
logic                              p8_ism_idle;
logic                              p8_cg_inprogress;
logic                              p8_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              island0_pok_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = cfg_sbr_b_cgctrl[15];
always_comb cfg_clkgatedef    = cfg_sbr_b_cgctrl[14];
always_comb cfg_idlecnt       = cfg_sbr_b_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = cfg_sbr_b_cgovrd[3];
always_comb jta_force_idle    = cfg_sbr_b_cgovrd[1];
always_comb jta_force_notidle = cfg_sbr_b_cgovrd[0];
always_comb jta_force_creditreq = cfg_sbr_b_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

// Asynchronous port signals
logic                              p6_clkgaten;
logic                              p6_clkgatedef;
logic                              p6_clkgate_ovrd;
logic                              p6_force_idle;
logic                              p6_force_notidle;
logic                              p6_force_creditreq;
logic                              p6_clken;
logic                              p6_gated_clk;
logic                              p6_agent_idle;
logic                              p6_eagent_idle;
logic                              p6_port_idle;
logic                              p6_ififo_idle;
logic                              p6_efifo_idle;
logic                              p6_pctrdy;
logic                              p6_pcirdy;
logic             [INTMAXPLDBIT:0] p6_pcdata;
logic                              p6_pceom;
logic                              p6_nptrdy;
logic                              p6_npirdy;
logic                              p6_npfence;
logic             [INTMAXPLDBIT:0] p6_npdata;
logic                              p6_npeom;
logic                              p6_enpstall;
logic                              p6_epctrdy;
logic                              p6_enptrdy;
logic                              p6_epcirdy;
logic                              p6_enpirdy;
logic                              p6_eom;
logic             [INTMAXPLDBIT:0] p6_data;

logic                              p8_clkgaten;
logic                              p8_clkgatedef;
logic                              p8_clkgate_ovrd;
logic                              p8_force_idle;
logic                              p8_force_notidle;
logic                              p8_force_creditreq;
logic                              p8_clken;
logic                              p8_gated_clk;
logic                              p8_agent_idle;
logic                              p8_eagent_idle;
logic                              p8_port_idle;
logic                              p8_ififo_idle;
logic                              p8_efifo_idle;
logic                              p8_pctrdy;
logic                              p8_pcirdy;
logic             [INTMAXPLDBIT:0] p8_pcdata;
logic                              p8_pceom;
logic                              p8_nptrdy;
logic                              p8_npirdy;
logic                              p8_npfence;
logic             [INTMAXPLDBIT:0] p8_npdata;
logic                              p8_npeom;
logic                              p8_enpstall;
logic                              p8_epctrdy;
logic                              p8_enptrdy;
logic                              p8_epcirdy;
logic                              p8_enpirdy;
logic                              p8_eom;
logic             [INTMAXPLDBIT:0] p8_data;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_b_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_b_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// Async clock reset synchronization
//
//------------------------------------------------------------------------------
logic clk_200_rst_b, clk_200_rst_b_pre;
sbc_doublesync sync_rst_clk_200 (
  .d     ( 1'b1 ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_200 ),
  .q     ( clk_200_rst_b_pre ));

always_comb clk_200_rst_b = fscan_rstbypen ? fscan_byprst_b : clk_200_rst_b_pre;


//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_creditreq               )
);

sbc_doublesync sync_p8_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_force_idle                 )
);

sbc_doublesync sync_p8_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_force_notidle              )
);

sbc_doublesync sync_p8_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_force_creditreq            )
);

sbc_doublesync sync_p6_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_force_idle                 )
);

sbc_doublesync sync_p6_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_force_notidle              )
);

sbc_doublesync sync_p6_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_force_creditreq            )
);

//------------------------------------------------------------------------------
//
// Asynchronous port local clock gating
//
//------------------------------------------------------------------------------
// Port 8
sbc_doublesync sync_p8_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_clkgaten                   )
);

sbc_doublesync sync_p8_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_clkgatedef                 )
);

sbc_doublesync sync_p8_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p8_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p8_clken <= '1;
  else
    p8_clken <= ~p8_clkgate_ovrd &
      (p8_clkgatedef | ~p8_clkgaten | ~p8_cg_inprogress |
       ((psf_0_north_sbr_b_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_b_psf_0_north_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (psf_0_north_sbr_b_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((psf_0_north_sbr_b_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_b_psf_0_north_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p8_clkgate  (
  .en                  ( p8_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p8_gated_clk                  )
);

// Port 6
sbc_doublesync sync_p6_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_clkgaten                   )
);

sbc_doublesync sync_p6_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_clkgatedef                 )
);

sbc_doublesync sync_p6_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p6_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p6_clken <= '1;
  else
    p6_clken <= ~p6_clkgate_ovrd &
      (p6_clkgatedef | ~p6_clkgaten | ~p6_cg_inprogress |
       ((psf_1_sbr_b_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_b_psf_1_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (psf_1_sbr_b_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((psf_1_sbr_b_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_b_psf_1_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p6_clkgate  (
  .en                  ( p6_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p6_gated_clk                  )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_island0_pok (
  .d                   ( island0_pok                   ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( island0_pok_ff2               )
);


always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          island0_pok_ff2
                        };

logic p0_gated_clk;
sbc_clock_gate p0_pwr_clkgate  (
  .en ( endpoint_pwrgd[0] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p0_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  p8_efifo_idle
                  &  (p7_ism_idle | ~endpoint_pwrgd[7])
                  &  p6_efifo_idle
                  &  (p5_ism_idle | ~endpoint_pwrgd[5])
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
logic p6_ism_idle_ff2, p6_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p6_ism_idle_pre <= '1;
  else
    p6_ism_idle_pre <= p6_ism_idle;

sbc_doublesync sync_idle_p6 (
  .d ( p6_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p6_ism_idle_ff2 ));

logic p8_ism_idle_ff2, p8_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p8_ism_idle_pre <= '1;
  else
    p8_ism_idle_pre <= p8_ism_idle;

sbc_doublesync sync_idle_p8 (
  .d ( p8_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p8_ism_idle_ff2 ));

// SBR_IDLE signal for PMU
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle &
                  p2_ism_idle &
                  p3_ism_idle &
                  p4_ism_idle &
                  p5_ism_idle &
                  p6_ism_idle_ff2 &
                  p7_ism_idle &
                  p8_ism_idle_ff2;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 1'b0,
                 p7_npfence,
                 1'b0,
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 pcirdy[8],
                 p7_pcdstvld,
                 pcirdy[6],
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 npirdy[8],
                 p7_npdstvld,
                 npirdy[6],
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_clk_100 = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk_100                       ),
  .side_rst_b          ( rst_b_100                     ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_clk_100 = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle & agent_idle[0] & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle & p0_side_clk_valid )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_clk_100 = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_clk_100 = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( p0_gated_clk                  ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( sbr_a_sbr_b_side_ism_agent    ),
  .side_ism_out        ( sbr_b_sbr_a_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_b_sbr_a_pccup             ),
  .tnpcup              ( sbr_b_sbr_a_npcup             ),
  .tpcput              ( sbr_a_sbr_b_pcput             ),
  .tnpput              ( sbr_a_sbr_b_npput             ),
  .teom                ( sbr_a_sbr_b_eom               ),
  .tpayload            ( sbr_a_sbr_b_payload           ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( sbr_a_sbr_b_pccup             ),
  .mnpcup              ( sbr_a_sbr_b_npcup             ),
  .mpcput              ( sbr_b_sbr_a_pcput             ),
  .mnpput              ( sbr_b_sbr_a_npput             ),
  .meom                ( sbr_b_sbr_a_eom               ),
  .mpayload            ( sbr_b_sbr_a_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit & p1_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle & (~agent_idle[1] || ~p1_idle_egress) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle & agent_idle[1] & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle & p1_side_clk_valid )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle )
          p1_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

  always_comb
    begin
      visa_p1_tier1_clk_100 = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_clk_100 = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( pcie_afe_sbr_b_side_ism_agent ),
  .side_ism_out        ( sbr_b_pcie_afe_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .idle_egress         ( p1_idle_egress                ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_b_pcie_afe_pccup          ),
  .tnpcup              ( sbr_b_pcie_afe_npcup          ),
  .tpcput              ( pcie_afe_sbr_b_pcput          ),
  .tnpput              ( pcie_afe_sbr_b_npput          ),
  .teom                ( pcie_afe_sbr_b_eom            ),
  .tpayload            ( pcie_afe_sbr_b_payload        ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( pcie_afe_sbr_b_pccup          ),
  .mnpcup              ( pcie_afe_sbr_b_npcup          ),
  .mpcput              ( sbr_b_pcie_afe_pcput          ),
  .mnpput              ( sbr_b_pcie_afe_npput          ),
  .meom                ( sbr_b_pcie_afe_eom            ),
  .mpayload            ( sbr_b_pcie_afe_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

// Port 2
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit & p2_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle & (~agent_idle[2] || ~p2_idle_egress) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle & agent_idle[2] & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle & p2_side_clk_valid )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle )
          p2_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

  always_comb
    begin
      visa_p2_tier1_clk_100 = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_clk_100 = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( sata_afe_sbr_b_side_ism_agent ),
  .side_ism_out        ( sbr_b_sata_afe_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .idle_egress         ( p2_idle_egress                ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_b_sata_afe_pccup          ),
  .tnpcup              ( sbr_b_sata_afe_npcup          ),
  .tpcput              ( sata_afe_sbr_b_pcput          ),
  .tnpput              ( sata_afe_sbr_b_npput          ),
  .teom                ( sata_afe_sbr_b_eom            ),
  .tpayload            ( sata_afe_sbr_b_payload        ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( sata_afe_sbr_b_pccup          ),
  .mnpcup              ( sata_afe_sbr_b_npcup          ),
  .mpcput              ( sbr_b_sata_afe_pcput          ),
  .mnpput              ( sbr_b_sata_afe_npput          ),
  .meom                ( sbr_b_sata_afe_eom            ),
  .mpayload            ( sbr_b_sata_afe_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

// Port 3
logic p3_side_clk_valid, p3_idle_egress, p3_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_rst_suppress <= 1'b1;
    else
      p3_rst_suppress <= p3_credit_reinit & p3_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p3_fab_init_idle_exit <= '1;
    else
      if ( ~p3_rst_suppress & (p3_ism_idle & (~agent_idle[3] || ~p3_idle_egress) & ~p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '1;
      else if ( ~p3_rst_suppress & (p3_ism_idle & agent_idle[3] & p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( p3_ism_idle & p3_side_clk_valid )
          p3_side_clk_valid <= '0;
        else if ( (p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack) || ~p3_ism_idle )
          p3_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

  always_comb
    begin
      visa_p3_tier1_clk_100 = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_clk_100 = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( usb_afe_sbr_b_side_ism_agent  ),
  .side_ism_out        ( sbr_b_usb_afe_side_ism_fabric ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .idle_egress         ( p3_idle_egress                ),
  .ism_idle            ( p3_ism_idle                   ),
  .credit_reinit       ( p3_credit_reinit              ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_b_usb_afe_pccup           ),
  .tnpcup              ( sbr_b_usb_afe_npcup           ),
  .tpcput              ( usb_afe_sbr_b_pcput           ),
  .tnpput              ( usb_afe_sbr_b_npput           ),
  .teom                ( usb_afe_sbr_b_eom             ),
  .tpayload            ( usb_afe_sbr_b_payload         ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( usb_afe_sbr_b_pccup           ),
  .mnpcup              ( usb_afe_sbr_b_npcup           ),
  .mpcput              ( sbr_b_usb_afe_pcput           ),
  .mnpput              ( sbr_b_usb_afe_npput           ),
  .meom                ( sbr_b_usb_afe_eom             ),
  .mpayload            ( sbr_b_usb_afe_payload         ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
logic p4_side_clk_valid, p4_idle_egress, p4_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_rst_suppress <= 1'b1;
    else
      p4_rst_suppress <= p4_credit_reinit & p4_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p4_fab_init_idle_exit <= '1;
    else
      if ( ~p4_rst_suppress & (p4_ism_idle & (~agent_idle[4] || ~p4_idle_egress) & ~p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '1;
      else if ( ~p4_rst_suppress & (p4_ism_idle & agent_idle[4] & p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( p4_ism_idle & p4_side_clk_valid )
          p4_side_clk_valid <= '0;
        else if ( (p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack) || ~p4_ism_idle )
          p4_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

  always_comb
    begin
      visa_p4_tier1_clk_100 = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_clk_100 = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( sata_ctrl_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_sata_ctrl_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .idle_egress         ( p4_idle_egress                ),
  .ism_idle            ( p4_ism_idle                   ),
  .credit_reinit       ( p4_credit_reinit              ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_b_sata_ctrl_pccup         ),
  .tnpcup              ( sbr_b_sata_ctrl_npcup         ),
  .tpcput              ( sata_ctrl_sbr_b_pcput         ),
  .tnpput              ( sata_ctrl_sbr_b_npput         ),
  .teom                ( sata_ctrl_sbr_b_eom           ),
  .tpayload            ( sata_ctrl_sbr_b_payload       ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( sata_ctrl_sbr_b_pccup         ),
  .mnpcup              ( sata_ctrl_sbr_b_npcup         ),
  .mpcput              ( sbr_b_sata_ctrl_pcput         ),
  .mnpput              ( sbr_b_sata_ctrl_npput         ),
  .meom                ( sbr_b_sata_ctrl_eom           ),
  .mpayload            ( sbr_b_sata_ctrl_payload       ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

// Port 5
logic p5_side_clk_valid, p5_idle_egress, p5_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p5_rst_suppress <= 1'b1;
    else
      p5_rst_suppress <= p5_credit_reinit & p5_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p5_fab_init_idle_exit <= '1;
    else
      if ( ~p5_rst_suppress & (p5_ism_idle & (~agent_idle[5] || ~p5_idle_egress) & ~p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '1;
      else if ( ~p5_rst_suppress & (p5_ism_idle & agent_idle[5] & p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p5_side_clk_valid <= 1'b0;
    else
      begin
        if ( p5_ism_idle & p5_side_clk_valid )
          p5_side_clk_valid <= '0;
        else if ( (p5_fab_init_idle_exit & p5_fab_init_idle_exit_ack) || ~p5_ism_idle )
          p5_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p5_dbgbus;

  always_comb
    begin
      visa_p5_tier1_clk_100 = { p5_dbgbus[31],
                            p5_dbgbus[27:24],
                            p5_dbgbus[21:19],
                            p5_dbgbus[15:12],
                            p5_dbgbus[7:4] };
      visa_p5_tier2_clk_100 = { p5_dbgbus[30:28],
                            p5_dbgbus[23:22],
                            p5_dbgbus[18:16],
                            p5_dbgbus[11:8],
                            p5_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport5 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( pcie_ctrl_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_pcie_ctrl_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[5] ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .idle_egress         ( p5_idle_egress                ),
  .ism_idle            ( p5_ism_idle                   ),
  .credit_reinit       ( p5_credit_reinit              ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr_b_pcie_ctrl_pccup         ),
  .tnpcup              ( sbr_b_pcie_ctrl_npcup         ),
  .tpcput              ( pcie_ctrl_sbr_b_pcput         ),
  .tnpput              ( pcie_ctrl_sbr_b_npput         ),
  .teom                ( pcie_ctrl_sbr_b_eom           ),
  .tpayload            ( pcie_ctrl_sbr_b_payload       ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( pcie_ctrl_sbr_b_pccup         ),
  .mnpcup              ( pcie_ctrl_sbr_b_npcup         ),
  .mpcput              ( sbr_b_pcie_ctrl_pcput         ),
  .mnpput              ( sbr_b_pcie_ctrl_npput         ),
  .meom                ( sbr_b_pcie_ctrl_eom           ),
  .mpayload            ( sbr_b_pcie_ctrl_payload       ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p5_dbgbus                     )
);

// Port 6 (Asynchronous port)
logic p6_side_clk_valid, p6_idle_egress, p6_rst_suppress;
  logic p6_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p6_rst_suppress <= 1'b1;
    else
      p6_rst_suppress <= p6_credit_reinit_ff2 & p6_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p6_fab_init_idle_exit <= '1;
    else
      if ( ~p6_rst_suppress & (p6_ism_idle_ff2 & (~agent_idle[6] || ~p6_efifo_idle) & ~p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '1;
      else if ( ~p6_rst_suppress & (p6_ism_idle_ff2 & agent_idle[6] & p6_efifo_idle & p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p6_side_clk_valid <= 1'b0;
    else
      begin
        if ( p6_ism_idle_ff2 & p6_side_clk_valid & ~p6_fab_init_idle_exit )
          p6_side_clk_valid <= '0;
        else if ( (p6_fab_init_idle_exit & p6_fab_init_idle_exit_ack) || ~p6_ism_idle_ff2 )
          p6_side_clk_valid <= '1;
      end

logic p6_side_clk_valid_ff2;
sbc_doublesync sync_p6_clk_valid (
  .d     ( p6_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p6_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p6_credit_reinit (
  .d     ( p6_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p6_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p6_dbgbus;

logic [15:0] p6_dbgbus_ing;
logic [15:0] p6_dbgbus_egr;
  always_comb
    begin
      visa_p6_tier1_clk_200 = { p6_dbgbus[31],
                            p6_dbgbus[27:24],
                            p6_dbgbus[21:19],
                            p6_dbgbus[15:12],
                            p6_dbgbus[7:4] };
      visa_p6_tier2_clk_200 = { p6_dbgbus[30:28],
                            p6_dbgbus[23:22],
                            p6_dbgbus[18:16],
                            p6_dbgbus[11:8],
                            p6_dbgbus[3:0] };
      visa_p6_ififo_tier1_clk_100 = { p6_dbgbus_ing[15:14],
                             p6_dbgbus_ing[5:0]};
      visa_p6_ififo_tier2_clk_100 = { p6_dbgbus_ing[13:6] };
      visa_p6_efifo_tier1_clk_100 = { p6_dbgbus_egr[7:0] };
      visa_p6_efifo_tier2_clk_100 = { p6_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport6 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p6_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p6_side_clk_valid_ff2         ),
  .side_ism_in         ( psf_1_sbr_b_side_ism_agent    ),
  .side_ism_out        ( sbr_b_psf_1_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[6] ),
  .agent_idle          ( p6_agent_idle                 ),
  .port_idle           ( p6_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p6_ism_idle                   ),
  .credit_reinit       ( p6_credit_reinit              ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr_b_psf_1_pccup             ),
  .tnpcup              ( sbr_b_psf_1_npcup             ),
  .tpcput              ( psf_1_sbr_b_pcput             ),
  .tnpput              ( psf_1_sbr_b_npput             ),
  .teom                ( psf_1_sbr_b_eom               ),
  .tpayload            ( psf_1_sbr_b_payload           ),
  .pctrdy              ( p6_pctrdy                     ),
  .pcirdy              ( p6_pcirdy                     ),
  .pcdata              ( p6_pcdata                     ),
  .pceom               ( p6_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p6_nptrdy                     ),
  .npirdy              ( p6_npirdy                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( p6_npdata                     ),
  .npeom               ( p6_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( psf_1_sbr_b_pccup             ),
  .mnpcup              ( psf_1_sbr_b_npcup             ),
  .mpcput              ( sbr_b_psf_1_pcput             ),
  .mnpput              ( sbr_b_psf_1_npput             ),
  .meom                ( sbr_b_psf_1_eom               ),
  .mpayload            ( sbr_b_psf_1_payload           ),
  .enpstall            ( p6_enpstall                   ),
  .epctrdy             ( p6_epctrdy                    ),
  .enptrdy             ( p6_enptrdy                    ),
  .epcirdy             ( p6_epcirdy                    ),
  .enpirdy             ( p6_enpirdy                    ),
  .data                ( p6_data                       ),
  .eom                 ( p6_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p6_clkgaten                   ),
  .force_idle          ( p6_force_idle                 ),
  .force_notidle       ( p6_force_notidle              ),
  .force_creditreq     ( p6_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p6_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress6 (
  .ing_side_clk        ( p6_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p6_port_idle                  ),
  .pcirdy              ( p6_pcirdy                     ),
  .npirdy              ( p6_npirdy                     ),
  .npfence             ( p6_npfence                    ),
  .pceom               ( p6_pceom                      ),
  .pcdata              ( p6_pcdata                     ),
  .npeom               ( p6_npeom                      ),
  .npdata              ( p6_npdata                     ),
  .pctrdy              ( p6_pctrdy                     ),
  .nptrdy              ( p6_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p6_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[6]                     ),
  .enptrdy             ( nptrdy[6]                     ),
  .epcirdy             ( pcirdy[6]                     ),
  .enpirdy             ( npirdy[6]                     ),
  .eom                 ( npeom[6]                      ),
  .data                ( npdata[6]                     ),
  .opceom              ( pceom[6]                      ),
  .opcdata             ( pcdata[6]                     ),
  .agent_idle          ( port_idle[6]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p6_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress6 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[6]                 ),
  .pcirdy              ( epcirdy[6]                    ),
  .npirdy              ( enpirdy[6]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[6]                    ),
  .nptrdy              ( enptrdy[6]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p6_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p6_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p6_enpstall                   ),
  .epctrdy             ( p6_epctrdy                    ),
  .enptrdy             ( p6_enptrdy                    ),
  .epcirdy             ( p6_epcirdy                    ),
  .enpirdy             ( p6_enpirdy                    ),
  .eom                 ( p6_eom                        ),
  .data                ( p6_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p6_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p6_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p6_agent_idle  = p6_eagent_idle & p6_ififo_idle;

// Port 7
logic p7_side_clk_valid, p7_idle_egress, p7_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p7_rst_suppress <= 1'b1;
    else
      p7_rst_suppress <= p7_credit_reinit & p7_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p7_fab_init_idle_exit <= '1;
    else
      if ( ~p7_rst_suppress & (p7_ism_idle & (~agent_idle[7] || ~p7_idle_egress) & ~p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '1;
      else if ( ~p7_rst_suppress & (p7_ism_idle & agent_idle[7] & p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p7_side_clk_valid <= 1'b0;
    else
      begin
        if ( p7_ism_idle & p7_side_clk_valid )
          p7_side_clk_valid <= '0;
        else if ( (p7_fab_init_idle_exit & p7_fab_init_idle_exit_ack) || ~p7_ism_idle )
          p7_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p7_dbgbus;

  always_comb
    begin
      visa_p7_tier1_clk_100 = { p7_dbgbus[31],
                            p7_dbgbus[27:24],
                            p7_dbgbus[21:19],
                            p7_dbgbus[15:12],
                            p7_dbgbus[7:4] };
      visa_p7_tier2_clk_100 = { p7_dbgbus[30:28],
                            p7_dbgbus[23:22],
                            p7_dbgbus[18:16],
                            p7_dbgbus[11:8],
                            p7_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport7 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( psf_0_south_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_psf_0_south_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[7] ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .idle_egress         ( p7_idle_egress                ),
  .ism_idle            ( p7_ism_idle                   ),
  .credit_reinit       ( p7_credit_reinit              ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr_b_psf_0_south_pccup       ),
  .tnpcup              ( sbr_b_psf_0_south_npcup       ),
  .tpcput              ( psf_0_south_sbr_b_pcput       ),
  .tnpput              ( psf_0_south_sbr_b_npput       ),
  .teom                ( psf_0_south_sbr_b_eom         ),
  .tpayload            ( psf_0_south_sbr_b_payload     ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( psf_0_south_sbr_b_pccup       ),
  .mnpcup              ( psf_0_south_sbr_b_npcup       ),
  .mpcput              ( sbr_b_psf_0_south_pcput       ),
  .mnpput              ( sbr_b_psf_0_south_npput       ),
  .meom                ( sbr_b_psf_0_south_eom         ),
  .mpayload            ( sbr_b_psf_0_south_payload     ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p7_dbgbus                     )
);

// Port 8 (Asynchronous port)
logic p8_side_clk_valid, p8_idle_egress, p8_rst_suppress;
  logic p8_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p8_rst_suppress <= 1'b1;
    else
      p8_rst_suppress <= p8_credit_reinit_ff2 & p8_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p8_fab_init_idle_exit <= '1;
    else
      if ( ~p8_rst_suppress & (p8_ism_idle_ff2 & (~agent_idle[8] || ~p8_efifo_idle) & ~p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '1;
      else if ( ~p8_rst_suppress & (p8_ism_idle_ff2 & agent_idle[8] & p8_efifo_idle & p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p8_side_clk_valid <= 1'b0;
    else
      begin
        if ( p8_ism_idle_ff2 & p8_side_clk_valid & ~p8_fab_init_idle_exit )
          p8_side_clk_valid <= '0;
        else if ( (p8_fab_init_idle_exit & p8_fab_init_idle_exit_ack) || ~p8_ism_idle_ff2 )
          p8_side_clk_valid <= '1;
      end

logic p8_side_clk_valid_ff2;
sbc_doublesync sync_p8_clk_valid (
  .d     ( p8_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p8_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p8_credit_reinit (
  .d     ( p8_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p8_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p8_dbgbus;

logic [15:0] p8_dbgbus_ing;
logic [15:0] p8_dbgbus_egr;
  always_comb
    begin
      visa_p8_tier1_clk_200 = { p8_dbgbus[31],
                            p8_dbgbus[27:24],
                            p8_dbgbus[21:19],
                            p8_dbgbus[15:12],
                            p8_dbgbus[7:4] };
      visa_p8_tier2_clk_200 = { p8_dbgbus[30:28],
                            p8_dbgbus[23:22],
                            p8_dbgbus[18:16],
                            p8_dbgbus[11:8],
                            p8_dbgbus[3:0] };
      visa_p8_ififo_tier1_clk_100 = { p8_dbgbus_ing[15:14],
                             p8_dbgbus_ing[5:0]};
      visa_p8_ififo_tier2_clk_100 = { p8_dbgbus_ing[13:6] };
      visa_p8_efifo_tier1_clk_100 = { p8_dbgbus_egr[7:0] };
      visa_p8_efifo_tier2_clk_100 = { p8_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport8 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p8_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p8_side_clk_valid_ff2         ),
  .side_ism_in         ( psf_0_north_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_psf_0_north_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[8] ),
  .agent_idle          ( p8_agent_idle                 ),
  .port_idle           ( p8_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p8_ism_idle                   ),
  .credit_reinit       ( p8_credit_reinit              ),
  .cg_inprogress       ( p8_cg_inprogress              ),
  .tpccup              ( sbr_b_psf_0_north_pccup       ),
  .tnpcup              ( sbr_b_psf_0_north_npcup       ),
  .tpcput              ( psf_0_north_sbr_b_pcput       ),
  .tnpput              ( psf_0_north_sbr_b_npput       ),
  .teom                ( psf_0_north_sbr_b_eom         ),
  .tpayload            ( psf_0_north_sbr_b_payload     ),
  .pctrdy              ( p8_pctrdy                     ),
  .pcirdy              ( p8_pcirdy                     ),
  .pcdata              ( p8_pcdata                     ),
  .pceom               ( p8_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p8_nptrdy                     ),
  .npirdy              ( p8_npirdy                     ),
  .npfence             ( p8_npfence                    ),
  .npdata              ( p8_npdata                     ),
  .npeom               ( p8_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( psf_0_north_sbr_b_pccup       ),
  .mnpcup              ( psf_0_north_sbr_b_npcup       ),
  .mpcput              ( sbr_b_psf_0_north_pcput       ),
  .mnpput              ( sbr_b_psf_0_north_npput       ),
  .meom                ( sbr_b_psf_0_north_eom         ),
  .mpayload            ( sbr_b_psf_0_north_payload     ),
  .enpstall            ( p8_enpstall                   ),
  .epctrdy             ( p8_epctrdy                    ),
  .enptrdy             ( p8_enptrdy                    ),
  .epcirdy             ( p8_epcirdy                    ),
  .enpirdy             ( p8_enpirdy                    ),
  .data                ( p8_data                       ),
  .eom                 ( p8_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p8_clkgaten                   ),
  .force_idle          ( p8_force_idle                 ),
  .force_notidle       ( p8_force_notidle              ),
  .force_creditreq     ( p8_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p8_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress8 (
  .ing_side_clk        ( p8_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p8_port_idle                  ),
  .pcirdy              ( p8_pcirdy                     ),
  .npirdy              ( p8_npirdy                     ),
  .npfence             ( p8_npfence                    ),
  .pceom               ( p8_pceom                      ),
  .pcdata              ( p8_pcdata                     ),
  .npeom               ( p8_npeom                      ),
  .npdata              ( p8_npdata                     ),
  .pctrdy              ( p8_pctrdy                     ),
  .nptrdy              ( p8_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p8_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[8]                     ),
  .enptrdy             ( nptrdy[8]                     ),
  .epcirdy             ( pcirdy[8]                     ),
  .enpirdy             ( npirdy[8]                     ),
  .eom                 ( npeom[8]                      ),
  .data                ( npdata[8]                     ),
  .opceom              ( pceom[8]                      ),
  .opcdata             ( pcdata[8]                     ),
  .agent_idle          ( port_idle[8]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p8_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress8 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[8]                 ),
  .pcirdy              ( epcirdy[8]                    ),
  .npirdy              ( enpirdy[8]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[8]                    ),
  .nptrdy              ( enptrdy[8]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p8_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p8_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p8_enpstall                   ),
  .epctrdy             ( p8_epctrdy                    ),
  .enptrdy             ( p8_enptrdy                    ),
  .epcirdy             ( p8_epcirdy                    ),
  .enpirdy             ( p8_enpirdy                    ),
  .eom                 ( p8_eom                        ),
  .data                ( p8_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p8_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p8_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p8_agent_idle  = p8_eagent_idle & p8_ififo_idle;

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_b_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_b_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk_100 or negedge rst_b_100)

      if (~rst_b_100) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 1, clk_100, rst_b_100, 0, , 5ns
ClockReset, 0, clk_200, rst_b_200, 0, , 2.5ns
ClockReset, 2, clk_27, rst_b_27, 0, , 18.5ns
Endpoint, SAPms,3, 1, 1, 0, 3, 3, 1, 65, 2, 2, 
Endpoint, adac,0, 1, 1, 0, 3, 3, 1, 129, 2, 2, 
Endpoint, apll,0, 1, 2, 0, 3, 3, 1, 139, 2, 2, 
Endpoint, bunit,2, 1, 0, 0, 3, 3, 1, 03, 2, 2, 
Endpoint, cpunit,2, 1, 1, 0, 3, 3, 1, 10, 2, 2, 
Endpoint, cunit,2, 1, 0, 0, 3, 3, 1, 07, 2, 2, 
Endpoint, ddrio,2, 1, 1, 0, 3, 3, 1, 80, 2, 2, 
Endpoint, dfx_jtag,2, 1, 1, 0, 3, 3, 1, 58, 2, 2, 
Endpoint, dfx_lakemore,2, 1, 1, 0, 3, 3, 1, 56, 2, 2, 
Endpoint, dfx_omar,2, 1, 1, 0, 3, 3, 1, 57, 2, 2, 
Endpoint, dpll,0, 1, 2, 0, 3, 3, 1, 138, 2, 2, 
Endpoint, fpll,0, 1, 2, 0, 3, 3, 1, 136, 2, 2, 
Endpoint, hdmi_rx,0, 1, 1, 0, 3, 3, 1, 131, 2, 2, 
Endpoint, hdmi_tx,0, 1, 1, 0, 3, 3, 1, 130, 2, 2, 
Endpoint, hpll,0, 1, 2, 0, 3, 3, 1, 137, 2, 2, 
Endpoint, hunit,2, 1, 0, 0, 3, 3, 1, 02, 2, 2, 
Endpoint, itunit,2, 1, 1, 0, 3, 3, 1, 64, 2, 2, 
Endpoint, itunit2,2, 1, 1, 0, 3, 3, 1, 66, 2, 2, 
Endpoint, legacy,2, 1, 1, 0, 3, 3, 10, 11,12,13,32,33,34,35,36,37,38, 2, 2, 
Endpoint, mcu,2, 1, 0, 0, 3, 3, 1, 01, 2, 2, 
Endpoint, pcie_afe,4, 1, 1, 0, 3, 3, 1, 17, 2, 2, 
Endpoint, pcie_ctrl,4, 1, 1, 0, 3, 3, 1, 16, 2, 2, 
Endpoint, psf_0_north,4, 1, 0, 0, 3, 3, 1, 50, 2, 2, 
Endpoint, psf_0_south,4, 1, 1, 0, 3, 3, 1, 144, 2, 2, 
Endpoint, psf_1,4, 1, 0, 0, 3, 3, 1, 145, 2, 2, 
Endpoint, psf_3,2, 1, 0, 0, 3, 3, 1, 147, 2, 2, 
Endpoint, punit,1, 1, 2, 0, 3, 3, 1, 04, 2, 2, 
Endpoint, reut_0,2, 1, 1, 0, 3, 3, 1, 84, 2, 2, 
Endpoint, reut_1,2, 1, 1, 0, 3, 3, 1, 85, 2, 2, 
Endpoint, sata_afe,4, 1, 1, 0, 3, 3, 1, 89, 2, 2, 
Endpoint, sata_ctrl,4, 1, 1, 0, 3, 3, 1, 88, 2, 2, 
SyncRouter, sbr_a, sbr_a,1, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 2, 8, sbr_e, sbr_b, sbr_c, dpll, apll, hpll, fpll, punit, , , , , , , , , 
RouterAgentPort, sbr_a, 0
RouterAgentPort, sbr_a, 1
RouterAgentPort, sbr_a, 2
RouterRange, sbr_a, 0, 48,49
SyncRouter, sbr_b, sbr_b,4, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 9, sbr_a, pcie_afe, sata_afe, usb_afe, sata_ctrl, pcie_ctrl, psf_1, psf_0_south, psf_0_north, , , , , , , , 
RouterRange, sbr_b, 0, 51,51
SyncRouter, sbr_c, sbr_c,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 15, sbr_a, sbr_d, vtunit, hunit, bunit, cunit, cpunit, legacy, dfx_lakemore, dfx_omar, dfx_jtag, itunit, psf_3, SAPms, itunit2, , 
RouterAgentPort, sbr_c, 1
RouterRange, sbr_c, 0, 52,52
SyncRouter, sbr_d, sbr_d,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_c, mcu, ddrio, reut_0, reut_1, , , , , , , , , , , , 
RouterRange, sbr_d, 0, 54,55
SyncRouter, sbr_e, sbr_e,5, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_a, vdac, adac, hdmi_tx, hdmi_rx, , , , , , , , , , , , 
Endpoint, usb_afe,4, 1, 1, 0, 3, 3, 1, 96, 2, 2, 
Endpoint, vdac,0, 1, 1, 0, 3, 3, 1, 128, 2, 2, 
Endpoint, vtunit,2, 1, 0, 0, 3, 3, 1, 00, 2, 2, 
AsyncPort, sbr_a, 0, 10, 4, 0, 
AsyncPort, sbr_a, 1, 10, 4, 0, 
AsyncPort, sbr_a, 2, 10, 4, 0, 
AsyncPort, sbr_b, 6, 4, 2, 0, 
AsyncPort, sbr_b, 8, 4, 2, 0, 
AsyncPort, sbr_c, 12, 4, 2, 0, 
AsyncPort, sbr_c, 2, 10, 4, 0, 
AsyncPort, sbr_c, 3, 10, 4, 0, 
AsyncPort, sbr_c, 4, 10, 4, 0, 
AsyncPort, sbr_c, 5, 10, 4, 0, 
AsyncPort, sbr_d, 1, 10, 4, 0, 
PowerWell, 0, 
PowerWell, 1, island0_pok
PowerWell, 2, island1_pok
PowerWell, 3, island2_pok
PowerWell, 4, island3_pok
PowerWell, 5, island8_pok
*/
//------------------------------------------------------------------------------
