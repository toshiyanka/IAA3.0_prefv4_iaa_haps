VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf096b256e1r1w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf096b256e1r1w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 43.2 BY 41.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 21.48 23.872 22.68 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 19.56 21.428 20.76 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 21.48 19.116 22.68 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 21.48 19.372 22.68 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 21.48 19.628 22.68 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 21.48 19.716 22.68 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 21.48 19.928 22.68 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 21.48 20.016 22.68 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 21.48 20.272 22.68 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 21.48 20.528 22.68 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 21.48 18.472 22.68 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 21.48 18.728 22.68 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 21.48 18.816 22.68 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 21.48 19.028 22.68 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 19.56 22.416 20.76 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 19.56 22.628 20.76 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 19.56 22.716 20.76 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 19.56 22.972 20.76 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 19.56 23.228 20.76 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 19.56 23.316 20.76 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.484 19.56 23.528 20.76 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 19.56 23.616 20.76 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 19.56 21.516 20.76 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 19.56 21.728 20.76 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 3.84 22.716 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 3.84 22.972 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 4.56 19.116 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 4.56 19.372 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 5.28 20.272 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 5.28 20.528 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 6 20.916 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 6 21.172 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 6.72 21.728 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 6.72 21.816 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 7.44 22.416 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 7.44 22.628 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 8.16 18.472 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 8.16 18.728 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 8.88 19.928 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 8.88 20.016 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 9.6 20.616 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 9.6 20.828 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 10.32 21.428 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 10.32 21.516 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 0.96 19.928 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 11.04 22.072 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 11.04 22.328 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 11.76 22.716 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 11.76 22.972 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 12.48 19.116 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 12.48 19.372 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 13.2 20.272 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 13.2 20.528 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 13.92 20.916 15.12 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 13.92 21.172 15.12 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 0.96 20.016 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 14.64 21.728 15.84 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 14.64 21.816 15.84 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 15.36 22.416 16.56 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 15.36 22.628 16.56 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 16.08 18.472 17.28 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 16.08 18.728 17.28 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 16.8 19.928 18 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 16.8 20.016 18 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 17.52 20.616 18.72 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 17.52 20.828 18.72 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.68 20.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 23.28 22.716 24.48 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 23.28 22.972 24.48 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 24 18.816 25.2 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 24 19.028 25.2 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 24.72 20.272 25.92 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 24.72 20.528 25.92 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 25.44 20.916 26.64 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 25.44 21.172 26.64 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 26.16 21.728 27.36 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 26.16 21.816 27.36 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 1.68 20.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 26.88 22.416 28.08 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 26.88 22.628 28.08 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 27.6 18.472 28.8 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 27.6 18.728 28.8 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 28.32 19.928 29.52 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 28.32 20.016 29.52 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 29.04 20.616 30.24 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 29.04 20.828 30.24 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 29.76 21.428 30.96 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 29.76 21.516 30.96 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 2.4 21.428 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 30.48 22.072 31.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 30.48 22.328 31.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 31.2 22.716 32.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 31.2 22.972 32.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 31.92 19.116 33.12 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 31.92 19.372 33.12 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 32.64 20.272 33.84 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 32.64 20.528 33.84 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 33.36 20.916 34.56 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 33.36 21.172 34.56 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 2.4 21.516 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 34.08 21.728 35.28 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 34.08 21.816 35.28 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 34.8 22.416 36 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 34.8 22.628 36 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 35.52 18.472 36.72 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 35.52 18.728 36.72 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 36.24 19.928 37.44 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 36.24 20.016 37.44 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 36.96 20.616 38.16 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 36.96 20.828 38.16 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 3.12 22.072 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 37.68 21.428 38.88 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 37.68 21.516 38.88 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 38.4 22.072 39.6 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 38.4 22.328 39.6 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 39.12 22.716 40.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 39.12 22.972 40.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 39.84 19.116 41.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 39.84 19.372 41.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 3.12 22.328 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 19.56 22.072 20.76 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 19.56 22.328 20.76 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 19.56 21.816 20.76 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 3.84 18.472 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 3.84 18.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 4.56 19.628 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 4.56 19.716 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 5.28 20.616 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 5.28 20.828 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 6 21.428 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 6 21.516 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 6.72 22.072 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 6.72 22.328 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 7.44 22.716 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 7.44 22.972 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.16 18.816 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.16 19.028 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 8.88 20.272 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 8.88 20.528 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 9.6 20.916 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 9.6 21.172 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 10.32 21.728 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 10.32 21.816 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 0.96 20.272 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 11.04 22.416 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 11.04 22.628 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 11.76 18.472 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.76 18.728 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 12.48 19.628 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 12.48 19.716 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 13.2 20.616 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 13.2 20.828 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 13.92 21.428 15.12 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 13.92 21.516 15.12 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 0.96 20.528 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 14.64 22.072 15.84 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 14.64 22.328 15.84 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 15.36 22.716 16.56 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 15.36 22.972 16.56 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 16.08 18.816 17.28 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 16.08 19.028 17.28 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 16.8 20.272 18 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 16.8 20.528 18 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 17.52 20.916 18.72 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 17.52 21.172 18.72 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 1.68 20.916 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 23.28 20.616 24.48 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 23.28 20.828 24.48 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 24 19.116 25.2 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 24 19.372 25.2 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 24.72 20.616 25.92 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 24.72 20.828 25.92 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 25.44 21.428 26.64 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 25.44 21.516 26.64 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 26.16 22.072 27.36 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 26.16 22.328 27.36 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 1.68 21.172 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 26.88 22.716 28.08 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 26.88 22.972 28.08 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 27.6 18.816 28.8 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 27.6 19.028 28.8 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 28.32 20.272 29.52 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 28.32 20.528 29.52 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 29.04 20.916 30.24 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 29.04 21.172 30.24 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 29.76 21.728 30.96 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 29.76 21.816 30.96 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 2.4 21.728 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 30.48 22.416 31.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 30.48 22.628 31.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 31.2 18.472 32.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 31.2 18.728 32.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 31.92 19.628 33.12 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 31.92 19.716 33.12 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 32.64 20.616 33.84 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 32.64 20.828 33.84 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 33.36 21.428 34.56 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 33.36 21.516 34.56 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.4 21.816 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 34.08 22.072 35.28 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 34.08 22.328 35.28 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 34.8 22.716 36 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 34.8 22.972 36 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 35.52 18.816 36.72 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 35.52 19.028 36.72 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 36.24 20.272 37.44 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 36.24 20.528 37.44 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 36.96 20.916 38.16 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 36.96 21.172 38.16 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 3.12 22.416 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 37.68 21.728 38.88 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 37.68 21.816 38.88 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 38.4 22.416 39.6 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 38.4 22.628 39.6 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 39.12 18.472 40.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 39.12 18.728 40.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 39.84 19.628 41.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 39.84 19.716 41.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 3.12 22.628 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 41.22 ;
        RECT 2.662 0.06 2.738 41.22 ;
        RECT 4.462 0.06 4.538 41.22 ;
        RECT 6.262 0.06 6.338 41.22 ;
        RECT 8.062 0.06 8.138 41.22 ;
        RECT 9.862 0.06 9.938 41.22 ;
        RECT 11.662 0.06 11.738 41.22 ;
        RECT 13.462 0.06 13.538 41.22 ;
        RECT 15.262 0.06 15.338 41.22 ;
        RECT 17.062 0.06 17.138 41.22 ;
        RECT 18.862 0.06 18.938 41.22 ;
        RECT 20.662 0.06 20.738 41.22 ;
        RECT 22.462 0.06 22.538 41.22 ;
        RECT 24.262 0.06 24.338 41.22 ;
        RECT 26.062 0.06 26.138 41.22 ;
        RECT 27.862 0.06 27.938 41.22 ;
        RECT 29.662 0.06 29.738 41.22 ;
        RECT 31.462 0.06 31.538 41.22 ;
        RECT 33.262 0.06 33.338 41.22 ;
        RECT 35.062 0.06 35.138 41.22 ;
        RECT 36.862 0.06 36.938 41.22 ;
        RECT 38.662 0.06 38.738 41.22 ;
        RECT 40.462 0.06 40.538 41.22 ;
        RECT 42.262 0.06 42.338 41.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 41.22 ;
        RECT 3.562 0.06 3.638 41.22 ;
        RECT 5.362 0.06 5.438 41.22 ;
        RECT 7.162 0.06 7.238 41.22 ;
        RECT 8.962 0.06 9.038 41.22 ;
        RECT 10.762 0.06 10.838 41.22 ;
        RECT 12.562 0.06 12.638 41.22 ;
        RECT 14.362 0.06 14.438 41.22 ;
        RECT 16.162 0.06 16.238 41.22 ;
        RECT 17.962 0.06 18.038 41.22 ;
        RECT 19.762 0.06 19.838 41.22 ;
        RECT 21.562 0.06 21.638 41.22 ;
        RECT 23.362 0.06 23.438 41.22 ;
        RECT 25.162 0.06 25.238 41.22 ;
        RECT 26.962 0.06 27.038 41.22 ;
        RECT 28.762 0.06 28.838 41.22 ;
        RECT 30.562 0.06 30.638 41.22 ;
        RECT 32.362 0.06 32.438 41.22 ;
        RECT 34.162 0.06 34.238 41.22 ;
        RECT 35.962 0.06 36.038 41.22 ;
        RECT 37.762 0.06 37.838 41.22 ;
        RECT 39.562 0.06 39.638 41.22 ;
        RECT 41.362 0.06 41.438 41.22 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 43.216 41.294 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 43.22 41.3 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 43.2705 41.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 43.235 41.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 43.27 41.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 43.259 41.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 43.29 41.342 ;
    LAYER m7 SPACING 0 ;
      RECT 42.338 41.34 43.24 41.4 ;
      RECT 42.338 -0.06 43.292 41.34 ;
      RECT 42.338 -0.12 43.24 -0.06 ;
      RECT 41.438 -0.12 42.262 41.4 ;
      RECT 40.538 -0.12 41.362 41.4 ;
      RECT 39.638 -0.12 40.462 41.4 ;
      RECT 38.738 -0.12 39.562 41.4 ;
      RECT 37.838 -0.12 38.662 41.4 ;
      RECT 36.938 -0.12 37.762 41.4 ;
      RECT 36.038 -0.12 36.862 41.4 ;
      RECT 35.138 -0.12 35.962 41.4 ;
      RECT 34.238 -0.12 35.062 41.4 ;
      RECT 33.338 -0.12 34.162 41.4 ;
      RECT 32.438 -0.12 33.262 41.4 ;
      RECT 31.538 -0.12 32.362 41.4 ;
      RECT 30.638 -0.12 31.462 41.4 ;
      RECT 29.738 -0.12 30.562 41.4 ;
      RECT 28.838 -0.12 29.662 41.4 ;
      RECT 27.938 -0.12 28.762 41.4 ;
      RECT 27.038 -0.12 27.862 41.4 ;
      RECT 26.138 -0.12 26.962 41.4 ;
      RECT 25.238 -0.12 26.062 41.4 ;
      RECT 24.338 -0.12 25.162 41.4 ;
      RECT 23.438 22.68 24.262 41.4 ;
      RECT 23.438 21.48 23.828 22.68 ;
      RECT 23.872 21.48 24.262 22.68 ;
      RECT 23.438 20.76 24.262 21.48 ;
      RECT 23.438 19.56 23.484 20.76 ;
      RECT 23.528 19.56 23.572 20.76 ;
      RECT 23.616 19.56 24.262 20.76 ;
      RECT 23.438 -0.12 24.262 19.56 ;
      RECT 22.538 40.32 23.362 41.4 ;
      RECT 22.538 39.6 22.672 40.32 ;
      RECT 22.716 39.12 22.928 40.32 ;
      RECT 22.972 39.12 23.362 40.32 ;
      RECT 22.628 39.12 22.672 39.6 ;
      RECT 22.538 38.4 22.584 39.6 ;
      RECT 22.628 38.4 23.362 39.12 ;
      RECT 22.538 36 23.362 38.4 ;
      RECT 22.538 34.8 22.584 36 ;
      RECT 22.628 34.8 22.672 36 ;
      RECT 22.716 34.8 22.928 36 ;
      RECT 22.972 34.8 23.362 36 ;
      RECT 22.538 32.4 23.362 34.8 ;
      RECT 22.538 31.68 22.672 32.4 ;
      RECT 22.716 31.2 22.928 32.4 ;
      RECT 22.972 31.2 23.362 32.4 ;
      RECT 22.628 31.2 22.672 31.68 ;
      RECT 22.538 30.48 22.584 31.68 ;
      RECT 22.628 30.48 23.362 31.2 ;
      RECT 22.538 28.08 23.362 30.48 ;
      RECT 22.538 26.88 22.584 28.08 ;
      RECT 22.628 26.88 22.672 28.08 ;
      RECT 22.716 26.88 22.928 28.08 ;
      RECT 22.972 26.88 23.362 28.08 ;
      RECT 22.538 24.48 23.362 26.88 ;
      RECT 22.538 23.28 22.672 24.48 ;
      RECT 22.716 23.28 22.928 24.48 ;
      RECT 22.972 23.28 23.362 24.48 ;
      RECT 22.538 20.76 23.362 23.28 ;
      RECT 22.538 19.56 22.584 20.76 ;
      RECT 22.628 19.56 22.672 20.76 ;
      RECT 22.716 19.56 22.928 20.76 ;
      RECT 22.972 19.56 23.184 20.76 ;
      RECT 23.228 19.56 23.272 20.76 ;
      RECT 23.316 19.56 23.362 20.76 ;
      RECT 22.538 16.56 23.362 19.56 ;
      RECT 22.538 15.36 22.584 16.56 ;
      RECT 22.628 15.36 22.672 16.56 ;
      RECT 22.716 15.36 22.928 16.56 ;
      RECT 22.972 15.36 23.362 16.56 ;
      RECT 22.538 12.96 23.362 15.36 ;
      RECT 22.538 12.24 22.672 12.96 ;
      RECT 22.716 11.76 22.928 12.96 ;
      RECT 22.972 11.76 23.362 12.96 ;
      RECT 22.628 11.76 22.672 12.24 ;
      RECT 22.538 11.04 22.584 12.24 ;
      RECT 22.628 11.04 23.362 11.76 ;
      RECT 22.538 8.64 23.362 11.04 ;
      RECT 22.538 7.44 22.584 8.64 ;
      RECT 22.628 7.44 22.672 8.64 ;
      RECT 22.716 7.44 22.928 8.64 ;
      RECT 22.972 7.44 23.362 8.64 ;
      RECT 22.538 5.04 23.362 7.44 ;
      RECT 22.538 4.32 22.672 5.04 ;
      RECT 22.716 3.84 22.928 5.04 ;
      RECT 22.972 3.84 23.362 5.04 ;
      RECT 22.628 3.84 22.672 4.32 ;
      RECT 22.538 3.12 22.584 4.32 ;
      RECT 22.628 3.12 23.362 3.84 ;
      RECT 22.538 -0.12 23.362 3.12 ;
      RECT 21.638 39.6 22.462 41.4 ;
      RECT 21.638 38.88 22.028 39.6 ;
      RECT 22.072 38.4 22.284 39.6 ;
      RECT 22.328 38.4 22.372 39.6 ;
      RECT 22.416 38.4 22.462 39.6 ;
      RECT 21.816 38.4 22.028 38.88 ;
      RECT 21.638 37.68 21.684 38.88 ;
      RECT 21.728 37.68 21.772 38.88 ;
      RECT 21.816 37.68 22.462 38.4 ;
      RECT 21.638 36 22.462 37.68 ;
      RECT 21.638 35.28 22.372 36 ;
      RECT 22.416 34.8 22.462 36 ;
      RECT 22.328 34.8 22.372 35.28 ;
      RECT 21.638 34.08 21.684 35.28 ;
      RECT 21.728 34.08 21.772 35.28 ;
      RECT 21.816 34.08 22.028 35.28 ;
      RECT 22.072 34.08 22.284 35.28 ;
      RECT 22.328 34.08 22.462 34.8 ;
      RECT 21.638 31.68 22.462 34.08 ;
      RECT 21.638 30.96 22.028 31.68 ;
      RECT 22.072 30.48 22.284 31.68 ;
      RECT 22.328 30.48 22.372 31.68 ;
      RECT 22.416 30.48 22.462 31.68 ;
      RECT 21.816 30.48 22.028 30.96 ;
      RECT 21.638 29.76 21.684 30.96 ;
      RECT 21.728 29.76 21.772 30.96 ;
      RECT 21.816 29.76 22.462 30.48 ;
      RECT 21.638 28.08 22.462 29.76 ;
      RECT 21.638 27.36 22.372 28.08 ;
      RECT 22.416 26.88 22.462 28.08 ;
      RECT 22.328 26.88 22.372 27.36 ;
      RECT 21.638 26.16 21.684 27.36 ;
      RECT 21.728 26.16 21.772 27.36 ;
      RECT 21.816 26.16 22.028 27.36 ;
      RECT 22.072 26.16 22.284 27.36 ;
      RECT 22.328 26.16 22.462 26.88 ;
      RECT 21.638 20.76 22.462 26.16 ;
      RECT 21.638 19.56 21.684 20.76 ;
      RECT 21.728 19.56 21.772 20.76 ;
      RECT 21.816 19.56 22.028 20.76 ;
      RECT 22.072 19.56 22.284 20.76 ;
      RECT 22.328 19.56 22.372 20.76 ;
      RECT 22.416 19.56 22.462 20.76 ;
      RECT 21.638 16.56 22.462 19.56 ;
      RECT 21.638 15.84 22.372 16.56 ;
      RECT 22.416 15.36 22.462 16.56 ;
      RECT 22.328 15.36 22.372 15.84 ;
      RECT 21.638 14.64 21.684 15.84 ;
      RECT 21.728 14.64 21.772 15.84 ;
      RECT 21.816 14.64 22.028 15.84 ;
      RECT 22.072 14.64 22.284 15.84 ;
      RECT 22.328 14.64 22.462 15.36 ;
      RECT 21.638 12.24 22.462 14.64 ;
      RECT 21.638 11.52 22.028 12.24 ;
      RECT 22.072 11.04 22.284 12.24 ;
      RECT 22.328 11.04 22.372 12.24 ;
      RECT 22.416 11.04 22.462 12.24 ;
      RECT 21.816 11.04 22.028 11.52 ;
      RECT 21.638 10.32 21.684 11.52 ;
      RECT 21.728 10.32 21.772 11.52 ;
      RECT 21.816 10.32 22.462 11.04 ;
      RECT 21.638 8.64 22.462 10.32 ;
      RECT 21.638 7.92 22.372 8.64 ;
      RECT 22.416 7.44 22.462 8.64 ;
      RECT 22.328 7.44 22.372 7.92 ;
      RECT 21.638 6.72 21.684 7.92 ;
      RECT 21.728 6.72 21.772 7.92 ;
      RECT 21.816 6.72 22.028 7.92 ;
      RECT 22.072 6.72 22.284 7.92 ;
      RECT 22.328 6.72 22.462 7.44 ;
      RECT 21.638 4.32 22.462 6.72 ;
      RECT 21.638 3.6 22.028 4.32 ;
      RECT 22.072 3.12 22.284 4.32 ;
      RECT 22.328 3.12 22.372 4.32 ;
      RECT 22.416 3.12 22.462 4.32 ;
      RECT 21.816 3.12 22.028 3.6 ;
      RECT 21.638 2.4 21.684 3.6 ;
      RECT 21.728 2.4 21.772 3.6 ;
      RECT 21.816 2.4 22.462 3.12 ;
      RECT 21.638 -0.12 22.462 2.4 ;
      RECT 20.738 38.88 21.562 41.4 ;
      RECT 20.738 38.16 21.384 38.88 ;
      RECT 21.428 37.68 21.472 38.88 ;
      RECT 21.516 37.68 21.562 38.88 ;
      RECT 21.172 37.68 21.384 38.16 ;
      RECT 20.738 36.96 20.784 38.16 ;
      RECT 20.828 36.96 20.872 38.16 ;
      RECT 20.916 36.96 21.128 38.16 ;
      RECT 21.172 36.96 21.562 37.68 ;
      RECT 20.738 34.56 21.562 36.96 ;
      RECT 20.738 33.84 20.872 34.56 ;
      RECT 20.916 33.36 21.128 34.56 ;
      RECT 21.172 33.36 21.384 34.56 ;
      RECT 21.428 33.36 21.472 34.56 ;
      RECT 21.516 33.36 21.562 34.56 ;
      RECT 20.828 33.36 20.872 33.84 ;
      RECT 20.738 32.64 20.784 33.84 ;
      RECT 20.828 32.64 21.562 33.36 ;
      RECT 20.738 30.96 21.562 32.64 ;
      RECT 20.738 30.24 21.384 30.96 ;
      RECT 21.428 29.76 21.472 30.96 ;
      RECT 21.516 29.76 21.562 30.96 ;
      RECT 21.172 29.76 21.384 30.24 ;
      RECT 20.738 29.04 20.784 30.24 ;
      RECT 20.828 29.04 20.872 30.24 ;
      RECT 20.916 29.04 21.128 30.24 ;
      RECT 21.172 29.04 21.562 29.76 ;
      RECT 20.738 26.64 21.562 29.04 ;
      RECT 20.738 25.92 20.872 26.64 ;
      RECT 20.916 25.44 21.128 26.64 ;
      RECT 21.172 25.44 21.384 26.64 ;
      RECT 21.428 25.44 21.472 26.64 ;
      RECT 21.516 25.44 21.562 26.64 ;
      RECT 20.828 25.44 20.872 25.92 ;
      RECT 20.738 24.72 20.784 25.92 ;
      RECT 20.828 24.72 21.562 25.44 ;
      RECT 20.738 24.48 21.562 24.72 ;
      RECT 20.738 23.28 20.784 24.48 ;
      RECT 20.828 23.28 21.562 24.48 ;
      RECT 20.738 20.76 21.562 23.28 ;
      RECT 20.738 19.56 21.384 20.76 ;
      RECT 21.428 19.56 21.472 20.76 ;
      RECT 21.516 19.56 21.562 20.76 ;
      RECT 20.738 18.72 21.562 19.56 ;
      RECT 20.738 17.52 20.784 18.72 ;
      RECT 20.828 17.52 20.872 18.72 ;
      RECT 20.916 17.52 21.128 18.72 ;
      RECT 21.172 17.52 21.562 18.72 ;
      RECT 20.738 15.12 21.562 17.52 ;
      RECT 20.738 14.4 20.872 15.12 ;
      RECT 20.916 13.92 21.128 15.12 ;
      RECT 21.172 13.92 21.384 15.12 ;
      RECT 21.428 13.92 21.472 15.12 ;
      RECT 21.516 13.92 21.562 15.12 ;
      RECT 20.828 13.92 20.872 14.4 ;
      RECT 20.738 13.2 20.784 14.4 ;
      RECT 20.828 13.2 21.562 13.92 ;
      RECT 20.738 11.52 21.562 13.2 ;
      RECT 20.738 10.8 21.384 11.52 ;
      RECT 21.428 10.32 21.472 11.52 ;
      RECT 21.516 10.32 21.562 11.52 ;
      RECT 21.172 10.32 21.384 10.8 ;
      RECT 20.738 9.6 20.784 10.8 ;
      RECT 20.828 9.6 20.872 10.8 ;
      RECT 20.916 9.6 21.128 10.8 ;
      RECT 21.172 9.6 21.562 10.32 ;
      RECT 20.738 7.2 21.562 9.6 ;
      RECT 20.738 6.48 20.872 7.2 ;
      RECT 20.916 6 21.128 7.2 ;
      RECT 21.172 6 21.384 7.2 ;
      RECT 21.428 6 21.472 7.2 ;
      RECT 21.516 6 21.562 7.2 ;
      RECT 20.828 6 20.872 6.48 ;
      RECT 20.738 5.28 20.784 6.48 ;
      RECT 20.828 5.28 21.562 6 ;
      RECT 20.738 3.6 21.562 5.28 ;
      RECT 20.738 2.88 21.384 3.6 ;
      RECT 21.428 2.4 21.472 3.6 ;
      RECT 21.516 2.4 21.562 3.6 ;
      RECT 21.172 2.4 21.384 2.88 ;
      RECT 20.738 1.68 20.784 2.88 ;
      RECT 20.828 1.68 20.872 2.88 ;
      RECT 20.916 1.68 21.128 2.88 ;
      RECT 21.172 1.68 21.562 2.4 ;
      RECT 20.738 -0.12 21.562 1.68 ;
      RECT 19.838 38.16 20.662 41.4 ;
      RECT 19.838 37.44 20.572 38.16 ;
      RECT 20.616 36.96 20.662 38.16 ;
      RECT 20.528 36.96 20.572 37.44 ;
      RECT 19.838 36.24 19.884 37.44 ;
      RECT 19.928 36.24 19.972 37.44 ;
      RECT 20.016 36.24 20.228 37.44 ;
      RECT 20.272 36.24 20.484 37.44 ;
      RECT 20.528 36.24 20.662 36.96 ;
      RECT 19.838 33.84 20.662 36.24 ;
      RECT 19.838 32.64 20.228 33.84 ;
      RECT 20.272 32.64 20.484 33.84 ;
      RECT 20.528 32.64 20.572 33.84 ;
      RECT 20.616 32.64 20.662 33.84 ;
      RECT 19.838 30.24 20.662 32.64 ;
      RECT 19.838 29.52 20.572 30.24 ;
      RECT 20.616 29.04 20.662 30.24 ;
      RECT 20.528 29.04 20.572 29.52 ;
      RECT 19.838 28.32 19.884 29.52 ;
      RECT 19.928 28.32 19.972 29.52 ;
      RECT 20.016 28.32 20.228 29.52 ;
      RECT 20.272 28.32 20.484 29.52 ;
      RECT 20.528 28.32 20.662 29.04 ;
      RECT 19.838 25.92 20.662 28.32 ;
      RECT 19.838 24.72 20.228 25.92 ;
      RECT 20.272 24.72 20.484 25.92 ;
      RECT 20.528 24.72 20.572 25.92 ;
      RECT 20.616 24.72 20.662 25.92 ;
      RECT 19.838 24.48 20.662 24.72 ;
      RECT 19.838 23.28 20.572 24.48 ;
      RECT 20.616 23.28 20.662 24.48 ;
      RECT 19.838 22.68 20.662 23.28 ;
      RECT 19.838 21.48 19.884 22.68 ;
      RECT 19.928 21.48 19.972 22.68 ;
      RECT 20.016 21.48 20.228 22.68 ;
      RECT 20.272 21.48 20.484 22.68 ;
      RECT 20.528 21.48 20.662 22.68 ;
      RECT 19.838 18.72 20.662 21.48 ;
      RECT 19.838 18 20.572 18.72 ;
      RECT 20.616 17.52 20.662 18.72 ;
      RECT 20.528 17.52 20.572 18 ;
      RECT 19.838 16.8 19.884 18 ;
      RECT 19.928 16.8 19.972 18 ;
      RECT 20.016 16.8 20.228 18 ;
      RECT 20.272 16.8 20.484 18 ;
      RECT 20.528 16.8 20.662 17.52 ;
      RECT 19.838 14.4 20.662 16.8 ;
      RECT 19.838 13.2 20.228 14.4 ;
      RECT 20.272 13.2 20.484 14.4 ;
      RECT 20.528 13.2 20.572 14.4 ;
      RECT 20.616 13.2 20.662 14.4 ;
      RECT 19.838 10.8 20.662 13.2 ;
      RECT 19.838 10.08 20.572 10.8 ;
      RECT 20.616 9.6 20.662 10.8 ;
      RECT 20.528 9.6 20.572 10.08 ;
      RECT 19.838 8.88 19.884 10.08 ;
      RECT 19.928 8.88 19.972 10.08 ;
      RECT 20.016 8.88 20.228 10.08 ;
      RECT 20.272 8.88 20.484 10.08 ;
      RECT 20.528 8.88 20.662 9.6 ;
      RECT 19.838 6.48 20.662 8.88 ;
      RECT 19.838 5.28 20.228 6.48 ;
      RECT 20.272 5.28 20.484 6.48 ;
      RECT 20.528 5.28 20.572 6.48 ;
      RECT 20.616 5.28 20.662 6.48 ;
      RECT 19.838 2.88 20.662 5.28 ;
      RECT 19.838 2.16 20.572 2.88 ;
      RECT 20.616 1.68 20.662 2.88 ;
      RECT 20.528 1.68 20.572 2.16 ;
      RECT 19.838 0.96 19.884 2.16 ;
      RECT 19.928 0.96 19.972 2.16 ;
      RECT 20.016 0.96 20.228 2.16 ;
      RECT 20.272 0.96 20.484 2.16 ;
      RECT 20.528 0.96 20.662 1.68 ;
      RECT 19.838 -0.12 20.662 0.96 ;
      RECT 18.938 41.04 19.762 41.4 ;
      RECT 18.938 39.84 19.072 41.04 ;
      RECT 19.116 39.84 19.328 41.04 ;
      RECT 19.372 39.84 19.584 41.04 ;
      RECT 19.628 39.84 19.672 41.04 ;
      RECT 19.716 39.84 19.762 41.04 ;
      RECT 18.938 36.72 19.762 39.84 ;
      RECT 18.938 35.52 18.984 36.72 ;
      RECT 19.028 35.52 19.762 36.72 ;
      RECT 18.938 33.12 19.762 35.52 ;
      RECT 18.938 31.92 19.072 33.12 ;
      RECT 19.116 31.92 19.328 33.12 ;
      RECT 19.372 31.92 19.584 33.12 ;
      RECT 19.628 31.92 19.672 33.12 ;
      RECT 19.716 31.92 19.762 33.12 ;
      RECT 18.938 28.8 19.762 31.92 ;
      RECT 18.938 27.6 18.984 28.8 ;
      RECT 19.028 27.6 19.762 28.8 ;
      RECT 18.938 25.2 19.762 27.6 ;
      RECT 18.938 24 18.984 25.2 ;
      RECT 19.028 24 19.072 25.2 ;
      RECT 19.116 24 19.328 25.2 ;
      RECT 19.372 24 19.762 25.2 ;
      RECT 18.938 22.68 19.762 24 ;
      RECT 18.938 21.48 18.984 22.68 ;
      RECT 19.028 21.48 19.072 22.68 ;
      RECT 19.116 21.48 19.328 22.68 ;
      RECT 19.372 21.48 19.584 22.68 ;
      RECT 19.628 21.48 19.672 22.68 ;
      RECT 19.716 21.48 19.762 22.68 ;
      RECT 18.938 17.28 19.762 21.48 ;
      RECT 18.938 16.08 18.984 17.28 ;
      RECT 19.028 16.08 19.762 17.28 ;
      RECT 18.938 13.68 19.762 16.08 ;
      RECT 18.938 12.48 19.072 13.68 ;
      RECT 19.116 12.48 19.328 13.68 ;
      RECT 19.372 12.48 19.584 13.68 ;
      RECT 19.628 12.48 19.672 13.68 ;
      RECT 19.716 12.48 19.762 13.68 ;
      RECT 18.938 9.36 19.762 12.48 ;
      RECT 18.938 8.16 18.984 9.36 ;
      RECT 19.028 8.16 19.762 9.36 ;
      RECT 18.938 5.76 19.762 8.16 ;
      RECT 18.938 4.56 19.072 5.76 ;
      RECT 19.116 4.56 19.328 5.76 ;
      RECT 19.372 4.56 19.584 5.76 ;
      RECT 19.628 4.56 19.672 5.76 ;
      RECT 19.716 4.56 19.762 5.76 ;
      RECT 18.938 1.44 19.762 4.56 ;
      RECT 18.938 0.24 18.984 1.44 ;
      RECT 19.028 0.24 19.762 1.44 ;
      RECT 18.938 -0.12 19.762 0.24 ;
      RECT 18.038 40.32 18.862 41.4 ;
      RECT 18.038 39.12 18.428 40.32 ;
      RECT 18.472 39.12 18.684 40.32 ;
      RECT 18.728 39.12 18.862 40.32 ;
      RECT 18.038 36.72 18.862 39.12 ;
      RECT 18.038 35.52 18.428 36.72 ;
      RECT 18.472 35.52 18.684 36.72 ;
      RECT 18.728 35.52 18.772 36.72 ;
      RECT 18.816 35.52 18.862 36.72 ;
      RECT 18.038 32.4 18.862 35.52 ;
      RECT 18.038 31.2 18.428 32.4 ;
      RECT 18.472 31.2 18.684 32.4 ;
      RECT 18.728 31.2 18.862 32.4 ;
      RECT 18.038 28.8 18.862 31.2 ;
      RECT 18.038 27.6 18.428 28.8 ;
      RECT 18.472 27.6 18.684 28.8 ;
      RECT 18.728 27.6 18.772 28.8 ;
      RECT 18.816 27.6 18.862 28.8 ;
      RECT 18.038 25.2 18.862 27.6 ;
      RECT 18.038 24 18.772 25.2 ;
      RECT 18.816 24 18.862 25.2 ;
      RECT 18.038 22.68 18.862 24 ;
      RECT 18.038 21.48 18.428 22.68 ;
      RECT 18.472 21.48 18.684 22.68 ;
      RECT 18.728 21.48 18.772 22.68 ;
      RECT 18.816 21.48 18.862 22.68 ;
      RECT 18.038 17.28 18.862 21.48 ;
      RECT 18.038 16.08 18.428 17.28 ;
      RECT 18.472 16.08 18.684 17.28 ;
      RECT 18.728 16.08 18.772 17.28 ;
      RECT 18.816 16.08 18.862 17.28 ;
      RECT 18.038 12.96 18.862 16.08 ;
      RECT 18.038 11.76 18.428 12.96 ;
      RECT 18.472 11.76 18.684 12.96 ;
      RECT 18.728 11.76 18.862 12.96 ;
      RECT 18.038 9.36 18.862 11.76 ;
      RECT 18.038 8.16 18.428 9.36 ;
      RECT 18.472 8.16 18.684 9.36 ;
      RECT 18.728 8.16 18.772 9.36 ;
      RECT 18.816 8.16 18.862 9.36 ;
      RECT 18.038 5.04 18.862 8.16 ;
      RECT 18.038 3.84 18.428 5.04 ;
      RECT 18.472 3.84 18.684 5.04 ;
      RECT 18.728 3.84 18.862 5.04 ;
      RECT 18.038 1.44 18.862 3.84 ;
      RECT 18.038 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.772 1.44 ;
      RECT 18.816 0.24 18.862 1.44 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 41.4 ;
      RECT 16.238 -0.12 17.062 41.4 ;
      RECT 15.338 -0.12 16.162 41.4 ;
      RECT 14.438 -0.12 15.262 41.4 ;
      RECT 13.538 -0.12 14.362 41.4 ;
      RECT 12.638 -0.12 13.462 41.4 ;
      RECT 11.738 -0.12 12.562 41.4 ;
      RECT 10.838 -0.12 11.662 41.4 ;
      RECT 9.938 -0.12 10.762 41.4 ;
      RECT 9.038 -0.12 9.862 41.4 ;
      RECT 8.138 -0.12 8.962 41.4 ;
      RECT 7.238 -0.12 8.062 41.4 ;
      RECT 6.338 -0.12 7.162 41.4 ;
      RECT 5.438 -0.12 6.262 41.4 ;
      RECT 4.538 -0.12 5.362 41.4 ;
      RECT 3.638 -0.12 4.462 41.4 ;
      RECT 2.738 -0.12 3.562 41.4 ;
      RECT 1.838 -0.12 2.662 41.4 ;
      RECT 0.938 -0.12 1.762 41.4 ;
      RECT -0.04 41.34 0.862 41.4 ;
      RECT -0.092 -0.06 0.862 41.34 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 42.458 0 43.12 41.28 ;
      RECT 41.558 0 42.142 41.28 ;
      RECT 40.658 0 41.242 41.28 ;
      RECT 39.758 0 40.342 41.28 ;
      RECT 38.858 0 39.442 41.28 ;
      RECT 37.958 0 38.542 41.28 ;
      RECT 37.058 0 37.642 41.28 ;
      RECT 36.158 0 36.742 41.28 ;
      RECT 35.258 0 35.842 41.28 ;
      RECT 34.358 0 34.942 41.28 ;
      RECT 33.458 0 34.042 41.28 ;
      RECT 32.558 0 33.142 41.28 ;
      RECT 31.658 0 32.242 41.28 ;
      RECT 30.758 0 31.342 41.28 ;
      RECT 29.858 0 30.442 41.28 ;
      RECT 28.958 0 29.542 41.28 ;
      RECT 28.058 0 28.642 41.28 ;
      RECT 27.158 0 27.742 41.28 ;
      RECT 26.258 0 26.842 41.28 ;
      RECT 25.358 0 25.942 41.28 ;
      RECT 24.458 0 25.042 41.28 ;
      RECT 23.558 22.8 24.142 41.28 ;
      RECT 23.558 21.36 23.708 22.8 ;
      RECT 23.992 21.36 24.142 22.8 ;
      RECT 23.558 20.88 24.142 21.36 ;
      RECT 23.736 19.44 24.142 20.88 ;
      RECT 23.558 0 24.142 19.44 ;
      RECT 22.658 40.44 23.242 41.28 ;
      RECT 23.092 39 23.242 40.44 ;
      RECT 22.748 38.28 23.242 39 ;
      RECT 22.658 36.12 23.242 38.28 ;
      RECT 23.092 34.68 23.242 36.12 ;
      RECT 22.658 32.52 23.242 34.68 ;
      RECT 23.092 31.08 23.242 32.52 ;
      RECT 22.748 30.36 23.242 31.08 ;
      RECT 22.658 28.2 23.242 30.36 ;
      RECT 23.092 26.76 23.242 28.2 ;
      RECT 22.658 24.6 23.242 26.76 ;
      RECT 23.092 23.16 23.242 24.6 ;
      RECT 22.658 20.88 23.242 23.16 ;
      RECT 21.758 39.72 22.342 41.28 ;
      RECT 21.758 39 21.908 39.72 ;
      RECT 20.858 39 21.442 41.28 ;
      RECT 20.858 38.28 21.264 39 ;
      RECT 19.958 38.28 20.542 41.28 ;
      RECT 19.958 37.56 20.452 38.28 ;
      RECT 19.058 41.16 19.642 41.28 ;
      RECT 18.158 40.44 18.742 41.28 ;
      RECT 18.158 39 18.308 40.44 ;
      RECT 18.158 36.84 18.742 39 ;
      RECT 18.158 35.4 18.308 36.84 ;
      RECT 18.158 32.52 18.742 35.4 ;
      RECT 18.158 31.08 18.308 32.52 ;
      RECT 18.158 28.92 18.742 31.08 ;
      RECT 18.158 27.48 18.308 28.92 ;
      RECT 18.158 25.32 18.742 27.48 ;
      RECT 18.158 23.88 18.652 25.32 ;
      RECT 18.158 22.8 18.742 23.88 ;
      RECT 18.158 21.36 18.308 22.8 ;
      RECT 18.158 17.4 18.742 21.36 ;
      RECT 18.158 15.96 18.308 17.4 ;
      RECT 18.158 13.08 18.742 15.96 ;
      RECT 18.158 11.64 18.308 13.08 ;
      RECT 18.158 9.48 18.742 11.64 ;
      RECT 18.158 8.04 18.308 9.48 ;
      RECT 18.158 5.16 18.742 8.04 ;
      RECT 18.158 3.72 18.308 5.16 ;
      RECT 18.158 1.56 18.742 3.72 ;
      RECT 18.158 0.12 18.308 1.56 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 41.28 ;
      RECT 16.358 0 16.942 41.28 ;
      RECT 15.458 0 16.042 41.28 ;
      RECT 14.558 0 15.142 41.28 ;
      RECT 13.658 0 14.242 41.28 ;
      RECT 12.758 0 13.342 41.28 ;
      RECT 11.858 0 12.442 41.28 ;
      RECT 10.958 0 11.542 41.28 ;
      RECT 10.058 0 10.642 41.28 ;
      RECT 9.158 0 9.742 41.28 ;
      RECT 8.258 0 8.842 41.28 ;
      RECT 7.358 0 7.942 41.28 ;
      RECT 6.458 0 7.042 41.28 ;
      RECT 5.558 0 6.142 41.28 ;
      RECT 4.658 0 5.242 41.28 ;
      RECT 3.758 0 4.342 41.28 ;
      RECT 2.858 0 3.442 41.28 ;
      RECT 1.958 0 2.542 41.28 ;
      RECT 1.058 0 1.642 41.28 ;
      RECT 0.08 0 0.742 41.28 ;
      RECT 19.058 36.84 19.642 39.72 ;
      RECT 19.148 35.4 19.642 36.84 ;
      RECT 19.058 33.24 19.642 35.4 ;
      RECT 21.936 37.56 22.342 38.28 ;
      RECT 21.758 36.12 22.342 37.56 ;
      RECT 21.758 35.4 22.252 36.12 ;
      RECT 21.292 36.84 21.442 37.56 ;
      RECT 20.858 34.68 21.442 36.84 ;
      RECT 19.958 33.96 20.542 36.12 ;
      RECT 19.958 32.52 20.108 33.96 ;
      RECT 19.958 30.36 20.542 32.52 ;
      RECT 19.958 29.64 20.452 30.36 ;
      RECT 21.758 31.8 22.342 33.96 ;
      RECT 21.758 31.08 21.908 31.8 ;
      RECT 20.948 32.52 21.442 33.24 ;
      RECT 20.858 31.08 21.442 32.52 ;
      RECT 20.858 30.36 21.264 31.08 ;
      RECT 19.058 28.92 19.642 31.8 ;
      RECT 19.148 27.48 19.642 28.92 ;
      RECT 19.058 25.32 19.642 27.48 ;
      RECT 19.492 23.88 19.642 25.32 ;
      RECT 19.058 22.8 19.642 23.88 ;
      RECT 21.936 29.64 22.342 30.36 ;
      RECT 21.758 28.2 22.342 29.64 ;
      RECT 21.758 27.48 22.252 28.2 ;
      RECT 21.292 28.92 21.442 29.64 ;
      RECT 20.858 26.76 21.442 28.92 ;
      RECT 19.958 26.04 20.542 28.2 ;
      RECT 19.958 24.6 20.108 26.04 ;
      RECT 19.958 23.16 20.452 24.6 ;
      RECT 19.958 22.8 20.542 23.16 ;
      RECT 21.758 20.88 22.342 26.04 ;
      RECT 20.948 23.16 21.442 25.32 ;
      RECT 20.858 20.88 21.442 23.16 ;
      RECT 20.858 19.44 21.264 20.88 ;
      RECT 20.858 18.84 21.442 19.44 ;
      RECT 21.292 17.4 21.442 18.84 ;
      RECT 20.858 15.24 21.442 17.4 ;
      RECT 19.958 18.84 20.542 21.36 ;
      RECT 19.958 18.12 20.452 18.84 ;
      RECT 19.058 17.4 19.642 21.36 ;
      RECT 19.148 15.96 19.642 17.4 ;
      RECT 19.058 13.8 19.642 15.96 ;
      RECT 22.658 16.68 23.242 19.44 ;
      RECT 23.092 15.24 23.242 16.68 ;
      RECT 22.658 13.08 23.242 15.24 ;
      RECT 23.092 11.64 23.242 13.08 ;
      RECT 22.748 10.92 23.242 11.64 ;
      RECT 22.658 8.76 23.242 10.92 ;
      RECT 23.092 7.32 23.242 8.76 ;
      RECT 22.658 5.16 23.242 7.32 ;
      RECT 23.092 3.72 23.242 5.16 ;
      RECT 22.748 3 23.242 3.72 ;
      RECT 22.658 0 23.242 3 ;
      RECT 21.758 16.68 22.342 19.44 ;
      RECT 21.758 15.96 22.252 16.68 ;
      RECT 19.958 14.52 20.542 16.68 ;
      RECT 19.958 13.08 20.108 14.52 ;
      RECT 19.958 10.92 20.542 13.08 ;
      RECT 19.958 10.2 20.452 10.92 ;
      RECT 21.758 12.36 22.342 14.52 ;
      RECT 21.758 11.64 21.908 12.36 ;
      RECT 20.948 13.08 21.442 13.8 ;
      RECT 20.858 11.64 21.442 13.08 ;
      RECT 20.858 10.92 21.264 11.64 ;
      RECT 19.058 9.48 19.642 12.36 ;
      RECT 19.148 8.04 19.642 9.48 ;
      RECT 19.058 5.88 19.642 8.04 ;
      RECT 21.936 10.2 22.342 10.92 ;
      RECT 21.758 8.76 22.342 10.2 ;
      RECT 21.758 8.04 22.252 8.76 ;
      RECT 21.292 9.48 21.442 10.2 ;
      RECT 20.858 7.32 21.442 9.48 ;
      RECT 19.958 6.6 20.542 8.76 ;
      RECT 19.958 5.16 20.108 6.6 ;
      RECT 19.958 3 20.542 5.16 ;
      RECT 19.958 2.28 20.452 3 ;
      RECT 21.758 4.44 22.342 6.6 ;
      RECT 21.758 3.72 21.908 4.44 ;
      RECT 20.948 5.16 21.442 5.88 ;
      RECT 20.858 3.72 21.442 5.16 ;
      RECT 20.858 3 21.264 3.72 ;
      RECT 19.058 1.56 19.642 4.44 ;
      RECT 19.148 0.12 19.642 1.56 ;
      RECT 19.058 0 19.642 0.12 ;
      RECT 21.936 2.28 22.342 3 ;
      RECT 21.758 0 22.342 2.28 ;
      RECT 21.292 1.56 21.442 2.28 ;
      RECT 20.858 0 21.442 1.56 ;
      RECT 19.958 0 20.542 0.84 ;
    LAYER m0 ;
      RECT 0 0.002 43.2 41.278 ;
    LAYER m1 ;
      RECT 0 0 43.2 41.28 ;
    LAYER m2 ;
      RECT 0 0.015 43.2 41.265 ;
    LAYER m3 ;
      RECT 0.015 0 43.185 41.28 ;
    LAYER m4 ;
      RECT 0 0.02 43.2 41.26 ;
    LAYER m5 ;
      RECT 0.012 0 43.188 41.28 ;
    LAYER m6 ;
      RECT 0 0.012 43.2 41.268 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf096b256e1r1w0cbbeheaa4acw

END LIBRARY
