VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf086b128e1r1w0cbbehsaa4acw
  CLASS BLOCK ;
  FOREIGN arf086b128e1r1w0cbbehsaa4acw ;
  ORIGIN 0 0 ;
  SIZE 23.4 BY 37.44 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 19.56 0.388 20.76 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 17.64 0.388 18.84 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 19.56 1.628 20.76 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 19.56 1.928 20.76 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 19.56 2.356 20.76 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.56 2.616 20.76 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 19.56 2.916 20.76 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 19.56 3.172 20.76 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 19.56 3.728 20.76 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 19.56 0.556 20.76 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 19.56 0.816 20.76 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 19.56 1.116 20.76 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 19.56 1.372 20.76 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 17.64 1.928 18.84 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 17.64 2.356 18.84 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 17.64 2.616 18.84 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 17.64 2.916 18.84 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 17.64 3.172 18.84 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 17.64 3.728 18.84 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 17.64 3.988 18.84 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 17.64 0.556 18.84 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 17.64 0.816 18.84 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.24 1.928 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 3.84 2.828 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 3.84 2.916 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 4.56 2.016 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 4.56 2.188 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.28 2.828 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 5.28 2.916 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 6 2.016 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 6 2.188 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 6.72 2.828 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 6.72 2.916 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 0.24 2.016 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 7.44 2.016 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 7.44 2.188 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 8.16 2.828 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 8.16 2.916 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 8.88 2.016 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 8.88 2.188 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 9.6 2.828 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 9.6 2.916 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 10.32 2.016 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 10.32 2.188 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 0.96 2.616 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 11.04 2.828 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 11.04 2.916 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 11.76 2.016 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 11.76 2.188 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12.48 2.828 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 12.48 2.916 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 13.2 2.016 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 13.2 2.188 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 13.92 2.828 15.12 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 13.92 2.916 15.12 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 0.96 2.828 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 14.64 2.016 15.84 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 14.64 2.188 15.84 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 15.36 2.828 16.56 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 15.36 2.916 16.56 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 16.08 2.016 17.28 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 16.08 2.188 17.28 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 21.6 2.188 22.8 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 21.6 2.272 22.8 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 22.32 2.828 23.52 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 22.32 2.916 23.52 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 1.68 2.016 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 23.04 2.016 24.24 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 23.04 2.188 24.24 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 23.76 2.828 24.96 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 23.76 2.916 24.96 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 24.48 2.016 25.68 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 24.48 2.188 25.68 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 25.2 2.828 26.4 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 25.2 2.916 26.4 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 25.92 2.016 27.12 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 25.92 2.188 27.12 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 1.68 2.188 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 26.64 2.828 27.84 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 26.64 2.916 27.84 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 27.36 2.016 28.56 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 27.36 2.188 28.56 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 28.08 2.828 29.28 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 28.08 2.916 29.28 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 28.8 2.016 30 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 28.8 2.188 30 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 29.52 2.828 30.72 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 29.52 2.916 30.72 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 2.4 2.828 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 30.24 2.016 31.44 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 30.24 2.188 31.44 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 30.96 2.828 32.16 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 30.96 2.916 32.16 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 31.68 2.016 32.88 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 31.68 2.188 32.88 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 32.4 2.828 33.6 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 32.4 2.916 33.6 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 33.12 2.016 34.32 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 33.12 2.188 34.32 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 2.4 2.916 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 33.84 2.828 35.04 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 33.84 2.916 35.04 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 34.56 2.016 35.76 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 34.56 2.188 35.76 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 35.28 2.828 36.48 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 35.28 2.916 36.48 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 36 2.016 37.2 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 36 2.188 37.2 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 3.12 2.016 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 3.12 2.188 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 17.64 1.372 18.84 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 17.64 1.628 18.84 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 17.64 1.116 18.84 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 0.24 3.256 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 3.84 4.156 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 3.84 4.328 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.56 3.428 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 4.56 3.516 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 5.28 4.156 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 5.28 4.328 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6 3.428 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 6 3.516 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 6.72 4.156 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6.72 4.328 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.24 3.428 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 7.44 3.428 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.44 3.516 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 8.16 4.156 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 8.16 4.328 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 8.88 3.428 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.88 3.516 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 9.6 4.156 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.6 4.328 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 10.32 3.428 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 10.32 3.516 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 0.96 4.072 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 11.04 4.156 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 11.04 4.328 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 11.76 3.428 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.76 3.516 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 12.48 4.156 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 12.48 4.328 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 13.2 3.428 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 13.2 3.516 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 13.92 4.156 15.12 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 13.92 4.328 15.12 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 0.96 4.156 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 14.64 3.428 15.84 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 14.64 3.516 15.84 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 15.36 4.156 16.56 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 15.36 4.328 16.56 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.08 3.428 17.28 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.08 3.516 17.28 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 21.6 3.516 22.8 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 21.6 3.816 22.8 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 22.32 4.156 23.52 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 22.32 4.328 23.52 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 1.68 3.428 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 23.04 3.428 24.24 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 23.04 3.516 24.24 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 23.76 4.156 24.96 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 23.76 4.328 24.96 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 24.48 3.428 25.68 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 24.48 3.516 25.68 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 25.2 4.156 26.4 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 25.2 4.328 26.4 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 25.92 3.428 27.12 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 25.92 3.516 27.12 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 1.68 3.516 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 26.64 4.156 27.84 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 26.64 4.328 27.84 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 27.36 3.428 28.56 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 27.36 3.516 28.56 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 28.08 4.156 29.28 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 28.08 4.328 29.28 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 28.8 3.428 30 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 28.8 3.516 30 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 29.52 4.156 30.72 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 29.52 4.328 30.72 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 2.4 4.156 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 30.24 3.428 31.44 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 30.24 3.516 31.44 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 30.96 4.156 32.16 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 30.96 4.328 32.16 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 31.68 3.428 32.88 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 31.68 3.516 32.88 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 32.4 4.156 33.6 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 32.4 4.328 33.6 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 33.12 3.428 34.32 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 33.12 3.516 34.32 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 2.4 4.328 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 33.84 4.156 35.04 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 33.84 4.328 35.04 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 34.56 3.428 35.76 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 34.56 3.516 35.76 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 35.28 4.156 36.48 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 35.28 4.328 36.48 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 36 3.428 37.2 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 36 3.516 37.2 ;
    END
  END rddatap0[87]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 3.12 3.428 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.12 3.516 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 37.38 ;
        RECT 2.662 0.06 2.738 37.38 ;
        RECT 4.462 0.06 4.538 37.38 ;
        RECT 6.262 0.06 6.338 37.38 ;
        RECT 8.062 0.06 8.138 37.38 ;
        RECT 9.862 0.06 9.938 37.38 ;
        RECT 11.662 0.06 11.738 37.38 ;
        RECT 13.462 0.06 13.538 37.38 ;
        RECT 15.262 0.06 15.338 37.38 ;
        RECT 17.062 0.06 17.138 37.38 ;
        RECT 18.862 0.06 18.938 37.38 ;
        RECT 20.662 0.06 20.738 37.38 ;
        RECT 22.462 0.06 22.538 37.38 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 37.38 ;
        RECT 3.562 0.06 3.638 37.38 ;
        RECT 5.362 0.06 5.438 37.38 ;
        RECT 7.162 0.06 7.238 37.38 ;
        RECT 8.962 0.06 9.038 37.38 ;
        RECT 10.762 0.06 10.838 37.38 ;
        RECT 12.562 0.06 12.638 37.38 ;
        RECT 14.362 0.06 14.438 37.38 ;
        RECT 16.162 0.06 16.238 37.38 ;
        RECT 17.962 0.06 18.038 37.38 ;
        RECT 19.762 0.06 19.838 37.38 ;
        RECT 21.562 0.06 21.638 37.38 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 23.416 37.454 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 23.42 37.46 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 23.4705 37.478 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 23.435 37.51 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 23.47 37.478 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 23.459 37.53 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 23.49 37.502 ;
    LAYER m7 SPACING 0 ;
      RECT 22.538 37.5 23.44 37.56 ;
      RECT 22.538 -0.06 23.492 37.5 ;
      RECT 22.538 -0.12 23.44 -0.06 ;
      RECT 21.638 -0.12 22.462 37.56 ;
      RECT 20.738 -0.12 21.562 37.56 ;
      RECT 19.838 -0.12 20.662 37.56 ;
      RECT 18.938 -0.12 19.762 37.56 ;
      RECT 18.038 -0.12 18.862 37.56 ;
      RECT 17.138 -0.12 17.962 37.56 ;
      RECT 16.238 -0.12 17.062 37.56 ;
      RECT 15.338 -0.12 16.162 37.56 ;
      RECT 14.438 -0.12 15.262 37.56 ;
      RECT 13.538 -0.12 14.362 37.56 ;
      RECT 12.638 -0.12 13.462 37.56 ;
      RECT 11.738 -0.12 12.562 37.56 ;
      RECT 10.838 -0.12 11.662 37.56 ;
      RECT 9.938 -0.12 10.762 37.56 ;
      RECT 9.038 -0.12 9.862 37.56 ;
      RECT 8.138 -0.12 8.962 37.56 ;
      RECT 7.238 -0.12 8.062 37.56 ;
      RECT 6.338 -0.12 7.162 37.56 ;
      RECT 5.438 -0.12 6.262 37.56 ;
      RECT 4.538 -0.12 5.362 37.56 ;
      RECT 3.638 36.48 4.462 37.56 ;
      RECT 3.638 35.28 4.112 36.48 ;
      RECT 4.156 35.28 4.284 36.48 ;
      RECT 4.328 35.28 4.462 36.48 ;
      RECT 3.638 35.04 4.462 35.28 ;
      RECT 3.638 33.84 4.112 35.04 ;
      RECT 4.156 33.84 4.284 35.04 ;
      RECT 4.328 33.84 4.462 35.04 ;
      RECT 3.638 33.6 4.462 33.84 ;
      RECT 3.638 32.4 4.112 33.6 ;
      RECT 4.156 32.4 4.284 33.6 ;
      RECT 4.328 32.4 4.462 33.6 ;
      RECT 3.638 32.16 4.462 32.4 ;
      RECT 3.638 30.96 4.112 32.16 ;
      RECT 4.156 30.96 4.284 32.16 ;
      RECT 4.328 30.96 4.462 32.16 ;
      RECT 3.638 30.72 4.462 30.96 ;
      RECT 3.638 29.52 4.112 30.72 ;
      RECT 4.156 29.52 4.284 30.72 ;
      RECT 4.328 29.52 4.462 30.72 ;
      RECT 3.638 29.28 4.462 29.52 ;
      RECT 3.638 28.08 4.112 29.28 ;
      RECT 4.156 28.08 4.284 29.28 ;
      RECT 4.328 28.08 4.462 29.28 ;
      RECT 3.638 27.84 4.462 28.08 ;
      RECT 3.638 26.64 4.112 27.84 ;
      RECT 4.156 26.64 4.284 27.84 ;
      RECT 4.328 26.64 4.462 27.84 ;
      RECT 3.638 26.4 4.462 26.64 ;
      RECT 3.638 25.2 4.112 26.4 ;
      RECT 4.156 25.2 4.284 26.4 ;
      RECT 4.328 25.2 4.462 26.4 ;
      RECT 3.638 24.96 4.462 25.2 ;
      RECT 3.638 23.76 4.112 24.96 ;
      RECT 4.156 23.76 4.284 24.96 ;
      RECT 4.328 23.76 4.462 24.96 ;
      RECT 3.638 23.52 4.462 23.76 ;
      RECT 3.638 22.8 4.112 23.52 ;
      RECT 4.156 22.32 4.284 23.52 ;
      RECT 4.328 22.32 4.462 23.52 ;
      RECT 3.816 22.32 4.112 22.8 ;
      RECT 3.638 21.6 3.772 22.8 ;
      RECT 3.816 21.6 4.462 22.32 ;
      RECT 3.638 20.76 4.462 21.6 ;
      RECT 3.638 19.56 3.684 20.76 ;
      RECT 3.728 19.56 4.462 20.76 ;
      RECT 3.638 18.84 4.462 19.56 ;
      RECT 3.638 17.64 3.684 18.84 ;
      RECT 3.728 17.64 3.944 18.84 ;
      RECT 3.988 17.64 4.462 18.84 ;
      RECT 3.638 16.56 4.462 17.64 ;
      RECT 3.638 15.36 4.112 16.56 ;
      RECT 4.156 15.36 4.284 16.56 ;
      RECT 4.328 15.36 4.462 16.56 ;
      RECT 3.638 15.12 4.462 15.36 ;
      RECT 3.638 13.92 4.112 15.12 ;
      RECT 4.156 13.92 4.284 15.12 ;
      RECT 4.328 13.92 4.462 15.12 ;
      RECT 3.638 13.68 4.462 13.92 ;
      RECT 3.638 12.48 4.112 13.68 ;
      RECT 4.156 12.48 4.284 13.68 ;
      RECT 4.328 12.48 4.462 13.68 ;
      RECT 3.638 12.24 4.462 12.48 ;
      RECT 3.638 11.04 4.112 12.24 ;
      RECT 4.156 11.04 4.284 12.24 ;
      RECT 4.328 11.04 4.462 12.24 ;
      RECT 3.638 10.8 4.462 11.04 ;
      RECT 3.638 9.6 4.112 10.8 ;
      RECT 4.156 9.6 4.284 10.8 ;
      RECT 4.328 9.6 4.462 10.8 ;
      RECT 3.638 9.36 4.462 9.6 ;
      RECT 3.638 8.16 4.112 9.36 ;
      RECT 4.156 8.16 4.284 9.36 ;
      RECT 4.328 8.16 4.462 9.36 ;
      RECT 3.638 7.92 4.462 8.16 ;
      RECT 3.638 6.72 4.112 7.92 ;
      RECT 4.156 6.72 4.284 7.92 ;
      RECT 4.328 6.72 4.462 7.92 ;
      RECT 3.638 6.48 4.462 6.72 ;
      RECT 3.638 5.28 4.112 6.48 ;
      RECT 4.156 5.28 4.284 6.48 ;
      RECT 4.328 5.28 4.462 6.48 ;
      RECT 3.638 5.04 4.462 5.28 ;
      RECT 3.638 3.84 4.112 5.04 ;
      RECT 4.156 3.84 4.284 5.04 ;
      RECT 4.328 3.84 4.462 5.04 ;
      RECT 3.638 3.6 4.462 3.84 ;
      RECT 3.638 2.4 4.112 3.6 ;
      RECT 4.156 2.4 4.284 3.6 ;
      RECT 4.328 2.4 4.462 3.6 ;
      RECT 3.638 2.16 4.462 2.4 ;
      RECT 3.638 0.96 4.028 2.16 ;
      RECT 4.072 0.96 4.112 2.16 ;
      RECT 4.156 0.96 4.462 2.16 ;
      RECT 3.638 -0.12 4.462 0.96 ;
      RECT 2.738 37.2 3.562 37.56 ;
      RECT 2.738 36.48 3.384 37.2 ;
      RECT 3.428 36 3.472 37.2 ;
      RECT 3.516 36 3.562 37.2 ;
      RECT 2.916 36 3.384 36.48 ;
      RECT 2.916 35.76 3.562 36 ;
      RECT 2.738 35.28 2.784 36.48 ;
      RECT 2.828 35.28 2.872 36.48 ;
      RECT 2.916 35.28 3.384 35.76 ;
      RECT 2.738 35.04 3.384 35.28 ;
      RECT 3.428 34.56 3.472 35.76 ;
      RECT 3.516 34.56 3.562 35.76 ;
      RECT 2.916 34.56 3.384 35.04 ;
      RECT 2.916 34.32 3.562 34.56 ;
      RECT 2.738 33.84 2.784 35.04 ;
      RECT 2.828 33.84 2.872 35.04 ;
      RECT 2.916 33.84 3.384 34.32 ;
      RECT 2.738 33.6 3.384 33.84 ;
      RECT 3.428 33.12 3.472 34.32 ;
      RECT 3.516 33.12 3.562 34.32 ;
      RECT 2.916 33.12 3.384 33.6 ;
      RECT 2.916 32.88 3.562 33.12 ;
      RECT 2.738 32.4 2.784 33.6 ;
      RECT 2.828 32.4 2.872 33.6 ;
      RECT 2.916 32.4 3.384 32.88 ;
      RECT 2.738 32.16 3.384 32.4 ;
      RECT 3.428 31.68 3.472 32.88 ;
      RECT 3.516 31.68 3.562 32.88 ;
      RECT 2.916 31.68 3.384 32.16 ;
      RECT 2.916 31.44 3.562 31.68 ;
      RECT 2.738 30.96 2.784 32.16 ;
      RECT 2.828 30.96 2.872 32.16 ;
      RECT 2.916 30.96 3.384 31.44 ;
      RECT 2.738 30.72 3.384 30.96 ;
      RECT 3.428 30.24 3.472 31.44 ;
      RECT 3.516 30.24 3.562 31.44 ;
      RECT 2.916 30.24 3.384 30.72 ;
      RECT 2.916 30 3.562 30.24 ;
      RECT 2.738 29.52 2.784 30.72 ;
      RECT 2.828 29.52 2.872 30.72 ;
      RECT 2.916 29.52 3.384 30 ;
      RECT 2.738 29.28 3.384 29.52 ;
      RECT 3.428 28.8 3.472 30 ;
      RECT 3.516 28.8 3.562 30 ;
      RECT 2.916 28.8 3.384 29.28 ;
      RECT 2.916 28.56 3.562 28.8 ;
      RECT 2.738 28.08 2.784 29.28 ;
      RECT 2.828 28.08 2.872 29.28 ;
      RECT 2.916 28.08 3.384 28.56 ;
      RECT 2.738 27.84 3.384 28.08 ;
      RECT 3.428 27.36 3.472 28.56 ;
      RECT 3.516 27.36 3.562 28.56 ;
      RECT 2.916 27.36 3.384 27.84 ;
      RECT 2.916 27.12 3.562 27.36 ;
      RECT 2.738 26.64 2.784 27.84 ;
      RECT 2.828 26.64 2.872 27.84 ;
      RECT 2.916 26.64 3.384 27.12 ;
      RECT 2.738 26.4 3.384 26.64 ;
      RECT 3.428 25.92 3.472 27.12 ;
      RECT 3.516 25.92 3.562 27.12 ;
      RECT 2.916 25.92 3.384 26.4 ;
      RECT 2.916 25.68 3.562 25.92 ;
      RECT 2.738 25.2 2.784 26.4 ;
      RECT 2.828 25.2 2.872 26.4 ;
      RECT 2.916 25.2 3.384 25.68 ;
      RECT 2.738 24.96 3.384 25.2 ;
      RECT 3.428 24.48 3.472 25.68 ;
      RECT 3.516 24.48 3.562 25.68 ;
      RECT 2.916 24.48 3.384 24.96 ;
      RECT 2.916 24.24 3.562 24.48 ;
      RECT 2.738 23.76 2.784 24.96 ;
      RECT 2.828 23.76 2.872 24.96 ;
      RECT 2.916 23.76 3.384 24.24 ;
      RECT 2.738 23.52 3.384 23.76 ;
      RECT 3.428 23.04 3.472 24.24 ;
      RECT 3.516 23.04 3.562 24.24 ;
      RECT 2.916 23.04 3.384 23.52 ;
      RECT 2.916 22.8 3.562 23.04 ;
      RECT 2.738 22.32 2.784 23.52 ;
      RECT 2.828 22.32 2.872 23.52 ;
      RECT 2.916 22.32 3.472 22.8 ;
      RECT 3.516 21.6 3.562 22.8 ;
      RECT 2.738 21.6 3.472 22.32 ;
      RECT 2.738 20.76 3.562 21.6 ;
      RECT 2.738 19.56 2.872 20.76 ;
      RECT 2.916 19.56 3.128 20.76 ;
      RECT 3.172 19.56 3.562 20.76 ;
      RECT 2.738 18.84 3.562 19.56 ;
      RECT 2.738 17.64 2.872 18.84 ;
      RECT 2.916 17.64 3.128 18.84 ;
      RECT 3.172 17.64 3.562 18.84 ;
      RECT 2.738 17.28 3.562 17.64 ;
      RECT 2.738 16.56 3.384 17.28 ;
      RECT 3.428 16.08 3.472 17.28 ;
      RECT 3.516 16.08 3.562 17.28 ;
      RECT 2.916 16.08 3.384 16.56 ;
      RECT 2.916 15.84 3.562 16.08 ;
      RECT 2.738 15.36 2.784 16.56 ;
      RECT 2.828 15.36 2.872 16.56 ;
      RECT 2.916 15.36 3.384 15.84 ;
      RECT 2.738 15.12 3.384 15.36 ;
      RECT 3.428 14.64 3.472 15.84 ;
      RECT 3.516 14.64 3.562 15.84 ;
      RECT 2.916 14.64 3.384 15.12 ;
      RECT 2.916 14.4 3.562 14.64 ;
      RECT 2.738 13.92 2.784 15.12 ;
      RECT 2.828 13.92 2.872 15.12 ;
      RECT 2.916 13.92 3.384 14.4 ;
      RECT 2.738 13.68 3.384 13.92 ;
      RECT 3.428 13.2 3.472 14.4 ;
      RECT 3.516 13.2 3.562 14.4 ;
      RECT 2.916 13.2 3.384 13.68 ;
      RECT 2.916 12.96 3.562 13.2 ;
      RECT 2.738 12.48 2.784 13.68 ;
      RECT 2.828 12.48 2.872 13.68 ;
      RECT 2.916 12.48 3.384 12.96 ;
      RECT 2.738 12.24 3.384 12.48 ;
      RECT 3.428 11.76 3.472 12.96 ;
      RECT 3.516 11.76 3.562 12.96 ;
      RECT 2.916 11.76 3.384 12.24 ;
      RECT 2.916 11.52 3.562 11.76 ;
      RECT 2.738 11.04 2.784 12.24 ;
      RECT 2.828 11.04 2.872 12.24 ;
      RECT 2.916 11.04 3.384 11.52 ;
      RECT 2.738 10.8 3.384 11.04 ;
      RECT 3.428 10.32 3.472 11.52 ;
      RECT 3.516 10.32 3.562 11.52 ;
      RECT 2.916 10.32 3.384 10.8 ;
      RECT 2.916 10.08 3.562 10.32 ;
      RECT 2.738 9.6 2.784 10.8 ;
      RECT 2.828 9.6 2.872 10.8 ;
      RECT 2.916 9.6 3.384 10.08 ;
      RECT 2.738 9.36 3.384 9.6 ;
      RECT 3.428 8.88 3.472 10.08 ;
      RECT 3.516 8.88 3.562 10.08 ;
      RECT 2.916 8.88 3.384 9.36 ;
      RECT 2.916 8.64 3.562 8.88 ;
      RECT 2.738 8.16 2.784 9.36 ;
      RECT 2.828 8.16 2.872 9.36 ;
      RECT 2.916 8.16 3.384 8.64 ;
      RECT 2.738 7.92 3.384 8.16 ;
      RECT 3.428 7.44 3.472 8.64 ;
      RECT 3.516 7.44 3.562 8.64 ;
      RECT 2.916 7.44 3.384 7.92 ;
      RECT 2.916 7.2 3.562 7.44 ;
      RECT 2.738 6.72 2.784 7.92 ;
      RECT 2.828 6.72 2.872 7.92 ;
      RECT 2.916 6.72 3.384 7.2 ;
      RECT 2.738 6.48 3.384 6.72 ;
      RECT 3.428 6 3.472 7.2 ;
      RECT 3.516 6 3.562 7.2 ;
      RECT 2.916 6 3.384 6.48 ;
      RECT 2.916 5.76 3.562 6 ;
      RECT 2.738 5.28 2.784 6.48 ;
      RECT 2.828 5.28 2.872 6.48 ;
      RECT 2.916 5.28 3.384 5.76 ;
      RECT 2.738 5.04 3.384 5.28 ;
      RECT 3.428 4.56 3.472 5.76 ;
      RECT 3.516 4.56 3.562 5.76 ;
      RECT 2.916 4.56 3.384 5.04 ;
      RECT 2.916 4.32 3.562 4.56 ;
      RECT 2.738 3.84 2.784 5.04 ;
      RECT 2.828 3.84 2.872 5.04 ;
      RECT 2.916 3.84 3.384 4.32 ;
      RECT 2.738 3.6 3.384 3.84 ;
      RECT 3.428 3.12 3.472 4.32 ;
      RECT 3.516 3.12 3.562 4.32 ;
      RECT 2.916 3.12 3.384 3.6 ;
      RECT 2.916 2.88 3.562 3.12 ;
      RECT 2.738 2.4 2.784 3.6 ;
      RECT 2.828 2.4 2.872 3.6 ;
      RECT 2.916 2.4 3.384 2.88 ;
      RECT 2.738 2.16 3.384 2.4 ;
      RECT 3.428 1.68 3.472 2.88 ;
      RECT 3.516 1.68 3.562 2.88 ;
      RECT 2.828 1.68 3.384 2.16 ;
      RECT 2.828 1.44 3.562 1.68 ;
      RECT 2.738 0.96 2.784 2.16 ;
      RECT 2.828 0.96 3.212 1.44 ;
      RECT 3.256 0.24 3.384 1.44 ;
      RECT 3.428 0.24 3.562 1.44 ;
      RECT 2.738 0.24 3.212 0.96 ;
      RECT 2.738 -0.12 3.562 0.24 ;
      RECT 1.838 37.2 2.662 37.56 ;
      RECT 1.838 36 1.972 37.2 ;
      RECT 2.016 36 2.144 37.2 ;
      RECT 2.188 36 2.662 37.2 ;
      RECT 1.838 35.76 2.662 36 ;
      RECT 1.838 34.56 1.972 35.76 ;
      RECT 2.016 34.56 2.144 35.76 ;
      RECT 2.188 34.56 2.662 35.76 ;
      RECT 1.838 34.32 2.662 34.56 ;
      RECT 1.838 33.12 1.972 34.32 ;
      RECT 2.016 33.12 2.144 34.32 ;
      RECT 2.188 33.12 2.662 34.32 ;
      RECT 1.838 32.88 2.662 33.12 ;
      RECT 1.838 31.68 1.972 32.88 ;
      RECT 2.016 31.68 2.144 32.88 ;
      RECT 2.188 31.68 2.662 32.88 ;
      RECT 1.838 31.44 2.662 31.68 ;
      RECT 1.838 30.24 1.972 31.44 ;
      RECT 2.016 30.24 2.144 31.44 ;
      RECT 2.188 30.24 2.662 31.44 ;
      RECT 1.838 30 2.662 30.24 ;
      RECT 1.838 28.8 1.972 30 ;
      RECT 2.016 28.8 2.144 30 ;
      RECT 2.188 28.8 2.662 30 ;
      RECT 1.838 28.56 2.662 28.8 ;
      RECT 1.838 27.36 1.972 28.56 ;
      RECT 2.016 27.36 2.144 28.56 ;
      RECT 2.188 27.36 2.662 28.56 ;
      RECT 1.838 27.12 2.662 27.36 ;
      RECT 1.838 25.92 1.972 27.12 ;
      RECT 2.016 25.92 2.144 27.12 ;
      RECT 2.188 25.92 2.662 27.12 ;
      RECT 1.838 25.68 2.662 25.92 ;
      RECT 1.838 24.48 1.972 25.68 ;
      RECT 2.016 24.48 2.144 25.68 ;
      RECT 2.188 24.48 2.662 25.68 ;
      RECT 1.838 24.24 2.662 24.48 ;
      RECT 1.838 23.04 1.972 24.24 ;
      RECT 2.016 23.04 2.144 24.24 ;
      RECT 2.188 23.04 2.662 24.24 ;
      RECT 1.838 22.8 2.662 23.04 ;
      RECT 1.838 21.6 2.144 22.8 ;
      RECT 2.188 21.6 2.228 22.8 ;
      RECT 2.272 21.6 2.662 22.8 ;
      RECT 1.838 20.76 2.662 21.6 ;
      RECT 1.838 19.56 1.884 20.76 ;
      RECT 1.928 19.56 2.312 20.76 ;
      RECT 2.356 19.56 2.572 20.76 ;
      RECT 2.616 19.56 2.662 20.76 ;
      RECT 1.838 18.84 2.662 19.56 ;
      RECT 1.838 17.64 1.884 18.84 ;
      RECT 1.928 17.64 2.312 18.84 ;
      RECT 2.356 17.64 2.572 18.84 ;
      RECT 2.616 17.64 2.662 18.84 ;
      RECT 1.838 17.28 2.662 17.64 ;
      RECT 1.838 16.08 1.972 17.28 ;
      RECT 2.016 16.08 2.144 17.28 ;
      RECT 2.188 16.08 2.662 17.28 ;
      RECT 1.838 15.84 2.662 16.08 ;
      RECT 1.838 14.64 1.972 15.84 ;
      RECT 2.016 14.64 2.144 15.84 ;
      RECT 2.188 14.64 2.662 15.84 ;
      RECT 1.838 14.4 2.662 14.64 ;
      RECT 1.838 13.2 1.972 14.4 ;
      RECT 2.016 13.2 2.144 14.4 ;
      RECT 2.188 13.2 2.662 14.4 ;
      RECT 1.838 12.96 2.662 13.2 ;
      RECT 1.838 11.76 1.972 12.96 ;
      RECT 2.016 11.76 2.144 12.96 ;
      RECT 2.188 11.76 2.662 12.96 ;
      RECT 1.838 11.52 2.662 11.76 ;
      RECT 1.838 10.32 1.972 11.52 ;
      RECT 2.016 10.32 2.144 11.52 ;
      RECT 2.188 10.32 2.662 11.52 ;
      RECT 1.838 10.08 2.662 10.32 ;
      RECT 1.838 8.88 1.972 10.08 ;
      RECT 2.016 8.88 2.144 10.08 ;
      RECT 2.188 8.88 2.662 10.08 ;
      RECT 1.838 8.64 2.662 8.88 ;
      RECT 1.838 7.44 1.972 8.64 ;
      RECT 2.016 7.44 2.144 8.64 ;
      RECT 2.188 7.44 2.662 8.64 ;
      RECT 1.838 7.2 2.662 7.44 ;
      RECT 1.838 6 1.972 7.2 ;
      RECT 2.016 6 2.144 7.2 ;
      RECT 2.188 6 2.662 7.2 ;
      RECT 1.838 5.76 2.662 6 ;
      RECT 1.838 4.56 1.972 5.76 ;
      RECT 2.016 4.56 2.144 5.76 ;
      RECT 2.188 4.56 2.662 5.76 ;
      RECT 1.838 4.32 2.662 4.56 ;
      RECT 1.838 3.12 1.972 4.32 ;
      RECT 2.016 3.12 2.144 4.32 ;
      RECT 2.188 3.12 2.662 4.32 ;
      RECT 1.838 2.88 2.662 3.12 ;
      RECT 2.188 2.16 2.662 2.88 ;
      RECT 1.838 1.68 1.972 2.88 ;
      RECT 2.016 1.68 2.144 2.88 ;
      RECT 2.188 1.68 2.572 2.16 ;
      RECT 1.838 1.44 2.572 1.68 ;
      RECT 2.616 0.96 2.662 2.16 ;
      RECT 2.016 0.96 2.572 1.44 ;
      RECT 1.838 0.24 1.884 1.44 ;
      RECT 1.928 0.24 1.972 1.44 ;
      RECT 2.016 0.24 2.662 0.96 ;
      RECT 1.838 -0.12 2.662 0.24 ;
      RECT 0.938 20.76 1.762 37.56 ;
      RECT 0.938 19.56 1.072 20.76 ;
      RECT 1.116 19.56 1.328 20.76 ;
      RECT 1.372 19.56 1.584 20.76 ;
      RECT 1.628 19.56 1.762 20.76 ;
      RECT 0.938 18.84 1.762 19.56 ;
      RECT 0.938 17.64 1.072 18.84 ;
      RECT 1.116 17.64 1.328 18.84 ;
      RECT 1.372 17.64 1.584 18.84 ;
      RECT 1.628 17.64 1.762 18.84 ;
      RECT 0.938 -0.12 1.762 17.64 ;
      RECT -0.04 37.5 0.862 37.56 ;
      RECT -0.092 20.76 0.862 37.5 ;
      RECT -0.092 19.56 0.344 20.76 ;
      RECT 0.388 19.56 0.512 20.76 ;
      RECT 0.556 19.56 0.772 20.76 ;
      RECT 0.816 19.56 0.862 20.76 ;
      RECT -0.092 18.84 0.862 19.56 ;
      RECT -0.092 17.64 0.344 18.84 ;
      RECT 0.388 17.64 0.512 18.84 ;
      RECT 0.556 17.64 0.772 18.84 ;
      RECT 0.816 17.64 0.862 18.84 ;
      RECT -0.092 -0.06 0.862 17.64 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 22.658 0 23.32 37.44 ;
      RECT 21.758 0 22.342 37.44 ;
      RECT 20.858 0 21.442 37.44 ;
      RECT 19.958 0 20.542 37.44 ;
      RECT 19.058 0 19.642 37.44 ;
      RECT 18.158 0 18.742 37.44 ;
      RECT 17.258 0 17.842 37.44 ;
      RECT 16.358 0 16.942 37.44 ;
      RECT 15.458 0 16.042 37.44 ;
      RECT 14.558 0 15.142 37.44 ;
      RECT 13.658 0 14.242 37.44 ;
      RECT 12.758 0 13.342 37.44 ;
      RECT 11.858 0 12.442 37.44 ;
      RECT 10.958 0 11.542 37.44 ;
      RECT 10.058 0 10.642 37.44 ;
      RECT 9.158 0 9.742 37.44 ;
      RECT 8.258 0 8.842 37.44 ;
      RECT 7.358 0 7.942 37.44 ;
      RECT 6.458 0 7.042 37.44 ;
      RECT 5.558 0 6.142 37.44 ;
      RECT 4.658 0 5.242 37.44 ;
      RECT 3.758 36.6 4.342 37.44 ;
      RECT 3.758 22.92 3.992 36.6 ;
      RECT 3.936 22.2 3.992 22.92 ;
      RECT 3.936 21.48 4.342 22.2 ;
      RECT 3.758 20.88 4.342 21.48 ;
      RECT 3.848 19.44 4.342 20.88 ;
      RECT 3.758 18.96 4.342 19.44 ;
      RECT 4.108 17.52 4.342 18.96 ;
      RECT 3.758 16.68 4.342 17.52 ;
      RECT 3.758 2.28 3.992 16.68 ;
      RECT 3.758 0.84 3.908 2.28 ;
      RECT 4.276 0.84 4.342 2.28 ;
      RECT 3.758 0 4.342 0.84 ;
      RECT 2.858 37.32 3.442 37.44 ;
      RECT 2.858 36.6 3.264 37.32 ;
      RECT 3.036 22.92 3.264 36.6 ;
      RECT 3.036 22.2 3.352 22.92 ;
      RECT 2.858 21.48 3.352 22.2 ;
      RECT 2.858 20.88 3.442 21.48 ;
      RECT 3.292 19.44 3.442 20.88 ;
      RECT 2.858 18.96 3.442 19.44 ;
      RECT 3.292 17.52 3.442 18.96 ;
      RECT 2.858 17.4 3.442 17.52 ;
      RECT 2.858 16.68 3.264 17.4 ;
      RECT 3.036 2.28 3.264 16.68 ;
      RECT 2.948 1.56 3.264 2.28 ;
      RECT 2.948 0.84 3.092 1.56 ;
      RECT 2.858 0.12 3.092 0.84 ;
      RECT 2.858 0 3.442 0.12 ;
      RECT 1.958 37.32 2.542 37.44 ;
      RECT 2.308 22.92 2.542 37.32 ;
      RECT 1.958 21.48 2.024 22.92 ;
      RECT 2.392 21.48 2.542 22.92 ;
      RECT 1.958 20.88 2.542 21.48 ;
      RECT 2.048 19.44 2.192 20.88 ;
      RECT 1.958 18.96 2.542 19.44 ;
      RECT 2.048 17.52 2.192 18.96 ;
      RECT 1.958 17.4 2.542 17.52 ;
      RECT 2.308 2.28 2.542 17.4 ;
      RECT 2.308 1.56 2.452 2.28 ;
      RECT 2.136 0.84 2.452 1.56 ;
      RECT 2.136 0.12 2.542 0.84 ;
      RECT 1.958 0 2.542 0.12 ;
      RECT 1.058 20.88 1.642 37.44 ;
      RECT 0.08 20.88 0.742 37.44 ;
      RECT 0.08 19.44 0.224 20.88 ;
      RECT 0.08 18.96 0.742 19.44 ;
      RECT 0.08 17.52 0.224 18.96 ;
      RECT 0.08 0 0.742 17.52 ;
      RECT 1.058 18.96 1.642 19.44 ;
      RECT 1.058 0 1.642 17.52 ;
    LAYER m0 ;
      RECT 0 0.002 23.4 37.438 ;
    LAYER m1 ;
      RECT 0 0 23.4 37.44 ;
    LAYER m2 ;
      RECT 0 0.015 23.4 37.425 ;
    LAYER m3 ;
      RECT 0.015 0 23.385 37.44 ;
    LAYER m4 ;
      RECT 0 0.02 23.4 37.42 ;
    LAYER m5 ;
      RECT 0.012 0 23.388 37.44 ;
    LAYER m6 ;
      RECT 0 0.012 23.4 37.428 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf086b128e1r1w0cbbehsaa4acw

END LIBRARY
