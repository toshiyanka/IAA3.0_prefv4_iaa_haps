//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr_b : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv rev -1.00
//
//------------------------------------------------------------------------------

`include "sbcglobal.vm"
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------

module sbr_b
(
  // Synchronous Clock/Reset
  input  logic        clk_200,
  input  logic        rst_b_200,

  // NOA Debug Signal/Clock Outputs
  output logic [31:0] sbr_b_visa_dbgbus_arb,
  output logic [31:0] sbr_b_visa_dbgbus_vp,
  output logic [31:0] sbr_b_visa_p0_dbgbus,
  output logic [31:0] sbr_b_visa_p1_dbgbus,
  output logic [31:0] sbr_b_visa_p2_dbgbus,
  output logic [31:0] sbr_b_visa_p3_dbgbus,
  output logic [31:0] sbr_b_visa_p4_dbgbus,
  output logic [31:0] sbr_b_visa_p5_dbgbus,
  output logic [31:0] sbr_b_visa_p6_dbgbus,
  output logic [31:0] sbr_b_visa_p7_dbgbus,
  output logic        sbr_b_visa_dbgclk,

  // Register wires
  input  logic [ 4:0] cfg_sbr_b_cgovrd,
  input  logic [15:0] cfg_sbr_b_cgctrl,

  input  logic        su_local_ugt,
  // Port 0 declarations
  input  logic [ 2:0] sbr_a_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_sbr_a_side_ism_fabric,
  input  logic        sbr_a_sbr_b_pccup,
  input  logic        sbr_a_sbr_b_npcup,
  output logic        sbr_b_sbr_a_pcput,
  output logic        sbr_b_sbr_a_npput,
  output logic        sbr_b_sbr_a_eom,
  output logic [31:0] sbr_b_sbr_a_payload,
  output logic        sbr_b_sbr_a_pccup,
  output logic        sbr_b_sbr_a_npcup,
  input  logic        sbr_a_sbr_b_pcput,
  input  logic        sbr_a_sbr_b_npput,
  input  logic        sbr_a_sbr_b_eom,
  input  logic [31:0] sbr_a_sbr_b_payload,

  // Port 1 declarations
  input  logic        pcie_afe_sbr_b_side_clkreq,
  output logic        sbr_b_pcie_afe_side_clkack,
  input  logic [ 2:0] pcie_afe_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_pcie_afe_side_ism_fabric,
  input  logic        pcie_afe_sbr_b_pccup,
  input  logic        pcie_afe_sbr_b_npcup,
  output logic        sbr_b_pcie_afe_pcput,
  output logic        sbr_b_pcie_afe_npput,
  output logic        sbr_b_pcie_afe_eom,
  output logic [ 7:0] sbr_b_pcie_afe_payload,
  output logic        sbr_b_pcie_afe_pccup,
  output logic        sbr_b_pcie_afe_npcup,
  input  logic        pcie_afe_sbr_b_pcput,
  input  logic        pcie_afe_sbr_b_npput,
  input  logic        pcie_afe_sbr_b_eom,
  input  logic [ 7:0] pcie_afe_sbr_b_payload,

  // Port 2 declarations
  input  logic        sata_afe_sbr_b_side_clkreq,
  output logic        sbr_b_sata_afe_side_clkack,
  input  logic [ 2:0] sata_afe_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_sata_afe_side_ism_fabric,
  input  logic        sata_afe_sbr_b_pccup,
  input  logic        sata_afe_sbr_b_npcup,
  output logic        sbr_b_sata_afe_pcput,
  output logic        sbr_b_sata_afe_npput,
  output logic        sbr_b_sata_afe_eom,
  output logic [ 7:0] sbr_b_sata_afe_payload,
  output logic        sbr_b_sata_afe_pccup,
  output logic        sbr_b_sata_afe_npcup,
  input  logic        sata_afe_sbr_b_pcput,
  input  logic        sata_afe_sbr_b_npput,
  input  logic        sata_afe_sbr_b_eom,
  input  logic [ 7:0] sata_afe_sbr_b_payload,

  // Port 3 declarations
  input  logic        usb_afe_sbr_b_side_clkreq,
  output logic        sbr_b_usb_afe_side_clkack,
  input  logic [ 2:0] usb_afe_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_usb_afe_side_ism_fabric,
  input  logic        usb_afe_sbr_b_pccup,
  input  logic        usb_afe_sbr_b_npcup,
  output logic        sbr_b_usb_afe_pcput,
  output logic        sbr_b_usb_afe_npput,
  output logic        sbr_b_usb_afe_eom,
  output logic [ 7:0] sbr_b_usb_afe_payload,
  output logic        sbr_b_usb_afe_pccup,
  output logic        sbr_b_usb_afe_npcup,
  input  logic        usb_afe_sbr_b_pcput,
  input  logic        usb_afe_sbr_b_npput,
  input  logic        usb_afe_sbr_b_eom,
  input  logic [ 7:0] usb_afe_sbr_b_payload,

  // Port 4 declarations
  input  logic        sata_ctrl_sbr_b_side_clkreq,
  output logic        sbr_b_sata_ctrl_side_clkack,
  input  logic [ 2:0] sata_ctrl_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_sata_ctrl_side_ism_fabric,
  input  logic        sata_ctrl_sbr_b_pccup,
  input  logic        sata_ctrl_sbr_b_npcup,
  output logic        sbr_b_sata_ctrl_pcput,
  output logic        sbr_b_sata_ctrl_npput,
  output logic        sbr_b_sata_ctrl_eom,
  output logic [ 7:0] sbr_b_sata_ctrl_payload,
  output logic        sbr_b_sata_ctrl_pccup,
  output logic        sbr_b_sata_ctrl_npcup,
  input  logic        sata_ctrl_sbr_b_pcput,
  input  logic        sata_ctrl_sbr_b_npput,
  input  logic        sata_ctrl_sbr_b_eom,
  input  logic [ 7:0] sata_ctrl_sbr_b_payload,

  // Port 5 declarations
  input  logic        pcie_ctrl_sbr_b_side_clkreq,
  output logic        sbr_b_pcie_ctrl_side_clkack,
  input  logic [ 2:0] pcie_ctrl_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_pcie_ctrl_side_ism_fabric,
  input  logic        pcie_ctrl_sbr_b_pccup,
  input  logic        pcie_ctrl_sbr_b_npcup,
  output logic        sbr_b_pcie_ctrl_pcput,
  output logic        sbr_b_pcie_ctrl_npput,
  output logic        sbr_b_pcie_ctrl_eom,
  output logic [ 7:0] sbr_b_pcie_ctrl_payload,
  output logic        sbr_b_pcie_ctrl_pccup,
  output logic        sbr_b_pcie_ctrl_npcup,
  input  logic        pcie_ctrl_sbr_b_pcput,
  input  logic        pcie_ctrl_sbr_b_npput,
  input  logic        pcie_ctrl_sbr_b_eom,
  input  logic [ 7:0] pcie_ctrl_sbr_b_payload,

  // Port 6 declarations
  input  logic        psf_1_sbr_b_side_clkreq,
  output logic        sbr_b_psf_1_side_clkack,
  input  logic [ 2:0] psf_1_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_psf_1_side_ism_fabric,
  input  logic        psf_1_sbr_b_pccup,
  input  logic        psf_1_sbr_b_npcup,
  output logic        sbr_b_psf_1_pcput,
  output logic        sbr_b_psf_1_npput,
  output logic        sbr_b_psf_1_eom,
  output logic [ 7:0] sbr_b_psf_1_payload,
  output logic        sbr_b_psf_1_pccup,
  output logic        sbr_b_psf_1_npcup,
  input  logic        psf_1_sbr_b_pcput,
  input  logic        psf_1_sbr_b_npput,
  input  logic        psf_1_sbr_b_eom,
  input  logic [ 7:0] psf_1_sbr_b_payload,

  // Port 7 declarations
  input  logic        spare_b_sbr_b_side_clkreq,
  output logic        sbr_b_spare_b_side_clkack,
  input  logic [ 2:0] spare_b_sbr_b_side_ism_agent,
  output logic [ 2:0] sbr_b_spare_b_side_ism_fabric,
  input  logic        spare_b_sbr_b_pccup,
  input  logic        spare_b_sbr_b_npcup,
  output logic        sbr_b_spare_b_pcput,
  output logic        sbr_b_spare_b_npput,
  output logic        sbr_b_spare_b_eom,
  output logic [ 7:0] sbr_b_spare_b_payload,
  output logic        sbr_b_spare_b_pccup,
  output logic        sbr_b_spare_b_npcup,
  input  logic        spare_b_sbr_b_pcput,
  input  logic        spare_b_sbr_b_npput,
  input  logic        spare_b_sbr_b_eom,
  input  logic [ 7:0] spare_b_sbr_b_payload
);


//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_b_sbcportmap;
always_comb sbr_b_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr_b (sbr_b)                                 SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  107 { 17'b0_0000_0000_0000_0000 }},   //   254:148      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //   147          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   146          SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //   145          SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0000 }},   //   144:140      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   139:136      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   135:132      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   131:128      SBCPORTMAPTABLE
      {   31 { 17'b0_0000_0000_0000_0000 }},   //   127: 97      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //    96          SBCPORTMAPTABLE
      {    6 { 17'b0_0000_0000_0000_0000 }},   //    95: 90      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //    89          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //    88          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    87: 86      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    85: 84      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0000 }},   //    83: 81      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    80          SBCPORTMAPTABLE
      {   14 { 17'b0_0000_0000_0000_0000 }},   //    79: 66      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    65: 64      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0000 }},   //    63: 59      SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_0000_0001 }},   //    58: 52      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_1000_0000 }},   //    51: 50      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    49: 48      SBCPORTMAPTABLE
      {    9 { 17'b0_0000_0000_0000_0000 }},   //    47: 39      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    38: 37      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //    36          SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //    35: 32      SBCPORTMAPTABLE
      {   14 { 17'b0_0000_0000_0000_0000 }},   //    31: 18      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //    17          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //    16          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    15: 14      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    13: 12      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //    11          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    10          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //     7          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     6:  5      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0001 }}    //     4:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  7;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;
logic                              p6_pcdstvld;
logic                              p7_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic                              p6_npfence;
logic                              p7_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;
logic                              p6_npdstvld;
logic                              p7_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              pms_request;
logic                              p0_pms_request;
logic                              p1_pms_request;
logic                              p2_pms_request;
logic                              p3_pms_request;
logic                              p4_pms_request;
logic                              p5_pms_request;
logic                              p6_pms_request;
logic                              p7_pms_request;
logic                              p0_ism_idle;
logic                              p1_ism_idle;
logic                              p2_ism_idle;
logic                              p3_ism_idle;
logic                              p4_ism_idle;
logic                              p5_ism_idle;
logic                              p6_ism_idle;
logic                              p7_ism_idle;
logic                              p0_cg_inprogress;
logic                              p1_cg_inprogress;
logic                              p2_cg_inprogress;
logic                              p3_cg_inprogress;
logic                              p4_cg_inprogress;
logic                              p5_cg_inprogress;
logic                              p6_cg_inprogress;
logic                              p7_cg_inprogress;
logic                              all_idle;
logic                              arbiter_idle;
logic                              p0_pms_leave_idle;
logic                              p1_pms_leave_idle;
logic                              p2_pms_leave_idle;
logic                              p3_pms_leave_idle;
logic                              p4_pms_leave_idle;
logic                              p5_pms_leave_idle;
logic                              p6_pms_leave_idle;
logic                              p7_pms_leave_idle;
logic                              block_pms_req;
logic                              gated_side_clk;
logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_clkreq;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = cfg_sbr_b_cgctrl[15];
always_comb cfg_clkgatedef    = cfg_sbr_b_cgctrl[14];
always_comb cfg_idlecnt       = cfg_sbr_b_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = cfg_sbr_b_cgovrd[3];
always_comb jta_force_clkreq  = cfg_sbr_b_cgovrd[2];
always_comb jta_force_idle    = cfg_sbr_b_cgovrd[1];
always_comb jta_force_notidle = cfg_sbr_b_cgovrd[0];
always_comb jta_force_creditreq = cfg_sbr_b_cgovrd[4];

logic                              dt_latchopen;
logic                              dt_latchclosed_b;

always_comb dt_latchopen     = '0;
always_comb dt_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_b_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_b_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rst_b_200                     ),
  .clk                 ( clk_200                       ),
  .q                   ( force_idle                    )
);

doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rst_b_200                     ),
  .clk                 ( clk_200                       ),
  .q                   ( force_notidle                 )
);

doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rst_b_200                     ),
  .clk                 ( clk_200                       ),
  .q                   ( force_creditreq               )
);

always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1
                        };

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p7_ism_idle | ~endpoint_pwrgd[7])
                  & ~p7_pms_leave_idle
                  &  (p6_ism_idle | ~endpoint_pwrgd[6])
                  & ~p6_pms_leave_idle
                  &  (p5_ism_idle | ~endpoint_pwrgd[5])
                  & ~p5_pms_leave_idle
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  & ~p4_pms_leave_idle
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  & ~p3_pms_leave_idle
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  & ~p2_pms_leave_idle
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  & ~p1_pms_leave_idle
                  &  (p0_ism_idle | ~endpoint_pwrgd[0])
                  & ~p0_pms_leave_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p7_npfence,
                 p6_npfence,
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p7_pcdstvld,
                 p6_pcdstvld,
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p7_npdstvld,
                 p6_npdstvld,
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .SBCPMUFLOPS         (  0                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk_200                       ),
  .side_rst_b          ( rst_b_200                     ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .block_pms_req       ( block_pms_req                 ),
  .arbiter_idle        ( arbiter_idle                  ),
  .pms_grant           ( pms_request                   ),
  .pms_request         ( pms_request                   ),
  .pms_gated           (                               ),
  .pms_gating          ( 1'b0                          ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( su_local_ugt                  ),
  .dbgbus              ( sbr_b_visa_dbgbus_arb         )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( sbr_b_visa_dbgbus_vp          )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
  logic        p0_side_clk_valid;
  always_comb  p0_side_clk_valid = 1'b1;

sbcport #(
  .EXTMAXPLDBIT        ( 31                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( sbr_a_sbr_b_side_ism_agent    ),
  .side_ism_out        ( sbr_b_sbr_a_side_ism_fabric   ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p0_pms_request                ),
  .pms_grant           ( p0_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .pms_leave_idle      ( p0_pms_leave_idle             ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .ism_idle            ( p0_ism_idle                   ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_b_sbr_a_pccup             ),
  .tnpcup              ( sbr_b_sbr_a_npcup             ),
  .tpcput              ( sbr_a_sbr_b_pcput             ),
  .tnpput              ( sbr_a_sbr_b_npput             ),
  .teom                ( sbr_a_sbr_b_eom               ),
  .tpayload            ( sbr_a_sbr_b_payload           ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( sbr_a_sbr_b_pccup             ),
  .mnpcup              ( sbr_a_sbr_b_npcup             ),
  .mpcput              ( sbr_b_sbr_a_pcput             ),
  .mnpput              ( sbr_b_sbr_a_npput             ),
  .meom                ( sbr_b_sbr_a_eom               ),
  .mpayload            ( sbr_b_sbr_a_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p0_dbgbus          )
);

// Port 1
// Temporary handling of clkack handshake.
logic p1_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_pcie_afe_side_clkack <= 1;
  else
    sbr_b_pcie_afe_side_clkack <= pcie_afe_sbr_b_side_clkreq;

always_comb
  p1_side_clk_valid = sbr_b_pcie_afe_side_clkack | p1_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( pcie_afe_sbr_b_side_ism_agent ),
  .side_ism_out        ( sbr_b_pcie_afe_side_ism_fabric),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p1_pms_request                ),
  .pms_grant           ( p1_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .pms_leave_idle      ( p1_pms_leave_idle             ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .ism_idle            ( p1_ism_idle                   ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_b_pcie_afe_pccup          ),
  .tnpcup              ( sbr_b_pcie_afe_npcup          ),
  .tpcput              ( pcie_afe_sbr_b_pcput          ),
  .tnpput              ( pcie_afe_sbr_b_npput          ),
  .teom                ( pcie_afe_sbr_b_eom            ),
  .tpayload            ( pcie_afe_sbr_b_payload        ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( pcie_afe_sbr_b_pccup          ),
  .mnpcup              ( pcie_afe_sbr_b_npcup          ),
  .mpcput              ( sbr_b_pcie_afe_pcput          ),
  .mnpput              ( sbr_b_pcie_afe_npput          ),
  .meom                ( sbr_b_pcie_afe_eom            ),
  .mpayload            ( sbr_b_pcie_afe_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p1_dbgbus          )
);

// Port 2
// Temporary handling of clkack handshake.
logic p2_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_sata_afe_side_clkack <= 1;
  else
    sbr_b_sata_afe_side_clkack <= sata_afe_sbr_b_side_clkreq;

always_comb
  p2_side_clk_valid = sbr_b_sata_afe_side_clkack | p2_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( sata_afe_sbr_b_side_ism_agent ),
  .side_ism_out        ( sbr_b_sata_afe_side_ism_fabric),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p2_pms_request                ),
  .pms_grant           ( p2_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .pms_leave_idle      ( p2_pms_leave_idle             ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .ism_idle            ( p2_ism_idle                   ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_b_sata_afe_pccup          ),
  .tnpcup              ( sbr_b_sata_afe_npcup          ),
  .tpcput              ( sata_afe_sbr_b_pcput          ),
  .tnpput              ( sata_afe_sbr_b_npput          ),
  .teom                ( sata_afe_sbr_b_eom            ),
  .tpayload            ( sata_afe_sbr_b_payload        ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( sata_afe_sbr_b_pccup          ),
  .mnpcup              ( sata_afe_sbr_b_npcup          ),
  .mpcput              ( sbr_b_sata_afe_pcput          ),
  .mnpput              ( sbr_b_sata_afe_npput          ),
  .meom                ( sbr_b_sata_afe_eom            ),
  .mpayload            ( sbr_b_sata_afe_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p2_dbgbus          )
);

// Port 3
// Temporary handling of clkack handshake.
logic p3_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_usb_afe_side_clkack <= 1;
  else
    sbr_b_usb_afe_side_clkack <= usb_afe_sbr_b_side_clkreq;

always_comb
  p3_side_clk_valid = sbr_b_usb_afe_side_clkack | p3_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( usb_afe_sbr_b_side_ism_agent  ),
  .side_ism_out        ( sbr_b_usb_afe_side_ism_fabric ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p3_pms_request                ),
  .pms_grant           ( p3_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .pms_leave_idle      ( p3_pms_leave_idle             ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .ism_idle            ( p3_ism_idle                   ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_b_usb_afe_pccup           ),
  .tnpcup              ( sbr_b_usb_afe_npcup           ),
  .tpcput              ( usb_afe_sbr_b_pcput           ),
  .tnpput              ( usb_afe_sbr_b_npput           ),
  .teom                ( usb_afe_sbr_b_eom             ),
  .tpayload            ( usb_afe_sbr_b_payload         ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( usb_afe_sbr_b_pccup           ),
  .mnpcup              ( usb_afe_sbr_b_npcup           ),
  .mpcput              ( sbr_b_usb_afe_pcput           ),
  .mnpput              ( sbr_b_usb_afe_npput           ),
  .meom                ( sbr_b_usb_afe_eom             ),
  .mpayload            ( sbr_b_usb_afe_payload         ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p3_dbgbus          )
);

// Port 4
// Temporary handling of clkack handshake.
logic p4_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_sata_ctrl_side_clkack <= 1;
  else
    sbr_b_sata_ctrl_side_clkack <= sata_ctrl_sbr_b_side_clkreq;

always_comb
  p4_side_clk_valid = sbr_b_sata_ctrl_side_clkack | p4_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( sata_ctrl_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_sata_ctrl_side_ism_fabric),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p4_pms_request                ),
  .pms_grant           ( p4_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .pms_leave_idle      ( p4_pms_leave_idle             ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .ism_idle            ( p4_ism_idle                   ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_b_sata_ctrl_pccup         ),
  .tnpcup              ( sbr_b_sata_ctrl_npcup         ),
  .tpcput              ( sata_ctrl_sbr_b_pcput         ),
  .tnpput              ( sata_ctrl_sbr_b_npput         ),
  .teom                ( sata_ctrl_sbr_b_eom           ),
  .tpayload            ( sata_ctrl_sbr_b_payload       ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( sata_ctrl_sbr_b_pccup         ),
  .mnpcup              ( sata_ctrl_sbr_b_npcup         ),
  .mpcput              ( sbr_b_sata_ctrl_pcput         ),
  .mnpput              ( sbr_b_sata_ctrl_npput         ),
  .meom                ( sbr_b_sata_ctrl_eom           ),
  .mpayload            ( sbr_b_sata_ctrl_payload       ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p4_dbgbus          )
);

// Port 5
// Temporary handling of clkack handshake.
logic p5_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_pcie_ctrl_side_clkack <= 1;
  else
    sbr_b_pcie_ctrl_side_clkack <= pcie_ctrl_sbr_b_side_clkreq;

always_comb
  p5_side_clk_valid = sbr_b_pcie_ctrl_side_clkack | p5_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport5 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( pcie_ctrl_sbr_b_side_ism_agent),
  .side_ism_out        ( sbr_b_pcie_ctrl_side_ism_fabric),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p5_pms_request                ),
  .pms_grant           ( p5_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[5] ),
  .pms_leave_idle      ( p5_pms_leave_idle             ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .ism_idle            ( p5_ism_idle                   ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr_b_pcie_ctrl_pccup         ),
  .tnpcup              ( sbr_b_pcie_ctrl_npcup         ),
  .tpcput              ( pcie_ctrl_sbr_b_pcput         ),
  .tnpput              ( pcie_ctrl_sbr_b_npput         ),
  .teom                ( pcie_ctrl_sbr_b_eom           ),
  .tpayload            ( pcie_ctrl_sbr_b_payload       ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( pcie_ctrl_sbr_b_pccup         ),
  .mnpcup              ( pcie_ctrl_sbr_b_npcup         ),
  .mpcput              ( sbr_b_pcie_ctrl_pcput         ),
  .mnpput              ( sbr_b_pcie_ctrl_npput         ),
  .meom                ( sbr_b_pcie_ctrl_eom           ),
  .mpayload            ( sbr_b_pcie_ctrl_payload       ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p5_dbgbus          )
);

// Port 6
// Temporary handling of clkack handshake.
logic p6_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_psf_1_side_clkack <= 1;
  else
    sbr_b_psf_1_side_clkack <= psf_1_sbr_b_side_clkreq;

always_comb
  p6_side_clk_valid = sbr_b_psf_1_side_clkack | p6_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport6 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p6_side_clk_valid             ),
  .side_ism_in         ( psf_1_sbr_b_side_ism_agent    ),
  .side_ism_out        ( sbr_b_psf_1_side_ism_fabric   ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p6_pms_request                ),
  .pms_grant           ( p6_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[6] ),
  .pms_leave_idle      ( p6_pms_leave_idle             ),
  .agent_idle          ( agent_idle[6]                 ),
  .port_idle           ( port_idle[6]                  ),
  .ism_idle            ( p6_ism_idle                   ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr_b_psf_1_pccup             ),
  .tnpcup              ( sbr_b_psf_1_npcup             ),
  .tpcput              ( psf_1_sbr_b_pcput             ),
  .tnpput              ( psf_1_sbr_b_npput             ),
  .teom                ( psf_1_sbr_b_eom               ),
  .tpayload            ( psf_1_sbr_b_payload           ),
  .pctrdy              ( pctrdy[6]                     ),
  .pcirdy              ( pcirdy[6]                     ),
  .pcdata              ( pcdata[6]                     ),
  .pceom               ( pceom[6]                      ),
  .pcdstvld            ( p6_pcdstvld                   ),
  .nptrdy              ( nptrdy[6]                     ),
  .npirdy              ( npirdy[6]                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( npdata[6]                     ),
  .npeom               ( npeom[6]                      ),
  .npdstvld            ( p6_npdstvld                   ),
  .mpccup              ( psf_1_sbr_b_pccup             ),
  .mnpcup              ( psf_1_sbr_b_npcup             ),
  .mpcput              ( sbr_b_psf_1_pcput             ),
  .mnpput              ( sbr_b_psf_1_npput             ),
  .meom                ( sbr_b_psf_1_eom               ),
  .mpayload            ( sbr_b_psf_1_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[6]                    ),
  .enptrdy             ( enptrdy[6]                    ),
  .epcirdy             ( epcirdy[6]                    ),
  .enpirdy             ( enpirdy[6]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p6_dbgbus          )
);

// Port 7
// Temporary handling of clkack handshake.
logic p7_side_clk_valid;
always_ff @(posedge clk_200 or negedge rst_b_200)
  if ( ~ rst_b_200 )
    sbr_b_spare_b_side_clkack <= 1;
  else
    sbr_b_spare_b_side_clkack <= spare_b_sbr_b_side_clkreq;

always_comb
  p7_side_clk_valid = sbr_b_spare_b_side_clkack | p7_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport7 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_200                     ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( spare_b_sbr_b_side_ism_agent  ),
  .side_ism_out        ( sbr_b_spare_b_side_ism_fabric ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p7_pms_request                ),
  .pms_grant           ( p7_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .int_pok             ( endpoint_pwrgd[7] ),
  .pms_leave_idle      ( p7_pms_leave_idle             ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .ism_idle            ( p7_ism_idle                   ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr_b_spare_b_pccup           ),
  .tnpcup              ( sbr_b_spare_b_npcup           ),
  .tpcput              ( spare_b_sbr_b_pcput           ),
  .tnpput              ( spare_b_sbr_b_npput           ),
  .teom                ( spare_b_sbr_b_eom             ),
  .tpayload            ( spare_b_sbr_b_payload         ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( spare_b_sbr_b_pccup           ),
  .mnpcup              ( spare_b_sbr_b_npcup           ),
  .mpcput              ( sbr_b_spare_b_pcput           ),
  .mnpput              ( sbr_b_spare_b_npput           ),
  .meom                ( sbr_b_spare_b_eom             ),
  .mpayload            ( sbr_b_spare_b_payload         ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( sbr_b_visa_p7_dbgbus          )
);

//------------------------------------------------------------------------------
//
// NOA output assignments
//
//------------------------------------------------------------------------------
always_comb sbr_b_visa_dbgclk = clk_200;


//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------

`ifndef IOSF_SB_ASSERT_OFF

 // synopsys translate_off
    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_b_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_b_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk_200 or negedge rst_b_200)

      if (~rst_b_200) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk_200) disable iff (~rst_b_200)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk_200) disable iff (~rst_b_200)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

 // synopsys translate_on
`endif

endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv
//
//------------------------------------------------------------------------------
/*
Endpoint, adac,0, 1, 0, 0, 1, 129, 
Endpoint, apll,0, 1, 0, 0, 1, 139, 
Endpoint, bunit,2, 1, 0, 0, 1, 03, 
Endpoint, cpunit,2, 1, 0, 0, 1, 10, 
Endpoint, cunit,2, 1, 0, 0, 1, 07, 
Endpoint, ddrio,2, 1, 0, 0, 1, 80, 
Endpoint, dfx_jtag,2, 1, 0, 0, 1, 58, 
Endpoint, dfx_lakemore,2, 1, 0, 0, 1, 56, 
Endpoint, dfx_omar,2, 1, 0, 0, 1, 57, 
Endpoint, dpll,0, 1, 0, 0, 1, 138, 
Endpoint, fpll,0, 1, 0, 0, 1, 136, 
Endpoint, hdmi_rx,0, 1, 0, 0, 1, 131, 
Endpoint, hdmi_tx,0, 1, 0, 0, 1, 130, 
Endpoint, hpll,0, 1, 0, 0, 1, 137, 
Endpoint, hunit,2, 1, 0, 0, 1, 02, 
Endpoint, itunit,2, 1, 0, 0, 1, 64, 
Endpoint, legacy,2, 1, 0, 0, 8, 12,13,32,33,34,35,37,38, 
Endpoint, mcu,2, 1, 0, 0, 1, 01, 
Endpoint, pcie_afe,4, 1, 0, 0, 1, 17, 
Endpoint, pcie_ctrl,4, 1, 0, 0, 1, 16, 
Endpoint, psf_1,4, 1, 0, 0, 1, 145, 
Endpoint, psf_3,2, 1, 0, 0, 1, 147, 
Endpoint, punit,1, 1, 0, 0, 1, 04, 
Endpoint, reut_0,2, 1, 0, 0, 1, 84, 
Endpoint, reut_1,2, 1, 0, 0, 1, 85, 
Endpoint, sata_afe,4, 1, 0, 0, 1, 89, 
Endpoint, sata_ctrl,4, 1, 0, 0, 1, 88, 
SyncRouter, sbr_a, sbr_a,0, 0, 0, 3, 4, 4, 0, visa, cfg, 0, 9, sbr_e, sbr_b, sbr_c, dpll, apll, hpll, fpll, punit, spare_a, , , , , , , , 
SyncRouter, sbr_b, sbr_b,4, 0, 0, 3, 4, 4, 0, visa, cfg, 0, 8, sbr_a, pcie_afe, sata_afe, usb_afe, sata_ctrl, pcie_ctrl, psf_1, spare_b, , , , , , , , , 
SyncRouter, sbr_c, sbr_c,2, 0, 0, 3, 4, 4, 0, visa, cfg, 0, 14, sbr_a, sbr_d, vtunit, hunit, bunit, cunit, cpunit, legacy, dfx_lakemore, dfx_omar, dfx_jtag, itunit, psf_3, spare_c, , , 
SyncRouter, sbr_d, sbr_d,2, 0, 0, 3, 4, 4, 0, visa, cfg, 0, 7, sbr_c, mcu, sec, ddrio, reut_0, reut_1, spare_d, , , , , , , , , , 
SyncRouter, sbr_e, sbr_e,5, 0, 0, 3, 4, 4, 0, visa, cfg, 0, 5, sbr_a, vdac, adac, hdmi_tx, hdmi_rx, , , , , , , , , , , , 
Endpoint, sec,3, 1, 0, 0, 1, 65, 
Endpoint, spare_a,0, 1, 0, 0, 2, 48,49, 
Endpoint, spare_b,0, 1, 0, 0, 2, 50,51, 
Endpoint, spare_c,0, 1, 0, 0, 2, 52,53, 
Endpoint, spare_d,0, 1, 0, 0, 2, 54,55, 
Endpoint, usb_afe,4, 1, 0, 0, 1, 96, 
Endpoint, vdac,0, 1, 0, 0, 1, 128, 
Endpoint, vtunit,2, 1, 0, 0, 1, 00, 
ClockReset, 1, clk_100, rst_b_100, 0, , 5ns
ClockReset, 0, clk_200, rst_b_200, 0, , 2.5ns
ClockReset, 2, clk_27, rst_b_27, 0, , 18.5ns
PowerWell, 0, 
PowerWell, 1, well1_pok
PowerWell, 2, well2_pok
PowerWell, 3, well3_pok
PowerWell, 4, well4_pok
PowerWell, 5, well5_pok
*/
//------------------------------------------------------------------------------
