//------------------------------------------------------------------------------------------------------------------------
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2023 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code ("Material") are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//

//------------------------------------------------------------------------------------------------------------------------
// Intel Proprietary        Intel Confidential        Intel Proprietary        Intel Confidential        Intel Proprietary
//------------------------------------------------------------------------------------------------------------------------
// Generated by                  : cudoming
// Generated on                  : April 19, 2023
//------------------------------------------------------------------------------------------------------------------------
// General Information:
// ------------------------------
// 2r2w0c standard array for SDG server designs.
// Behavioral modeling of a parameterized register file core with no DFX features.
// RTL is written in SystemVerilog.
//------------------------------------------------------------------------------------------------------------------------
// Detail Information:
// ------------------------------
// Addresses        : RD/WR addresses are encoded.
//                    Input addresses will be valid at the array in 1 phases after being driven.
//                    Address latency of 1 is corresponding to a B-latch.
// Enables          : RD/WR enables are used to condition the clock and wordlines.
//                  : Input enables will be valid at the array in 1 phases after being driven.
//                    Enable latency of 1 is corresponding to a B-latch.
// Write Data       : Write data will be valid at the array 2 phases after being driven.
//                    Write data latency of 2 is corresponding to a rising-edge flop. 
// Read Data        : Read data will be valid at the output of a SDL 1 phase after being read.
//                    Read data latency of 1 is corresponding to a B-latch.
// Address Offset   : 
//------------------------------------------------------------------------------------------------------------------------

//------------------------------------------------------------------------------------------------------------------------
// Other Information:
// ------------------------------
// SDG RFIP RTL Release Path:
// /p/hdk/rtl/ip_releases/shdk74/array_macro_module
//
//------------------------------------------------------------------------------------------------------------------------


/// Parent Module    : arf028b032e2r2w0cbbehraa4acw_dfx_wrapper
/// Child Module     : array_generic_rwx_std

`ifndef ARF028B032E2R2W0CBBEHRAA4ACW_SV
`define ARF028B032E2R2W0CBBEHRAA4ACW_SV

//------------------------------------------------------------------------------------------------------------------------
// module arf028b032e2r2w0cbbehraa4acw
//------------------------------------------------------------------------------------------------------------------------
module arf028b032e2r2w0cbbehraa4acw #(

//------------------------------------------------------------------------------------------------------------------------
// local parameters
//------------------------------------------------------------------------------------------------------------------------
  localparam MODULE                 = "arf028b032e2r2w0cbbehraa4acw",
  localparam BITS                   = 30,
  localparam ENTRIES                = 32,
  localparam DWIDTH                 = 30,
  localparam AWIDTH                 = 5,
  localparam RD_PORTS               = 2,
  localparam WR_PORTS               = 2,
  localparam CM_PORTS               = 0,
  localparam BPHASE_RD              = 0,
  localparam BPHASE_WR              = 0,
  localparam BPHASE_CM              = 0,
  localparam SEGMENTS               = 0,
  localparam BITS_PER_SEGMENT       = 0,
  localparam SDL_INITVAL            = {1'b0,1'b0},
  localparam ADDRESS_OFFSET         = 0,
  localparam NO_CAM_LATENCY         = 0,
  localparam NO_CAM_LSB             = 0
)
(

//------------------------------------------------------------------------------------------------------------------------
// interfaces
//------------------------------------------------------------------------------------------------------------------------

  //------------------------------
  // read interfaces
  //------------------------------
  input   wire                            ckrdp0,
  input   wire                            rdenp0,
  input   wire    [AWIDTH-1:0]            rdaddrp0,
  output  wire    [DWIDTH-1:0]            rddatap0,
  input   wire                            sdl_initp0,
  input   wire                            ckrdp1,
  input   wire                            rdenp1,
  input   wire    [AWIDTH-1:0]            rdaddrp1,
  output  wire    [DWIDTH-1:0]            rddatap1,
  input   wire                            sdl_initp1,

  //------------------------------
  // write interfaces
  //------------------------------
  input   wire                            ckwrp0,
  input   wire                            wrenp0,
  input   wire    [AWIDTH-1:0]            wraddrp0,
  input   wire    [DWIDTH-1:0]            wrdatap0,
  input   wire                            ckwrp1,
  input   wire                            wrenp1,
  input   wire    [AWIDTH-1:0]            wraddrp1,
  input   wire    [DWIDTH-1:0]            wrdatap1,



  //------------------------------
  // rcb interfaces
  //------------------------------
  input   wire                            rdaddrp0_fd,
  input   wire                            rdaddrp0_rd,
  input   wire                            rdaddrp1_fd,
  input   wire                            rdaddrp1_rd,
  input   wire                            wraddrp0_fd,
  input   wire                            wraddrp0_rd,
  input   wire                            wrdatap0_fd,
  input   wire                            wrdatap0_rd,
  input   wire                            wraddrp1_fd,
  input   wire                            wraddrp1_rd,
  input   wire                            wrdatap1_fd,
  input   wire                            wrdatap1_rd

);



//------------------------------------------------------------------------------------------------------------------------
// instantiation array_generic_rwx_std
//------------------------------------------------------------------------------------------------------------------------
arf028b032e2r2w0cbbehraa4acw_array_generic_rwx_std #
(

  .MODULE                     (MODULE),
  .BITS                       (BITS),
  .ENTRIES                    (ENTRIES),
  .AWIDTH                     (AWIDTH),
  .DWIDTH                     (DWIDTH),
  .RD_PORTS                   (RD_PORTS),
  .WR_PORTS                   (WR_PORTS),
  .CM_PORTS                   (CM_PORTS),
  .BPHASE_RD                  (BPHASE_RD),
  .BPHASE_WR                  (BPHASE_WR),
  .BPHASE_CM                  (BPHASE_CM),
  .SEGMENTS                   (SEGMENTS),
  .BITS_PER_SEGMENT           (BITS_PER_SEGMENT),
  .SDL_INITVAL                (SDL_INITVAL),
  .ADDRESS_OFFSET             (ADDRESS_OFFSET),
  .NO_CAM_LATENCY             (NO_CAM_LATENCY),
  .NO_CAM_LSB                 (NO_CAM_LSB)

)
array_generic
(

  //------------------------------
  // read interfaces
  //------------------------------
  .ckrd             ( {>>{ ckrdp0, ckrdp1  }} ),
  .rden             ( {>>{ rdenp0, rdenp1 }} ),
  .rdaddr           ( {>>{ rdaddrp0, rdaddrp1 }} ),
  .rddata           ( {>>{ rddatap0, rddatap1 }} ),
  .sdl_init         ( {>>{ sdl_initp0, sdl_initp1 }} ),

  //------------------------------
  // write interfaces
  //------------------------------
  .ckwr             ( {>>{ ckwrp0, ckwrp1 }} ),
  .wren             ( {>>{ wrenp0, wrenp1 }} ),
  .wraddr           ( {>>{ wraddrp0, wraddrp1 }} ),
  .wrdata           ( {>>{ wrdatap0, wrdatap1 }} ),



  //------------------------------
  // rcb interfaces
  //------------------------------
  .rdaddr_fd        ( {>>{ rdaddrp0_fd, rdaddrp1_fd }} ),
  .rdaddr_rd        ( {>>{ rdaddrp0_rd, rdaddrp1_rd }} ),
  .wraddr_fd        ( {>>{ wraddrp0_fd, wraddrp1_fd }} ),
  .wraddr_rd        ( {>>{ wraddrp0_rd, wraddrp1_rd }} ),
  .wrdata_fd        ( {>>{ wrdatap0_fd, wrdatap1_fd }} ),
  .wrdata_rd        ( {>>{ wrdatap0_rd, wrdatap1_rd }} )


);

`ifdef INTC_MEM_GLS

  //err variables
  logic errSDL_INITP0, errSDL_INITP1;
  logic errsdl_initp0, errsdl_initp1;
  logic errRDENP0, errRDENP1;
  logic errrdenp0, errrdenp1;
  logic errRDADDRP0, errRDADDRP1;
  logic errrdaddrp0, errrdaddrp1;
  
  logic errWRENP0, errWRENP1;
  logic errwrenp0, errwrenp1;
  logic errWRADDRP0, errWRADDRP1;
  logic errwraddrp0, errwraddrp1;
  logic errWRDATAP0, errWRDATAP1;
  logic errwrdatap0, errwrdatap1;


  always @(errSDL_INITP0) errsdl_initp0 = 1'b1;
  always @(errRDENP0) errrdenp0 = 1'b1;
  always @(errRDADDRP0) errrdaddrp0 = 1'b1;

  always @(errSDL_INITP1) errsdl_initp1 = 1'b1;
  always @(errRDENP1) errrdenp1 = 1'b1;
  always @(errRDADDRP1) errrdaddrp1 = 1'b1;

  always @(errWRENP0) errwrenp0 = 1'b1;
  always @(errWRADDRP0) errwraddrp0 = 1'b1;
  always @(errWRDATAP0) errwrdatap0 = 1'b1;

  always @(errWRENP1) errwrenp1 = 1'b1;
  always @(errWRADDRP1) errwraddrp1 = 1'b1;
  always @(errWRDATAP1) errwrdatap1 = 1'b1;

  always @(negedge ckrdp0) begin
    errsdl_initp0 = 1'b0;
    errrdenp0 = 1'b0;
    errrdaddrp0 = 1'b0;
  end

  always @(negedge ckrdp1) begin
    errsdl_initp1 = 1'b0;
    errrdenp1 = 1'b0;
    errrdaddrp1 = 1'b0;
  end

  always @(negedge ckwrp0) begin
    errwrenp0 = 1'b0;
    errwraddrp0 = 1'b0;
    errwrdatap0 = 1'b0;
  end

  always @(negedge ckwrp1) begin
    errwrenp1 = 1'b0;
    errwraddrp1 = 1'b0;
    errwrdatap1 = 1'b0;
  end


specify
  specparam trddatap0_r = 0.00:0.00:0.00;
  specparam trddatap0_f = 0.00:0.00:0.00;

  specparam trddatap1_r = 0.00:0.00:0.00;
  specparam trddatap1_f = 0.00:0.00:0.00;

  specparam tsdl_initp0_sr = 0.00:0.00:0.00;
  specparam tsdl_initp0_sf = 0.00:0.00:0.00;
  specparam tsdl_initp0_hr = 0.00:0.00:0.00;
  specparam tsdl_initp0_hf = 0.00:0.00:0.00;

  specparam tsdl_initp1_sr = 0.00:0.00:0.00;
  specparam tsdl_initp1_sf = 0.00:0.00:0.00;
  specparam tsdl_initp1_hr = 0.00:0.00:0.00;
  specparam tsdl_initp1_hf = 0.00:0.00:0.00;

  specparam trdenp0_sr = 0.00:0.00:0.00;
  specparam trdenp0_sf = 0.00:0.00:0.00;
  specparam trdenp0_hr = 0.00:0.00:0.00;
  specparam trdenp0_hf = 0.00:0.00:0.00;

  specparam trdenp1_sr = 0.00:0.00:0.00;
  specparam trdenp1_sf = 0.00:0.00:0.00;
  specparam trdenp1_hr = 0.00:0.00:0.00;
  specparam trdenp1_hf = 0.00:0.00:0.00;

  specparam trdaddrp0_sr = 0.00:0.00:0.00;
  specparam trdaddrp0_sf = 0.00:0.00:0.00;
  specparam trdaddrp0_hr = 0.00:0.00:0.00;
  specparam trdaddrp0_hf = 0.00:0.00:0.00;

  specparam trdaddrp1_sr = 0.00:0.00:0.00;
  specparam trdaddrp1_sf = 0.00:0.00:0.00;
  specparam trdaddrp1_hr = 0.00:0.00:0.00;
  specparam trdaddrp1_hf = 0.00:0.00:0.00;

  specparam twrenp0_sr = 0.00:0.00:0.00;
  specparam twrenp0_sf = 0.00:0.00:0.00;
  specparam twrenp0_hr = 0.00:0.00:0.00;
  specparam twrenp0_hf = 0.00:0.00:0.00;

  specparam twrenp1_sr = 0.00:0.00:0.00;
  specparam twrenp1_sf = 0.00:0.00:0.00;
  specparam twrenp1_hr = 0.00:0.00:0.00;
  specparam twrenp1_hf = 0.00:0.00:0.00;

  specparam twraddrp0_sr = 0.00:0.00:0.00;
  specparam twraddrp0_sf = 0.00:0.00:0.00;
  specparam twraddrp0_hr = 0.00:0.00:0.00;
  specparam twraddrp0_hf = 0.00:0.00:0.00;
  specparam twraddrp1_sr = 0.00:0.00:0.00;
  specparam twraddrp1_sf = 0.00:0.00:0.00;
  specparam twraddrp1_hr = 0.00:0.00:0.00;
  specparam twraddrp1_hf = 0.00:0.00:0.00;
  
  specparam twrdatap0_sr = 0.00:0.00:0.00;
  specparam twrdatap0_sf = 0.00:0.00:0.00;
  specparam twrdatap0_hr = 0.00:0.00:0.00;
  specparam twrdatap0_hf = 0.00:0.00:0.00;  
  specparam twrdatap1_sr = 0.00:0.00:0.00;
  specparam twrdatap1_sf = 0.00:0.00:0.00;
  specparam twrdatap1_hr = 0.00:0.00:0.00;
  specparam twrdatap1_hf = 0.00:0.00:0.00;

  //sdl_init
  $setuphold(posedge ckrdp0, posedge sdl_initp0, tsdl_initp0_sr, tsdl_initp0_hr, errSDL_INITP0);
  $setuphold(posedge ckrdp0, negedge sdl_initp0, tsdl_initp0_sf, tsdl_initp0_hf, errSDL_INITP0);

  $setuphold(posedge ckrdp1, posedge sdl_initp1, tsdl_initp1_sr, tsdl_initp1_hr, errSDL_INITP1);
  $setuphold(posedge ckrdp1, negedge sdl_initp1, tsdl_initp1_sf, tsdl_initp1_hf, errSDL_INITP1);


  //rden
  $setuphold(posedge ckrdp0, posedge rdenp0, trdenp0_sr, trdenp0_hr, errRDENP0);
  $setuphold(posedge ckrdp0, negedge rdenp0, trdenp0_sf, trdenp0_hf, errRDENP0);

  $setuphold(posedge ckrdp1, posedge rdenp1, trdenp1_sr, trdenp1_hr, errRDENP1);
  $setuphold(posedge ckrdp1, negedge rdenp1, trdenp1_sf, trdenp1_hf, errRDENP1);

  
  //rdaddr
  $setuphold(posedge ckrdp0, posedge rdaddrp0[4], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[4], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[3], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[3], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[2], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[2], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[1], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[1], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[0], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[0], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);

  $setuphold(posedge ckrdp1, posedge rdaddrp1[4], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[4], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[3], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[3], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[2], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[2], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[1], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[1], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[0], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[0], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);


  //wren
  $setuphold(posedge ckwrp0, posedge wrenp0, twrenp0_sr, twrenp0_hr, errWRENP0);
  $setuphold(posedge ckwrp0, negedge wrenp0, twrenp0_sf, twrenp0_hf, errWRENP0);

  $setuphold(posedge ckwrp1, posedge wrenp1, twrenp1_sr, twrenp1_hr, errWRENP1);
  $setuphold(posedge ckwrp1, negedge wrenp1, twrenp1_sf, twrenp1_hf, errWRENP1);

 
  //wraddr
  $setuphold(posedge ckwrp0, posedge wraddrp0[4], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[4], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[3], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[3], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[2], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[2], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[1], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[1], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[0], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[0], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);

  $setuphold(posedge ckwrp1, posedge wraddrp1[4], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[4], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[3], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[3], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[2], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[2], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[1], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[1], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[0], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[0], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);

  
  //wrdata
  $setuphold(posedge ckwrp0, posedge wrdatap0[29], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[29], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[28], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[28], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[27], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[27], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[26], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[26], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[25], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[25], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[24], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[24], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[23], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[23], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[22], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[22], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[21], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[21], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[20], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[20], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[19], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[19], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[18], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[18], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[17], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[17], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[16], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[16], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[15], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[15], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[14], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[14], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[13], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[13], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[12], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[12], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[11], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[11], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[10], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[10], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[9], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[9], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[8], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[8], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[7], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[7], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[6], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[6], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[5], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[5], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[4], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[4], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[3], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[3], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[2], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[2], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[1], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[1], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[0], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[0], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);

  $setuphold(posedge ckwrp1, posedge wrdatap1[29], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[29], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[28], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[28], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[27], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[27], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[26], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[26], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[25], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[25], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[24], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[24], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[23], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[23], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[22], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[22], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[21], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[21], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[20], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[20], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[19], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[19], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[18], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[18], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[17], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[17], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[16], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[16], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[15], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[15], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[14], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[14], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[13], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[13], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[12], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[12], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[11], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[11], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[10], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[10], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[9], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[9], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[8], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[8], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[7], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[7], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[6], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[6], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[5], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[5], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[4], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[4], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[3], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[3], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[2], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[2], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[1], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[1], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[0], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[0], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);


  //q 
  (posedge ckrdp0 => rddatap0[29]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[28]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[27]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[26]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[25]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[24]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[23]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[22]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[21]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[20]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[19]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[18]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[17]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[16]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[15]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[14]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[13]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[12]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[11]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[10]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[9]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[8]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[7]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[6]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[5]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[4]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[3]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[2]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[1]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[0]) = (trddatap0_r, trddatap0_f);
 
  (posedge ckrdp1 => rddatap1[29]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[28]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[27]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[26]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[25]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[24]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[23]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[22]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[21]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[20]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[19]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[18]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[17]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[16]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[15]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[14]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[13]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[12]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[11]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[10]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[9]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[8]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[7]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[6]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[5]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[4]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[3]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[2]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[1]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[0]) = (trddatap1_r, trddatap1_f);

endspecify

`endif



endmodule // end module arf028b032e2r2w0cbbehraa4acw
`endif // endif ifndef ARF028B032E2R2W0CBBEHRAA4ACW_SV
