
///
///  INTEL CONFIDENTIAL
///
///  Copyright 2015 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
module hqm_rcfwl_gclk_iclk_clkdiv 
 (
    input  logic clk,
    input  logic rst_b,
    input  logic [3:0] div,

    output logic clkdiv
);

//NON_POR DIRECTIVE
//`ifdef EMULATION

hqm_rcfwl_gclk_iclk_clkdiv_emulation iclk_clkdiv_emulation (
   .clk,
   .rst_b,
   .div,
   .clkdiv
);   

//`else

hqm_rcfwl_gclk_iclk_clkpostdiv clkdiv_div (
   .predivout(clk),
   .ratiom3(div),
   .postdiven(rst_b),
   .dutycyc_50p_en(1'b1),

   .clkdivout(clkdiv)
);

//`endif


endmodule
