//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../gen/sbccfg rev 0.61
//  Fabric configuration file:  generated_code/lv0_sbr_cfg_1/lv0_sbr_cfg_1.csv rev -1.00
//
//------------------------------------------------------------------------------

`include "sbcglobal.vm"
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------

module sbr
(
  // Synchronous Clock/Reset
  input  logic        clk,
  input  logic        rstb,

  // Power Well Isolation Input Signals
  input  logic        pd1_pwrgd,

  // DFx signals
  input  logic        dt_latchopen,
  input  logic        dt_latchclosed_b,

  input  logic        su_local_ugt,
  // Port 0 declarations
  input  logic        ep0_sbr_side_clkreq,
  output logic        sbr_ep0_side_clkack,
  input  logic [ 2:0] ep0_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep0_side_ism_fabric,
  input  logic        ep0_sbr_pccup,
  input  logic        ep0_sbr_npcup,
  output logic        sbr_ep0_pcput,
  output logic        sbr_ep0_npput,
  output logic        sbr_ep0_eom,
  output logic [ 7:0] sbr_ep0_payload,
  output logic        sbr_ep0_pccup,
  output logic        sbr_ep0_npcup,
  input  logic        ep0_sbr_pcput,
  input  logic        ep0_sbr_npput,
  input  logic        ep0_sbr_eom,
  input  logic [ 7:0] ep0_sbr_payload,

  // Port 1 declarations
  input  logic        ep1_sbr_side_clkreq,
  output logic        sbr_ep1_side_clkack,
  input  logic [ 2:0] ep1_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep1_side_ism_fabric,
  input  logic        ep1_sbr_pccup,
  input  logic        ep1_sbr_npcup,
  output logic        sbr_ep1_pcput,
  output logic        sbr_ep1_npput,
  output logic        sbr_ep1_eom,
  output logic [ 7:0] sbr_ep1_payload,
  output logic        sbr_ep1_pccup,
  output logic        sbr_ep1_npcup,
  input  logic        ep1_sbr_pcput,
  input  logic        ep1_sbr_npput,
  input  logic        ep1_sbr_eom,
  input  logic [ 7:0] ep1_sbr_payload,

  // Port 2 declarations
  input  logic        ep2_sbr_side_clkreq,
  output logic        sbr_ep2_side_clkack,
  input  logic [ 2:0] ep2_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep2_side_ism_fabric,
  input  logic        ep2_sbr_pccup,
  input  logic        ep2_sbr_npcup,
  output logic        sbr_ep2_pcput,
  output logic        sbr_ep2_npput,
  output logic        sbr_ep2_eom,
  output logic [15:0] sbr_ep2_payload,
  output logic        sbr_ep2_pccup,
  output logic        sbr_ep2_npcup,
  input  logic        ep2_sbr_pcput,
  input  logic        ep2_sbr_npput,
  input  logic        ep2_sbr_eom,
  input  logic [15:0] ep2_sbr_payload,

  // Port 3 declarations
  input  logic        ep3_sbr_side_clkreq,
  output logic        sbr_ep3_side_clkack,
  input  logic [ 2:0] ep3_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep3_side_ism_fabric,
  input  logic        ep3_sbr_pccup,
  input  logic        ep3_sbr_npcup,
  output logic        sbr_ep3_pcput,
  output logic        sbr_ep3_npput,
  output logic        sbr_ep3_eom,
  output logic [15:0] sbr_ep3_payload,
  output logic        sbr_ep3_pccup,
  output logic        sbr_ep3_npcup,
  input  logic        ep3_sbr_pcput,
  input  logic        ep3_sbr_npput,
  input  logic        ep3_sbr_eom,
  input  logic [15:0] ep3_sbr_payload,

  // Port 4 declarations
  input  logic        ep4_sbr_side_clkreq,
  output logic        sbr_ep4_side_clkack,
  input  logic [ 2:0] ep4_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep4_side_ism_fabric,
  input  logic        ep4_sbr_pccup,
  input  logic        ep4_sbr_npcup,
  output logic        sbr_ep4_pcput,
  output logic        sbr_ep4_npput,
  output logic        sbr_ep4_eom,
  output logic [ 7:0] sbr_ep4_payload,
  output logic        sbr_ep4_pccup,
  output logic        sbr_ep4_npcup,
  input  logic        ep4_sbr_pcput,
  input  logic        ep4_sbr_npput,
  input  logic        ep4_sbr_eom,
  input  logic [ 7:0] ep4_sbr_payload,

  // Port 5 declarations
  input  logic        ep5_sbr_side_clkreq,
  output logic        sbr_ep5_side_clkack,
  input  logic [ 2:0] ep5_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep5_side_ism_fabric,
  input  logic        ep5_sbr_pccup,
  input  logic        ep5_sbr_npcup,
  output logic        sbr_ep5_pcput,
  output logic        sbr_ep5_npput,
  output logic        sbr_ep5_eom,
  output logic [ 7:0] sbr_ep5_payload,
  output logic        sbr_ep5_pccup,
  output logic        sbr_ep5_npcup,
  input  logic        ep5_sbr_pcput,
  input  logic        ep5_sbr_npput,
  input  logic        ep5_sbr_eom,
  input  logic [ 7:0] ep5_sbr_payload,

  // Port 6 declarations
  input  logic        ep6_sbr_side_clkreq,
  output logic        sbr_ep6_side_clkack,
  input  logic [ 2:0] ep6_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep6_side_ism_fabric,
  input  logic        ep6_sbr_pccup,
  input  logic        ep6_sbr_npcup,
  output logic        sbr_ep6_pcput,
  output logic        sbr_ep6_npput,
  output logic        sbr_ep6_eom,
  output logic [15:0] sbr_ep6_payload,
  output logic        sbr_ep6_pccup,
  output logic        sbr_ep6_npcup,
  input  logic        ep6_sbr_pcput,
  input  logic        ep6_sbr_npput,
  input  logic        ep6_sbr_eom,
  input  logic [15:0] ep6_sbr_payload,

  // Port 7 declarations
  input  logic        ep7_sbr_side_clkreq,
  output logic        sbr_ep7_side_clkack,
  input  logic [ 2:0] ep7_sbr_side_ism_agent,
  output logic [ 2:0] sbr_ep7_side_ism_fabric,
  input  logic        ep7_sbr_pccup,
  input  logic        ep7_sbr_npcup,
  output logic        sbr_ep7_pcput,
  output logic        sbr_ep7_npput,
  output logic        sbr_ep7_eom,
  output logic [15:0] sbr_ep7_payload,
  output logic        sbr_ep7_pccup,
  output logic        sbr_ep7_npcup,
  input  logic        ep7_sbr_pcput,
  input  logic        ep7_sbr_npput,
  input  logic        ep7_sbr_eom,
  input  logic [15:0] ep7_sbr_payload
);


//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_sbcportmap;
always_comb sbr_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr (sbr)                                     SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  222 { 17'b0_0000_0000_0000_0000 }},   //   254: 33      SBCPORTMAPTABLE
               17'b1_0000_0000_0000_1111,      //    32          SBCPORTMAPTABLE
      {   18 { 17'b0_0000_0000_0000_0000 }},   //    31: 14      SBCPORTMAPTABLE
               17'b0_0000_0000_1000_0000,      //    13          SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //    12          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //    11          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //    10          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //     9          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //     8          SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0010 }},   //     7:  4      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }}    //     3:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  7;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;
logic                              p6_pcdstvld;
logic                              p7_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic                              p6_npfence;
logic                              p7_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;
logic                              p6_npdstvld;
logic                              p7_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              pms_request;
logic                              p0_pms_request;
logic                              p1_pms_request;
logic                              p2_pms_request;
logic                              p3_pms_request;
logic                              p4_pms_request;
logic                              p5_pms_request;
logic                              p6_pms_request;
logic                              p7_pms_request;
logic                              p0_ism_idle;
logic                              p1_ism_idle;
logic                              p2_ism_idle;
logic                              p3_ism_idle;
logic                              p4_ism_idle;
logic                              p5_ism_idle;
logic                              p6_ism_idle;
logic                              p7_ism_idle;
logic                              p0_cg_inprogress;
logic                              p1_cg_inprogress;
logic                              p2_cg_inprogress;
logic                              p3_cg_inprogress;
logic                              p4_cg_inprogress;
logic                              p5_cg_inprogress;
logic                              p6_cg_inprogress;
logic                              p7_cg_inprogress;
logic                              all_idle;
logic                              arbiter_idle;
logic                              p0_pms_leave_idle;
logic                              p1_pms_leave_idle;
logic                              p2_pms_leave_idle;
logic                              p3_pms_leave_idle;
logic                              p4_pms_leave_idle;
logic                              p5_pms_leave_idle;
logic                              p6_pms_leave_idle;
logic                              p7_pms_leave_idle;
logic                              block_pms_req;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                       [31:0] p0_dbgbus;
logic                       [31:0] p1_dbgbus;
logic                       [31:0] p2_dbgbus;
logic                       [31:0] p3_dbgbus;
logic                       [31:0] p4_dbgbus;
logic                       [31:0] p5_dbgbus;
logic                       [31:0] p6_dbgbus;
logic                       [31:0] p7_dbgbus;
logic                              pd1_pwrgd_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_clkreq;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              force_idle;
logic                              force_notidle;

always_comb cfg_clkgaten      = '1;
always_comb cfg_clkgatedef    = '0;
always_comb cfg_idlecnt       = 8'h10;
always_comb jta_clkgate_ovrd  = '0;
always_comb jta_force_clkreq  = '0;
always_comb jta_force_idle    = '0;
always_comb jta_force_notidle = '0;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_idle                    )
);

doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_notidle                 )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
doublesync sync_pd1_pwrgd (
  .d                   ( pd1_pwrgd                     ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( pd1_pwrgd_ff2                 )
);


always_comb endpoint_pwrgd = { pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1
                        };

logic p7_gated_clk;
clock_gate p7_pwr_clkgate  (
  .en ( endpoint_pwrgd[7] ),
  .te                  ( su_local_ugt                  ),
  .clk                 ( clk                           ),
  .enclk ( p7_gated_clk )
);

logic p5_gated_clk;
clock_gate p5_pwr_clkgate  (
  .en ( endpoint_pwrgd[5] ),
  .te                  ( su_local_ugt                  ),
  .clk                 ( clk                           ),
  .enclk ( p5_gated_clk )
);

logic p3_gated_clk;
clock_gate p3_pwr_clkgate  (
  .en ( endpoint_pwrgd[3] ),
  .te                  ( su_local_ugt                  ),
  .clk                 ( clk                           ),
  .enclk ( p3_gated_clk )
);

logic p1_gated_clk;
clock_gate p1_pwr_clkgate  (
  .en ( endpoint_pwrgd[1] ),
  .te                  ( su_local_ugt                  ),
  .clk                 ( clk                           ),
  .enclk ( p1_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &port_idle
                  &  p7_ism_idle
                  & ~p7_pms_leave_idle
                  &  p6_ism_idle
                  & ~p6_pms_leave_idle
                  &  p5_ism_idle
                  & ~p5_pms_leave_idle
                  &  p4_ism_idle
                  & ~p4_pms_leave_idle
                  &  p3_ism_idle
                  & ~p3_pms_leave_idle
                  &  p2_ism_idle
                  & ~p2_pms_leave_idle
                  &  p1_ism_idle
                  & ~p1_pms_leave_idle
                  &  p0_ism_idle
                  & ~p0_pms_leave_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p7_npfence,
                 p6_npfence,
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p7_pcdstvld,
                 p6_pcdstvld,
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p7_npdstvld,
                 p6_npdstvld,
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .SBCPMUFLOPS         (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk                           ),
  .side_rst_b          ( rstb                          ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .block_pms_req       ( block_pms_req                 ),
  .arbiter_idle        ( arbiter_idle                  ),
  .pms_grant           ( pms_request                   ),
  .pms_request         ( pms_request                   ),
  .pms_gated           (                               ),
  .pms_gating          ( 1'b0                          ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( su_local_ugt                  ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
// Temporary handling of clkack handshake.
logic p0_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep0_side_clkack <= 0;
  else
    sbr_ep0_side_clkack <= ep0_sbr_side_clkreq;

always_comb
  p0_side_clk_valid = sbr_ep0_side_clkack | p0_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport0 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( ep0_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep0_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p0_pms_request                ),
  .pms_grant           ( p0_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .int_pok  ( 1'b1 ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p0_pms_leave_idle             ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .ism_idle            ( p0_ism_idle                   ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_ep0_pccup                 ),
  .tnpcup              ( sbr_ep0_npcup                 ),
  .tpcput              ( ep0_sbr_pcput                 ),
  .tnpput              ( ep0_sbr_npput                 ),
  .teom                ( ep0_sbr_eom                   ),
  .tpayload            ( ep0_sbr_payload               ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( ep0_sbr_pccup                 ),
  .mnpcup              ( ep0_sbr_npcup                 ),
  .mpcput              ( sbr_ep0_pcput                 ),
  .mnpput              ( sbr_ep0_npput                 ),
  .meom                ( sbr_ep0_eom                   ),
  .mpayload            ( sbr_ep0_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_creditreq (1'b0),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
// Temporary handling of clkack handshake.
logic p1_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep1_side_clkack <= 0;
  else
    sbr_ep1_side_clkack <= ep1_sbr_side_clkreq;

always_comb
  p1_side_clk_valid = sbr_ep1_side_clkack | p1_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport1 (
  .int_pok  ( 1'b1 ),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( ep1_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep1_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p1_pms_request                ),
  .pms_grant           ( p1_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p1_pms_leave_idle             ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .ism_idle            ( p1_ism_idle                   ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_ep1_pccup                 ),
  .tnpcup              ( sbr_ep1_npcup                 ),
  .tpcput              ( ep1_sbr_pcput                 ),
  .tnpput              ( ep1_sbr_npput                 ),
  .teom                ( ep1_sbr_eom                   ),
  .tpayload            ( ep1_sbr_payload               ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( ep1_sbr_pccup                 ),
  .mnpcup              ( ep1_sbr_npcup                 ),
  .mpcput              ( sbr_ep1_pcput                 ),
  .mnpput              ( sbr_ep1_npput                 ),
  .meom                ( sbr_ep1_eom                   ),
  .mpayload            ( sbr_ep1_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq (1'b0),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p1_dbgbus                     )
);

// Port 2
// Temporary handling of clkack handshake.
logic p2_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep2_side_clkack <= 0;
  else
    sbr_ep2_side_clkack <= ep2_sbr_side_clkreq;

always_comb
  p2_side_clk_valid = sbr_ep2_side_clkack | p2_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport2 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( ep2_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep2_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p2_pms_request                ),
  .pms_grant           ( p2_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p2_pms_leave_idle             ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .ism_idle            ( p2_ism_idle                   ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_ep2_pccup                 ),
  .tnpcup              ( sbr_ep2_npcup                 ),
  .tpcput              ( ep2_sbr_pcput                 ),
  .tnpput              ( ep2_sbr_npput                 ),
  .teom                ( ep2_sbr_eom                   ),
  .tpayload            ( ep2_sbr_payload               ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( ep2_sbr_pccup                 ),
  .mnpcup              ( ep2_sbr_npcup                 ),
  .mpcput              ( sbr_ep2_pcput                 ),
  .mnpput              ( sbr_ep2_npput                 ),
  .meom                ( sbr_ep2_eom                   ),
  .mpayload            ( sbr_ep2_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p2_dbgbus                     )
);

// Port 3
// Temporary handling of clkack handshake.
logic p3_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep3_side_clkack <= 0;
  else
    sbr_ep3_side_clkack <= ep3_sbr_side_clkreq;

always_comb
  p3_side_clk_valid = sbr_ep3_side_clkack | p3_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport3 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p3_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( ep3_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep3_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p3_pms_request                ),
  .pms_grant           ( p3_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p3_pms_leave_idle             ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .ism_idle            ( p3_ism_idle                   ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_ep3_pccup                 ),
  .tnpcup              ( sbr_ep3_npcup                 ),
  .tpcput              ( ep3_sbr_pcput                 ),
  .tnpput              ( ep3_sbr_npput                 ),
  .teom                ( ep3_sbr_eom                   ),
  .tpayload            ( ep3_sbr_payload               ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( ep3_sbr_pccup                 ),
  .mnpcup              ( ep3_sbr_npcup                 ),
  .mpcput              ( sbr_ep3_pcput                 ),
  .mnpput              ( sbr_ep3_npput                 ),
  .meom                ( sbr_ep3_eom                   ),
  .mpayload            ( sbr_ep3_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
// Temporary handling of clkack handshake.
logic p4_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep4_side_clkack <= 0;
  else
    sbr_ep4_side_clkack <= ep4_sbr_side_clkreq;

always_comb
  p4_side_clk_valid = sbr_ep4_side_clkack | p4_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport4 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( ep4_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep4_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p4_pms_request                ),
  .pms_grant           ( p4_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p4_pms_leave_idle             ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .ism_idle            ( p4_ism_idle                   ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_ep4_pccup                 ),
  .tnpcup              ( sbr_ep4_npcup                 ),
  .tpcput              ( ep4_sbr_pcput                 ),
  .tnpput              ( ep4_sbr_npput                 ),
  .teom                ( ep4_sbr_eom                   ),
  .tpayload            ( ep4_sbr_payload               ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( ep4_sbr_pccup                 ),
  .mnpcup              ( ep4_sbr_npcup                 ),
  .mpcput              ( sbr_ep4_pcput                 ),
  .mnpput              ( sbr_ep4_npput                 ),
  .meom                ( sbr_ep4_eom                   ),
  .mpayload            ( sbr_ep4_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p4_dbgbus                     )
);

// Port 5
// Temporary handling of clkack handshake.
logic p5_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep5_side_clkack <= 0;
  else
    sbr_ep5_side_clkack <= ep5_sbr_side_clkreq;

always_comb
  p5_side_clk_valid = sbr_ep5_side_clkack | p5_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport5 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p5_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( ep5_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep5_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p5_pms_request                ),
  .pms_grant           ( p5_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p5_pms_leave_idle             ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .ism_idle            ( p5_ism_idle                   ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr_ep5_pccup                 ),
  .tnpcup              ( sbr_ep5_npcup                 ),
  .tpcput              ( ep5_sbr_pcput                 ),
  .tnpput              ( ep5_sbr_npput                 ),
  .teom                ( ep5_sbr_eom                   ),
  .tpayload            ( ep5_sbr_payload               ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( ep5_sbr_pccup                 ),
  .mnpcup              ( ep5_sbr_npcup                 ),
  .mpcput              ( sbr_ep5_pcput                 ),
  .mnpput              ( sbr_ep5_npput                 ),
  .meom                ( sbr_ep5_eom                   ),
  .mpayload            ( sbr_ep5_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p5_dbgbus                     )
);

// Port 6
// Temporary handling of clkack handshake.
logic p6_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep6_side_clkack <= 0;
  else
    sbr_ep6_side_clkack <= ep6_sbr_side_clkreq;

always_comb
  p6_side_clk_valid = sbr_ep6_side_clkack | p6_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport6 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p6_side_clk_valid             ),
  .side_ism_in         ( ep6_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep6_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p6_pms_request                ),
  .pms_grant           ( p6_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p6_pms_leave_idle             ),
  .agent_idle          ( agent_idle[6]                 ),
  .port_idle           ( port_idle[6]                  ),
  .ism_idle            ( p6_ism_idle                   ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr_ep6_pccup                 ),
  .tnpcup              ( sbr_ep6_npcup                 ),
  .tpcput              ( ep6_sbr_pcput                 ),
  .tnpput              ( ep6_sbr_npput                 ),
  .teom                ( ep6_sbr_eom                   ),
  .tpayload            ( ep6_sbr_payload               ),
  .pctrdy              ( pctrdy[6]                     ),
  .pcirdy              ( pcirdy[6]                     ),
  .pcdata              ( pcdata[6]                     ),
  .pceom               ( pceom[6]                      ),
  .pcdstvld            ( p6_pcdstvld                   ),
  .nptrdy              ( nptrdy[6]                     ),
  .npirdy              ( npirdy[6]                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( npdata[6]                     ),
  .npeom               ( npeom[6]                      ),
  .npdstvld            ( p6_npdstvld                   ),
  .mpccup              ( ep6_sbr_pccup                 ),
  .mnpcup              ( ep6_sbr_npcup                 ),
  .mpcput              ( sbr_ep6_pcput                 ),
  .mnpput              ( sbr_ep6_npput                 ),
  .meom                ( sbr_ep6_eom                   ),
  .mpayload            ( sbr_ep6_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[6]                    ),
  .enptrdy             ( enptrdy[6]                    ),
  .epcirdy             ( epcirdy[6]                    ),
  .enpirdy             ( enpirdy[6]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p6_dbgbus                     )
);

// Port 7
// Temporary handling of clkack handshake.
logic p7_side_clk_valid;
always_ff @(posedge clk or negedge rstb)
  if ( ~ rstb )
    sbr_ep7_side_clkack <= 0;
  else
    sbr_ep7_side_clkack <= ep7_sbr_side_clkreq;

always_comb
  p7_side_clk_valid = sbr_ep7_side_clkack | p7_pms_leave_idle;

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .QUEUEDEPTH          (  2                            ),
  .SBCISMISAGENT       (  0                            ),
  .SBCPMUFLOPS         (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport7 (
  .int_pok  ( 1'b1 ),
  .force_creditreq (1'b0),
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p7_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( ep7_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep7_side_ism_fabric       ),
  .block_pms_req       ( block_pms_req                 ),
  .pms_request         ( p7_pms_request                ),
  .pms_grant           ( p7_pms_request                ),
  .pms_gating          ( 1'b0                          ),
  .pms_gated           (                               ),
  .pms_leave_idle      ( p7_pms_leave_idle             ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .ism_idle            ( p7_ism_idle                   ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr_ep7_pccup                 ),
  .tnpcup              ( sbr_ep7_npcup                 ),
  .tpcput              ( ep7_sbr_pcput                 ),
  .tnpput              ( ep7_sbr_npput                 ),
  .teom                ( ep7_sbr_eom                   ),
  .tpayload            ( ep7_sbr_payload               ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( ep7_sbr_pccup                 ),
  .mnpcup              ( ep7_sbr_npcup                 ),
  .mpcput              ( sbr_ep7_pcput                 ),
  .mnpput              ( sbr_ep7_npput                 ),
  .meom                ( sbr_ep7_eom                   ),
  .mpayload            ( sbr_ep7_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .dt_latchopen        ( dt_latchopen                  ),
  .dt_latchclosed_b    ( dt_latchclosed_b              ),
  .dbgbus              ( p7_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------

`ifndef IOSF_SB_ASSERT_OFF

 // synopsys translate_off
    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk or negedge rstb)

      if (~rstb) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (~rstb)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (~rstb)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

 // synopsys translate_on
`endif

endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: generated_code/lv0_sbr_cfg_1/lv0_sbr_cfg_1.csv
//
//------------------------------------------------------------------------------
/*
Endpoint, ep0,0, 1, 0, 1, 4, 0,1,2,3, 
Endpoint, ep1,1, 1, 0, 1, 4, 4,5,6,7, 
Endpoint, ep2,0, 2, 0, 1, 1, 8, 
Endpoint, ep3,1, 2, 0, 1, 1, 9, 
Endpoint, ep4,0, 1, 0, 1, 1, 10, 
Endpoint, ep5,1, 1, 0, 1, 1, 11, 
Endpoint, ep6,0, 2, 0, 1, 1, 12, 
Endpoint, ep7,1, 2, 0, 1, 1, 13, 
SyncRouter, sbr, sbr,0, 1, 0, 3, 4, 4, 0, , , 0, 8, ep0, ep1, ep2, ep3, ep4, ep5, ep6, ep7, , , , , , , , , 
Multicast, 32, 4, 0,4,8,9
ClockReset, 0, clk, rstb, 0, , 1ns
PowerWell, 0, 
PowerWell, 1, pd1_pwrgd
*/
//------------------------------------------------------------------------------
