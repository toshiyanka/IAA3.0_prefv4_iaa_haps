`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

,
    (* inserted_by="VISA IT" *) output logic [29:0] visaRt_probe_from_i_hqm_system_visa_probe


`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
