//------------------------------------------------------------------------------
//  INTEL CONFIDENTIAL
//
//  Copyright 2020 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//  Collateral Description:
//  dteg-stap
//
//  Source organization:
//  DTEG Engineering Group (DTEG)
//
//  Support Information:
//  HSD: https://hsdes.intel.com/appstore/article/#/dft_services.bugeco/create
//
//  Revision:
//  DTEG_sTAP_2020WW05_RTL1P0_PIC6_V1
//
//  Module <sTAP> :  < put your functional description here in plain text >
//
//------------------------------------------------------------------------------

//----------------------------------------------------------------------
// Intel Proprietary -- Copyright 2020 Intel -- All rights reserved
//----------------------------------------------------------------------
// NOTE: Log history is at end of file.
//----------------------------------------------------------------------
//
//    FILENAME    : stap_irdecoder.sv
//    DESIGNER    : B.S.Adithya
//    PROJECT     : sTAP
//
//    PURPOSE     : sTAP IR Decoder Logic
//    DESCRIPTION :
//       This module generated decoder enable signals. This is generated by
//       comparing instruction address with address defined by parameter.
//----------------------------------------------------------------------
//    LOCAL PARAMETERS:
//
//    HIGH
//       This is 1 bit one value
//
//    LOW
//       This is 1 bit zero value
//
//    ONE
//       This is number 1 to and is declared just to avoid lint warnings
//
//    IRDECODER_STAP_SIZE_OF_POLICY_OPCODE
//       This parameter specifies MSB STAP_SIZE_OF_EACH_INSTRUCTION number of 
//       bits for address opcodes and concatinated with LSB 2 bits for 
//       security color code.
//----------------------------------------------------------------------
module stap_irdecoder
   #(
   parameter IRDECODER_STAP_SWCOMP_ACTIVE                  = 1,
   parameter IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION       = 8,
   parameter IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS      = 0,
   parameter IRDECODER_STAP_INSTRUCTION_FOR_DATA_REGISTERS = 0,
   parameter IRDECODER_STAP_ADDRESS_OF_CLAMP               = 0,
   parameter IRDECODER_STAP_MINIMUM_SIZEOF_INSTRUCTION     = 0,
   parameter IRDECODER_STAP_ENABLE_BSCAN                   = 0,
   parameter IRDECODER_STAP_SECURE_GREEN                   = 2'b00,
   parameter IRDECODER_STAP_SECURE_ORANGE                  = 2'b01,
   parameter IRDECODER_STAP_SECURE_RED                     = 2'b10
   )
   (
   input  logic                                                    powergood_rst_trst_b, //kbbhagwa cdc fix
   input  logic [(IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  stap_irreg_ireg,
   input  logic [(IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  stap_irreg_ireg_nxt,//kbbhagwa cdc fix
   input  logic                                                    ftap_tck, //kbbhagwa cdc fix
   input  logic                                                    feature_green_en,
   input  logic                                                    feature_orange_en,
   input  logic                                                    feature_red_en,
   input  logic                                                    stap_isol_en_b, //badithya edit for SWCOMP implementation: PCR 1604263740

   output logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] stap_irdecoder_drselect,
   output logic                                                    tap_swcomp_active, //badithya edit for SWCOMP implementation
   output logic                                                    stap_and_all_bits_irreg
   );

   // *********************************************************************
   // Local parameters
   // *********************************************************************
   localparam HIGH                               = 1'b1;
   localparam LOW                                = 1'b0;
   localparam ONE                                = 1;
   localparam IRDECODER_STAP_POSITION_OF_HIGHZ   = 2;
   localparam IRDECODER_STAP_POSITION_OF_SLVIDCODE = (IRDECODER_STAP_ENABLE_BSCAN == 1) ? 4 : 1; //kbbhagwa cdc fix
   localparam IRDECODER_STAP_SIZE_OF_POLICY_OPCODE = IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION + 2;  

   // *********************************************************************
   // Internal signals
   // *********************************************************************
   logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] decoder_drselect;
   logic                                                    decode_clamp;

   logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] irdecoder_drselect_nxt; //kbbhagwa cdc fix
   logic                                                    and_all_bits_irreg_nxt; //kbbhagwa cdc fix

   logic                                                    bypass_enable ; //badithya fix for SWCOMP

   // *********************************************************************
   // Generate construct is used to generate number of decoded output lines
   // which is equal to IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS
   // *********************************************************************
   generate
      for (genvar k = 0; k < IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS; k = k + 1)
      begin:generate_decoder
         stap_decoder #(
                        .DECODER_INSTRUCTION_TO_DECODE
                             (IRDECODER_STAP_INSTRUCTION_FOR_DATA_REGISTERS[
                               ((IRDECODER_STAP_SIZE_OF_POLICY_OPCODE + 
                                (IRDECODER_STAP_SIZE_OF_POLICY_OPCODE * k)) - 1) :
                               ((IRDECODER_STAP_SIZE_OF_POLICY_OPCODE * k) + 2)]),
                        .DECODER_STAP_SIZE_OF_EACH_INSTRUCTION
                           (IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION),
                        .DECODER_STAP_DFX_SECURE_POLICY_OPCODE
                             (IRDECODER_STAP_INSTRUCTION_FOR_DATA_REGISTERS[
                                (((IRDECODER_STAP_SIZE_OF_POLICY_OPCODE + 
                                  (IRDECODER_STAP_SIZE_OF_POLICY_OPCODE * k)) -
                                   IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION) - 1) :
                                  (IRDECODER_STAP_SIZE_OF_POLICY_OPCODE * k)]),
                        .DECODER_STAP_SECURE_GREEN  (IRDECODER_STAP_SECURE_GREEN),
                        .DECODER_STAP_SECURE_ORANGE (IRDECODER_STAP_SECURE_ORANGE),
                        .DECODER_STAP_SECURE_RED    (IRDECODER_STAP_SECURE_RED)
                       )
         i_stap_decoder (
                         .stap_irreg_ireg  (stap_irreg_ireg_nxt), //kbbhagwa cdc fix
                         .decoder_drselect (decoder_drselect[k]),
                         .feature_green_en (feature_green_en),
                         .feature_orange_en(feature_orange_en),
                         .feature_red_en   (feature_red_en)
                        );
      end
   endgenerate

always_ff @(negedge ftap_tck or negedge powergood_rst_trst_b)
  if (~ powergood_rst_trst_b)
      for (integer count = 0; count <= (IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1); count++)
      begin
         if (count == IRDECODER_STAP_POSITION_OF_SLVIDCODE)
             stap_irdecoder_drselect[IRDECODER_STAP_POSITION_OF_SLVIDCODE] <= 1'b1;
         else
             stap_irdecoder_drselect[count] <= 1'b0;
      end
  else
      stap_irdecoder_drselect <= irdecoder_drselect_nxt;

   // *********************************************************************
   // Decoding of some of the Instructions
   // *********************************************************************
   assign stap_and_all_bits_irreg = &(stap_irreg_ireg);
   assign and_all_bits_irreg_nxt  = &(stap_irreg_ireg_nxt) | bypass_enable ; //kbbhagwa cdc fix //badithya fix for making IRREG go to bypass whenever bypass_enable is 1. 

   assign decode_clamp = (stap_irreg_ireg_nxt == IRDECODER_STAP_ADDRESS_OF_CLAMP) ? HIGH : LOW;

   generate
     if(IRDECODER_STAP_SWCOMP_ACTIVE == 1)
     begin:generate_enable

//      always_comb begin
//            if(((stap_irreg_ireg == 'h20) | (stap_irreg_ireg == 'h21))  && (stap_isol_en_b == 1'b0) ) //Whenever SWCOMP registers are selected and SWCOMP is powered down, bypass register should be selected.
//            begin
//                bypass_enable = 1'b1;
//            end
//            else
//            begin 
//                bypass_enable = 1'b0;
//            end
//        
//            if(bypass_enable == 1'b0)  // Whenever bypass enable = 0 and SWCOMP registers are selected, tap_swcomp_active should be high
//              begin
//               if((stap_irreg_ireg == 'h20 | stap_irreg_ireg == 'h21))
//                   tap_swcomp_active = 1'b1;
//               else
//                   tap_swcomp_active = 1'b0;
//              end
//            else 
//            begin
//                   tap_swcomp_active = 1'b1 ;
//            end 
//          end
//
  always_comb begin
	  if(stap_isol_en_b == 1'b0)
	  begin
          if((stap_irreg_ireg == 'h20) | (stap_irreg_ireg == 'h21))
			  begin
                   bypass_enable = 1'b1;
                   tap_swcomp_active = 1'b1;
		      end
         else 
		      begin
                   bypass_enable = 1'b0;
                   tap_swcomp_active = 1'b1;
		      end
	  end
	  else
	  begin
          if((stap_irreg_ireg == 'h20) | (stap_irreg_ireg == 'h21))
			  begin
                   bypass_enable = 1'b0;
                  tap_swcomp_active = 1'b1;
			  end
          else
              begin
                   bypass_enable = 1'b0;
				  tap_swcomp_active = 1'b0;
			  end    
      end
  end
		  
     end
     else
     begin:generate_enable
        assign  bypass_enable = 1'b0;
        assign  tap_swcomp_active = 1'b1;
     end
     endgenerate


   generate
      if (IRDECODER_STAP_ENABLE_BSCAN == 1)
      begin:generate_irdec
         assign irdecoder_drselect_nxt = (and_all_bits_irreg_nxt == HIGH) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} : (decode_clamp == HIGH) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} :
            (decoder_drselect == {IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS{LOW}}) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} :
            (decoder_drselect[IRDECODER_STAP_POSITION_OF_HIGHZ] == HIGH) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} : decoder_drselect;
      end
      else
      begin:generate_irdec
         assign irdecoder_drselect_nxt = (and_all_bits_irreg_nxt == HIGH) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} :
            (decoder_drselect == {IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS{LOW}}) ?
            {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH} : decoder_drselect;

   end
   endgenerate

endmodule
