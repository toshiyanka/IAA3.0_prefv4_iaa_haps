module ctech_lib_msff_meta_hard (o,d,clk);
   input logic d,clk;
   output logic o;
   d04hgn10ld0b0 ctech_lib_dcszo (.clk(clk), .d(d), .o(o));
endmodule
