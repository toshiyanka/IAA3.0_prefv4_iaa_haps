mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dir_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_rop_dp_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_dir.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_dqed.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_dir.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_dp_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rop_dp_enq_ro.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_rfw.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_pgcb_rfw.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_wu_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_dir_tok_lim_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_tok_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_enq_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atq_enqueue_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_inflight_limit_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2priov_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_replay_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_aqed_active_limit_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dir_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_max_depth_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_dir_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_1_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_inflight_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_atm_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_atm_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_uno_atm_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_sel_nalb_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq2qid_0_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_ldb_token_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_aqed_lsp_deq_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_ldb_token_rtn_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_atm_active_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_aqed_active_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_dir_max_depth_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_qid_ldb_replay_count_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_nalb_qid_dpth_thrsh_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_rw_cfg_cq_ldb_token_depth_select_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_nalb_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_list_sel_pipe_rfw.i_rf_cq_nalb_pri_arbindex_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_nalb_qed_data.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_rx_sync_dp_dqed_data.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_rfw.i_rf_qed_chp_sch_data.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_srw.i_sr_nalb_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_0.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_7.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_5.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_2.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_3.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_1.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_6.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_qed_pipe_srw.i_sr_qed_4.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_unoord.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_unoord.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_tp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_lsp_enq_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_qed.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rofrag_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_replay_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_nalb_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_atq_hp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rx_sync_rop_nalb_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_rop_nalb_enq_ro.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_nalb_pipe_rfw.i_rf_lsp_nalb_sch_unoord.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_6.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_hist_list.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_4.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_0.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_7.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_5.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_3.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_2.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_srw.i_sr_freelist_1.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hcw_enq_w_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_depth.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_tok_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_outbound_hcw_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_hist_list_minmax.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_hist_list_ptr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_wptr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_wptr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_to_cq_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_intr_thresh.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ord_qid_sn_map.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_dir_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_cmp_id_chk_enbl_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_dir_cq_depth.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_ldb_cq_token_depth_select.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_count_rmw_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_aqed_chp_sch_rx_sync_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_qed_chp_sch_rx_sync_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_credit_hist_pipe_rfw.i_rf_rw_threshold_r_pipe_ldb_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b2.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b3.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_qed_pipe.i_hqm_dir_pipe_srw.i_sr_dir_nxthp.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rx_sync_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_freelist_return.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_qid_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_qed_aqed_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_rw_aqed_qid_fid_limit.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fid_cnt.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_cnt_pri1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_fifo_aqed_chp_sch.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_rfw.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_phdr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_nphdr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_npdata.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_pdata_rxq.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ph_req_fifo.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_ri_tlq_fifo_pdata.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_rfw.i_iosf_rf_cpldata_rxq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_aqed_ap_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_lsp_enq.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b2.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin3.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin3.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rlst_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_atm_fifo_ap_aqed.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b3.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_rw_aqed_qid2cqidix.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin3.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin3.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_slst_cnt.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hp_bin2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_tp_bin0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_fid2cqqidix.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_sch_cnt_dup1.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_tp_bin1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_qid_rdylst_clamp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_schlst_hp_bin2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_lsp_atm_pipe_rfw.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_st_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbtp_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_ldb_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirhp_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_cnt_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_lbhp_mem.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_lsp_reordercmp_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_dir_rply_req_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn0_order_shft_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_ordered_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_reord_dirtp_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn_complete_fifo_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_sn1_order_shft_mem.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_reorder_pipe_rfw.i_rf_chp_rop_hcw_fifo_mem.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_pd_fifo.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.hqm_system_aon_wrap.i_hqm_iosf_dc_rfw.i_ti_trn_ph_fifo.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_dc_rfw.i_hcw_enq_fifo.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_l.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_u.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_pasid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b1.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_pp2vas.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_data.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid2qid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp2pp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_isr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vpp2pp.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vpp_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_data.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_isr.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_ldb_wb0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_ldb_vqid_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd0.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_ai_addr_u.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_qid2vqid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_pasid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_vasqid_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_dir_wb1.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_alarm_vf_synd2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_addr_u.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_sch_out_fifo.i_rf_b0.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_vasqid_v.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq2vf_pf.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_msix_tbl_word2.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_vf_dir_vqid2qid.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_dir_cq_addr_l.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_cq_ai_addr_l.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_rf_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_rfw.i_lut_ldb_pp2vas.i_rf.FUSE_MISC_RF_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_system.i_hqm_system_srw.i_system_csr_ram0.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_freelist.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed_ll_qe_hpnxt.i_sram.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b1.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b0.FUSE_MISC_SSA_IN[19]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[0]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[0]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[1]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[1]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[2]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[2]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[3]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[3]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[4]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[4]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[5]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[5]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[6]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[6]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[9]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[9]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[10]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[10]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[11]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[11]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[12]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[12]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[13]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[13]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[14]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[14]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[15]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[15]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[16]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[16]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[17]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[17]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[18]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[18]");
mem_trim_fuse_ip_bit_q.push_back("hqm_tb_top.u_hqm.fary_ffuse_ssa_trim[19]");
mem_trim_fuse_op_bit_q.push_back("hqm_tb_top.u_hqm.par_hqm_list_sel_pipe.i_hqm_aqed_pipe_srw.i_sr_aqed.i_sram_b2.FUSE_MISC_SSA_IN[19]");
