// File output was printed on: Saturday, January 19, 2013 2:59:29 PM
// Chassis TAP Tool version: 0.6.0.0
//----------------------------------------------------------------------
// ENUM DECLARATIONS
//------------------------------------------------------------------------
typedef enum int {
   IPLEVEL_STAP   =  'd0,
   NOTAP          =  'hFFFF_FFFF
} Tap_t;


