VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf028b032e2r2w0cbbehraa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf028b032e2r2w0cbbehraa4acw 0 0 ;
  SIZE 18 BY 20.16 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 3.24 0.388 4.44 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 3.24 2.916 4.44 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 0.84 0.388 2.04 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 0.84 3.172 2.04 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 3.24 1.628 4.44 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 3.24 1.928 4.44 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 3.24 2.188 4.44 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 3.24 2.356 4.44 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.24 2.616 4.44 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 3.24 0.556 4.44 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 3.24 0.816 4.44 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 3.24 4.156 4.44 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 3.24 4.416 4.44 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 3.24 4.716 4.44 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 3.24 4.972 4.44 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 3.24 5.228 4.44 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 3.24 3.172 4.44 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 3.24 3.428 4.44 ;
    END
  END rdaddrp1_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 5.16 5.956 6.36 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 9.96 5.616 11.16 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 9.96 5.788 11.16 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 10.92 5.316 12.12 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 10.92 5.528 12.12 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 11.88 6.856 13.08 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 11.88 7.028 13.08 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 12.84 6.428 14.04 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 12.84 6.516 14.04 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 13.8 5.788 15 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 13.8 5.872 15 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 5.16 6.128 6.36 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 14.76 5.316 15.96 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 14.76 5.528 15.96 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 15.72 6.856 16.92 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 15.72 7.028 16.92 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 16.68 6.428 17.88 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 16.68 6.516 17.88 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 17.64 5.788 18.84 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 17.64 5.872 18.84 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 18.6 5.316 19.8 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 18.6 5.528 19.8 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 6.12 5.528 7.32 ;
    END
  END rddatap0[2]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 6.12 5.616 7.32 ;
    END
  END rddatap0[3]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 7.08 7.028 8.28 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 7.08 5.316 8.28 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 8.04 6.688 9.24 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 8.04 6.772 9.24 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 9 6.128 10.2 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 9 6.216 10.2 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 5.16 6.216 6.36 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 9.96 5.872 11.16 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 9.96 5.956 11.16 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 10.92 6.128 12.12 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 10.92 6.216 12.12 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 11.88 5.616 13.08 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 11.88 5.788 13.08 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 12.84 6.688 14.04 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 12.84 6.772 14.04 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 13.8 5.956 15 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 13.8 6.128 15 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 5.16 6.428 6.36 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 14.76 5.616 15.96 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 14.76 6.216 15.96 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 15.72 5.788 16.92 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 15.72 5.872 16.92 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 16.68 6.688 17.88 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 16.68 6.772 17.88 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 17.64 5.956 18.84 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 17.64 6.128 18.84 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 18.6 5.616 19.8 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 18.6 6.216 19.8 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 6.12 5.788 7.32 ;
    END
  END rddatap1[2]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 6.12 5.872 7.32 ;
    END
  END rddatap1[3]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 7.08 5.956 8.28 ;
    END
  END rddatap1[4]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 7.08 6.128 8.28 ;
    END
  END rddatap1[5]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 8.04 6.856 9.24 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 8.04 5.528 9.24 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 9 6.428 10.2 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 9 6.516 10.2 ;
    END
  END rddatap1[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 3.24 1.116 4.44 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.24 3.728 4.44 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 3.24 1.372 4.44 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 3.24 3.988 4.44 ;
    END
  END sdl_initp1
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 17.062 0.06 17.138 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.262 0.06 15.338 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 20.1 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 16.162 0.06 16.238 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.362 0.06 14.438 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 20.1 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 20.1 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.84 1.928 2.04 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 0.84 2.188 2.04 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 0.84 2.356 2.04 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 0.84 2.616 2.04 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.84 2.916 2.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 0.84 0.556 2.04 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 0.84 0.816 2.04 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 0.84 4.716 2.04 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 0.84 4.972 2.04 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 0.84 5.228 2.04 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 0.84 5.528 2.04 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 0.84 5.788 2.04 ;
    END
  END wraddrp1[4]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.84 3.428 2.04 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.84 3.728 2.04 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 5.16 3.256 6.36 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 9.96 4.888 11.16 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 9.96 4.972 11.16 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 10.92 4.156 12.12 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 10.92 4.328 12.12 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 11.88 3.728 13.08 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 11.88 3.816 13.08 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 12.84 3.428 14.04 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.84 3.516 14.04 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 13.8 4.972 15 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 13.8 3.172 15 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.16 3.516 6.36 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 14.76 4.416 15.96 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 14.76 4.628 15.96 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 15.72 3.728 16.92 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 15.72 3.816 16.92 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.68 3.428 17.88 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.68 3.516 17.88 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 17.64 4.972 18.84 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 17.64 3.172 18.84 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 18.6 4.416 19.8 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 18.6 4.628 19.8 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 6.12 4.716 7.32 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 6.12 4.888 7.32 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 7.08 3.988 8.28 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 7.08 4.072 8.28 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.04 3.516 9.24 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 8.04 3.728 9.24 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 9 3.256 10.2 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9 3.428 10.2 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 0.84 1.372 2.04 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 0.84 1.628 2.04 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 5.16 3.816 6.36 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 9.96 3.172 11.16 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 9.96 3.516 11.16 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 10.92 4.416 12.12 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 10.92 4.628 12.12 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 11.88 3.988 13.08 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 11.88 4.072 13.08 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 12.84 4.156 14.04 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 12.84 4.328 14.04 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 13.8 3.256 15 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 13.8 3.728 15 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 5.16 4.072 6.36 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 14.76 4.716 15.96 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 14.76 4.888 15.96 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 15.72 3.988 16.92 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 15.72 4.072 16.92 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 16.68 4.156 17.88 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 16.68 4.328 17.88 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 17.64 3.256 18.84 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 17.64 3.728 18.84 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 18.6 4.716 19.8 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 18.6 4.888 19.8 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 6.12 4.972 7.32 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 6.12 3.172 7.32 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 7.08 4.156 8.28 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 7.08 4.328 8.28 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 8.04 3.816 9.24 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 8.04 4.416 9.24 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 9 3.988 10.2 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 9 4.072 10.2 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 0.84 4.156 2.04 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 0.84 4.416 2.04 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 0.84 1.116 2.04 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 0.84 3.988 2.04 ;
    END
  END wrenp1
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 18 20.16 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 18 20.16 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 18.0705 20.198 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 18.035 20.23 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 18.07 20.198 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 18.059 20.25 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 18.09 20.222 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 18.092 20.22 ;
  END
END arf028b032e2r2w0cbbehraa4acw
END LIBRARY
