module ctech_lib_msff_clkb (
   input logic clkb,
   input logic d,
   output logic o
);
   d04fkn80ld0b0 ctech_lib_dcszo (.clkb(clkb), .d(d), .o(o));
endmodule
