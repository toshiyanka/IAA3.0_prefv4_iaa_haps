VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO ip764hduspsr1024x52m4b2s0r2p0d0
  CLASS BLOCK ;
  FIXEDMASK ;
  FOREIGN ip764hduspsr1024x52m4b2s0r2p0d0 ;
  ORIGIN 0 0 ;
  SIZE 36.3 BY 72.72 ;
  SYMMETRY X Y ;
  SITE ip764hduspsr1024x52m4b2s0r2p0d0 ;
  PIN adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.344 34.902 17.384 34.938 ;
      LAYER m5 ;
        RECT 17.344 34.18 17.384 35.14 ;
    END
  END adr[0]
  PIN adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.48 34.6005 17.52 34.6365 ;
      LAYER m5 ;
        RECT 17.48 34.3 17.52 35.26 ;
    END
  END adr[1]
  PIN adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.48 34.0035 17.52 34.0395 ;
      LAYER m5 ;
        RECT 17.48 33.3 17.52 34.26 ;
    END
  END adr[2]
  PIN adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 34.902 17.176 34.938 ;
      LAYER m5 ;
        RECT 17.136 34.3 17.176 35.26 ;
    END
  END adr[3]
  PIN adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.284 33.942 18.328 33.978 ;
      LAYER m5 ;
        RECT 18.284 33.18 18.328 34.14 ;
    END
  END adr[4]
  PIN adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 33.942 17.176 33.978 ;
      LAYER m5 ;
        RECT 17.136 33.3 17.176 34.26 ;
    END
  END adr[5]
  PIN adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.944 33.222 17.984 33.258 ;
      LAYER m5 ;
        RECT 17.944 33.18 17.984 34.14 ;
    END
  END adr[6]
  PIN adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.284 34.902 18.328 34.938 ;
      LAYER m5 ;
        RECT 18.284 34.18 18.328 35.14 ;
    END
  END adr[7]
  PIN adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.272 34.2435 17.316 34.2795 ;
      LAYER m5 ;
        RECT 17.272 34.18 17.316 35.14 ;
    END
  END adr[8]
  PIN adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.616 34.3605 17.656 34.3965 ;
      LAYER m5 ;
        RECT 17.616 34.18 17.656 35.14 ;
    END
  END adr[9]
  PIN arysleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.344 32.2005 17.384 32.2365 ;
      LAYER m5 ;
        RECT 17.344 32.18 17.384 33.14 ;
    END
  END arysleep
  PIN async_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.616 32.3235 17.656 32.3595 ;
      LAYER m5 ;
        RECT 17.616 32.18 17.656 33.14 ;
    END
  END async_reset
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 36.342 17.176 36.378 ;
      LAYER m5 ;
        RECT 17.136 35.85 17.176 36.81 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 1.558 17.452 1.594 ;
      LAYER m5 ;
        RECT 17.412 0.62 17.452 1.78 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 13.558 17.452 13.594 ;
      LAYER m5 ;
        RECT 17.412 12.62 17.452 13.78 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 14.758 17.452 14.794 ;
      LAYER m5 ;
        RECT 17.412 13.82 17.452 14.98 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 15.958 17.452 15.994 ;
      LAYER m5 ;
        RECT 17.412 15.02 17.452 16.18 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 17.158 17.452 17.194 ;
      LAYER m5 ;
        RECT 17.412 16.22 17.452 17.38 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 18.358 17.452 18.394 ;
      LAYER m5 ;
        RECT 17.412 17.42 17.452 18.58 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 19.558 17.452 19.594 ;
      LAYER m5 ;
        RECT 17.412 18.62 17.452 19.78 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 20.758 17.452 20.794 ;
      LAYER m5 ;
        RECT 17.412 19.82 17.452 20.98 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 21.958 17.452 21.994 ;
      LAYER m5 ;
        RECT 17.412 21.02 17.452 22.18 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 23.158 17.452 23.194 ;
      LAYER m5 ;
        RECT 17.412 22.22 17.452 23.38 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 24.358 17.452 24.394 ;
      LAYER m5 ;
        RECT 17.412 23.42 17.452 24.58 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 2.758 17.452 2.794 ;
      LAYER m5 ;
        RECT 17.412 1.82 17.452 2.98 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 25.558 17.452 25.594 ;
      LAYER m5 ;
        RECT 17.412 24.62 17.452 25.78 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 26.758 17.452 26.794 ;
      LAYER m5 ;
        RECT 17.412 25.82 17.452 26.98 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 27.958 17.452 27.994 ;
      LAYER m5 ;
        RECT 17.412 27.02 17.452 28.18 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 29.158 17.452 29.194 ;
      LAYER m5 ;
        RECT 17.412 28.22 17.452 29.38 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 30.358 17.452 30.394 ;
      LAYER m5 ;
        RECT 17.412 29.42 17.452 30.58 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 31.558 17.452 31.594 ;
      LAYER m5 ;
        RECT 17.412 30.62 17.452 31.78 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 40.678 17.452 40.714 ;
      LAYER m5 ;
        RECT 17.412 39.74 17.452 40.9 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 41.878 17.452 41.914 ;
      LAYER m5 ;
        RECT 17.412 40.94 17.452 42.1 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 43.078 17.452 43.114 ;
      LAYER m5 ;
        RECT 17.412 42.14 17.452 43.3 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 44.278 17.452 44.314 ;
      LAYER m5 ;
        RECT 17.412 43.34 17.452 44.5 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 3.958 17.452 3.994 ;
      LAYER m5 ;
        RECT 17.412 3.02 17.452 4.18 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 45.478 17.452 45.514 ;
      LAYER m5 ;
        RECT 17.412 44.54 17.452 45.7 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 46.678 17.452 46.714 ;
      LAYER m5 ;
        RECT 17.412 45.74 17.452 46.9 ;
    END
  END din[31]
  PIN din[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 47.878 17.452 47.914 ;
      LAYER m5 ;
        RECT 17.412 46.94 17.452 48.1 ;
    END
  END din[32]
  PIN din[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 49.078 17.452 49.114 ;
      LAYER m5 ;
        RECT 17.412 48.14 17.452 49.3 ;
    END
  END din[33]
  PIN din[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 50.278 17.452 50.314 ;
      LAYER m5 ;
        RECT 17.412 49.34 17.452 50.5 ;
    END
  END din[34]
  PIN din[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 51.478 17.452 51.514 ;
      LAYER m5 ;
        RECT 17.412 50.54 17.452 51.7 ;
    END
  END din[35]
  PIN din[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 52.678 17.452 52.714 ;
      LAYER m5 ;
        RECT 17.412 51.74 17.452 52.9 ;
    END
  END din[36]
  PIN din[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 53.878 17.452 53.914 ;
      LAYER m5 ;
        RECT 17.412 52.94 17.452 54.1 ;
    END
  END din[37]
  PIN din[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 55.078 17.452 55.114 ;
      LAYER m5 ;
        RECT 17.412 54.14 17.452 55.3 ;
    END
  END din[38]
  PIN din[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 56.278 17.452 56.314 ;
      LAYER m5 ;
        RECT 17.412 55.34 17.452 56.5 ;
    END
  END din[39]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 5.158 17.452 5.194 ;
      LAYER m5 ;
        RECT 17.412 4.22 17.452 5.38 ;
    END
  END din[3]
  PIN din[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 57.478 17.452 57.514 ;
      LAYER m5 ;
        RECT 17.412 56.54 17.452 57.7 ;
    END
  END din[40]
  PIN din[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 58.678 17.452 58.714 ;
      LAYER m5 ;
        RECT 17.412 57.74 17.452 58.9 ;
    END
  END din[41]
  PIN din[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 59.878 17.452 59.914 ;
      LAYER m5 ;
        RECT 17.412 58.94 17.452 60.1 ;
    END
  END din[42]
  PIN din[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 61.078 17.452 61.114 ;
      LAYER m5 ;
        RECT 17.412 60.14 17.452 61.3 ;
    END
  END din[43]
  PIN din[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 62.278 17.452 62.314 ;
      LAYER m5 ;
        RECT 17.412 61.34 17.452 62.5 ;
    END
  END din[44]
  PIN din[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 63.478 17.452 63.514 ;
      LAYER m5 ;
        RECT 17.412 62.54 17.452 63.7 ;
    END
  END din[45]
  PIN din[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 64.678 17.452 64.714 ;
      LAYER m5 ;
        RECT 17.412 63.74 17.452 64.9 ;
    END
  END din[46]
  PIN din[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 65.878 17.452 65.914 ;
      LAYER m5 ;
        RECT 17.412 64.94 17.452 66.1 ;
    END
  END din[47]
  PIN din[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 67.078 17.452 67.114 ;
      LAYER m5 ;
        RECT 17.412 66.14 17.452 67.3 ;
    END
  END din[48]
  PIN din[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 68.278 17.452 68.314 ;
      LAYER m5 ;
        RECT 17.412 67.34 17.452 68.5 ;
    END
  END din[49]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 6.358 17.452 6.394 ;
      LAYER m5 ;
        RECT 17.412 5.42 17.452 6.58 ;
    END
  END din[4]
  PIN din[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 69.478 17.452 69.514 ;
      LAYER m5 ;
        RECT 17.412 68.54 17.452 69.7 ;
    END
  END din[50]
  PIN din[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 70.678 17.452 70.714 ;
      LAYER m5 ;
        RECT 17.412 69.74 17.452 70.9 ;
    END
  END din[51]
  PIN din[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 71.878 17.452 71.914 ;
      LAYER m5 ;
        RECT 17.412 70.94 17.452 72.1 ;
    END
  END din[52]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 7.558 17.452 7.594 ;
      LAYER m5 ;
        RECT 17.412 6.62 17.452 7.78 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 8.758 17.452 8.794 ;
      LAYER m5 ;
        RECT 17.412 7.82 17.452 8.98 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 9.958 17.452 9.994 ;
      LAYER m5 ;
        RECT 17.412 9.02 17.452 10.18 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 11.158 17.452 11.194 ;
      LAYER m5 ;
        RECT 17.412 10.22 17.452 11.38 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.412 12.358 17.452 12.394 ;
      LAYER m5 ;
        RECT 17.412 11.42 17.452 12.58 ;
    END
  END din[9]
  PIN mce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 38.022 17.176 38.058 ;
      LAYER m5 ;
        RECT 17.136 37.85 17.176 38.81 ;
    END
  END mce
  PIN ra[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.424 37.7205 18.464 37.7565 ;
      LAYER m5 ;
        RECT 18.424 36.85 18.464 37.81 ;
    END
  END ra[0]
  PIN ra[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.012 37.542 18.052 37.578 ;
      LAYER m5 ;
        RECT 18.012 36.85 18.052 37.81 ;
    END
  END ra[1]
  PIN redrowen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.616 36.102 17.656 36.138 ;
      LAYER m5 ;
        RECT 17.616 35.85 17.656 36.81 ;
    END
  END redrowen[0]
  PIN redrowen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.012 33.462 18.052 33.498 ;
      LAYER m5 ;
        RECT 18.012 33.18 18.052 34.14 ;
    END
  END redrowen[1]
  PIN ren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.064 34.422 17.108 34.458 ;
      LAYER m5 ;
        RECT 17.064 34.18 17.108 35.14 ;
    END
  END ren
  PIN rmce[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.616 38.502 17.656 38.538 ;
      LAYER m5 ;
        RECT 17.616 37.85 17.656 38.81 ;
    END
  END rmce[0]
  PIN rmce[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.548 38.2005 17.588 38.2365 ;
      LAYER m5 ;
        RECT 17.548 37.85 17.588 38.81 ;
    END
  END rmce[1]
  PIN rmce[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.344 37.9605 17.384 37.9965 ;
      LAYER m5 ;
        RECT 17.344 37.85 17.384 38.81 ;
    END
  END rmce[2]
  PIN rmce[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.48 38.3235 17.52 38.3595 ;
      LAYER m5 ;
        RECT 17.48 37.97 17.52 38.93 ;
    END
  END rmce[3]
  PIN sbc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.284 32.262 18.328 32.298 ;
      LAYER m5 ;
        RECT 18.284 32.18 18.328 33.14 ;
    END
  END sbc[0]
  PIN sbc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.548 32.4405 17.588 32.4765 ;
      LAYER m5 ;
        RECT 17.548 32.18 17.588 33.14 ;
    END
  END sbc[1]
  PIN stbyp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.012 34.662 18.052 34.698 ;
      LAYER m5 ;
        RECT 18.012 34.18 18.052 35.14 ;
    END
  END stbyp
  PIN wa[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.616 37.302 17.656 37.338 ;
      LAYER m5 ;
        RECT 17.616 36.85 17.656 37.81 ;
    END
  END wa[0]
  PIN wa[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.344 36.342 17.384 36.378 ;
      LAYER m5 ;
        RECT 17.344 35.85 17.384 36.81 ;
    END
  END wa[1]
  PIN wa[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 18.08 36.8835 18.12 36.9195 ;
      LAYER m5 ;
        RECT 18.08 36.85 18.12 37.81 ;
    END
  END wa[2]
  PIN wen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.272 33.7635 17.316 33.7995 ;
      LAYER m5 ;
        RECT 17.272 33.18 17.316 34.14 ;
    END
  END wen
  PIN wmce[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.48 37.3635 17.52 37.3995 ;
      LAYER m5 ;
        RECT 17.48 36.97 17.52 37.93 ;
    END
  END wmce[0]
  PIN wmce[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.344 36.8835 17.384 36.9195 ;
      LAYER m5 ;
        RECT 17.344 36.85 17.384 37.81 ;
    END
  END wmce[1]
  PIN wpulse[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.548 37.4805 17.588 37.5165 ;
      LAYER m5 ;
        RECT 17.548 36.85 17.588 37.81 ;
    END
  END wpulse[0]
  PIN wpulse[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 37.2405 17.176 37.2765 ;
      LAYER m5 ;
        RECT 17.136 36.85 17.176 37.81 ;
    END
  END wpulse[1]
  PIN wpulse[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.944 37.2405 17.984 37.2765 ;
      LAYER m5 ;
        RECT 17.944 36.85 17.984 37.81 ;
    END
  END wpulse[2]
  PIN q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 1.329 17.176 1.365 ;
      LAYER m5 ;
        RECT 17.136 0.62 17.176 1.78 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 13.329 17.176 13.365 ;
      LAYER m5 ;
        RECT 17.136 12.62 17.176 13.78 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 14.529 17.176 14.565 ;
      LAYER m5 ;
        RECT 17.136 13.82 17.176 14.98 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 15.729 17.176 15.765 ;
      LAYER m5 ;
        RECT 17.136 15.02 17.176 16.18 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 16.929 17.176 16.965 ;
      LAYER m5 ;
        RECT 17.136 16.22 17.176 17.38 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 18.129 17.176 18.165 ;
      LAYER m5 ;
        RECT 17.136 17.42 17.176 18.58 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 19.329 17.176 19.365 ;
      LAYER m5 ;
        RECT 17.136 18.62 17.176 19.78 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 20.529 17.176 20.565 ;
      LAYER m5 ;
        RECT 17.136 19.82 17.176 20.98 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 21.729 17.176 21.765 ;
      LAYER m5 ;
        RECT 17.136 21.02 17.176 22.18 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 22.929 17.176 22.965 ;
      LAYER m5 ;
        RECT 17.136 22.22 17.176 23.38 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 24.129 17.176 24.165 ;
      LAYER m5 ;
        RECT 17.136 23.42 17.176 24.58 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 2.529 17.176 2.565 ;
      LAYER m5 ;
        RECT 17.136 1.82 17.176 2.98 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 25.329 17.176 25.365 ;
      LAYER m5 ;
        RECT 17.136 24.62 17.176 25.78 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 26.529 17.176 26.565 ;
      LAYER m5 ;
        RECT 17.136 25.82 17.176 26.98 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 27.729 17.176 27.765 ;
      LAYER m5 ;
        RECT 17.136 27.02 17.176 28.18 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 28.929 17.176 28.965 ;
      LAYER m5 ;
        RECT 17.136 28.22 17.176 29.38 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 30.129 17.176 30.165 ;
      LAYER m5 ;
        RECT 17.136 29.42 17.176 30.58 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 31.329 17.176 31.365 ;
      LAYER m5 ;
        RECT 17.136 30.62 17.176 31.78 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 40.449 17.176 40.485 ;
      LAYER m5 ;
        RECT 17.136 39.74 17.176 40.9 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 41.649 17.176 41.685 ;
      LAYER m5 ;
        RECT 17.136 40.94 17.176 42.1 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 42.849 17.176 42.885 ;
      LAYER m5 ;
        RECT 17.136 42.14 17.176 43.3 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 44.049 17.176 44.085 ;
      LAYER m5 ;
        RECT 17.136 43.34 17.176 44.5 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 3.729 17.176 3.765 ;
      LAYER m5 ;
        RECT 17.136 3.02 17.176 4.18 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 45.249 17.176 45.285 ;
      LAYER m5 ;
        RECT 17.136 44.54 17.176 45.7 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 46.449 17.176 46.485 ;
      LAYER m5 ;
        RECT 17.136 45.74 17.176 46.9 ;
    END
  END q[31]
  PIN q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 47.649 17.176 47.685 ;
      LAYER m5 ;
        RECT 17.136 46.94 17.176 48.1 ;
    END
  END q[32]
  PIN q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 48.849 17.176 48.885 ;
      LAYER m5 ;
        RECT 17.136 48.14 17.176 49.3 ;
    END
  END q[33]
  PIN q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 50.049 17.176 50.085 ;
      LAYER m5 ;
        RECT 17.136 49.34 17.176 50.5 ;
    END
  END q[34]
  PIN q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 51.249 17.176 51.285 ;
      LAYER m5 ;
        RECT 17.136 50.54 17.176 51.7 ;
    END
  END q[35]
  PIN q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 52.449 17.176 52.485 ;
      LAYER m5 ;
        RECT 17.136 51.74 17.176 52.9 ;
    END
  END q[36]
  PIN q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 53.649 17.176 53.685 ;
      LAYER m5 ;
        RECT 17.136 52.94 17.176 54.1 ;
    END
  END q[37]
  PIN q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 54.849 17.176 54.885 ;
      LAYER m5 ;
        RECT 17.136 54.14 17.176 55.3 ;
    END
  END q[38]
  PIN q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 56.049 17.176 56.085 ;
      LAYER m5 ;
        RECT 17.136 55.34 17.176 56.5 ;
    END
  END q[39]
  PIN q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 4.929 17.176 4.965 ;
      LAYER m5 ;
        RECT 17.136 4.22 17.176 5.38 ;
    END
  END q[3]
  PIN q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 57.249 17.176 57.285 ;
      LAYER m5 ;
        RECT 17.136 56.54 17.176 57.7 ;
    END
  END q[40]
  PIN q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 58.449 17.176 58.485 ;
      LAYER m5 ;
        RECT 17.136 57.74 17.176 58.9 ;
    END
  END q[41]
  PIN q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 59.649 17.176 59.685 ;
      LAYER m5 ;
        RECT 17.136 58.94 17.176 60.1 ;
    END
  END q[42]
  PIN q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 60.849 17.176 60.885 ;
      LAYER m5 ;
        RECT 17.136 60.14 17.176 61.3 ;
    END
  END q[43]
  PIN q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 62.049 17.176 62.085 ;
      LAYER m5 ;
        RECT 17.136 61.34 17.176 62.5 ;
    END
  END q[44]
  PIN q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 63.249 17.176 63.285 ;
      LAYER m5 ;
        RECT 17.136 62.54 17.176 63.7 ;
    END
  END q[45]
  PIN q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 64.449 17.176 64.485 ;
      LAYER m5 ;
        RECT 17.136 63.74 17.176 64.9 ;
    END
  END q[46]
  PIN q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 65.649 17.176 65.685 ;
      LAYER m5 ;
        RECT 17.136 64.94 17.176 66.1 ;
    END
  END q[47]
  PIN q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 66.849 17.176 66.885 ;
      LAYER m5 ;
        RECT 17.136 66.14 17.176 67.3 ;
    END
  END q[48]
  PIN q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 68.049 17.176 68.085 ;
      LAYER m5 ;
        RECT 17.136 67.34 17.176 68.5 ;
    END
  END q[49]
  PIN q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 6.129 17.176 6.165 ;
      LAYER m5 ;
        RECT 17.136 5.42 17.176 6.58 ;
    END
  END q[4]
  PIN q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 69.249 17.176 69.285 ;
      LAYER m5 ;
        RECT 17.136 68.54 17.176 69.7 ;
    END
  END q[50]
  PIN q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 70.449 17.176 70.485 ;
      LAYER m5 ;
        RECT 17.136 69.74 17.176 70.9 ;
    END
  END q[51]
  PIN q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 71.649 17.176 71.685 ;
      LAYER m5 ;
        RECT 17.136 70.94 17.176 72.1 ;
    END
  END q[52]
  PIN q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 7.329 17.176 7.365 ;
      LAYER m5 ;
        RECT 17.136 6.62 17.176 7.78 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 8.529 17.176 8.565 ;
      LAYER m5 ;
        RECT 17.136 7.82 17.176 8.98 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 9.729 17.176 9.765 ;
      LAYER m5 ;
        RECT 17.136 9.02 17.176 10.18 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 10.929 17.176 10.965 ;
      LAYER m5 ;
        RECT 17.136 10.22 17.176 11.38 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER v4 ;
        RECT 17.136 12.129 17.176 12.165 ;
      LAYER m5 ;
        RECT 17.136 11.42 17.176 12.58 ;
    END
  END q[9]
  PIN vddp
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER v4 ;
        RECT 16.964 0.7345 17.036 0.7595 ;
        RECT 17.844 0.7345 17.916 0.7595 ;
        RECT 18.664 0.7345 18.736 0.7595 ;
        RECT 18.964 0.7345 19.036 0.7595 ;
        RECT 14.05 0.729 14.104 0.765 ;
        RECT 14.932 0.729 14.986 0.765 ;
        RECT 15.318 0.729 15.37 0.765 ;
        RECT 15.478 0.729 15.53 0.765 ;
        RECT 15.874 0.729 15.926 0.765 ;
        RECT 16.034 0.729 16.086 0.765 ;
        RECT 16.8 0.729 16.854 0.765 ;
        RECT 18.148 0.729 18.188 0.765 ;
        RECT 18.356 0.729 18.396 0.765 ;
        RECT 19.914 0.729 19.966 0.765 ;
        RECT 20.074 0.729 20.126 0.765 ;
        RECT 20.47 0.729 20.522 0.765 ;
        RECT 20.63 0.729 20.682 0.765 ;
        RECT 21.014 0.729 21.068 0.765 ;
        RECT 21.896 0.729 21.95 0.765 ;
        RECT 16.964 0.9635 17.036 0.9885 ;
        RECT 18.664 0.9635 18.736 0.9885 ;
        RECT 18.964 0.9635 19.036 0.9885 ;
        RECT 14.05 0.958 14.104 0.994 ;
        RECT 14.296 0.958 14.35 0.994 ;
        RECT 14.932 0.958 14.986 0.994 ;
        RECT 15.318 0.958 15.37 0.994 ;
        RECT 15.478 0.958 15.53 0.994 ;
        RECT 15.874 0.958 15.926 0.994 ;
        RECT 16.034 0.958 16.086 0.994 ;
        RECT 16.8 0.958 16.854 0.994 ;
        RECT 18.148 0.958 18.188 0.994 ;
        RECT 19.914 0.958 19.966 0.994 ;
        RECT 20.074 0.958 20.126 0.994 ;
        RECT 20.47 0.958 20.522 0.994 ;
        RECT 20.63 0.958 20.682 0.994 ;
        RECT 21.014 0.958 21.068 0.994 ;
        RECT 21.65 0.958 21.704 0.994 ;
        RECT 21.896 0.958 21.95 0.994 ;
        RECT 17.844 1.0405 17.916 1.0655 ;
        RECT 18.356 1.035 18.396 1.071 ;
        RECT 16.964 1.4115 17.036 1.4365 ;
        RECT 17.844 1.4115 17.916 1.4365 ;
        RECT 18.964 1.4115 19.036 1.4365 ;
        RECT 14.05 1.406 14.104 1.442 ;
        RECT 14.296 1.406 14.35 1.442 ;
        RECT 14.932 1.406 14.986 1.442 ;
        RECT 15.318 1.406 15.37 1.442 ;
        RECT 15.874 1.406 15.926 1.442 ;
        RECT 16.034 1.406 16.086 1.442 ;
        RECT 18.356 1.406 18.396 1.442 ;
        RECT 19.914 1.406 19.966 1.442 ;
        RECT 20.074 1.406 20.126 1.442 ;
        RECT 20.63 1.406 20.682 1.442 ;
        RECT 21.014 1.406 21.068 1.442 ;
        RECT 21.65 1.406 21.704 1.442 ;
        RECT 21.896 1.406 21.95 1.442 ;
        RECT 17.844 1.5635 17.916 1.5885 ;
        RECT 18.356 1.558 18.396 1.594 ;
        RECT 18.664 1.6405 18.736 1.6655 ;
        RECT 18.964 1.6405 19.036 1.6655 ;
        RECT 14.296 1.635 14.35 1.671 ;
        RECT 14.932 1.635 14.986 1.671 ;
        RECT 15.318 1.635 15.37 1.671 ;
        RECT 15.478 1.635 15.53 1.671 ;
        RECT 15.874 1.635 15.926 1.671 ;
        RECT 18.148 1.635 18.188 1.671 ;
        RECT 20.074 1.635 20.126 1.671 ;
        RECT 20.47 1.635 20.522 1.671 ;
        RECT 20.63 1.635 20.682 1.671 ;
        RECT 21.014 1.635 21.068 1.671 ;
        RECT 21.65 1.635 21.704 1.671 ;
        RECT 16.964 1.9345 17.036 1.9595 ;
        RECT 17.844 1.9345 17.916 1.9595 ;
        RECT 18.664 1.9345 18.736 1.9595 ;
        RECT 18.964 1.9345 19.036 1.9595 ;
        RECT 14.05 1.929 14.104 1.965 ;
        RECT 14.932 1.929 14.986 1.965 ;
        RECT 15.318 1.929 15.37 1.965 ;
        RECT 15.478 1.929 15.53 1.965 ;
        RECT 15.874 1.929 15.926 1.965 ;
        RECT 16.034 1.929 16.086 1.965 ;
        RECT 16.8 1.929 16.854 1.965 ;
        RECT 18.148 1.929 18.188 1.965 ;
        RECT 18.356 1.929 18.396 1.965 ;
        RECT 19.914 1.929 19.966 1.965 ;
        RECT 20.074 1.929 20.126 1.965 ;
        RECT 20.47 1.929 20.522 1.965 ;
        RECT 20.63 1.929 20.682 1.965 ;
        RECT 21.014 1.929 21.068 1.965 ;
        RECT 21.896 1.929 21.95 1.965 ;
        RECT 16.964 2.1635 17.036 2.1885 ;
        RECT 18.664 2.1635 18.736 2.1885 ;
        RECT 18.964 2.1635 19.036 2.1885 ;
        RECT 14.05 2.158 14.104 2.194 ;
        RECT 14.296 2.158 14.35 2.194 ;
        RECT 14.932 2.158 14.986 2.194 ;
        RECT 15.318 2.158 15.37 2.194 ;
        RECT 15.478 2.158 15.53 2.194 ;
        RECT 15.874 2.158 15.926 2.194 ;
        RECT 16.034 2.158 16.086 2.194 ;
        RECT 16.8 2.158 16.854 2.194 ;
        RECT 18.148 2.158 18.188 2.194 ;
        RECT 19.914 2.158 19.966 2.194 ;
        RECT 20.074 2.158 20.126 2.194 ;
        RECT 20.47 2.158 20.522 2.194 ;
        RECT 20.63 2.158 20.682 2.194 ;
        RECT 21.014 2.158 21.068 2.194 ;
        RECT 21.65 2.158 21.704 2.194 ;
        RECT 21.896 2.158 21.95 2.194 ;
        RECT 17.844 2.2405 17.916 2.2655 ;
        RECT 18.356 2.235 18.396 2.271 ;
        RECT 16.964 2.6115 17.036 2.6365 ;
        RECT 17.844 2.6115 17.916 2.6365 ;
        RECT 18.964 2.6115 19.036 2.6365 ;
        RECT 14.05 2.606 14.104 2.642 ;
        RECT 14.296 2.606 14.35 2.642 ;
        RECT 14.932 2.606 14.986 2.642 ;
        RECT 15.318 2.606 15.37 2.642 ;
        RECT 15.874 2.606 15.926 2.642 ;
        RECT 16.034 2.606 16.086 2.642 ;
        RECT 18.356 2.606 18.396 2.642 ;
        RECT 19.914 2.606 19.966 2.642 ;
        RECT 20.074 2.606 20.126 2.642 ;
        RECT 20.63 2.606 20.682 2.642 ;
        RECT 21.014 2.606 21.068 2.642 ;
        RECT 21.65 2.606 21.704 2.642 ;
        RECT 21.896 2.606 21.95 2.642 ;
        RECT 17.844 2.7635 17.916 2.7885 ;
        RECT 18.356 2.758 18.396 2.794 ;
        RECT 18.664 2.8405 18.736 2.8655 ;
        RECT 18.964 2.8405 19.036 2.8655 ;
        RECT 14.296 2.835 14.35 2.871 ;
        RECT 14.932 2.835 14.986 2.871 ;
        RECT 15.318 2.835 15.37 2.871 ;
        RECT 15.478 2.835 15.53 2.871 ;
        RECT 15.874 2.835 15.926 2.871 ;
        RECT 18.148 2.835 18.188 2.871 ;
        RECT 20.074 2.835 20.126 2.871 ;
        RECT 20.47 2.835 20.522 2.871 ;
        RECT 20.63 2.835 20.682 2.871 ;
        RECT 21.014 2.835 21.068 2.871 ;
        RECT 21.65 2.835 21.704 2.871 ;
        RECT 16.964 3.1345 17.036 3.1595 ;
        RECT 17.844 3.1345 17.916 3.1595 ;
        RECT 18.664 3.1345 18.736 3.1595 ;
        RECT 18.964 3.1345 19.036 3.1595 ;
        RECT 14.05 3.129 14.104 3.165 ;
        RECT 14.932 3.129 14.986 3.165 ;
        RECT 15.318 3.129 15.37 3.165 ;
        RECT 15.478 3.129 15.53 3.165 ;
        RECT 15.874 3.129 15.926 3.165 ;
        RECT 16.034 3.129 16.086 3.165 ;
        RECT 16.8 3.129 16.854 3.165 ;
        RECT 18.148 3.129 18.188 3.165 ;
        RECT 18.356 3.129 18.396 3.165 ;
        RECT 19.914 3.129 19.966 3.165 ;
        RECT 20.074 3.129 20.126 3.165 ;
        RECT 20.47 3.129 20.522 3.165 ;
        RECT 20.63 3.129 20.682 3.165 ;
        RECT 21.014 3.129 21.068 3.165 ;
        RECT 21.896 3.129 21.95 3.165 ;
        RECT 16.964 3.3635 17.036 3.3885 ;
        RECT 18.664 3.3635 18.736 3.3885 ;
        RECT 18.964 3.3635 19.036 3.3885 ;
        RECT 14.05 3.358 14.104 3.394 ;
        RECT 14.296 3.358 14.35 3.394 ;
        RECT 14.932 3.358 14.986 3.394 ;
        RECT 15.318 3.358 15.37 3.394 ;
        RECT 15.478 3.358 15.53 3.394 ;
        RECT 15.874 3.358 15.926 3.394 ;
        RECT 16.034 3.358 16.086 3.394 ;
        RECT 16.8 3.358 16.854 3.394 ;
        RECT 18.148 3.358 18.188 3.394 ;
        RECT 19.914 3.358 19.966 3.394 ;
        RECT 20.074 3.358 20.126 3.394 ;
        RECT 20.47 3.358 20.522 3.394 ;
        RECT 20.63 3.358 20.682 3.394 ;
        RECT 21.014 3.358 21.068 3.394 ;
        RECT 21.65 3.358 21.704 3.394 ;
        RECT 21.896 3.358 21.95 3.394 ;
        RECT 17.844 3.4405 17.916 3.4655 ;
        RECT 18.356 3.435 18.396 3.471 ;
        RECT 16.964 3.8115 17.036 3.8365 ;
        RECT 17.844 3.8115 17.916 3.8365 ;
        RECT 18.964 3.8115 19.036 3.8365 ;
        RECT 14.05 3.806 14.104 3.842 ;
        RECT 14.296 3.806 14.35 3.842 ;
        RECT 14.932 3.806 14.986 3.842 ;
        RECT 15.318 3.806 15.37 3.842 ;
        RECT 15.874 3.806 15.926 3.842 ;
        RECT 16.034 3.806 16.086 3.842 ;
        RECT 18.356 3.806 18.396 3.842 ;
        RECT 19.914 3.806 19.966 3.842 ;
        RECT 20.074 3.806 20.126 3.842 ;
        RECT 20.63 3.806 20.682 3.842 ;
        RECT 21.014 3.806 21.068 3.842 ;
        RECT 21.65 3.806 21.704 3.842 ;
        RECT 21.896 3.806 21.95 3.842 ;
        RECT 17.844 3.9635 17.916 3.9885 ;
        RECT 18.356 3.958 18.396 3.994 ;
        RECT 18.664 4.0405 18.736 4.0655 ;
        RECT 18.964 4.0405 19.036 4.0655 ;
        RECT 14.296 4.035 14.35 4.071 ;
        RECT 14.932 4.035 14.986 4.071 ;
        RECT 15.318 4.035 15.37 4.071 ;
        RECT 15.478 4.035 15.53 4.071 ;
        RECT 15.874 4.035 15.926 4.071 ;
        RECT 18.148 4.035 18.188 4.071 ;
        RECT 20.074 4.035 20.126 4.071 ;
        RECT 20.47 4.035 20.522 4.071 ;
        RECT 20.63 4.035 20.682 4.071 ;
        RECT 21.014 4.035 21.068 4.071 ;
        RECT 21.65 4.035 21.704 4.071 ;
        RECT 16.964 4.3345 17.036 4.3595 ;
        RECT 17.844 4.3345 17.916 4.3595 ;
        RECT 18.664 4.3345 18.736 4.3595 ;
        RECT 18.964 4.3345 19.036 4.3595 ;
        RECT 14.05 4.329 14.104 4.365 ;
        RECT 14.932 4.329 14.986 4.365 ;
        RECT 15.318 4.329 15.37 4.365 ;
        RECT 15.478 4.329 15.53 4.365 ;
        RECT 15.874 4.329 15.926 4.365 ;
        RECT 16.034 4.329 16.086 4.365 ;
        RECT 16.8 4.329 16.854 4.365 ;
        RECT 18.148 4.329 18.188 4.365 ;
        RECT 18.356 4.329 18.396 4.365 ;
        RECT 19.914 4.329 19.966 4.365 ;
        RECT 20.074 4.329 20.126 4.365 ;
        RECT 20.47 4.329 20.522 4.365 ;
        RECT 20.63 4.329 20.682 4.365 ;
        RECT 21.014 4.329 21.068 4.365 ;
        RECT 21.896 4.329 21.95 4.365 ;
        RECT 16.964 4.5635 17.036 4.5885 ;
        RECT 18.664 4.5635 18.736 4.5885 ;
        RECT 18.964 4.5635 19.036 4.5885 ;
        RECT 14.05 4.558 14.104 4.594 ;
        RECT 14.296 4.558 14.35 4.594 ;
        RECT 14.932 4.558 14.986 4.594 ;
        RECT 15.318 4.558 15.37 4.594 ;
        RECT 15.478 4.558 15.53 4.594 ;
        RECT 15.874 4.558 15.926 4.594 ;
        RECT 16.034 4.558 16.086 4.594 ;
        RECT 16.8 4.558 16.854 4.594 ;
        RECT 18.148 4.558 18.188 4.594 ;
        RECT 19.914 4.558 19.966 4.594 ;
        RECT 20.074 4.558 20.126 4.594 ;
        RECT 20.47 4.558 20.522 4.594 ;
        RECT 20.63 4.558 20.682 4.594 ;
        RECT 21.014 4.558 21.068 4.594 ;
        RECT 21.65 4.558 21.704 4.594 ;
        RECT 21.896 4.558 21.95 4.594 ;
        RECT 17.844 4.6405 17.916 4.6655 ;
        RECT 18.356 4.635 18.396 4.671 ;
        RECT 16.964 5.0115 17.036 5.0365 ;
        RECT 17.844 5.0115 17.916 5.0365 ;
        RECT 18.964 5.0115 19.036 5.0365 ;
        RECT 14.05 5.006 14.104 5.042 ;
        RECT 14.296 5.006 14.35 5.042 ;
        RECT 14.932 5.006 14.986 5.042 ;
        RECT 15.318 5.006 15.37 5.042 ;
        RECT 15.874 5.006 15.926 5.042 ;
        RECT 16.034 5.006 16.086 5.042 ;
        RECT 18.356 5.006 18.396 5.042 ;
        RECT 19.914 5.006 19.966 5.042 ;
        RECT 20.074 5.006 20.126 5.042 ;
        RECT 20.63 5.006 20.682 5.042 ;
        RECT 21.014 5.006 21.068 5.042 ;
        RECT 21.65 5.006 21.704 5.042 ;
        RECT 21.896 5.006 21.95 5.042 ;
        RECT 17.844 5.1635 17.916 5.1885 ;
        RECT 18.356 5.158 18.396 5.194 ;
        RECT 18.664 5.2405 18.736 5.2655 ;
        RECT 18.964 5.2405 19.036 5.2655 ;
        RECT 14.296 5.235 14.35 5.271 ;
        RECT 14.932 5.235 14.986 5.271 ;
        RECT 15.318 5.235 15.37 5.271 ;
        RECT 15.478 5.235 15.53 5.271 ;
        RECT 15.874 5.235 15.926 5.271 ;
        RECT 18.148 5.235 18.188 5.271 ;
        RECT 20.074 5.235 20.126 5.271 ;
        RECT 20.47 5.235 20.522 5.271 ;
        RECT 20.63 5.235 20.682 5.271 ;
        RECT 21.014 5.235 21.068 5.271 ;
        RECT 21.65 5.235 21.704 5.271 ;
        RECT 16.964 5.5345 17.036 5.5595 ;
        RECT 17.844 5.5345 17.916 5.5595 ;
        RECT 18.664 5.5345 18.736 5.5595 ;
        RECT 18.964 5.5345 19.036 5.5595 ;
        RECT 14.05 5.529 14.104 5.565 ;
        RECT 14.932 5.529 14.986 5.565 ;
        RECT 15.318 5.529 15.37 5.565 ;
        RECT 15.478 5.529 15.53 5.565 ;
        RECT 15.874 5.529 15.926 5.565 ;
        RECT 16.034 5.529 16.086 5.565 ;
        RECT 16.8 5.529 16.854 5.565 ;
        RECT 18.148 5.529 18.188 5.565 ;
        RECT 18.356 5.529 18.396 5.565 ;
        RECT 19.914 5.529 19.966 5.565 ;
        RECT 20.074 5.529 20.126 5.565 ;
        RECT 20.47 5.529 20.522 5.565 ;
        RECT 20.63 5.529 20.682 5.565 ;
        RECT 21.014 5.529 21.068 5.565 ;
        RECT 21.896 5.529 21.95 5.565 ;
        RECT 16.964 5.7635 17.036 5.7885 ;
        RECT 18.664 5.7635 18.736 5.7885 ;
        RECT 18.964 5.7635 19.036 5.7885 ;
        RECT 14.05 5.758 14.104 5.794 ;
        RECT 14.296 5.758 14.35 5.794 ;
        RECT 14.932 5.758 14.986 5.794 ;
        RECT 15.318 5.758 15.37 5.794 ;
        RECT 15.478 5.758 15.53 5.794 ;
        RECT 15.874 5.758 15.926 5.794 ;
        RECT 16.034 5.758 16.086 5.794 ;
        RECT 16.8 5.758 16.854 5.794 ;
        RECT 18.148 5.758 18.188 5.794 ;
        RECT 19.914 5.758 19.966 5.794 ;
        RECT 20.074 5.758 20.126 5.794 ;
        RECT 20.47 5.758 20.522 5.794 ;
        RECT 20.63 5.758 20.682 5.794 ;
        RECT 21.014 5.758 21.068 5.794 ;
        RECT 21.65 5.758 21.704 5.794 ;
        RECT 21.896 5.758 21.95 5.794 ;
        RECT 17.844 5.8405 17.916 5.8655 ;
        RECT 18.356 5.835 18.396 5.871 ;
        RECT 16.964 6.2115 17.036 6.2365 ;
        RECT 17.844 6.2115 17.916 6.2365 ;
        RECT 18.964 6.2115 19.036 6.2365 ;
        RECT 14.05 6.206 14.104 6.242 ;
        RECT 14.296 6.206 14.35 6.242 ;
        RECT 14.932 6.206 14.986 6.242 ;
        RECT 15.318 6.206 15.37 6.242 ;
        RECT 15.874 6.206 15.926 6.242 ;
        RECT 16.034 6.206 16.086 6.242 ;
        RECT 18.356 6.206 18.396 6.242 ;
        RECT 19.914 6.206 19.966 6.242 ;
        RECT 20.074 6.206 20.126 6.242 ;
        RECT 20.63 6.206 20.682 6.242 ;
        RECT 21.014 6.206 21.068 6.242 ;
        RECT 21.65 6.206 21.704 6.242 ;
        RECT 21.896 6.206 21.95 6.242 ;
        RECT 17.844 6.3635 17.916 6.3885 ;
        RECT 18.356 6.358 18.396 6.394 ;
        RECT 18.664 6.4405 18.736 6.4655 ;
        RECT 18.964 6.4405 19.036 6.4655 ;
        RECT 14.296 6.435 14.35 6.471 ;
        RECT 14.932 6.435 14.986 6.471 ;
        RECT 15.318 6.435 15.37 6.471 ;
        RECT 15.478 6.435 15.53 6.471 ;
        RECT 15.874 6.435 15.926 6.471 ;
        RECT 18.148 6.435 18.188 6.471 ;
        RECT 20.074 6.435 20.126 6.471 ;
        RECT 20.47 6.435 20.522 6.471 ;
        RECT 20.63 6.435 20.682 6.471 ;
        RECT 21.014 6.435 21.068 6.471 ;
        RECT 21.65 6.435 21.704 6.471 ;
        RECT 16.964 6.7345 17.036 6.7595 ;
        RECT 17.844 6.7345 17.916 6.7595 ;
        RECT 18.664 6.7345 18.736 6.7595 ;
        RECT 18.964 6.7345 19.036 6.7595 ;
        RECT 14.05 6.729 14.104 6.765 ;
        RECT 14.932 6.729 14.986 6.765 ;
        RECT 15.318 6.729 15.37 6.765 ;
        RECT 15.478 6.729 15.53 6.765 ;
        RECT 15.874 6.729 15.926 6.765 ;
        RECT 16.034 6.729 16.086 6.765 ;
        RECT 16.8 6.729 16.854 6.765 ;
        RECT 18.148 6.729 18.188 6.765 ;
        RECT 18.356 6.729 18.396 6.765 ;
        RECT 19.914 6.729 19.966 6.765 ;
        RECT 20.074 6.729 20.126 6.765 ;
        RECT 20.47 6.729 20.522 6.765 ;
        RECT 20.63 6.729 20.682 6.765 ;
        RECT 21.014 6.729 21.068 6.765 ;
        RECT 21.896 6.729 21.95 6.765 ;
        RECT 16.964 6.9635 17.036 6.9885 ;
        RECT 18.664 6.9635 18.736 6.9885 ;
        RECT 18.964 6.9635 19.036 6.9885 ;
        RECT 14.05 6.958 14.104 6.994 ;
        RECT 14.296 6.958 14.35 6.994 ;
        RECT 14.932 6.958 14.986 6.994 ;
        RECT 15.318 6.958 15.37 6.994 ;
        RECT 15.478 6.958 15.53 6.994 ;
        RECT 15.874 6.958 15.926 6.994 ;
        RECT 16.034 6.958 16.086 6.994 ;
        RECT 16.8 6.958 16.854 6.994 ;
        RECT 18.148 6.958 18.188 6.994 ;
        RECT 19.914 6.958 19.966 6.994 ;
        RECT 20.074 6.958 20.126 6.994 ;
        RECT 20.47 6.958 20.522 6.994 ;
        RECT 20.63 6.958 20.682 6.994 ;
        RECT 21.014 6.958 21.068 6.994 ;
        RECT 21.65 6.958 21.704 6.994 ;
        RECT 21.896 6.958 21.95 6.994 ;
        RECT 17.844 7.0405 17.916 7.0655 ;
        RECT 18.356 7.035 18.396 7.071 ;
        RECT 16.964 7.4115 17.036 7.4365 ;
        RECT 17.844 7.4115 17.916 7.4365 ;
        RECT 18.964 7.4115 19.036 7.4365 ;
        RECT 14.05 7.406 14.104 7.442 ;
        RECT 14.296 7.406 14.35 7.442 ;
        RECT 14.932 7.406 14.986 7.442 ;
        RECT 15.318 7.406 15.37 7.442 ;
        RECT 15.874 7.406 15.926 7.442 ;
        RECT 16.034 7.406 16.086 7.442 ;
        RECT 18.356 7.406 18.396 7.442 ;
        RECT 19.914 7.406 19.966 7.442 ;
        RECT 20.074 7.406 20.126 7.442 ;
        RECT 20.63 7.406 20.682 7.442 ;
        RECT 21.014 7.406 21.068 7.442 ;
        RECT 21.65 7.406 21.704 7.442 ;
        RECT 21.896 7.406 21.95 7.442 ;
        RECT 17.844 7.5635 17.916 7.5885 ;
        RECT 18.356 7.558 18.396 7.594 ;
        RECT 18.664 7.6405 18.736 7.6655 ;
        RECT 18.964 7.6405 19.036 7.6655 ;
        RECT 14.296 7.635 14.35 7.671 ;
        RECT 14.932 7.635 14.986 7.671 ;
        RECT 15.318 7.635 15.37 7.671 ;
        RECT 15.478 7.635 15.53 7.671 ;
        RECT 15.874 7.635 15.926 7.671 ;
        RECT 18.148 7.635 18.188 7.671 ;
        RECT 20.074 7.635 20.126 7.671 ;
        RECT 20.47 7.635 20.522 7.671 ;
        RECT 20.63 7.635 20.682 7.671 ;
        RECT 21.014 7.635 21.068 7.671 ;
        RECT 21.65 7.635 21.704 7.671 ;
        RECT 16.964 7.9345 17.036 7.9595 ;
        RECT 17.844 7.9345 17.916 7.9595 ;
        RECT 18.664 7.9345 18.736 7.9595 ;
        RECT 18.964 7.9345 19.036 7.9595 ;
        RECT 14.05 7.929 14.104 7.965 ;
        RECT 14.932 7.929 14.986 7.965 ;
        RECT 15.318 7.929 15.37 7.965 ;
        RECT 15.478 7.929 15.53 7.965 ;
        RECT 15.874 7.929 15.926 7.965 ;
        RECT 16.034 7.929 16.086 7.965 ;
        RECT 16.8 7.929 16.854 7.965 ;
        RECT 18.148 7.929 18.188 7.965 ;
        RECT 18.356 7.929 18.396 7.965 ;
        RECT 19.914 7.929 19.966 7.965 ;
        RECT 20.074 7.929 20.126 7.965 ;
        RECT 20.47 7.929 20.522 7.965 ;
        RECT 20.63 7.929 20.682 7.965 ;
        RECT 21.014 7.929 21.068 7.965 ;
        RECT 21.896 7.929 21.95 7.965 ;
        RECT 16.964 8.1635 17.036 8.1885 ;
        RECT 18.664 8.1635 18.736 8.1885 ;
        RECT 18.964 8.1635 19.036 8.1885 ;
        RECT 14.05 8.158 14.104 8.194 ;
        RECT 14.296 8.158 14.35 8.194 ;
        RECT 14.932 8.158 14.986 8.194 ;
        RECT 15.318 8.158 15.37 8.194 ;
        RECT 15.478 8.158 15.53 8.194 ;
        RECT 15.874 8.158 15.926 8.194 ;
        RECT 16.034 8.158 16.086 8.194 ;
        RECT 16.8 8.158 16.854 8.194 ;
        RECT 18.148 8.158 18.188 8.194 ;
        RECT 19.914 8.158 19.966 8.194 ;
        RECT 20.074 8.158 20.126 8.194 ;
        RECT 20.47 8.158 20.522 8.194 ;
        RECT 20.63 8.158 20.682 8.194 ;
        RECT 21.014 8.158 21.068 8.194 ;
        RECT 21.65 8.158 21.704 8.194 ;
        RECT 21.896 8.158 21.95 8.194 ;
        RECT 17.844 8.2405 17.916 8.2655 ;
        RECT 18.356 8.235 18.396 8.271 ;
        RECT 16.964 8.6115 17.036 8.6365 ;
        RECT 17.844 8.6115 17.916 8.6365 ;
        RECT 18.964 8.6115 19.036 8.6365 ;
        RECT 14.05 8.606 14.104 8.642 ;
        RECT 14.296 8.606 14.35 8.642 ;
        RECT 14.932 8.606 14.986 8.642 ;
        RECT 15.318 8.606 15.37 8.642 ;
        RECT 15.874 8.606 15.926 8.642 ;
        RECT 16.034 8.606 16.086 8.642 ;
        RECT 18.356 8.606 18.396 8.642 ;
        RECT 19.914 8.606 19.966 8.642 ;
        RECT 20.074 8.606 20.126 8.642 ;
        RECT 20.63 8.606 20.682 8.642 ;
        RECT 21.014 8.606 21.068 8.642 ;
        RECT 21.65 8.606 21.704 8.642 ;
        RECT 21.896 8.606 21.95 8.642 ;
        RECT 17.844 8.7635 17.916 8.7885 ;
        RECT 18.356 8.758 18.396 8.794 ;
        RECT 18.664 8.8405 18.736 8.8655 ;
        RECT 18.964 8.8405 19.036 8.8655 ;
        RECT 14.296 8.835 14.35 8.871 ;
        RECT 14.932 8.835 14.986 8.871 ;
        RECT 15.318 8.835 15.37 8.871 ;
        RECT 15.478 8.835 15.53 8.871 ;
        RECT 15.874 8.835 15.926 8.871 ;
        RECT 18.148 8.835 18.188 8.871 ;
        RECT 20.074 8.835 20.126 8.871 ;
        RECT 20.47 8.835 20.522 8.871 ;
        RECT 20.63 8.835 20.682 8.871 ;
        RECT 21.014 8.835 21.068 8.871 ;
        RECT 21.65 8.835 21.704 8.871 ;
        RECT 16.964 9.1345 17.036 9.1595 ;
        RECT 17.844 9.1345 17.916 9.1595 ;
        RECT 18.664 9.1345 18.736 9.1595 ;
        RECT 18.964 9.1345 19.036 9.1595 ;
        RECT 14.05 9.129 14.104 9.165 ;
        RECT 14.932 9.129 14.986 9.165 ;
        RECT 15.318 9.129 15.37 9.165 ;
        RECT 15.478 9.129 15.53 9.165 ;
        RECT 15.874 9.129 15.926 9.165 ;
        RECT 16.034 9.129 16.086 9.165 ;
        RECT 16.8 9.129 16.854 9.165 ;
        RECT 18.148 9.129 18.188 9.165 ;
        RECT 18.356 9.129 18.396 9.165 ;
        RECT 19.914 9.129 19.966 9.165 ;
        RECT 20.074 9.129 20.126 9.165 ;
        RECT 20.47 9.129 20.522 9.165 ;
        RECT 20.63 9.129 20.682 9.165 ;
        RECT 21.014 9.129 21.068 9.165 ;
        RECT 21.896 9.129 21.95 9.165 ;
        RECT 16.964 9.3635 17.036 9.3885 ;
        RECT 18.664 9.3635 18.736 9.3885 ;
        RECT 18.964 9.3635 19.036 9.3885 ;
        RECT 14.05 9.358 14.104 9.394 ;
        RECT 14.296 9.358 14.35 9.394 ;
        RECT 14.932 9.358 14.986 9.394 ;
        RECT 15.318 9.358 15.37 9.394 ;
        RECT 15.478 9.358 15.53 9.394 ;
        RECT 15.874 9.358 15.926 9.394 ;
        RECT 16.034 9.358 16.086 9.394 ;
        RECT 16.8 9.358 16.854 9.394 ;
        RECT 18.148 9.358 18.188 9.394 ;
        RECT 19.914 9.358 19.966 9.394 ;
        RECT 20.074 9.358 20.126 9.394 ;
        RECT 20.47 9.358 20.522 9.394 ;
        RECT 20.63 9.358 20.682 9.394 ;
        RECT 21.014 9.358 21.068 9.394 ;
        RECT 21.65 9.358 21.704 9.394 ;
        RECT 21.896 9.358 21.95 9.394 ;
        RECT 17.844 9.4405 17.916 9.4655 ;
        RECT 18.356 9.435 18.396 9.471 ;
        RECT 16.964 9.8115 17.036 9.8365 ;
        RECT 17.844 9.8115 17.916 9.8365 ;
        RECT 18.964 9.8115 19.036 9.8365 ;
        RECT 14.05 9.806 14.104 9.842 ;
        RECT 14.296 9.806 14.35 9.842 ;
        RECT 14.932 9.806 14.986 9.842 ;
        RECT 15.318 9.806 15.37 9.842 ;
        RECT 15.874 9.806 15.926 9.842 ;
        RECT 16.034 9.806 16.086 9.842 ;
        RECT 18.356 9.806 18.396 9.842 ;
        RECT 19.914 9.806 19.966 9.842 ;
        RECT 20.074 9.806 20.126 9.842 ;
        RECT 20.63 9.806 20.682 9.842 ;
        RECT 21.014 9.806 21.068 9.842 ;
        RECT 21.65 9.806 21.704 9.842 ;
        RECT 21.896 9.806 21.95 9.842 ;
        RECT 17.844 9.9635 17.916 9.9885 ;
        RECT 18.356 9.958 18.396 9.994 ;
        RECT 18.664 10.0405 18.736 10.0655 ;
        RECT 18.964 10.0405 19.036 10.0655 ;
        RECT 14.296 10.035 14.35 10.071 ;
        RECT 14.932 10.035 14.986 10.071 ;
        RECT 15.318 10.035 15.37 10.071 ;
        RECT 15.478 10.035 15.53 10.071 ;
        RECT 15.874 10.035 15.926 10.071 ;
        RECT 18.148 10.035 18.188 10.071 ;
        RECT 20.074 10.035 20.126 10.071 ;
        RECT 20.47 10.035 20.522 10.071 ;
        RECT 20.63 10.035 20.682 10.071 ;
        RECT 21.014 10.035 21.068 10.071 ;
        RECT 21.65 10.035 21.704 10.071 ;
        RECT 16.964 10.3345 17.036 10.3595 ;
        RECT 17.844 10.3345 17.916 10.3595 ;
        RECT 18.664 10.3345 18.736 10.3595 ;
        RECT 18.964 10.3345 19.036 10.3595 ;
        RECT 14.05 10.329 14.104 10.365 ;
        RECT 14.932 10.329 14.986 10.365 ;
        RECT 15.318 10.329 15.37 10.365 ;
        RECT 15.478 10.329 15.53 10.365 ;
        RECT 15.874 10.329 15.926 10.365 ;
        RECT 16.034 10.329 16.086 10.365 ;
        RECT 16.8 10.329 16.854 10.365 ;
        RECT 18.148 10.329 18.188 10.365 ;
        RECT 18.356 10.329 18.396 10.365 ;
        RECT 19.914 10.329 19.966 10.365 ;
        RECT 20.074 10.329 20.126 10.365 ;
        RECT 20.47 10.329 20.522 10.365 ;
        RECT 20.63 10.329 20.682 10.365 ;
        RECT 21.014 10.329 21.068 10.365 ;
        RECT 21.896 10.329 21.95 10.365 ;
        RECT 16.964 10.5635 17.036 10.5885 ;
        RECT 18.664 10.5635 18.736 10.5885 ;
        RECT 18.964 10.5635 19.036 10.5885 ;
        RECT 14.05 10.558 14.104 10.594 ;
        RECT 14.296 10.558 14.35 10.594 ;
        RECT 14.932 10.558 14.986 10.594 ;
        RECT 15.318 10.558 15.37 10.594 ;
        RECT 15.478 10.558 15.53 10.594 ;
        RECT 15.874 10.558 15.926 10.594 ;
        RECT 16.034 10.558 16.086 10.594 ;
        RECT 16.8 10.558 16.854 10.594 ;
        RECT 18.148 10.558 18.188 10.594 ;
        RECT 19.914 10.558 19.966 10.594 ;
        RECT 20.074 10.558 20.126 10.594 ;
        RECT 20.47 10.558 20.522 10.594 ;
        RECT 20.63 10.558 20.682 10.594 ;
        RECT 21.014 10.558 21.068 10.594 ;
        RECT 21.65 10.558 21.704 10.594 ;
        RECT 21.896 10.558 21.95 10.594 ;
        RECT 17.844 10.6405 17.916 10.6655 ;
        RECT 18.356 10.635 18.396 10.671 ;
        RECT 16.964 11.0115 17.036 11.0365 ;
        RECT 17.844 11.0115 17.916 11.0365 ;
        RECT 18.964 11.0115 19.036 11.0365 ;
        RECT 14.05 11.006 14.104 11.042 ;
        RECT 14.296 11.006 14.35 11.042 ;
        RECT 14.932 11.006 14.986 11.042 ;
        RECT 15.318 11.006 15.37 11.042 ;
        RECT 15.874 11.006 15.926 11.042 ;
        RECT 16.034 11.006 16.086 11.042 ;
        RECT 18.356 11.006 18.396 11.042 ;
        RECT 19.914 11.006 19.966 11.042 ;
        RECT 20.074 11.006 20.126 11.042 ;
        RECT 20.63 11.006 20.682 11.042 ;
        RECT 21.014 11.006 21.068 11.042 ;
        RECT 21.65 11.006 21.704 11.042 ;
        RECT 21.896 11.006 21.95 11.042 ;
        RECT 17.844 11.1635 17.916 11.1885 ;
        RECT 18.356 11.158 18.396 11.194 ;
        RECT 18.664 11.2405 18.736 11.2655 ;
        RECT 18.964 11.2405 19.036 11.2655 ;
        RECT 14.296 11.235 14.35 11.271 ;
        RECT 14.932 11.235 14.986 11.271 ;
        RECT 15.318 11.235 15.37 11.271 ;
        RECT 15.478 11.235 15.53 11.271 ;
        RECT 15.874 11.235 15.926 11.271 ;
        RECT 18.148 11.235 18.188 11.271 ;
        RECT 20.074 11.235 20.126 11.271 ;
        RECT 20.47 11.235 20.522 11.271 ;
        RECT 20.63 11.235 20.682 11.271 ;
        RECT 21.014 11.235 21.068 11.271 ;
        RECT 21.65 11.235 21.704 11.271 ;
        RECT 16.964 11.5345 17.036 11.5595 ;
        RECT 17.844 11.5345 17.916 11.5595 ;
        RECT 18.664 11.5345 18.736 11.5595 ;
        RECT 18.964 11.5345 19.036 11.5595 ;
        RECT 14.05 11.529 14.104 11.565 ;
        RECT 14.932 11.529 14.986 11.565 ;
        RECT 15.318 11.529 15.37 11.565 ;
        RECT 15.478 11.529 15.53 11.565 ;
        RECT 15.874 11.529 15.926 11.565 ;
        RECT 16.034 11.529 16.086 11.565 ;
        RECT 16.8 11.529 16.854 11.565 ;
        RECT 18.148 11.529 18.188 11.565 ;
        RECT 18.356 11.529 18.396 11.565 ;
        RECT 19.914 11.529 19.966 11.565 ;
        RECT 20.074 11.529 20.126 11.565 ;
        RECT 20.47 11.529 20.522 11.565 ;
        RECT 20.63 11.529 20.682 11.565 ;
        RECT 21.014 11.529 21.068 11.565 ;
        RECT 21.896 11.529 21.95 11.565 ;
        RECT 16.964 11.7635 17.036 11.7885 ;
        RECT 18.664 11.7635 18.736 11.7885 ;
        RECT 18.964 11.7635 19.036 11.7885 ;
        RECT 14.05 11.758 14.104 11.794 ;
        RECT 14.296 11.758 14.35 11.794 ;
        RECT 14.932 11.758 14.986 11.794 ;
        RECT 15.318 11.758 15.37 11.794 ;
        RECT 15.478 11.758 15.53 11.794 ;
        RECT 15.874 11.758 15.926 11.794 ;
        RECT 16.034 11.758 16.086 11.794 ;
        RECT 16.8 11.758 16.854 11.794 ;
        RECT 18.148 11.758 18.188 11.794 ;
        RECT 19.914 11.758 19.966 11.794 ;
        RECT 20.074 11.758 20.126 11.794 ;
        RECT 20.47 11.758 20.522 11.794 ;
        RECT 20.63 11.758 20.682 11.794 ;
        RECT 21.014 11.758 21.068 11.794 ;
        RECT 21.65 11.758 21.704 11.794 ;
        RECT 21.896 11.758 21.95 11.794 ;
        RECT 17.844 11.8405 17.916 11.8655 ;
        RECT 18.356 11.835 18.396 11.871 ;
        RECT 16.964 12.2115 17.036 12.2365 ;
        RECT 17.844 12.2115 17.916 12.2365 ;
        RECT 18.964 12.2115 19.036 12.2365 ;
        RECT 14.05 12.206 14.104 12.242 ;
        RECT 14.296 12.206 14.35 12.242 ;
        RECT 14.932 12.206 14.986 12.242 ;
        RECT 15.318 12.206 15.37 12.242 ;
        RECT 15.874 12.206 15.926 12.242 ;
        RECT 16.034 12.206 16.086 12.242 ;
        RECT 18.356 12.206 18.396 12.242 ;
        RECT 19.914 12.206 19.966 12.242 ;
        RECT 20.074 12.206 20.126 12.242 ;
        RECT 20.63 12.206 20.682 12.242 ;
        RECT 21.014 12.206 21.068 12.242 ;
        RECT 21.65 12.206 21.704 12.242 ;
        RECT 21.896 12.206 21.95 12.242 ;
        RECT 17.844 12.3635 17.916 12.3885 ;
        RECT 18.356 12.358 18.396 12.394 ;
        RECT 18.664 12.4405 18.736 12.4655 ;
        RECT 18.964 12.4405 19.036 12.4655 ;
        RECT 14.296 12.435 14.35 12.471 ;
        RECT 14.932 12.435 14.986 12.471 ;
        RECT 15.318 12.435 15.37 12.471 ;
        RECT 15.478 12.435 15.53 12.471 ;
        RECT 15.874 12.435 15.926 12.471 ;
        RECT 18.148 12.435 18.188 12.471 ;
        RECT 20.074 12.435 20.126 12.471 ;
        RECT 20.47 12.435 20.522 12.471 ;
        RECT 20.63 12.435 20.682 12.471 ;
        RECT 21.014 12.435 21.068 12.471 ;
        RECT 21.65 12.435 21.704 12.471 ;
        RECT 16.964 12.7345 17.036 12.7595 ;
        RECT 17.844 12.7345 17.916 12.7595 ;
        RECT 18.664 12.7345 18.736 12.7595 ;
        RECT 18.964 12.7345 19.036 12.7595 ;
        RECT 14.05 12.729 14.104 12.765 ;
        RECT 14.932 12.729 14.986 12.765 ;
        RECT 15.318 12.729 15.37 12.765 ;
        RECT 15.478 12.729 15.53 12.765 ;
        RECT 15.874 12.729 15.926 12.765 ;
        RECT 16.034 12.729 16.086 12.765 ;
        RECT 16.8 12.729 16.854 12.765 ;
        RECT 18.148 12.729 18.188 12.765 ;
        RECT 18.356 12.729 18.396 12.765 ;
        RECT 19.914 12.729 19.966 12.765 ;
        RECT 20.074 12.729 20.126 12.765 ;
        RECT 20.47 12.729 20.522 12.765 ;
        RECT 20.63 12.729 20.682 12.765 ;
        RECT 21.014 12.729 21.068 12.765 ;
        RECT 21.896 12.729 21.95 12.765 ;
        RECT 16.964 12.9635 17.036 12.9885 ;
        RECT 18.664 12.9635 18.736 12.9885 ;
        RECT 18.964 12.9635 19.036 12.9885 ;
        RECT 14.05 12.958 14.104 12.994 ;
        RECT 14.296 12.958 14.35 12.994 ;
        RECT 14.932 12.958 14.986 12.994 ;
        RECT 15.318 12.958 15.37 12.994 ;
        RECT 15.478 12.958 15.53 12.994 ;
        RECT 15.874 12.958 15.926 12.994 ;
        RECT 16.034 12.958 16.086 12.994 ;
        RECT 16.8 12.958 16.854 12.994 ;
        RECT 18.148 12.958 18.188 12.994 ;
        RECT 19.914 12.958 19.966 12.994 ;
        RECT 20.074 12.958 20.126 12.994 ;
        RECT 20.47 12.958 20.522 12.994 ;
        RECT 20.63 12.958 20.682 12.994 ;
        RECT 21.014 12.958 21.068 12.994 ;
        RECT 21.65 12.958 21.704 12.994 ;
        RECT 21.896 12.958 21.95 12.994 ;
        RECT 17.844 13.0405 17.916 13.0655 ;
        RECT 18.356 13.035 18.396 13.071 ;
        RECT 16.964 13.4115 17.036 13.4365 ;
        RECT 17.844 13.4115 17.916 13.4365 ;
        RECT 18.964 13.4115 19.036 13.4365 ;
        RECT 14.05 13.406 14.104 13.442 ;
        RECT 14.296 13.406 14.35 13.442 ;
        RECT 14.932 13.406 14.986 13.442 ;
        RECT 15.318 13.406 15.37 13.442 ;
        RECT 15.874 13.406 15.926 13.442 ;
        RECT 16.034 13.406 16.086 13.442 ;
        RECT 18.356 13.406 18.396 13.442 ;
        RECT 19.914 13.406 19.966 13.442 ;
        RECT 20.074 13.406 20.126 13.442 ;
        RECT 20.63 13.406 20.682 13.442 ;
        RECT 21.014 13.406 21.068 13.442 ;
        RECT 21.65 13.406 21.704 13.442 ;
        RECT 21.896 13.406 21.95 13.442 ;
        RECT 17.844 13.5635 17.916 13.5885 ;
        RECT 18.356 13.558 18.396 13.594 ;
        RECT 18.664 13.6405 18.736 13.6655 ;
        RECT 18.964 13.6405 19.036 13.6655 ;
        RECT 14.296 13.635 14.35 13.671 ;
        RECT 14.932 13.635 14.986 13.671 ;
        RECT 15.318 13.635 15.37 13.671 ;
        RECT 15.478 13.635 15.53 13.671 ;
        RECT 15.874 13.635 15.926 13.671 ;
        RECT 18.148 13.635 18.188 13.671 ;
        RECT 20.074 13.635 20.126 13.671 ;
        RECT 20.47 13.635 20.522 13.671 ;
        RECT 20.63 13.635 20.682 13.671 ;
        RECT 21.014 13.635 21.068 13.671 ;
        RECT 21.65 13.635 21.704 13.671 ;
        RECT 16.964 13.9345 17.036 13.9595 ;
        RECT 17.844 13.9345 17.916 13.9595 ;
        RECT 18.664 13.9345 18.736 13.9595 ;
        RECT 18.964 13.9345 19.036 13.9595 ;
        RECT 14.05 13.929 14.104 13.965 ;
        RECT 14.932 13.929 14.986 13.965 ;
        RECT 15.318 13.929 15.37 13.965 ;
        RECT 15.478 13.929 15.53 13.965 ;
        RECT 15.874 13.929 15.926 13.965 ;
        RECT 16.034 13.929 16.086 13.965 ;
        RECT 16.8 13.929 16.854 13.965 ;
        RECT 18.148 13.929 18.188 13.965 ;
        RECT 18.356 13.929 18.396 13.965 ;
        RECT 19.914 13.929 19.966 13.965 ;
        RECT 20.074 13.929 20.126 13.965 ;
        RECT 20.47 13.929 20.522 13.965 ;
        RECT 20.63 13.929 20.682 13.965 ;
        RECT 21.014 13.929 21.068 13.965 ;
        RECT 21.896 13.929 21.95 13.965 ;
        RECT 16.964 14.1635 17.036 14.1885 ;
        RECT 18.664 14.1635 18.736 14.1885 ;
        RECT 18.964 14.1635 19.036 14.1885 ;
        RECT 14.05 14.158 14.104 14.194 ;
        RECT 14.296 14.158 14.35 14.194 ;
        RECT 14.932 14.158 14.986 14.194 ;
        RECT 15.318 14.158 15.37 14.194 ;
        RECT 15.478 14.158 15.53 14.194 ;
        RECT 15.874 14.158 15.926 14.194 ;
        RECT 16.034 14.158 16.086 14.194 ;
        RECT 16.8 14.158 16.854 14.194 ;
        RECT 18.148 14.158 18.188 14.194 ;
        RECT 19.914 14.158 19.966 14.194 ;
        RECT 20.074 14.158 20.126 14.194 ;
        RECT 20.47 14.158 20.522 14.194 ;
        RECT 20.63 14.158 20.682 14.194 ;
        RECT 21.014 14.158 21.068 14.194 ;
        RECT 21.65 14.158 21.704 14.194 ;
        RECT 21.896 14.158 21.95 14.194 ;
        RECT 17.844 14.2405 17.916 14.2655 ;
        RECT 18.356 14.235 18.396 14.271 ;
        RECT 16.964 14.6115 17.036 14.6365 ;
        RECT 17.844 14.6115 17.916 14.6365 ;
        RECT 18.964 14.6115 19.036 14.6365 ;
        RECT 14.05 14.606 14.104 14.642 ;
        RECT 14.296 14.606 14.35 14.642 ;
        RECT 14.932 14.606 14.986 14.642 ;
        RECT 15.318 14.606 15.37 14.642 ;
        RECT 15.874 14.606 15.926 14.642 ;
        RECT 16.034 14.606 16.086 14.642 ;
        RECT 18.356 14.606 18.396 14.642 ;
        RECT 19.914 14.606 19.966 14.642 ;
        RECT 20.074 14.606 20.126 14.642 ;
        RECT 20.63 14.606 20.682 14.642 ;
        RECT 21.014 14.606 21.068 14.642 ;
        RECT 21.65 14.606 21.704 14.642 ;
        RECT 21.896 14.606 21.95 14.642 ;
        RECT 17.844 14.7635 17.916 14.7885 ;
        RECT 18.356 14.758 18.396 14.794 ;
        RECT 18.664 14.8405 18.736 14.8655 ;
        RECT 18.964 14.8405 19.036 14.8655 ;
        RECT 14.296 14.835 14.35 14.871 ;
        RECT 14.932 14.835 14.986 14.871 ;
        RECT 15.318 14.835 15.37 14.871 ;
        RECT 15.478 14.835 15.53 14.871 ;
        RECT 15.874 14.835 15.926 14.871 ;
        RECT 18.148 14.835 18.188 14.871 ;
        RECT 20.074 14.835 20.126 14.871 ;
        RECT 20.47 14.835 20.522 14.871 ;
        RECT 20.63 14.835 20.682 14.871 ;
        RECT 21.014 14.835 21.068 14.871 ;
        RECT 21.65 14.835 21.704 14.871 ;
        RECT 16.964 15.1345 17.036 15.1595 ;
        RECT 17.844 15.1345 17.916 15.1595 ;
        RECT 18.664 15.1345 18.736 15.1595 ;
        RECT 18.964 15.1345 19.036 15.1595 ;
        RECT 14.05 15.129 14.104 15.165 ;
        RECT 14.932 15.129 14.986 15.165 ;
        RECT 15.318 15.129 15.37 15.165 ;
        RECT 15.478 15.129 15.53 15.165 ;
        RECT 15.874 15.129 15.926 15.165 ;
        RECT 16.034 15.129 16.086 15.165 ;
        RECT 16.8 15.129 16.854 15.165 ;
        RECT 18.148 15.129 18.188 15.165 ;
        RECT 18.356 15.129 18.396 15.165 ;
        RECT 19.914 15.129 19.966 15.165 ;
        RECT 20.074 15.129 20.126 15.165 ;
        RECT 20.47 15.129 20.522 15.165 ;
        RECT 20.63 15.129 20.682 15.165 ;
        RECT 21.014 15.129 21.068 15.165 ;
        RECT 21.896 15.129 21.95 15.165 ;
        RECT 16.964 15.3635 17.036 15.3885 ;
        RECT 18.664 15.3635 18.736 15.3885 ;
        RECT 18.964 15.3635 19.036 15.3885 ;
        RECT 14.05 15.358 14.104 15.394 ;
        RECT 14.296 15.358 14.35 15.394 ;
        RECT 14.932 15.358 14.986 15.394 ;
        RECT 15.318 15.358 15.37 15.394 ;
        RECT 15.478 15.358 15.53 15.394 ;
        RECT 15.874 15.358 15.926 15.394 ;
        RECT 16.034 15.358 16.086 15.394 ;
        RECT 16.8 15.358 16.854 15.394 ;
        RECT 18.148 15.358 18.188 15.394 ;
        RECT 19.914 15.358 19.966 15.394 ;
        RECT 20.074 15.358 20.126 15.394 ;
        RECT 20.47 15.358 20.522 15.394 ;
        RECT 20.63 15.358 20.682 15.394 ;
        RECT 21.014 15.358 21.068 15.394 ;
        RECT 21.65 15.358 21.704 15.394 ;
        RECT 21.896 15.358 21.95 15.394 ;
        RECT 17.844 15.4405 17.916 15.4655 ;
        RECT 18.356 15.435 18.396 15.471 ;
        RECT 16.964 15.8115 17.036 15.8365 ;
        RECT 17.844 15.8115 17.916 15.8365 ;
        RECT 18.964 15.8115 19.036 15.8365 ;
        RECT 14.05 15.806 14.104 15.842 ;
        RECT 14.296 15.806 14.35 15.842 ;
        RECT 14.932 15.806 14.986 15.842 ;
        RECT 15.318 15.806 15.37 15.842 ;
        RECT 15.874 15.806 15.926 15.842 ;
        RECT 16.034 15.806 16.086 15.842 ;
        RECT 18.356 15.806 18.396 15.842 ;
        RECT 19.914 15.806 19.966 15.842 ;
        RECT 20.074 15.806 20.126 15.842 ;
        RECT 20.63 15.806 20.682 15.842 ;
        RECT 21.014 15.806 21.068 15.842 ;
        RECT 21.65 15.806 21.704 15.842 ;
        RECT 21.896 15.806 21.95 15.842 ;
        RECT 17.844 15.9635 17.916 15.9885 ;
        RECT 18.356 15.958 18.396 15.994 ;
        RECT 18.664 16.0405 18.736 16.0655 ;
        RECT 18.964 16.0405 19.036 16.0655 ;
        RECT 14.296 16.035 14.35 16.071 ;
        RECT 14.932 16.035 14.986 16.071 ;
        RECT 15.318 16.035 15.37 16.071 ;
        RECT 15.478 16.035 15.53 16.071 ;
        RECT 15.874 16.035 15.926 16.071 ;
        RECT 18.148 16.035 18.188 16.071 ;
        RECT 20.074 16.035 20.126 16.071 ;
        RECT 20.47 16.035 20.522 16.071 ;
        RECT 20.63 16.035 20.682 16.071 ;
        RECT 21.014 16.035 21.068 16.071 ;
        RECT 21.65 16.035 21.704 16.071 ;
        RECT 16.964 16.3345 17.036 16.3595 ;
        RECT 17.844 16.3345 17.916 16.3595 ;
        RECT 18.664 16.3345 18.736 16.3595 ;
        RECT 18.964 16.3345 19.036 16.3595 ;
        RECT 14.05 16.329 14.104 16.365 ;
        RECT 14.932 16.329 14.986 16.365 ;
        RECT 15.318 16.329 15.37 16.365 ;
        RECT 15.478 16.329 15.53 16.365 ;
        RECT 15.874 16.329 15.926 16.365 ;
        RECT 16.034 16.329 16.086 16.365 ;
        RECT 16.8 16.329 16.854 16.365 ;
        RECT 18.148 16.329 18.188 16.365 ;
        RECT 18.356 16.329 18.396 16.365 ;
        RECT 19.914 16.329 19.966 16.365 ;
        RECT 20.074 16.329 20.126 16.365 ;
        RECT 20.47 16.329 20.522 16.365 ;
        RECT 20.63 16.329 20.682 16.365 ;
        RECT 21.014 16.329 21.068 16.365 ;
        RECT 21.896 16.329 21.95 16.365 ;
        RECT 16.964 16.5635 17.036 16.5885 ;
        RECT 18.664 16.5635 18.736 16.5885 ;
        RECT 18.964 16.5635 19.036 16.5885 ;
        RECT 14.05 16.558 14.104 16.594 ;
        RECT 14.296 16.558 14.35 16.594 ;
        RECT 14.932 16.558 14.986 16.594 ;
        RECT 15.318 16.558 15.37 16.594 ;
        RECT 15.478 16.558 15.53 16.594 ;
        RECT 15.874 16.558 15.926 16.594 ;
        RECT 16.034 16.558 16.086 16.594 ;
        RECT 16.8 16.558 16.854 16.594 ;
        RECT 18.148 16.558 18.188 16.594 ;
        RECT 19.914 16.558 19.966 16.594 ;
        RECT 20.074 16.558 20.126 16.594 ;
        RECT 20.47 16.558 20.522 16.594 ;
        RECT 20.63 16.558 20.682 16.594 ;
        RECT 21.014 16.558 21.068 16.594 ;
        RECT 21.65 16.558 21.704 16.594 ;
        RECT 21.896 16.558 21.95 16.594 ;
        RECT 17.844 16.6405 17.916 16.6655 ;
        RECT 18.356 16.635 18.396 16.671 ;
        RECT 16.964 17.0115 17.036 17.0365 ;
        RECT 17.844 17.0115 17.916 17.0365 ;
        RECT 18.964 17.0115 19.036 17.0365 ;
        RECT 14.05 17.006 14.104 17.042 ;
        RECT 14.296 17.006 14.35 17.042 ;
        RECT 14.932 17.006 14.986 17.042 ;
        RECT 15.318 17.006 15.37 17.042 ;
        RECT 15.874 17.006 15.926 17.042 ;
        RECT 16.034 17.006 16.086 17.042 ;
        RECT 18.356 17.006 18.396 17.042 ;
        RECT 19.914 17.006 19.966 17.042 ;
        RECT 20.074 17.006 20.126 17.042 ;
        RECT 20.63 17.006 20.682 17.042 ;
        RECT 21.014 17.006 21.068 17.042 ;
        RECT 21.65 17.006 21.704 17.042 ;
        RECT 21.896 17.006 21.95 17.042 ;
        RECT 17.844 17.1635 17.916 17.1885 ;
        RECT 18.356 17.158 18.396 17.194 ;
        RECT 18.664 17.2405 18.736 17.2655 ;
        RECT 18.964 17.2405 19.036 17.2655 ;
        RECT 14.296 17.235 14.35 17.271 ;
        RECT 14.932 17.235 14.986 17.271 ;
        RECT 15.318 17.235 15.37 17.271 ;
        RECT 15.478 17.235 15.53 17.271 ;
        RECT 15.874 17.235 15.926 17.271 ;
        RECT 18.148 17.235 18.188 17.271 ;
        RECT 20.074 17.235 20.126 17.271 ;
        RECT 20.47 17.235 20.522 17.271 ;
        RECT 20.63 17.235 20.682 17.271 ;
        RECT 21.014 17.235 21.068 17.271 ;
        RECT 21.65 17.235 21.704 17.271 ;
        RECT 16.964 17.5345 17.036 17.5595 ;
        RECT 17.844 17.5345 17.916 17.5595 ;
        RECT 18.664 17.5345 18.736 17.5595 ;
        RECT 18.964 17.5345 19.036 17.5595 ;
        RECT 14.05 17.529 14.104 17.565 ;
        RECT 14.932 17.529 14.986 17.565 ;
        RECT 15.318 17.529 15.37 17.565 ;
        RECT 15.478 17.529 15.53 17.565 ;
        RECT 15.874 17.529 15.926 17.565 ;
        RECT 16.034 17.529 16.086 17.565 ;
        RECT 16.8 17.529 16.854 17.565 ;
        RECT 18.148 17.529 18.188 17.565 ;
        RECT 18.356 17.529 18.396 17.565 ;
        RECT 19.914 17.529 19.966 17.565 ;
        RECT 20.074 17.529 20.126 17.565 ;
        RECT 20.47 17.529 20.522 17.565 ;
        RECT 20.63 17.529 20.682 17.565 ;
        RECT 21.014 17.529 21.068 17.565 ;
        RECT 21.896 17.529 21.95 17.565 ;
        RECT 16.964 17.7635 17.036 17.7885 ;
        RECT 18.664 17.7635 18.736 17.7885 ;
        RECT 18.964 17.7635 19.036 17.7885 ;
        RECT 14.05 17.758 14.104 17.794 ;
        RECT 14.296 17.758 14.35 17.794 ;
        RECT 14.932 17.758 14.986 17.794 ;
        RECT 15.318 17.758 15.37 17.794 ;
        RECT 15.478 17.758 15.53 17.794 ;
        RECT 15.874 17.758 15.926 17.794 ;
        RECT 16.034 17.758 16.086 17.794 ;
        RECT 16.8 17.758 16.854 17.794 ;
        RECT 18.148 17.758 18.188 17.794 ;
        RECT 19.914 17.758 19.966 17.794 ;
        RECT 20.074 17.758 20.126 17.794 ;
        RECT 20.47 17.758 20.522 17.794 ;
        RECT 20.63 17.758 20.682 17.794 ;
        RECT 21.014 17.758 21.068 17.794 ;
        RECT 21.65 17.758 21.704 17.794 ;
        RECT 21.896 17.758 21.95 17.794 ;
        RECT 17.844 17.8405 17.916 17.8655 ;
        RECT 18.356 17.835 18.396 17.871 ;
        RECT 16.964 18.2115 17.036 18.2365 ;
        RECT 17.844 18.2115 17.916 18.2365 ;
        RECT 18.964 18.2115 19.036 18.2365 ;
        RECT 14.05 18.206 14.104 18.242 ;
        RECT 14.296 18.206 14.35 18.242 ;
        RECT 14.932 18.206 14.986 18.242 ;
        RECT 15.318 18.206 15.37 18.242 ;
        RECT 15.874 18.206 15.926 18.242 ;
        RECT 16.034 18.206 16.086 18.242 ;
        RECT 18.356 18.206 18.396 18.242 ;
        RECT 19.914 18.206 19.966 18.242 ;
        RECT 20.074 18.206 20.126 18.242 ;
        RECT 20.63 18.206 20.682 18.242 ;
        RECT 21.014 18.206 21.068 18.242 ;
        RECT 21.65 18.206 21.704 18.242 ;
        RECT 21.896 18.206 21.95 18.242 ;
        RECT 17.844 18.3635 17.916 18.3885 ;
        RECT 18.356 18.358 18.396 18.394 ;
        RECT 18.664 18.4405 18.736 18.4655 ;
        RECT 18.964 18.4405 19.036 18.4655 ;
        RECT 14.296 18.435 14.35 18.471 ;
        RECT 14.932 18.435 14.986 18.471 ;
        RECT 15.318 18.435 15.37 18.471 ;
        RECT 15.478 18.435 15.53 18.471 ;
        RECT 15.874 18.435 15.926 18.471 ;
        RECT 18.148 18.435 18.188 18.471 ;
        RECT 20.074 18.435 20.126 18.471 ;
        RECT 20.47 18.435 20.522 18.471 ;
        RECT 20.63 18.435 20.682 18.471 ;
        RECT 21.014 18.435 21.068 18.471 ;
        RECT 21.65 18.435 21.704 18.471 ;
        RECT 16.964 18.7345 17.036 18.7595 ;
        RECT 17.844 18.7345 17.916 18.7595 ;
        RECT 18.664 18.7345 18.736 18.7595 ;
        RECT 18.964 18.7345 19.036 18.7595 ;
        RECT 14.05 18.729 14.104 18.765 ;
        RECT 14.932 18.729 14.986 18.765 ;
        RECT 15.318 18.729 15.37 18.765 ;
        RECT 15.478 18.729 15.53 18.765 ;
        RECT 15.874 18.729 15.926 18.765 ;
        RECT 16.034 18.729 16.086 18.765 ;
        RECT 16.8 18.729 16.854 18.765 ;
        RECT 18.148 18.729 18.188 18.765 ;
        RECT 18.356 18.729 18.396 18.765 ;
        RECT 19.914 18.729 19.966 18.765 ;
        RECT 20.074 18.729 20.126 18.765 ;
        RECT 20.47 18.729 20.522 18.765 ;
        RECT 20.63 18.729 20.682 18.765 ;
        RECT 21.014 18.729 21.068 18.765 ;
        RECT 21.896 18.729 21.95 18.765 ;
        RECT 16.964 18.9635 17.036 18.9885 ;
        RECT 18.664 18.9635 18.736 18.9885 ;
        RECT 18.964 18.9635 19.036 18.9885 ;
        RECT 14.05 18.958 14.104 18.994 ;
        RECT 14.296 18.958 14.35 18.994 ;
        RECT 14.932 18.958 14.986 18.994 ;
        RECT 15.318 18.958 15.37 18.994 ;
        RECT 15.478 18.958 15.53 18.994 ;
        RECT 15.874 18.958 15.926 18.994 ;
        RECT 16.034 18.958 16.086 18.994 ;
        RECT 16.8 18.958 16.854 18.994 ;
        RECT 18.148 18.958 18.188 18.994 ;
        RECT 19.914 18.958 19.966 18.994 ;
        RECT 20.074 18.958 20.126 18.994 ;
        RECT 20.47 18.958 20.522 18.994 ;
        RECT 20.63 18.958 20.682 18.994 ;
        RECT 21.014 18.958 21.068 18.994 ;
        RECT 21.65 18.958 21.704 18.994 ;
        RECT 21.896 18.958 21.95 18.994 ;
        RECT 17.844 19.0405 17.916 19.0655 ;
        RECT 18.356 19.035 18.396 19.071 ;
        RECT 16.964 19.4115 17.036 19.4365 ;
        RECT 17.844 19.4115 17.916 19.4365 ;
        RECT 18.964 19.4115 19.036 19.4365 ;
        RECT 14.05 19.406 14.104 19.442 ;
        RECT 14.296 19.406 14.35 19.442 ;
        RECT 14.932 19.406 14.986 19.442 ;
        RECT 15.318 19.406 15.37 19.442 ;
        RECT 15.874 19.406 15.926 19.442 ;
        RECT 16.034 19.406 16.086 19.442 ;
        RECT 18.356 19.406 18.396 19.442 ;
        RECT 19.914 19.406 19.966 19.442 ;
        RECT 20.074 19.406 20.126 19.442 ;
        RECT 20.63 19.406 20.682 19.442 ;
        RECT 21.014 19.406 21.068 19.442 ;
        RECT 21.65 19.406 21.704 19.442 ;
        RECT 21.896 19.406 21.95 19.442 ;
        RECT 17.844 19.5635 17.916 19.5885 ;
        RECT 18.356 19.558 18.396 19.594 ;
        RECT 18.664 19.6405 18.736 19.6655 ;
        RECT 18.964 19.6405 19.036 19.6655 ;
        RECT 14.296 19.635 14.35 19.671 ;
        RECT 14.932 19.635 14.986 19.671 ;
        RECT 15.318 19.635 15.37 19.671 ;
        RECT 15.478 19.635 15.53 19.671 ;
        RECT 15.874 19.635 15.926 19.671 ;
        RECT 18.148 19.635 18.188 19.671 ;
        RECT 20.074 19.635 20.126 19.671 ;
        RECT 20.47 19.635 20.522 19.671 ;
        RECT 20.63 19.635 20.682 19.671 ;
        RECT 21.014 19.635 21.068 19.671 ;
        RECT 21.65 19.635 21.704 19.671 ;
        RECT 16.964 19.9345 17.036 19.9595 ;
        RECT 17.844 19.9345 17.916 19.9595 ;
        RECT 18.664 19.9345 18.736 19.9595 ;
        RECT 18.964 19.9345 19.036 19.9595 ;
        RECT 14.05 19.929 14.104 19.965 ;
        RECT 14.932 19.929 14.986 19.965 ;
        RECT 15.318 19.929 15.37 19.965 ;
        RECT 15.478 19.929 15.53 19.965 ;
        RECT 15.874 19.929 15.926 19.965 ;
        RECT 16.034 19.929 16.086 19.965 ;
        RECT 16.8 19.929 16.854 19.965 ;
        RECT 18.148 19.929 18.188 19.965 ;
        RECT 18.356 19.929 18.396 19.965 ;
        RECT 19.914 19.929 19.966 19.965 ;
        RECT 20.074 19.929 20.126 19.965 ;
        RECT 20.47 19.929 20.522 19.965 ;
        RECT 20.63 19.929 20.682 19.965 ;
        RECT 21.014 19.929 21.068 19.965 ;
        RECT 21.896 19.929 21.95 19.965 ;
        RECT 16.964 20.1635 17.036 20.1885 ;
        RECT 18.664 20.1635 18.736 20.1885 ;
        RECT 18.964 20.1635 19.036 20.1885 ;
        RECT 14.05 20.158 14.104 20.194 ;
        RECT 14.296 20.158 14.35 20.194 ;
        RECT 14.932 20.158 14.986 20.194 ;
        RECT 15.318 20.158 15.37 20.194 ;
        RECT 15.478 20.158 15.53 20.194 ;
        RECT 15.874 20.158 15.926 20.194 ;
        RECT 16.034 20.158 16.086 20.194 ;
        RECT 16.8 20.158 16.854 20.194 ;
        RECT 18.148 20.158 18.188 20.194 ;
        RECT 19.914 20.158 19.966 20.194 ;
        RECT 20.074 20.158 20.126 20.194 ;
        RECT 20.47 20.158 20.522 20.194 ;
        RECT 20.63 20.158 20.682 20.194 ;
        RECT 21.014 20.158 21.068 20.194 ;
        RECT 21.65 20.158 21.704 20.194 ;
        RECT 21.896 20.158 21.95 20.194 ;
        RECT 17.844 20.2405 17.916 20.2655 ;
        RECT 18.356 20.235 18.396 20.271 ;
        RECT 16.964 20.6115 17.036 20.6365 ;
        RECT 17.844 20.6115 17.916 20.6365 ;
        RECT 18.964 20.6115 19.036 20.6365 ;
        RECT 14.05 20.606 14.104 20.642 ;
        RECT 14.296 20.606 14.35 20.642 ;
        RECT 14.932 20.606 14.986 20.642 ;
        RECT 15.318 20.606 15.37 20.642 ;
        RECT 15.874 20.606 15.926 20.642 ;
        RECT 16.034 20.606 16.086 20.642 ;
        RECT 18.356 20.606 18.396 20.642 ;
        RECT 19.914 20.606 19.966 20.642 ;
        RECT 20.074 20.606 20.126 20.642 ;
        RECT 20.63 20.606 20.682 20.642 ;
        RECT 21.014 20.606 21.068 20.642 ;
        RECT 21.65 20.606 21.704 20.642 ;
        RECT 21.896 20.606 21.95 20.642 ;
        RECT 17.844 20.7635 17.916 20.7885 ;
        RECT 18.356 20.758 18.396 20.794 ;
        RECT 18.664 20.8405 18.736 20.8655 ;
        RECT 18.964 20.8405 19.036 20.8655 ;
        RECT 14.296 20.835 14.35 20.871 ;
        RECT 14.932 20.835 14.986 20.871 ;
        RECT 15.318 20.835 15.37 20.871 ;
        RECT 15.478 20.835 15.53 20.871 ;
        RECT 15.874 20.835 15.926 20.871 ;
        RECT 18.148 20.835 18.188 20.871 ;
        RECT 20.074 20.835 20.126 20.871 ;
        RECT 20.47 20.835 20.522 20.871 ;
        RECT 20.63 20.835 20.682 20.871 ;
        RECT 21.014 20.835 21.068 20.871 ;
        RECT 21.65 20.835 21.704 20.871 ;
        RECT 16.964 21.1345 17.036 21.1595 ;
        RECT 17.844 21.1345 17.916 21.1595 ;
        RECT 18.664 21.1345 18.736 21.1595 ;
        RECT 18.964 21.1345 19.036 21.1595 ;
        RECT 14.05 21.129 14.104 21.165 ;
        RECT 14.932 21.129 14.986 21.165 ;
        RECT 15.318 21.129 15.37 21.165 ;
        RECT 15.478 21.129 15.53 21.165 ;
        RECT 15.874 21.129 15.926 21.165 ;
        RECT 16.034 21.129 16.086 21.165 ;
        RECT 16.8 21.129 16.854 21.165 ;
        RECT 18.148 21.129 18.188 21.165 ;
        RECT 18.356 21.129 18.396 21.165 ;
        RECT 19.914 21.129 19.966 21.165 ;
        RECT 20.074 21.129 20.126 21.165 ;
        RECT 20.47 21.129 20.522 21.165 ;
        RECT 20.63 21.129 20.682 21.165 ;
        RECT 21.014 21.129 21.068 21.165 ;
        RECT 21.896 21.129 21.95 21.165 ;
        RECT 16.964 21.3635 17.036 21.3885 ;
        RECT 18.664 21.3635 18.736 21.3885 ;
        RECT 18.964 21.3635 19.036 21.3885 ;
        RECT 14.05 21.358 14.104 21.394 ;
        RECT 14.296 21.358 14.35 21.394 ;
        RECT 14.932 21.358 14.986 21.394 ;
        RECT 15.318 21.358 15.37 21.394 ;
        RECT 15.478 21.358 15.53 21.394 ;
        RECT 15.874 21.358 15.926 21.394 ;
        RECT 16.034 21.358 16.086 21.394 ;
        RECT 16.8 21.358 16.854 21.394 ;
        RECT 18.148 21.358 18.188 21.394 ;
        RECT 19.914 21.358 19.966 21.394 ;
        RECT 20.074 21.358 20.126 21.394 ;
        RECT 20.47 21.358 20.522 21.394 ;
        RECT 20.63 21.358 20.682 21.394 ;
        RECT 21.014 21.358 21.068 21.394 ;
        RECT 21.65 21.358 21.704 21.394 ;
        RECT 21.896 21.358 21.95 21.394 ;
        RECT 17.844 21.4405 17.916 21.4655 ;
        RECT 18.356 21.435 18.396 21.471 ;
        RECT 16.964 21.8115 17.036 21.8365 ;
        RECT 17.844 21.8115 17.916 21.8365 ;
        RECT 18.964 21.8115 19.036 21.8365 ;
        RECT 14.05 21.806 14.104 21.842 ;
        RECT 14.296 21.806 14.35 21.842 ;
        RECT 14.932 21.806 14.986 21.842 ;
        RECT 15.318 21.806 15.37 21.842 ;
        RECT 15.874 21.806 15.926 21.842 ;
        RECT 16.034 21.806 16.086 21.842 ;
        RECT 18.356 21.806 18.396 21.842 ;
        RECT 19.914 21.806 19.966 21.842 ;
        RECT 20.074 21.806 20.126 21.842 ;
        RECT 20.63 21.806 20.682 21.842 ;
        RECT 21.014 21.806 21.068 21.842 ;
        RECT 21.65 21.806 21.704 21.842 ;
        RECT 21.896 21.806 21.95 21.842 ;
        RECT 17.844 21.9635 17.916 21.9885 ;
        RECT 18.356 21.958 18.396 21.994 ;
        RECT 18.664 22.0405 18.736 22.0655 ;
        RECT 18.964 22.0405 19.036 22.0655 ;
        RECT 14.296 22.035 14.35 22.071 ;
        RECT 14.932 22.035 14.986 22.071 ;
        RECT 15.318 22.035 15.37 22.071 ;
        RECT 15.478 22.035 15.53 22.071 ;
        RECT 15.874 22.035 15.926 22.071 ;
        RECT 18.148 22.035 18.188 22.071 ;
        RECT 20.074 22.035 20.126 22.071 ;
        RECT 20.47 22.035 20.522 22.071 ;
        RECT 20.63 22.035 20.682 22.071 ;
        RECT 21.014 22.035 21.068 22.071 ;
        RECT 21.65 22.035 21.704 22.071 ;
        RECT 16.964 22.3345 17.036 22.3595 ;
        RECT 17.844 22.3345 17.916 22.3595 ;
        RECT 18.664 22.3345 18.736 22.3595 ;
        RECT 18.964 22.3345 19.036 22.3595 ;
        RECT 14.05 22.329 14.104 22.365 ;
        RECT 14.932 22.329 14.986 22.365 ;
        RECT 15.318 22.329 15.37 22.365 ;
        RECT 15.478 22.329 15.53 22.365 ;
        RECT 15.874 22.329 15.926 22.365 ;
        RECT 16.034 22.329 16.086 22.365 ;
        RECT 16.8 22.329 16.854 22.365 ;
        RECT 18.148 22.329 18.188 22.365 ;
        RECT 18.356 22.329 18.396 22.365 ;
        RECT 19.914 22.329 19.966 22.365 ;
        RECT 20.074 22.329 20.126 22.365 ;
        RECT 20.47 22.329 20.522 22.365 ;
        RECT 20.63 22.329 20.682 22.365 ;
        RECT 21.014 22.329 21.068 22.365 ;
        RECT 21.896 22.329 21.95 22.365 ;
        RECT 16.964 22.5635 17.036 22.5885 ;
        RECT 18.664 22.5635 18.736 22.5885 ;
        RECT 18.964 22.5635 19.036 22.5885 ;
        RECT 14.05 22.558 14.104 22.594 ;
        RECT 14.296 22.558 14.35 22.594 ;
        RECT 14.932 22.558 14.986 22.594 ;
        RECT 15.318 22.558 15.37 22.594 ;
        RECT 15.478 22.558 15.53 22.594 ;
        RECT 15.874 22.558 15.926 22.594 ;
        RECT 16.034 22.558 16.086 22.594 ;
        RECT 16.8 22.558 16.854 22.594 ;
        RECT 18.148 22.558 18.188 22.594 ;
        RECT 19.914 22.558 19.966 22.594 ;
        RECT 20.074 22.558 20.126 22.594 ;
        RECT 20.47 22.558 20.522 22.594 ;
        RECT 20.63 22.558 20.682 22.594 ;
        RECT 21.014 22.558 21.068 22.594 ;
        RECT 21.65 22.558 21.704 22.594 ;
        RECT 21.896 22.558 21.95 22.594 ;
        RECT 17.844 22.6405 17.916 22.6655 ;
        RECT 18.356 22.635 18.396 22.671 ;
        RECT 16.964 23.0115 17.036 23.0365 ;
        RECT 17.844 23.0115 17.916 23.0365 ;
        RECT 18.964 23.0115 19.036 23.0365 ;
        RECT 14.05 23.006 14.104 23.042 ;
        RECT 14.296 23.006 14.35 23.042 ;
        RECT 14.932 23.006 14.986 23.042 ;
        RECT 15.318 23.006 15.37 23.042 ;
        RECT 15.874 23.006 15.926 23.042 ;
        RECT 16.034 23.006 16.086 23.042 ;
        RECT 18.356 23.006 18.396 23.042 ;
        RECT 19.914 23.006 19.966 23.042 ;
        RECT 20.074 23.006 20.126 23.042 ;
        RECT 20.63 23.006 20.682 23.042 ;
        RECT 21.014 23.006 21.068 23.042 ;
        RECT 21.65 23.006 21.704 23.042 ;
        RECT 21.896 23.006 21.95 23.042 ;
        RECT 17.844 23.1635 17.916 23.1885 ;
        RECT 18.356 23.158 18.396 23.194 ;
        RECT 18.664 23.2405 18.736 23.2655 ;
        RECT 18.964 23.2405 19.036 23.2655 ;
        RECT 14.296 23.235 14.35 23.271 ;
        RECT 14.932 23.235 14.986 23.271 ;
        RECT 15.318 23.235 15.37 23.271 ;
        RECT 15.478 23.235 15.53 23.271 ;
        RECT 15.874 23.235 15.926 23.271 ;
        RECT 18.148 23.235 18.188 23.271 ;
        RECT 20.074 23.235 20.126 23.271 ;
        RECT 20.47 23.235 20.522 23.271 ;
        RECT 20.63 23.235 20.682 23.271 ;
        RECT 21.014 23.235 21.068 23.271 ;
        RECT 21.65 23.235 21.704 23.271 ;
        RECT 16.964 23.5345 17.036 23.5595 ;
        RECT 17.844 23.5345 17.916 23.5595 ;
        RECT 18.664 23.5345 18.736 23.5595 ;
        RECT 18.964 23.5345 19.036 23.5595 ;
        RECT 14.05 23.529 14.104 23.565 ;
        RECT 14.932 23.529 14.986 23.565 ;
        RECT 15.318 23.529 15.37 23.565 ;
        RECT 15.478 23.529 15.53 23.565 ;
        RECT 15.874 23.529 15.926 23.565 ;
        RECT 16.034 23.529 16.086 23.565 ;
        RECT 16.8 23.529 16.854 23.565 ;
        RECT 18.148 23.529 18.188 23.565 ;
        RECT 18.356 23.529 18.396 23.565 ;
        RECT 19.914 23.529 19.966 23.565 ;
        RECT 20.074 23.529 20.126 23.565 ;
        RECT 20.47 23.529 20.522 23.565 ;
        RECT 20.63 23.529 20.682 23.565 ;
        RECT 21.014 23.529 21.068 23.565 ;
        RECT 21.896 23.529 21.95 23.565 ;
        RECT 16.964 23.7635 17.036 23.7885 ;
        RECT 18.664 23.7635 18.736 23.7885 ;
        RECT 18.964 23.7635 19.036 23.7885 ;
        RECT 14.05 23.758 14.104 23.794 ;
        RECT 14.296 23.758 14.35 23.794 ;
        RECT 14.932 23.758 14.986 23.794 ;
        RECT 15.318 23.758 15.37 23.794 ;
        RECT 15.478 23.758 15.53 23.794 ;
        RECT 15.874 23.758 15.926 23.794 ;
        RECT 16.034 23.758 16.086 23.794 ;
        RECT 16.8 23.758 16.854 23.794 ;
        RECT 18.148 23.758 18.188 23.794 ;
        RECT 19.914 23.758 19.966 23.794 ;
        RECT 20.074 23.758 20.126 23.794 ;
        RECT 20.47 23.758 20.522 23.794 ;
        RECT 20.63 23.758 20.682 23.794 ;
        RECT 21.014 23.758 21.068 23.794 ;
        RECT 21.65 23.758 21.704 23.794 ;
        RECT 21.896 23.758 21.95 23.794 ;
        RECT 17.844 23.8405 17.916 23.8655 ;
        RECT 18.356 23.835 18.396 23.871 ;
        RECT 16.964 24.2115 17.036 24.2365 ;
        RECT 17.844 24.2115 17.916 24.2365 ;
        RECT 18.964 24.2115 19.036 24.2365 ;
        RECT 14.05 24.206 14.104 24.242 ;
        RECT 14.296 24.206 14.35 24.242 ;
        RECT 14.932 24.206 14.986 24.242 ;
        RECT 15.318 24.206 15.37 24.242 ;
        RECT 15.874 24.206 15.926 24.242 ;
        RECT 16.034 24.206 16.086 24.242 ;
        RECT 18.356 24.206 18.396 24.242 ;
        RECT 19.914 24.206 19.966 24.242 ;
        RECT 20.074 24.206 20.126 24.242 ;
        RECT 20.63 24.206 20.682 24.242 ;
        RECT 21.014 24.206 21.068 24.242 ;
        RECT 21.65 24.206 21.704 24.242 ;
        RECT 21.896 24.206 21.95 24.242 ;
        RECT 17.844 24.3635 17.916 24.3885 ;
        RECT 18.356 24.358 18.396 24.394 ;
        RECT 18.664 24.4405 18.736 24.4655 ;
        RECT 18.964 24.4405 19.036 24.4655 ;
        RECT 14.296 24.435 14.35 24.471 ;
        RECT 14.932 24.435 14.986 24.471 ;
        RECT 15.318 24.435 15.37 24.471 ;
        RECT 15.478 24.435 15.53 24.471 ;
        RECT 15.874 24.435 15.926 24.471 ;
        RECT 18.148 24.435 18.188 24.471 ;
        RECT 20.074 24.435 20.126 24.471 ;
        RECT 20.47 24.435 20.522 24.471 ;
        RECT 20.63 24.435 20.682 24.471 ;
        RECT 21.014 24.435 21.068 24.471 ;
        RECT 21.65 24.435 21.704 24.471 ;
        RECT 16.964 24.7345 17.036 24.7595 ;
        RECT 17.844 24.7345 17.916 24.7595 ;
        RECT 18.664 24.7345 18.736 24.7595 ;
        RECT 18.964 24.7345 19.036 24.7595 ;
        RECT 14.05 24.729 14.104 24.765 ;
        RECT 14.932 24.729 14.986 24.765 ;
        RECT 15.318 24.729 15.37 24.765 ;
        RECT 15.478 24.729 15.53 24.765 ;
        RECT 15.874 24.729 15.926 24.765 ;
        RECT 16.034 24.729 16.086 24.765 ;
        RECT 16.8 24.729 16.854 24.765 ;
        RECT 18.148 24.729 18.188 24.765 ;
        RECT 18.356 24.729 18.396 24.765 ;
        RECT 19.914 24.729 19.966 24.765 ;
        RECT 20.074 24.729 20.126 24.765 ;
        RECT 20.47 24.729 20.522 24.765 ;
        RECT 20.63 24.729 20.682 24.765 ;
        RECT 21.014 24.729 21.068 24.765 ;
        RECT 21.896 24.729 21.95 24.765 ;
        RECT 16.964 24.9635 17.036 24.9885 ;
        RECT 18.664 24.9635 18.736 24.9885 ;
        RECT 18.964 24.9635 19.036 24.9885 ;
        RECT 14.05 24.958 14.104 24.994 ;
        RECT 14.296 24.958 14.35 24.994 ;
        RECT 14.932 24.958 14.986 24.994 ;
        RECT 15.318 24.958 15.37 24.994 ;
        RECT 15.478 24.958 15.53 24.994 ;
        RECT 15.874 24.958 15.926 24.994 ;
        RECT 16.034 24.958 16.086 24.994 ;
        RECT 16.8 24.958 16.854 24.994 ;
        RECT 18.148 24.958 18.188 24.994 ;
        RECT 19.914 24.958 19.966 24.994 ;
        RECT 20.074 24.958 20.126 24.994 ;
        RECT 20.47 24.958 20.522 24.994 ;
        RECT 20.63 24.958 20.682 24.994 ;
        RECT 21.014 24.958 21.068 24.994 ;
        RECT 21.65 24.958 21.704 24.994 ;
        RECT 21.896 24.958 21.95 24.994 ;
        RECT 17.844 25.0405 17.916 25.0655 ;
        RECT 18.356 25.035 18.396 25.071 ;
        RECT 16.964 25.4115 17.036 25.4365 ;
        RECT 17.844 25.4115 17.916 25.4365 ;
        RECT 18.964 25.4115 19.036 25.4365 ;
        RECT 14.05 25.406 14.104 25.442 ;
        RECT 14.296 25.406 14.35 25.442 ;
        RECT 14.932 25.406 14.986 25.442 ;
        RECT 15.318 25.406 15.37 25.442 ;
        RECT 15.874 25.406 15.926 25.442 ;
        RECT 16.034 25.406 16.086 25.442 ;
        RECT 18.356 25.406 18.396 25.442 ;
        RECT 19.914 25.406 19.966 25.442 ;
        RECT 20.074 25.406 20.126 25.442 ;
        RECT 20.63 25.406 20.682 25.442 ;
        RECT 21.014 25.406 21.068 25.442 ;
        RECT 21.65 25.406 21.704 25.442 ;
        RECT 21.896 25.406 21.95 25.442 ;
        RECT 17.844 25.5635 17.916 25.5885 ;
        RECT 18.356 25.558 18.396 25.594 ;
        RECT 18.664 25.6405 18.736 25.6655 ;
        RECT 18.964 25.6405 19.036 25.6655 ;
        RECT 14.296 25.635 14.35 25.671 ;
        RECT 14.932 25.635 14.986 25.671 ;
        RECT 15.318 25.635 15.37 25.671 ;
        RECT 15.478 25.635 15.53 25.671 ;
        RECT 15.874 25.635 15.926 25.671 ;
        RECT 18.148 25.635 18.188 25.671 ;
        RECT 20.074 25.635 20.126 25.671 ;
        RECT 20.47 25.635 20.522 25.671 ;
        RECT 20.63 25.635 20.682 25.671 ;
        RECT 21.014 25.635 21.068 25.671 ;
        RECT 21.65 25.635 21.704 25.671 ;
        RECT 16.964 25.9345 17.036 25.9595 ;
        RECT 17.844 25.9345 17.916 25.9595 ;
        RECT 18.664 25.9345 18.736 25.9595 ;
        RECT 18.964 25.9345 19.036 25.9595 ;
        RECT 14.05 25.929 14.104 25.965 ;
        RECT 14.932 25.929 14.986 25.965 ;
        RECT 15.318 25.929 15.37 25.965 ;
        RECT 15.478 25.929 15.53 25.965 ;
        RECT 15.874 25.929 15.926 25.965 ;
        RECT 16.034 25.929 16.086 25.965 ;
        RECT 16.8 25.929 16.854 25.965 ;
        RECT 18.148 25.929 18.188 25.965 ;
        RECT 18.356 25.929 18.396 25.965 ;
        RECT 19.914 25.929 19.966 25.965 ;
        RECT 20.074 25.929 20.126 25.965 ;
        RECT 20.47 25.929 20.522 25.965 ;
        RECT 20.63 25.929 20.682 25.965 ;
        RECT 21.014 25.929 21.068 25.965 ;
        RECT 21.896 25.929 21.95 25.965 ;
        RECT 16.964 26.1635 17.036 26.1885 ;
        RECT 18.664 26.1635 18.736 26.1885 ;
        RECT 18.964 26.1635 19.036 26.1885 ;
        RECT 14.05 26.158 14.104 26.194 ;
        RECT 14.296 26.158 14.35 26.194 ;
        RECT 14.932 26.158 14.986 26.194 ;
        RECT 15.318 26.158 15.37 26.194 ;
        RECT 15.478 26.158 15.53 26.194 ;
        RECT 15.874 26.158 15.926 26.194 ;
        RECT 16.034 26.158 16.086 26.194 ;
        RECT 16.8 26.158 16.854 26.194 ;
        RECT 18.148 26.158 18.188 26.194 ;
        RECT 19.914 26.158 19.966 26.194 ;
        RECT 20.074 26.158 20.126 26.194 ;
        RECT 20.47 26.158 20.522 26.194 ;
        RECT 20.63 26.158 20.682 26.194 ;
        RECT 21.014 26.158 21.068 26.194 ;
        RECT 21.65 26.158 21.704 26.194 ;
        RECT 21.896 26.158 21.95 26.194 ;
        RECT 17.844 26.2405 17.916 26.2655 ;
        RECT 18.356 26.235 18.396 26.271 ;
        RECT 16.964 26.6115 17.036 26.6365 ;
        RECT 17.844 26.6115 17.916 26.6365 ;
        RECT 18.964 26.6115 19.036 26.6365 ;
        RECT 14.05 26.606 14.104 26.642 ;
        RECT 14.296 26.606 14.35 26.642 ;
        RECT 14.932 26.606 14.986 26.642 ;
        RECT 15.318 26.606 15.37 26.642 ;
        RECT 15.874 26.606 15.926 26.642 ;
        RECT 16.034 26.606 16.086 26.642 ;
        RECT 18.356 26.606 18.396 26.642 ;
        RECT 19.914 26.606 19.966 26.642 ;
        RECT 20.074 26.606 20.126 26.642 ;
        RECT 20.63 26.606 20.682 26.642 ;
        RECT 21.014 26.606 21.068 26.642 ;
        RECT 21.65 26.606 21.704 26.642 ;
        RECT 21.896 26.606 21.95 26.642 ;
        RECT 17.844 26.7635 17.916 26.7885 ;
        RECT 18.356 26.758 18.396 26.794 ;
        RECT 18.664 26.8405 18.736 26.8655 ;
        RECT 18.964 26.8405 19.036 26.8655 ;
        RECT 14.296 26.835 14.35 26.871 ;
        RECT 14.932 26.835 14.986 26.871 ;
        RECT 15.318 26.835 15.37 26.871 ;
        RECT 15.478 26.835 15.53 26.871 ;
        RECT 15.874 26.835 15.926 26.871 ;
        RECT 18.148 26.835 18.188 26.871 ;
        RECT 20.074 26.835 20.126 26.871 ;
        RECT 20.47 26.835 20.522 26.871 ;
        RECT 20.63 26.835 20.682 26.871 ;
        RECT 21.014 26.835 21.068 26.871 ;
        RECT 21.65 26.835 21.704 26.871 ;
        RECT 16.964 27.1345 17.036 27.1595 ;
        RECT 17.844 27.1345 17.916 27.1595 ;
        RECT 18.664 27.1345 18.736 27.1595 ;
        RECT 18.964 27.1345 19.036 27.1595 ;
        RECT 14.05 27.129 14.104 27.165 ;
        RECT 14.932 27.129 14.986 27.165 ;
        RECT 15.318 27.129 15.37 27.165 ;
        RECT 15.478 27.129 15.53 27.165 ;
        RECT 15.874 27.129 15.926 27.165 ;
        RECT 16.034 27.129 16.086 27.165 ;
        RECT 16.8 27.129 16.854 27.165 ;
        RECT 18.148 27.129 18.188 27.165 ;
        RECT 18.356 27.129 18.396 27.165 ;
        RECT 19.914 27.129 19.966 27.165 ;
        RECT 20.074 27.129 20.126 27.165 ;
        RECT 20.47 27.129 20.522 27.165 ;
        RECT 20.63 27.129 20.682 27.165 ;
        RECT 21.014 27.129 21.068 27.165 ;
        RECT 21.896 27.129 21.95 27.165 ;
        RECT 16.964 27.3635 17.036 27.3885 ;
        RECT 18.664 27.3635 18.736 27.3885 ;
        RECT 18.964 27.3635 19.036 27.3885 ;
        RECT 14.05 27.358 14.104 27.394 ;
        RECT 14.296 27.358 14.35 27.394 ;
        RECT 14.932 27.358 14.986 27.394 ;
        RECT 15.318 27.358 15.37 27.394 ;
        RECT 15.478 27.358 15.53 27.394 ;
        RECT 15.874 27.358 15.926 27.394 ;
        RECT 16.034 27.358 16.086 27.394 ;
        RECT 16.8 27.358 16.854 27.394 ;
        RECT 18.148 27.358 18.188 27.394 ;
        RECT 19.914 27.358 19.966 27.394 ;
        RECT 20.074 27.358 20.126 27.394 ;
        RECT 20.47 27.358 20.522 27.394 ;
        RECT 20.63 27.358 20.682 27.394 ;
        RECT 21.014 27.358 21.068 27.394 ;
        RECT 21.65 27.358 21.704 27.394 ;
        RECT 21.896 27.358 21.95 27.394 ;
        RECT 17.844 27.4405 17.916 27.4655 ;
        RECT 18.356 27.435 18.396 27.471 ;
        RECT 16.964 27.8115 17.036 27.8365 ;
        RECT 17.844 27.8115 17.916 27.8365 ;
        RECT 18.964 27.8115 19.036 27.8365 ;
        RECT 14.05 27.806 14.104 27.842 ;
        RECT 14.296 27.806 14.35 27.842 ;
        RECT 14.932 27.806 14.986 27.842 ;
        RECT 15.318 27.806 15.37 27.842 ;
        RECT 15.874 27.806 15.926 27.842 ;
        RECT 16.034 27.806 16.086 27.842 ;
        RECT 18.356 27.806 18.396 27.842 ;
        RECT 19.914 27.806 19.966 27.842 ;
        RECT 20.074 27.806 20.126 27.842 ;
        RECT 20.63 27.806 20.682 27.842 ;
        RECT 21.014 27.806 21.068 27.842 ;
        RECT 21.65 27.806 21.704 27.842 ;
        RECT 21.896 27.806 21.95 27.842 ;
        RECT 17.844 27.9635 17.916 27.9885 ;
        RECT 18.356 27.958 18.396 27.994 ;
        RECT 18.664 28.0405 18.736 28.0655 ;
        RECT 18.964 28.0405 19.036 28.0655 ;
        RECT 14.296 28.035 14.35 28.071 ;
        RECT 14.932 28.035 14.986 28.071 ;
        RECT 15.318 28.035 15.37 28.071 ;
        RECT 15.478 28.035 15.53 28.071 ;
        RECT 15.874 28.035 15.926 28.071 ;
        RECT 18.148 28.035 18.188 28.071 ;
        RECT 20.074 28.035 20.126 28.071 ;
        RECT 20.47 28.035 20.522 28.071 ;
        RECT 20.63 28.035 20.682 28.071 ;
        RECT 21.014 28.035 21.068 28.071 ;
        RECT 21.65 28.035 21.704 28.071 ;
        RECT 16.964 28.3345 17.036 28.3595 ;
        RECT 17.844 28.3345 17.916 28.3595 ;
        RECT 18.664 28.3345 18.736 28.3595 ;
        RECT 18.964 28.3345 19.036 28.3595 ;
        RECT 14.05 28.329 14.104 28.365 ;
        RECT 14.932 28.329 14.986 28.365 ;
        RECT 15.318 28.329 15.37 28.365 ;
        RECT 15.478 28.329 15.53 28.365 ;
        RECT 15.874 28.329 15.926 28.365 ;
        RECT 16.034 28.329 16.086 28.365 ;
        RECT 16.8 28.329 16.854 28.365 ;
        RECT 18.148 28.329 18.188 28.365 ;
        RECT 18.356 28.329 18.396 28.365 ;
        RECT 19.914 28.329 19.966 28.365 ;
        RECT 20.074 28.329 20.126 28.365 ;
        RECT 20.47 28.329 20.522 28.365 ;
        RECT 20.63 28.329 20.682 28.365 ;
        RECT 21.014 28.329 21.068 28.365 ;
        RECT 21.896 28.329 21.95 28.365 ;
        RECT 16.964 28.5635 17.036 28.5885 ;
        RECT 18.664 28.5635 18.736 28.5885 ;
        RECT 18.964 28.5635 19.036 28.5885 ;
        RECT 14.05 28.558 14.104 28.594 ;
        RECT 14.296 28.558 14.35 28.594 ;
        RECT 14.932 28.558 14.986 28.594 ;
        RECT 15.318 28.558 15.37 28.594 ;
        RECT 15.478 28.558 15.53 28.594 ;
        RECT 15.874 28.558 15.926 28.594 ;
        RECT 16.034 28.558 16.086 28.594 ;
        RECT 16.8 28.558 16.854 28.594 ;
        RECT 18.148 28.558 18.188 28.594 ;
        RECT 19.914 28.558 19.966 28.594 ;
        RECT 20.074 28.558 20.126 28.594 ;
        RECT 20.47 28.558 20.522 28.594 ;
        RECT 20.63 28.558 20.682 28.594 ;
        RECT 21.014 28.558 21.068 28.594 ;
        RECT 21.65 28.558 21.704 28.594 ;
        RECT 21.896 28.558 21.95 28.594 ;
        RECT 17.844 28.6405 17.916 28.6655 ;
        RECT 18.356 28.635 18.396 28.671 ;
        RECT 16.964 29.0115 17.036 29.0365 ;
        RECT 17.844 29.0115 17.916 29.0365 ;
        RECT 18.964 29.0115 19.036 29.0365 ;
        RECT 14.05 29.006 14.104 29.042 ;
        RECT 14.296 29.006 14.35 29.042 ;
        RECT 14.932 29.006 14.986 29.042 ;
        RECT 15.318 29.006 15.37 29.042 ;
        RECT 15.874 29.006 15.926 29.042 ;
        RECT 16.034 29.006 16.086 29.042 ;
        RECT 18.356 29.006 18.396 29.042 ;
        RECT 19.914 29.006 19.966 29.042 ;
        RECT 20.074 29.006 20.126 29.042 ;
        RECT 20.63 29.006 20.682 29.042 ;
        RECT 21.014 29.006 21.068 29.042 ;
        RECT 21.65 29.006 21.704 29.042 ;
        RECT 21.896 29.006 21.95 29.042 ;
        RECT 17.844 29.1635 17.916 29.1885 ;
        RECT 18.356 29.158 18.396 29.194 ;
        RECT 18.664 29.2405 18.736 29.2655 ;
        RECT 18.964 29.2405 19.036 29.2655 ;
        RECT 14.296 29.235 14.35 29.271 ;
        RECT 14.932 29.235 14.986 29.271 ;
        RECT 15.318 29.235 15.37 29.271 ;
        RECT 15.478 29.235 15.53 29.271 ;
        RECT 15.874 29.235 15.926 29.271 ;
        RECT 18.148 29.235 18.188 29.271 ;
        RECT 20.074 29.235 20.126 29.271 ;
        RECT 20.47 29.235 20.522 29.271 ;
        RECT 20.63 29.235 20.682 29.271 ;
        RECT 21.014 29.235 21.068 29.271 ;
        RECT 21.65 29.235 21.704 29.271 ;
        RECT 16.964 29.5345 17.036 29.5595 ;
        RECT 17.844 29.5345 17.916 29.5595 ;
        RECT 18.664 29.5345 18.736 29.5595 ;
        RECT 18.964 29.5345 19.036 29.5595 ;
        RECT 14.05 29.529 14.104 29.565 ;
        RECT 14.932 29.529 14.986 29.565 ;
        RECT 15.318 29.529 15.37 29.565 ;
        RECT 15.478 29.529 15.53 29.565 ;
        RECT 15.874 29.529 15.926 29.565 ;
        RECT 16.034 29.529 16.086 29.565 ;
        RECT 16.8 29.529 16.854 29.565 ;
        RECT 18.148 29.529 18.188 29.565 ;
        RECT 18.356 29.529 18.396 29.565 ;
        RECT 19.914 29.529 19.966 29.565 ;
        RECT 20.074 29.529 20.126 29.565 ;
        RECT 20.47 29.529 20.522 29.565 ;
        RECT 20.63 29.529 20.682 29.565 ;
        RECT 21.014 29.529 21.068 29.565 ;
        RECT 21.896 29.529 21.95 29.565 ;
        RECT 16.964 29.7635 17.036 29.7885 ;
        RECT 18.664 29.7635 18.736 29.7885 ;
        RECT 18.964 29.7635 19.036 29.7885 ;
        RECT 14.05 29.758 14.104 29.794 ;
        RECT 14.296 29.758 14.35 29.794 ;
        RECT 14.932 29.758 14.986 29.794 ;
        RECT 15.318 29.758 15.37 29.794 ;
        RECT 15.478 29.758 15.53 29.794 ;
        RECT 15.874 29.758 15.926 29.794 ;
        RECT 16.034 29.758 16.086 29.794 ;
        RECT 16.8 29.758 16.854 29.794 ;
        RECT 18.148 29.758 18.188 29.794 ;
        RECT 19.914 29.758 19.966 29.794 ;
        RECT 20.074 29.758 20.126 29.794 ;
        RECT 20.47 29.758 20.522 29.794 ;
        RECT 20.63 29.758 20.682 29.794 ;
        RECT 21.014 29.758 21.068 29.794 ;
        RECT 21.65 29.758 21.704 29.794 ;
        RECT 21.896 29.758 21.95 29.794 ;
        RECT 17.844 29.8405 17.916 29.8655 ;
        RECT 18.356 29.835 18.396 29.871 ;
        RECT 16.964 30.2115 17.036 30.2365 ;
        RECT 17.844 30.2115 17.916 30.2365 ;
        RECT 18.964 30.2115 19.036 30.2365 ;
        RECT 14.05 30.206 14.104 30.242 ;
        RECT 14.296 30.206 14.35 30.242 ;
        RECT 14.932 30.206 14.986 30.242 ;
        RECT 15.318 30.206 15.37 30.242 ;
        RECT 15.874 30.206 15.926 30.242 ;
        RECT 16.034 30.206 16.086 30.242 ;
        RECT 18.356 30.206 18.396 30.242 ;
        RECT 19.914 30.206 19.966 30.242 ;
        RECT 20.074 30.206 20.126 30.242 ;
        RECT 20.63 30.206 20.682 30.242 ;
        RECT 21.014 30.206 21.068 30.242 ;
        RECT 21.65 30.206 21.704 30.242 ;
        RECT 21.896 30.206 21.95 30.242 ;
        RECT 17.844 30.3635 17.916 30.3885 ;
        RECT 18.356 30.358 18.396 30.394 ;
        RECT 18.664 30.4405 18.736 30.4655 ;
        RECT 18.964 30.4405 19.036 30.4655 ;
        RECT 14.296 30.435 14.35 30.471 ;
        RECT 14.932 30.435 14.986 30.471 ;
        RECT 15.318 30.435 15.37 30.471 ;
        RECT 15.478 30.435 15.53 30.471 ;
        RECT 15.874 30.435 15.926 30.471 ;
        RECT 18.148 30.435 18.188 30.471 ;
        RECT 20.074 30.435 20.126 30.471 ;
        RECT 20.47 30.435 20.522 30.471 ;
        RECT 20.63 30.435 20.682 30.471 ;
        RECT 21.014 30.435 21.068 30.471 ;
        RECT 21.65 30.435 21.704 30.471 ;
        RECT 16.964 30.7345 17.036 30.7595 ;
        RECT 17.844 30.7345 17.916 30.7595 ;
        RECT 18.664 30.7345 18.736 30.7595 ;
        RECT 18.964 30.7345 19.036 30.7595 ;
        RECT 14.05 30.729 14.104 30.765 ;
        RECT 14.932 30.729 14.986 30.765 ;
        RECT 15.318 30.729 15.37 30.765 ;
        RECT 15.478 30.729 15.53 30.765 ;
        RECT 15.874 30.729 15.926 30.765 ;
        RECT 16.034 30.729 16.086 30.765 ;
        RECT 16.8 30.729 16.854 30.765 ;
        RECT 18.148 30.729 18.188 30.765 ;
        RECT 18.356 30.729 18.396 30.765 ;
        RECT 19.914 30.729 19.966 30.765 ;
        RECT 20.074 30.729 20.126 30.765 ;
        RECT 20.47 30.729 20.522 30.765 ;
        RECT 20.63 30.729 20.682 30.765 ;
        RECT 21.014 30.729 21.068 30.765 ;
        RECT 21.896 30.729 21.95 30.765 ;
        RECT 16.964 30.9635 17.036 30.9885 ;
        RECT 18.664 30.9635 18.736 30.9885 ;
        RECT 18.964 30.9635 19.036 30.9885 ;
        RECT 14.05 30.958 14.104 30.994 ;
        RECT 14.296 30.958 14.35 30.994 ;
        RECT 14.932 30.958 14.986 30.994 ;
        RECT 15.318 30.958 15.37 30.994 ;
        RECT 15.478 30.958 15.53 30.994 ;
        RECT 15.874 30.958 15.926 30.994 ;
        RECT 16.034 30.958 16.086 30.994 ;
        RECT 16.8 30.958 16.854 30.994 ;
        RECT 18.148 30.958 18.188 30.994 ;
        RECT 19.914 30.958 19.966 30.994 ;
        RECT 20.074 30.958 20.126 30.994 ;
        RECT 20.47 30.958 20.522 30.994 ;
        RECT 20.63 30.958 20.682 30.994 ;
        RECT 21.014 30.958 21.068 30.994 ;
        RECT 21.65 30.958 21.704 30.994 ;
        RECT 21.896 30.958 21.95 30.994 ;
        RECT 17.844 31.0405 17.916 31.0655 ;
        RECT 18.356 31.035 18.396 31.071 ;
        RECT 16.964 31.4115 17.036 31.4365 ;
        RECT 17.844 31.4115 17.916 31.4365 ;
        RECT 18.964 31.4115 19.036 31.4365 ;
        RECT 14.05 31.406 14.104 31.442 ;
        RECT 14.296 31.406 14.35 31.442 ;
        RECT 14.932 31.406 14.986 31.442 ;
        RECT 15.318 31.406 15.37 31.442 ;
        RECT 15.874 31.406 15.926 31.442 ;
        RECT 16.034 31.406 16.086 31.442 ;
        RECT 18.356 31.406 18.396 31.442 ;
        RECT 19.914 31.406 19.966 31.442 ;
        RECT 20.074 31.406 20.126 31.442 ;
        RECT 20.63 31.406 20.682 31.442 ;
        RECT 21.014 31.406 21.068 31.442 ;
        RECT 21.65 31.406 21.704 31.442 ;
        RECT 21.896 31.406 21.95 31.442 ;
        RECT 17.844 31.5635 17.916 31.5885 ;
        RECT 18.356 31.558 18.396 31.594 ;
        RECT 18.664 31.6405 18.736 31.6655 ;
        RECT 18.964 31.6405 19.036 31.6655 ;
        RECT 14.296 31.635 14.35 31.671 ;
        RECT 14.932 31.635 14.986 31.671 ;
        RECT 15.318 31.635 15.37 31.671 ;
        RECT 15.478 31.635 15.53 31.671 ;
        RECT 15.874 31.635 15.926 31.671 ;
        RECT 18.148 31.635 18.188 31.671 ;
        RECT 20.074 31.635 20.126 31.671 ;
        RECT 20.47 31.635 20.522 31.671 ;
        RECT 20.63 31.635 20.682 31.671 ;
        RECT 21.014 31.635 21.068 31.671 ;
        RECT 21.65 31.635 21.704 31.671 ;
        RECT 14.05 32.262 14.104 32.298 ;
        RECT 14.296 32.262 14.35 32.298 ;
        RECT 14.932 32.262 14.986 32.298 ;
        RECT 21.014 32.262 21.068 32.298 ;
        RECT 21.65 32.262 21.704 32.298 ;
        RECT 21.896 32.262 21.95 32.298 ;
        RECT 14.296 32.3875 14.35 32.4125 ;
        RECT 16.964 32.3875 17.036 32.4125 ;
        RECT 17.844 32.3875 17.916 32.4125 ;
        RECT 18.664 32.3875 18.736 32.4125 ;
        RECT 18.964 32.3875 19.036 32.4125 ;
        RECT 21.65 32.3875 21.704 32.4125 ;
        RECT 14.05 32.382 14.104 32.418 ;
        RECT 14.932 32.382 14.986 32.418 ;
        RECT 15.318 32.382 15.37 32.418 ;
        RECT 15.478 32.382 15.53 32.418 ;
        RECT 15.874 32.382 15.926 32.418 ;
        RECT 16.034 32.382 16.086 32.418 ;
        RECT 16.8 32.382 16.854 32.418 ;
        RECT 17.412 32.382 17.452 32.418 ;
        RECT 18.148 32.382 18.188 32.418 ;
        RECT 18.356 32.382 18.396 32.418 ;
        RECT 19.31 32.382 19.35 32.418 ;
        RECT 19.914 32.382 19.966 32.418 ;
        RECT 20.074 32.382 20.126 32.418 ;
        RECT 20.47 32.382 20.522 32.418 ;
        RECT 20.63 32.382 20.682 32.418 ;
        RECT 21.014 32.382 21.068 32.418 ;
        RECT 21.896 32.382 21.95 32.418 ;
        RECT 0.974 32.742 1.026 32.778 ;
        RECT 1.774 32.742 1.826 32.778 ;
        RECT 2.574 32.742 2.626 32.778 ;
        RECT 3.374 32.742 3.426 32.778 ;
        RECT 4.174 32.742 4.226 32.778 ;
        RECT 4.974 32.742 5.026 32.778 ;
        RECT 5.774 32.742 5.826 32.778 ;
        RECT 6.574 32.742 6.626 32.778 ;
        RECT 7.374 32.742 7.426 32.778 ;
        RECT 8.174 32.742 8.226 32.778 ;
        RECT 8.974 32.742 9.026 32.778 ;
        RECT 9.774 32.742 9.826 32.778 ;
        RECT 10.574 32.742 10.626 32.778 ;
        RECT 11.374 32.742 11.426 32.778 ;
        RECT 12.174 32.742 12.226 32.778 ;
        RECT 12.974 32.742 13.026 32.778 ;
        RECT 14.05 32.742 14.104 32.778 ;
        RECT 14.296 32.742 14.35 32.778 ;
        RECT 14.932 32.742 14.986 32.778 ;
        RECT 21.014 32.742 21.068 32.778 ;
        RECT 21.65 32.742 21.704 32.778 ;
        RECT 21.896 32.742 21.95 32.778 ;
        RECT 23.174 32.742 23.226 32.778 ;
        RECT 23.974 32.742 24.026 32.778 ;
        RECT 24.774 32.742 24.826 32.778 ;
        RECT 25.574 32.742 25.626 32.778 ;
        RECT 26.374 32.742 26.426 32.778 ;
        RECT 27.174 32.742 27.226 32.778 ;
        RECT 27.974 32.742 28.026 32.778 ;
        RECT 28.774 32.742 28.826 32.778 ;
        RECT 29.574 32.742 29.626 32.778 ;
        RECT 30.374 32.742 30.426 32.778 ;
        RECT 31.174 32.742 31.226 32.778 ;
        RECT 31.974 32.742 32.026 32.778 ;
        RECT 32.774 32.742 32.826 32.778 ;
        RECT 33.574 32.742 33.626 32.778 ;
        RECT 34.374 32.742 34.426 32.778 ;
        RECT 35.174 32.742 35.226 32.778 ;
        RECT 16.964 32.8675 17.036 32.8925 ;
        RECT 18.356 32.8675 18.396 32.8925 ;
        RECT 18.664 32.8675 18.736 32.8925 ;
        RECT 18.964 32.8675 19.036 32.8925 ;
        RECT 14.05 32.862 14.104 32.898 ;
        RECT 14.296 32.862 14.35 32.898 ;
        RECT 14.932 32.862 14.986 32.898 ;
        RECT 15.318 32.862 15.37 32.898 ;
        RECT 15.874 32.862 15.926 32.898 ;
        RECT 16.034 32.862 16.086 32.898 ;
        RECT 16.8 32.862 16.854 32.898 ;
        RECT 17.412 32.862 17.452 32.898 ;
        RECT 18.148 32.862 18.188 32.898 ;
        RECT 19.31 32.862 19.35 32.898 ;
        RECT 19.914 32.862 19.966 32.898 ;
        RECT 20.074 32.862 20.126 32.898 ;
        RECT 20.63 32.862 20.682 32.898 ;
        RECT 21.014 32.862 21.068 32.898 ;
        RECT 21.65 32.862 21.704 32.898 ;
        RECT 21.896 32.862 21.95 32.898 ;
        RECT 0.654 32.982 0.706 33.018 ;
        RECT 0.974 32.982 1.026 33.018 ;
        RECT 1.454 32.982 1.506 33.018 ;
        RECT 1.774 32.982 1.826 33.018 ;
        RECT 2.254 32.982 2.306 33.018 ;
        RECT 2.574 32.982 2.626 33.018 ;
        RECT 3.054 32.982 3.106 33.018 ;
        RECT 3.374 32.982 3.426 33.018 ;
        RECT 3.854 32.982 3.906 33.018 ;
        RECT 4.174 32.982 4.226 33.018 ;
        RECT 4.654 32.982 4.706 33.018 ;
        RECT 4.974 32.982 5.026 33.018 ;
        RECT 5.454 32.982 5.506 33.018 ;
        RECT 5.774 32.982 5.826 33.018 ;
        RECT 6.254 32.982 6.306 33.018 ;
        RECT 6.574 32.982 6.626 33.018 ;
        RECT 7.054 32.982 7.106 33.018 ;
        RECT 7.374 32.982 7.426 33.018 ;
        RECT 7.854 32.982 7.906 33.018 ;
        RECT 8.174 32.982 8.226 33.018 ;
        RECT 8.654 32.982 8.706 33.018 ;
        RECT 8.974 32.982 9.026 33.018 ;
        RECT 9.454 32.982 9.506 33.018 ;
        RECT 9.774 32.982 9.826 33.018 ;
        RECT 10.254 32.982 10.306 33.018 ;
        RECT 10.574 32.982 10.626 33.018 ;
        RECT 11.054 32.982 11.106 33.018 ;
        RECT 11.374 32.982 11.426 33.018 ;
        RECT 11.854 32.982 11.906 33.018 ;
        RECT 12.174 32.982 12.226 33.018 ;
        RECT 12.654 32.982 12.706 33.018 ;
        RECT 12.974 32.982 13.026 33.018 ;
        RECT 14.05 32.982 14.104 33.018 ;
        RECT 14.296 32.982 14.35 33.018 ;
        RECT 14.932 32.982 14.986 33.018 ;
        RECT 21.014 32.982 21.068 33.018 ;
        RECT 21.65 32.982 21.704 33.018 ;
        RECT 21.896 32.982 21.95 33.018 ;
        RECT 22.854 32.982 22.906 33.018 ;
        RECT 23.174 32.982 23.226 33.018 ;
        RECT 23.654 32.982 23.706 33.018 ;
        RECT 23.974 32.982 24.026 33.018 ;
        RECT 24.454 32.982 24.506 33.018 ;
        RECT 24.774 32.982 24.826 33.018 ;
        RECT 25.254 32.982 25.306 33.018 ;
        RECT 25.574 32.982 25.626 33.018 ;
        RECT 26.054 32.982 26.106 33.018 ;
        RECT 26.374 32.982 26.426 33.018 ;
        RECT 26.854 32.982 26.906 33.018 ;
        RECT 27.174 32.982 27.226 33.018 ;
        RECT 27.654 32.982 27.706 33.018 ;
        RECT 27.974 32.982 28.026 33.018 ;
        RECT 28.454 32.982 28.506 33.018 ;
        RECT 28.774 32.982 28.826 33.018 ;
        RECT 29.254 32.982 29.306 33.018 ;
        RECT 29.574 32.982 29.626 33.018 ;
        RECT 30.054 32.982 30.106 33.018 ;
        RECT 30.374 32.982 30.426 33.018 ;
        RECT 30.854 32.982 30.906 33.018 ;
        RECT 31.174 32.982 31.226 33.018 ;
        RECT 31.654 32.982 31.706 33.018 ;
        RECT 31.974 32.982 32.026 33.018 ;
        RECT 32.454 32.982 32.506 33.018 ;
        RECT 32.774 32.982 32.826 33.018 ;
        RECT 33.254 32.982 33.306 33.018 ;
        RECT 33.574 32.982 33.626 33.018 ;
        RECT 34.054 32.982 34.106 33.018 ;
        RECT 34.374 32.982 34.426 33.018 ;
        RECT 34.854 32.982 34.906 33.018 ;
        RECT 35.174 32.982 35.226 33.018 ;
        RECT 16.964 33.049 17.036 33.074 ;
        RECT 17.844 33.049 17.916 33.074 ;
        RECT 18.664 33.049 18.736 33.074 ;
        RECT 15.318 33.0435 15.37 33.0795 ;
        RECT 16.8 33.0435 16.854 33.0795 ;
        RECT 17.412 33.0435 17.452 33.0795 ;
        RECT 18.356 33.0435 18.396 33.0795 ;
        RECT 20.63 33.0435 20.682 33.0795 ;
        RECT 16.964 33.3475 17.036 33.3725 ;
        RECT 17.844 33.3475 17.916 33.3725 ;
        RECT 18.664 33.3475 18.736 33.3725 ;
        RECT 18.964 33.3475 19.036 33.3725 ;
        RECT 14.05 33.342 14.104 33.378 ;
        RECT 14.296 33.342 14.35 33.378 ;
        RECT 15.318 33.342 15.37 33.378 ;
        RECT 15.874 33.342 15.926 33.378 ;
        RECT 16.034 33.342 16.086 33.378 ;
        RECT 16.8 33.342 16.854 33.378 ;
        RECT 17.412 33.342 17.452 33.378 ;
        RECT 18.148 33.342 18.188 33.378 ;
        RECT 18.356 33.342 18.396 33.378 ;
        RECT 19.31 33.342 19.35 33.378 ;
        RECT 19.914 33.342 19.966 33.378 ;
        RECT 20.074 33.342 20.126 33.378 ;
        RECT 20.63 33.342 20.682 33.378 ;
        RECT 21.65 33.342 21.704 33.378 ;
        RECT 21.896 33.342 21.95 33.378 ;
        RECT 0.654 33.462 0.706 33.498 ;
        RECT 0.974 33.462 1.026 33.498 ;
        RECT 1.454 33.462 1.506 33.498 ;
        RECT 1.774 33.462 1.826 33.498 ;
        RECT 2.254 33.462 2.306 33.498 ;
        RECT 2.574 33.462 2.626 33.498 ;
        RECT 3.054 33.462 3.106 33.498 ;
        RECT 3.374 33.462 3.426 33.498 ;
        RECT 3.854 33.462 3.906 33.498 ;
        RECT 4.174 33.462 4.226 33.498 ;
        RECT 4.654 33.462 4.706 33.498 ;
        RECT 4.974 33.462 5.026 33.498 ;
        RECT 5.454 33.462 5.506 33.498 ;
        RECT 5.774 33.462 5.826 33.498 ;
        RECT 6.254 33.462 6.306 33.498 ;
        RECT 6.574 33.462 6.626 33.498 ;
        RECT 7.054 33.462 7.106 33.498 ;
        RECT 7.374 33.462 7.426 33.498 ;
        RECT 7.854 33.462 7.906 33.498 ;
        RECT 8.174 33.462 8.226 33.498 ;
        RECT 8.654 33.462 8.706 33.498 ;
        RECT 8.974 33.462 9.026 33.498 ;
        RECT 9.454 33.462 9.506 33.498 ;
        RECT 9.774 33.462 9.826 33.498 ;
        RECT 10.254 33.462 10.306 33.498 ;
        RECT 10.574 33.462 10.626 33.498 ;
        RECT 11.054 33.462 11.106 33.498 ;
        RECT 11.374 33.462 11.426 33.498 ;
        RECT 11.854 33.462 11.906 33.498 ;
        RECT 12.174 33.462 12.226 33.498 ;
        RECT 12.654 33.462 12.706 33.498 ;
        RECT 12.974 33.462 13.026 33.498 ;
        RECT 14.05 33.462 14.104 33.498 ;
        RECT 14.296 33.462 14.35 33.498 ;
        RECT 14.932 33.462 14.986 33.498 ;
        RECT 21.014 33.462 21.068 33.498 ;
        RECT 21.65 33.462 21.704 33.498 ;
        RECT 21.896 33.462 21.95 33.498 ;
        RECT 22.854 33.462 22.906 33.498 ;
        RECT 23.174 33.462 23.226 33.498 ;
        RECT 23.654 33.462 23.706 33.498 ;
        RECT 23.974 33.462 24.026 33.498 ;
        RECT 24.454 33.462 24.506 33.498 ;
        RECT 24.774 33.462 24.826 33.498 ;
        RECT 25.254 33.462 25.306 33.498 ;
        RECT 25.574 33.462 25.626 33.498 ;
        RECT 26.054 33.462 26.106 33.498 ;
        RECT 26.374 33.462 26.426 33.498 ;
        RECT 26.854 33.462 26.906 33.498 ;
        RECT 27.174 33.462 27.226 33.498 ;
        RECT 27.654 33.462 27.706 33.498 ;
        RECT 27.974 33.462 28.026 33.498 ;
        RECT 28.454 33.462 28.506 33.498 ;
        RECT 28.774 33.462 28.826 33.498 ;
        RECT 29.254 33.462 29.306 33.498 ;
        RECT 29.574 33.462 29.626 33.498 ;
        RECT 30.054 33.462 30.106 33.498 ;
        RECT 30.374 33.462 30.426 33.498 ;
        RECT 30.854 33.462 30.906 33.498 ;
        RECT 31.174 33.462 31.226 33.498 ;
        RECT 31.654 33.462 31.706 33.498 ;
        RECT 31.974 33.462 32.026 33.498 ;
        RECT 32.454 33.462 32.506 33.498 ;
        RECT 32.774 33.462 32.826 33.498 ;
        RECT 33.254 33.462 33.306 33.498 ;
        RECT 33.574 33.462 33.626 33.498 ;
        RECT 34.054 33.462 34.106 33.498 ;
        RECT 34.374 33.462 34.426 33.498 ;
        RECT 34.854 33.462 34.906 33.498 ;
        RECT 35.174 33.462 35.226 33.498 ;
        RECT 0.654 33.702 0.706 33.738 ;
        RECT 0.974 33.702 1.026 33.738 ;
        RECT 1.454 33.702 1.506 33.738 ;
        RECT 1.774 33.702 1.826 33.738 ;
        RECT 2.254 33.702 2.306 33.738 ;
        RECT 2.574 33.702 2.626 33.738 ;
        RECT 3.054 33.702 3.106 33.738 ;
        RECT 3.374 33.702 3.426 33.738 ;
        RECT 3.854 33.702 3.906 33.738 ;
        RECT 4.174 33.702 4.226 33.738 ;
        RECT 4.654 33.702 4.706 33.738 ;
        RECT 4.974 33.702 5.026 33.738 ;
        RECT 5.454 33.702 5.506 33.738 ;
        RECT 5.774 33.702 5.826 33.738 ;
        RECT 6.254 33.702 6.306 33.738 ;
        RECT 6.574 33.702 6.626 33.738 ;
        RECT 7.054 33.702 7.106 33.738 ;
        RECT 7.374 33.702 7.426 33.738 ;
        RECT 7.854 33.702 7.906 33.738 ;
        RECT 8.174 33.702 8.226 33.738 ;
        RECT 8.654 33.702 8.706 33.738 ;
        RECT 8.974 33.702 9.026 33.738 ;
        RECT 9.454 33.702 9.506 33.738 ;
        RECT 9.774 33.702 9.826 33.738 ;
        RECT 10.254 33.702 10.306 33.738 ;
        RECT 10.574 33.702 10.626 33.738 ;
        RECT 11.054 33.702 11.106 33.738 ;
        RECT 11.374 33.702 11.426 33.738 ;
        RECT 11.854 33.702 11.906 33.738 ;
        RECT 12.174 33.702 12.226 33.738 ;
        RECT 12.654 33.702 12.706 33.738 ;
        RECT 12.974 33.702 13.026 33.738 ;
        RECT 22.854 33.702 22.906 33.738 ;
        RECT 23.174 33.702 23.226 33.738 ;
        RECT 23.654 33.702 23.706 33.738 ;
        RECT 23.974 33.702 24.026 33.738 ;
        RECT 24.454 33.702 24.506 33.738 ;
        RECT 24.774 33.702 24.826 33.738 ;
        RECT 25.254 33.702 25.306 33.738 ;
        RECT 25.574 33.702 25.626 33.738 ;
        RECT 26.054 33.702 26.106 33.738 ;
        RECT 26.374 33.702 26.426 33.738 ;
        RECT 26.854 33.702 26.906 33.738 ;
        RECT 27.174 33.702 27.226 33.738 ;
        RECT 27.654 33.702 27.706 33.738 ;
        RECT 27.974 33.702 28.026 33.738 ;
        RECT 28.454 33.702 28.506 33.738 ;
        RECT 28.774 33.702 28.826 33.738 ;
        RECT 29.254 33.702 29.306 33.738 ;
        RECT 29.574 33.702 29.626 33.738 ;
        RECT 30.054 33.702 30.106 33.738 ;
        RECT 30.374 33.702 30.426 33.738 ;
        RECT 30.854 33.702 30.906 33.738 ;
        RECT 31.174 33.702 31.226 33.738 ;
        RECT 31.654 33.702 31.706 33.738 ;
        RECT 31.974 33.702 32.026 33.738 ;
        RECT 32.454 33.702 32.506 33.738 ;
        RECT 32.774 33.702 32.826 33.738 ;
        RECT 33.254 33.702 33.306 33.738 ;
        RECT 33.574 33.702 33.626 33.738 ;
        RECT 34.054 33.702 34.106 33.738 ;
        RECT 34.374 33.702 34.426 33.738 ;
        RECT 34.854 33.702 34.906 33.738 ;
        RECT 35.174 33.702 35.226 33.738 ;
        RECT 16.964 33.8275 17.036 33.8525 ;
        RECT 17.844 33.8275 17.916 33.8525 ;
        RECT 18.664 33.8275 18.736 33.8525 ;
        RECT 18.964 33.8275 19.036 33.8525 ;
        RECT 14.05 33.822 14.104 33.858 ;
        RECT 14.296 33.822 14.35 33.858 ;
        RECT 14.932 33.822 14.986 33.858 ;
        RECT 15.318 33.822 15.37 33.858 ;
        RECT 15.874 33.822 15.926 33.858 ;
        RECT 16.034 33.822 16.086 33.858 ;
        RECT 16.8 33.822 16.854 33.858 ;
        RECT 17.412 33.822 17.452 33.858 ;
        RECT 18.148 33.822 18.188 33.858 ;
        RECT 18.356 33.822 18.396 33.858 ;
        RECT 19.31 33.822 19.35 33.858 ;
        RECT 19.914 33.822 19.966 33.858 ;
        RECT 20.074 33.822 20.126 33.858 ;
        RECT 20.63 33.822 20.682 33.858 ;
        RECT 21.014 33.822 21.068 33.858 ;
        RECT 21.65 33.822 21.704 33.858 ;
        RECT 21.896 33.822 21.95 33.858 ;
        RECT 0.654 34.182 0.706 34.218 ;
        RECT 0.974 34.182 1.026 34.218 ;
        RECT 1.454 34.182 1.506 34.218 ;
        RECT 1.774 34.182 1.826 34.218 ;
        RECT 2.254 34.182 2.306 34.218 ;
        RECT 2.574 34.182 2.626 34.218 ;
        RECT 3.054 34.182 3.106 34.218 ;
        RECT 3.374 34.182 3.426 34.218 ;
        RECT 3.854 34.182 3.906 34.218 ;
        RECT 4.174 34.182 4.226 34.218 ;
        RECT 4.654 34.182 4.706 34.218 ;
        RECT 4.974 34.182 5.026 34.218 ;
        RECT 5.454 34.182 5.506 34.218 ;
        RECT 5.774 34.182 5.826 34.218 ;
        RECT 6.254 34.182 6.306 34.218 ;
        RECT 6.574 34.182 6.626 34.218 ;
        RECT 7.054 34.182 7.106 34.218 ;
        RECT 7.374 34.182 7.426 34.218 ;
        RECT 7.854 34.182 7.906 34.218 ;
        RECT 8.174 34.182 8.226 34.218 ;
        RECT 8.654 34.182 8.706 34.218 ;
        RECT 8.974 34.182 9.026 34.218 ;
        RECT 9.454 34.182 9.506 34.218 ;
        RECT 9.774 34.182 9.826 34.218 ;
        RECT 10.254 34.182 10.306 34.218 ;
        RECT 10.574 34.182 10.626 34.218 ;
        RECT 11.054 34.182 11.106 34.218 ;
        RECT 11.374 34.182 11.426 34.218 ;
        RECT 11.854 34.182 11.906 34.218 ;
        RECT 12.174 34.182 12.226 34.218 ;
        RECT 12.654 34.182 12.706 34.218 ;
        RECT 12.974 34.182 13.026 34.218 ;
        RECT 22.854 34.182 22.906 34.218 ;
        RECT 23.174 34.182 23.226 34.218 ;
        RECT 23.654 34.182 23.706 34.218 ;
        RECT 23.974 34.182 24.026 34.218 ;
        RECT 24.454 34.182 24.506 34.218 ;
        RECT 24.774 34.182 24.826 34.218 ;
        RECT 25.254 34.182 25.306 34.218 ;
        RECT 25.574 34.182 25.626 34.218 ;
        RECT 26.054 34.182 26.106 34.218 ;
        RECT 26.374 34.182 26.426 34.218 ;
        RECT 26.854 34.182 26.906 34.218 ;
        RECT 27.174 34.182 27.226 34.218 ;
        RECT 27.654 34.182 27.706 34.218 ;
        RECT 27.974 34.182 28.026 34.218 ;
        RECT 28.454 34.182 28.506 34.218 ;
        RECT 28.774 34.182 28.826 34.218 ;
        RECT 29.254 34.182 29.306 34.218 ;
        RECT 29.574 34.182 29.626 34.218 ;
        RECT 30.054 34.182 30.106 34.218 ;
        RECT 30.374 34.182 30.426 34.218 ;
        RECT 30.854 34.182 30.906 34.218 ;
        RECT 31.174 34.182 31.226 34.218 ;
        RECT 31.654 34.182 31.706 34.218 ;
        RECT 31.974 34.182 32.026 34.218 ;
        RECT 32.454 34.182 32.506 34.218 ;
        RECT 32.774 34.182 32.826 34.218 ;
        RECT 33.254 34.182 33.306 34.218 ;
        RECT 33.574 34.182 33.626 34.218 ;
        RECT 34.054 34.182 34.106 34.218 ;
        RECT 34.374 34.182 34.426 34.218 ;
        RECT 34.854 34.182 34.906 34.218 ;
        RECT 35.174 34.182 35.226 34.218 ;
        RECT 16.034 34.3075 16.086 34.3325 ;
        RECT 16.964 34.3075 17.036 34.3325 ;
        RECT 17.844 34.3075 17.916 34.3325 ;
        RECT 18.664 34.3075 18.736 34.3325 ;
        RECT 18.964 34.3075 19.036 34.3325 ;
        RECT 19.914 34.3075 19.966 34.3325 ;
        RECT 0.654 34.302 0.706 34.338 ;
        RECT 0.974 34.302 1.026 34.338 ;
        RECT 1.454 34.302 1.506 34.338 ;
        RECT 1.774 34.302 1.826 34.338 ;
        RECT 2.254 34.302 2.306 34.338 ;
        RECT 2.574 34.302 2.626 34.338 ;
        RECT 3.054 34.302 3.106 34.338 ;
        RECT 3.374 34.302 3.426 34.338 ;
        RECT 3.854 34.302 3.906 34.338 ;
        RECT 4.174 34.302 4.226 34.338 ;
        RECT 4.654 34.302 4.706 34.338 ;
        RECT 4.974 34.302 5.026 34.338 ;
        RECT 5.454 34.302 5.506 34.338 ;
        RECT 5.774 34.302 5.826 34.338 ;
        RECT 6.254 34.302 6.306 34.338 ;
        RECT 6.574 34.302 6.626 34.338 ;
        RECT 7.054 34.302 7.106 34.338 ;
        RECT 7.374 34.302 7.426 34.338 ;
        RECT 7.854 34.302 7.906 34.338 ;
        RECT 8.174 34.302 8.226 34.338 ;
        RECT 8.654 34.302 8.706 34.338 ;
        RECT 8.974 34.302 9.026 34.338 ;
        RECT 9.454 34.302 9.506 34.338 ;
        RECT 9.774 34.302 9.826 34.338 ;
        RECT 10.254 34.302 10.306 34.338 ;
        RECT 10.574 34.302 10.626 34.338 ;
        RECT 11.054 34.302 11.106 34.338 ;
        RECT 11.374 34.302 11.426 34.338 ;
        RECT 11.854 34.302 11.906 34.338 ;
        RECT 12.174 34.302 12.226 34.338 ;
        RECT 12.654 34.302 12.706 34.338 ;
        RECT 12.974 34.302 13.026 34.338 ;
        RECT 14.296 34.302 14.35 34.338 ;
        RECT 14.932 34.302 14.986 34.338 ;
        RECT 15.318 34.302 15.37 34.338 ;
        RECT 15.874 34.302 15.926 34.338 ;
        RECT 16.8 34.302 16.854 34.338 ;
        RECT 17.412 34.302 17.452 34.338 ;
        RECT 18.148 34.302 18.188 34.338 ;
        RECT 18.356 34.302 18.396 34.338 ;
        RECT 19.31 34.302 19.35 34.338 ;
        RECT 20.074 34.302 20.126 34.338 ;
        RECT 20.63 34.302 20.682 34.338 ;
        RECT 21.014 34.302 21.068 34.338 ;
        RECT 21.65 34.302 21.704 34.338 ;
        RECT 22.854 34.302 22.906 34.338 ;
        RECT 23.174 34.302 23.226 34.338 ;
        RECT 23.654 34.302 23.706 34.338 ;
        RECT 23.974 34.302 24.026 34.338 ;
        RECT 24.454 34.302 24.506 34.338 ;
        RECT 24.774 34.302 24.826 34.338 ;
        RECT 25.254 34.302 25.306 34.338 ;
        RECT 25.574 34.302 25.626 34.338 ;
        RECT 26.054 34.302 26.106 34.338 ;
        RECT 26.374 34.302 26.426 34.338 ;
        RECT 26.854 34.302 26.906 34.338 ;
        RECT 27.174 34.302 27.226 34.338 ;
        RECT 27.654 34.302 27.706 34.338 ;
        RECT 27.974 34.302 28.026 34.338 ;
        RECT 28.454 34.302 28.506 34.338 ;
        RECT 28.774 34.302 28.826 34.338 ;
        RECT 29.254 34.302 29.306 34.338 ;
        RECT 29.574 34.302 29.626 34.338 ;
        RECT 30.054 34.302 30.106 34.338 ;
        RECT 30.374 34.302 30.426 34.338 ;
        RECT 30.854 34.302 30.906 34.338 ;
        RECT 31.174 34.302 31.226 34.338 ;
        RECT 31.654 34.302 31.706 34.338 ;
        RECT 31.974 34.302 32.026 34.338 ;
        RECT 32.454 34.302 32.506 34.338 ;
        RECT 32.774 34.302 32.826 34.338 ;
        RECT 33.254 34.302 33.306 34.338 ;
        RECT 33.574 34.302 33.626 34.338 ;
        RECT 34.054 34.302 34.106 34.338 ;
        RECT 34.374 34.302 34.426 34.338 ;
        RECT 34.854 34.302 34.906 34.338 ;
        RECT 35.174 34.302 35.226 34.338 ;
        RECT 14.05 34.7875 14.104 34.8125 ;
        RECT 16.964 34.7875 17.036 34.8125 ;
        RECT 17.844 34.7875 17.916 34.8125 ;
        RECT 18.664 34.7875 18.736 34.8125 ;
        RECT 18.964 34.7875 19.036 34.8125 ;
        RECT 21.896 34.7875 21.95 34.8125 ;
        RECT 0.654 34.782 0.706 34.818 ;
        RECT 0.974 34.782 1.026 34.818 ;
        RECT 1.454 34.782 1.506 34.818 ;
        RECT 1.774 34.782 1.826 34.818 ;
        RECT 2.254 34.782 2.306 34.818 ;
        RECT 2.574 34.782 2.626 34.818 ;
        RECT 3.054 34.782 3.106 34.818 ;
        RECT 3.374 34.782 3.426 34.818 ;
        RECT 3.854 34.782 3.906 34.818 ;
        RECT 4.174 34.782 4.226 34.818 ;
        RECT 4.654 34.782 4.706 34.818 ;
        RECT 4.974 34.782 5.026 34.818 ;
        RECT 5.454 34.782 5.506 34.818 ;
        RECT 5.774 34.782 5.826 34.818 ;
        RECT 6.254 34.782 6.306 34.818 ;
        RECT 6.574 34.782 6.626 34.818 ;
        RECT 7.054 34.782 7.106 34.818 ;
        RECT 7.374 34.782 7.426 34.818 ;
        RECT 7.854 34.782 7.906 34.818 ;
        RECT 8.174 34.782 8.226 34.818 ;
        RECT 8.654 34.782 8.706 34.818 ;
        RECT 8.974 34.782 9.026 34.818 ;
        RECT 9.454 34.782 9.506 34.818 ;
        RECT 9.774 34.782 9.826 34.818 ;
        RECT 10.254 34.782 10.306 34.818 ;
        RECT 10.574 34.782 10.626 34.818 ;
        RECT 11.054 34.782 11.106 34.818 ;
        RECT 11.374 34.782 11.426 34.818 ;
        RECT 11.854 34.782 11.906 34.818 ;
        RECT 12.174 34.782 12.226 34.818 ;
        RECT 12.654 34.782 12.706 34.818 ;
        RECT 12.974 34.782 13.026 34.818 ;
        RECT 14.296 34.782 14.35 34.818 ;
        RECT 14.932 34.782 14.986 34.818 ;
        RECT 15.318 34.782 15.37 34.818 ;
        RECT 15.874 34.782 15.926 34.818 ;
        RECT 16.034 34.782 16.086 34.818 ;
        RECT 16.8 34.782 16.854 34.818 ;
        RECT 17.412 34.782 17.452 34.818 ;
        RECT 18.148 34.782 18.188 34.818 ;
        RECT 18.356 34.782 18.396 34.818 ;
        RECT 19.31 34.782 19.35 34.818 ;
        RECT 19.914 34.782 19.966 34.818 ;
        RECT 20.074 34.782 20.126 34.818 ;
        RECT 20.63 34.782 20.682 34.818 ;
        RECT 21.014 34.782 21.068 34.818 ;
        RECT 21.65 34.782 21.704 34.818 ;
        RECT 22.854 34.782 22.906 34.818 ;
        RECT 23.174 34.782 23.226 34.818 ;
        RECT 23.654 34.782 23.706 34.818 ;
        RECT 23.974 34.782 24.026 34.818 ;
        RECT 24.454 34.782 24.506 34.818 ;
        RECT 24.774 34.782 24.826 34.818 ;
        RECT 25.254 34.782 25.306 34.818 ;
        RECT 25.574 34.782 25.626 34.818 ;
        RECT 26.054 34.782 26.106 34.818 ;
        RECT 26.374 34.782 26.426 34.818 ;
        RECT 26.854 34.782 26.906 34.818 ;
        RECT 27.174 34.782 27.226 34.818 ;
        RECT 27.654 34.782 27.706 34.818 ;
        RECT 27.974 34.782 28.026 34.818 ;
        RECT 28.454 34.782 28.506 34.818 ;
        RECT 28.774 34.782 28.826 34.818 ;
        RECT 29.254 34.782 29.306 34.818 ;
        RECT 29.574 34.782 29.626 34.818 ;
        RECT 30.054 34.782 30.106 34.818 ;
        RECT 30.374 34.782 30.426 34.818 ;
        RECT 30.854 34.782 30.906 34.818 ;
        RECT 31.174 34.782 31.226 34.818 ;
        RECT 31.654 34.782 31.706 34.818 ;
        RECT 31.974 34.782 32.026 34.818 ;
        RECT 32.454 34.782 32.506 34.818 ;
        RECT 32.774 34.782 32.826 34.818 ;
        RECT 33.254 34.782 33.306 34.818 ;
        RECT 33.574 34.782 33.626 34.818 ;
        RECT 34.054 34.782 34.106 34.818 ;
        RECT 34.374 34.782 34.426 34.818 ;
        RECT 34.854 34.782 34.906 34.818 ;
        RECT 35.174 34.782 35.226 34.818 ;
        RECT 16.964 35.2675 17.036 35.2925 ;
        RECT 17.844 35.2675 17.916 35.2925 ;
        RECT 18.664 35.2675 18.736 35.2925 ;
        RECT 18.964 35.2675 19.036 35.2925 ;
        RECT 0.654 35.262 0.706 35.298 ;
        RECT 0.974 35.262 1.026 35.298 ;
        RECT 1.454 35.262 1.506 35.298 ;
        RECT 1.774 35.262 1.826 35.298 ;
        RECT 2.254 35.262 2.306 35.298 ;
        RECT 2.574 35.262 2.626 35.298 ;
        RECT 3.054 35.262 3.106 35.298 ;
        RECT 3.374 35.262 3.426 35.298 ;
        RECT 3.854 35.262 3.906 35.298 ;
        RECT 4.174 35.262 4.226 35.298 ;
        RECT 4.654 35.262 4.706 35.298 ;
        RECT 4.974 35.262 5.026 35.298 ;
        RECT 5.454 35.262 5.506 35.298 ;
        RECT 5.774 35.262 5.826 35.298 ;
        RECT 6.254 35.262 6.306 35.298 ;
        RECT 6.574 35.262 6.626 35.298 ;
        RECT 7.054 35.262 7.106 35.298 ;
        RECT 7.374 35.262 7.426 35.298 ;
        RECT 7.854 35.262 7.906 35.298 ;
        RECT 8.174 35.262 8.226 35.298 ;
        RECT 8.654 35.262 8.706 35.298 ;
        RECT 8.974 35.262 9.026 35.298 ;
        RECT 9.454 35.262 9.506 35.298 ;
        RECT 9.774 35.262 9.826 35.298 ;
        RECT 10.254 35.262 10.306 35.298 ;
        RECT 10.574 35.262 10.626 35.298 ;
        RECT 11.054 35.262 11.106 35.298 ;
        RECT 11.374 35.262 11.426 35.298 ;
        RECT 11.854 35.262 11.906 35.298 ;
        RECT 12.174 35.262 12.226 35.298 ;
        RECT 12.654 35.262 12.706 35.298 ;
        RECT 12.974 35.262 13.026 35.298 ;
        RECT 14.05 35.262 14.104 35.298 ;
        RECT 14.296 35.262 14.35 35.298 ;
        RECT 14.932 35.262 14.986 35.298 ;
        RECT 15.318 35.262 15.37 35.298 ;
        RECT 15.874 35.262 15.926 35.298 ;
        RECT 16.034 35.262 16.086 35.298 ;
        RECT 16.8 35.262 16.854 35.298 ;
        RECT 17.412 35.262 17.452 35.298 ;
        RECT 18.148 35.262 18.188 35.298 ;
        RECT 18.356 35.262 18.396 35.298 ;
        RECT 19.31 35.262 19.35 35.298 ;
        RECT 19.914 35.262 19.966 35.298 ;
        RECT 20.074 35.262 20.126 35.298 ;
        RECT 20.63 35.262 20.682 35.298 ;
        RECT 21.014 35.262 21.068 35.298 ;
        RECT 21.65 35.262 21.704 35.298 ;
        RECT 21.896 35.262 21.95 35.298 ;
        RECT 22.854 35.262 22.906 35.298 ;
        RECT 23.174 35.262 23.226 35.298 ;
        RECT 23.654 35.262 23.706 35.298 ;
        RECT 23.974 35.262 24.026 35.298 ;
        RECT 24.454 35.262 24.506 35.298 ;
        RECT 24.774 35.262 24.826 35.298 ;
        RECT 25.254 35.262 25.306 35.298 ;
        RECT 25.574 35.262 25.626 35.298 ;
        RECT 26.054 35.262 26.106 35.298 ;
        RECT 26.374 35.262 26.426 35.298 ;
        RECT 26.854 35.262 26.906 35.298 ;
        RECT 27.174 35.262 27.226 35.298 ;
        RECT 27.654 35.262 27.706 35.298 ;
        RECT 27.974 35.262 28.026 35.298 ;
        RECT 28.454 35.262 28.506 35.298 ;
        RECT 28.774 35.262 28.826 35.298 ;
        RECT 29.254 35.262 29.306 35.298 ;
        RECT 29.574 35.262 29.626 35.298 ;
        RECT 30.054 35.262 30.106 35.298 ;
        RECT 30.374 35.262 30.426 35.298 ;
        RECT 30.854 35.262 30.906 35.298 ;
        RECT 31.174 35.262 31.226 35.298 ;
        RECT 31.654 35.262 31.706 35.298 ;
        RECT 31.974 35.262 32.026 35.298 ;
        RECT 32.454 35.262 32.506 35.298 ;
        RECT 32.774 35.262 32.826 35.298 ;
        RECT 33.254 35.262 33.306 35.298 ;
        RECT 33.574 35.262 33.626 35.298 ;
        RECT 34.054 35.262 34.106 35.298 ;
        RECT 34.374 35.262 34.426 35.298 ;
        RECT 34.854 35.262 34.906 35.298 ;
        RECT 35.174 35.262 35.226 35.298 ;
        RECT 0.654 35.382 0.706 35.418 ;
        RECT 0.974 35.382 1.026 35.418 ;
        RECT 1.454 35.382 1.506 35.418 ;
        RECT 1.774 35.382 1.826 35.418 ;
        RECT 2.254 35.382 2.306 35.418 ;
        RECT 2.574 35.382 2.626 35.418 ;
        RECT 3.054 35.382 3.106 35.418 ;
        RECT 3.374 35.382 3.426 35.418 ;
        RECT 3.854 35.382 3.906 35.418 ;
        RECT 4.174 35.382 4.226 35.418 ;
        RECT 4.654 35.382 4.706 35.418 ;
        RECT 4.974 35.382 5.026 35.418 ;
        RECT 5.454 35.382 5.506 35.418 ;
        RECT 5.774 35.382 5.826 35.418 ;
        RECT 6.254 35.382 6.306 35.418 ;
        RECT 6.574 35.382 6.626 35.418 ;
        RECT 7.054 35.382 7.106 35.418 ;
        RECT 7.374 35.382 7.426 35.418 ;
        RECT 7.854 35.382 7.906 35.418 ;
        RECT 8.174 35.382 8.226 35.418 ;
        RECT 8.654 35.382 8.706 35.418 ;
        RECT 8.974 35.382 9.026 35.418 ;
        RECT 9.454 35.382 9.506 35.418 ;
        RECT 9.774 35.382 9.826 35.418 ;
        RECT 10.254 35.382 10.306 35.418 ;
        RECT 10.574 35.382 10.626 35.418 ;
        RECT 11.054 35.382 11.106 35.418 ;
        RECT 11.374 35.382 11.426 35.418 ;
        RECT 11.854 35.382 11.906 35.418 ;
        RECT 12.174 35.382 12.226 35.418 ;
        RECT 12.654 35.382 12.706 35.418 ;
        RECT 12.974 35.382 13.026 35.418 ;
        RECT 14.05 35.382 14.104 35.418 ;
        RECT 14.296 35.382 14.35 35.418 ;
        RECT 14.932 35.382 14.986 35.418 ;
        RECT 21.014 35.382 21.068 35.418 ;
        RECT 21.65 35.382 21.704 35.418 ;
        RECT 21.896 35.382 21.95 35.418 ;
        RECT 22.854 35.382 22.906 35.418 ;
        RECT 23.174 35.382 23.226 35.418 ;
        RECT 23.654 35.382 23.706 35.418 ;
        RECT 23.974 35.382 24.026 35.418 ;
        RECT 24.454 35.382 24.506 35.418 ;
        RECT 24.774 35.382 24.826 35.418 ;
        RECT 25.254 35.382 25.306 35.418 ;
        RECT 25.574 35.382 25.626 35.418 ;
        RECT 26.054 35.382 26.106 35.418 ;
        RECT 26.374 35.382 26.426 35.418 ;
        RECT 26.854 35.382 26.906 35.418 ;
        RECT 27.174 35.382 27.226 35.418 ;
        RECT 27.654 35.382 27.706 35.418 ;
        RECT 27.974 35.382 28.026 35.418 ;
        RECT 28.454 35.382 28.506 35.418 ;
        RECT 28.774 35.382 28.826 35.418 ;
        RECT 29.254 35.382 29.306 35.418 ;
        RECT 29.574 35.382 29.626 35.418 ;
        RECT 30.054 35.382 30.106 35.418 ;
        RECT 30.374 35.382 30.426 35.418 ;
        RECT 30.854 35.382 30.906 35.418 ;
        RECT 31.174 35.382 31.226 35.418 ;
        RECT 31.654 35.382 31.706 35.418 ;
        RECT 31.974 35.382 32.026 35.418 ;
        RECT 32.454 35.382 32.506 35.418 ;
        RECT 32.774 35.382 32.826 35.418 ;
        RECT 33.254 35.382 33.306 35.418 ;
        RECT 33.574 35.382 33.626 35.418 ;
        RECT 34.054 35.382 34.106 35.418 ;
        RECT 34.374 35.382 34.426 35.418 ;
        RECT 34.854 35.382 34.906 35.418 ;
        RECT 35.174 35.382 35.226 35.418 ;
        RECT 16.964 35.7475 17.036 35.7725 ;
        RECT 17.844 35.7475 17.916 35.7725 ;
        RECT 18.664 35.7475 18.736 35.7725 ;
        RECT 18.964 35.7475 19.036 35.7725 ;
        RECT 0.654 35.742 0.706 35.778 ;
        RECT 0.974 35.742 1.026 35.778 ;
        RECT 1.454 35.742 1.506 35.778 ;
        RECT 1.774 35.742 1.826 35.778 ;
        RECT 2.254 35.742 2.306 35.778 ;
        RECT 2.574 35.742 2.626 35.778 ;
        RECT 3.054 35.742 3.106 35.778 ;
        RECT 3.374 35.742 3.426 35.778 ;
        RECT 3.854 35.742 3.906 35.778 ;
        RECT 4.174 35.742 4.226 35.778 ;
        RECT 4.654 35.742 4.706 35.778 ;
        RECT 4.974 35.742 5.026 35.778 ;
        RECT 5.454 35.742 5.506 35.778 ;
        RECT 5.774 35.742 5.826 35.778 ;
        RECT 6.254 35.742 6.306 35.778 ;
        RECT 6.574 35.742 6.626 35.778 ;
        RECT 7.054 35.742 7.106 35.778 ;
        RECT 7.374 35.742 7.426 35.778 ;
        RECT 7.854 35.742 7.906 35.778 ;
        RECT 8.174 35.742 8.226 35.778 ;
        RECT 8.654 35.742 8.706 35.778 ;
        RECT 8.974 35.742 9.026 35.778 ;
        RECT 9.454 35.742 9.506 35.778 ;
        RECT 9.774 35.742 9.826 35.778 ;
        RECT 10.254 35.742 10.306 35.778 ;
        RECT 10.574 35.742 10.626 35.778 ;
        RECT 11.054 35.742 11.106 35.778 ;
        RECT 11.374 35.742 11.426 35.778 ;
        RECT 11.854 35.742 11.906 35.778 ;
        RECT 12.174 35.742 12.226 35.778 ;
        RECT 12.654 35.742 12.706 35.778 ;
        RECT 12.974 35.742 13.026 35.778 ;
        RECT 14.05 35.742 14.104 35.778 ;
        RECT 14.296 35.742 14.35 35.778 ;
        RECT 14.932 35.742 14.986 35.778 ;
        RECT 15.318 35.742 15.37 35.778 ;
        RECT 15.874 35.742 15.926 35.778 ;
        RECT 16.034 35.742 16.086 35.778 ;
        RECT 16.8 35.742 16.854 35.778 ;
        RECT 17.412 35.742 17.452 35.778 ;
        RECT 18.148 35.742 18.188 35.778 ;
        RECT 18.356 35.742 18.396 35.778 ;
        RECT 19.31 35.742 19.35 35.778 ;
        RECT 19.914 35.742 19.966 35.778 ;
        RECT 20.074 35.742 20.126 35.778 ;
        RECT 20.63 35.742 20.682 35.778 ;
        RECT 21.014 35.742 21.068 35.778 ;
        RECT 21.65 35.742 21.704 35.778 ;
        RECT 21.896 35.742 21.95 35.778 ;
        RECT 22.854 35.742 22.906 35.778 ;
        RECT 23.174 35.742 23.226 35.778 ;
        RECT 23.654 35.742 23.706 35.778 ;
        RECT 23.974 35.742 24.026 35.778 ;
        RECT 24.454 35.742 24.506 35.778 ;
        RECT 24.774 35.742 24.826 35.778 ;
        RECT 25.254 35.742 25.306 35.778 ;
        RECT 25.574 35.742 25.626 35.778 ;
        RECT 26.054 35.742 26.106 35.778 ;
        RECT 26.374 35.742 26.426 35.778 ;
        RECT 26.854 35.742 26.906 35.778 ;
        RECT 27.174 35.742 27.226 35.778 ;
        RECT 27.654 35.742 27.706 35.778 ;
        RECT 27.974 35.742 28.026 35.778 ;
        RECT 28.454 35.742 28.506 35.778 ;
        RECT 28.774 35.742 28.826 35.778 ;
        RECT 29.254 35.742 29.306 35.778 ;
        RECT 29.574 35.742 29.626 35.778 ;
        RECT 30.054 35.742 30.106 35.778 ;
        RECT 30.374 35.742 30.426 35.778 ;
        RECT 30.854 35.742 30.906 35.778 ;
        RECT 31.174 35.742 31.226 35.778 ;
        RECT 31.654 35.742 31.706 35.778 ;
        RECT 31.974 35.742 32.026 35.778 ;
        RECT 32.454 35.742 32.506 35.778 ;
        RECT 32.774 35.742 32.826 35.778 ;
        RECT 33.254 35.742 33.306 35.778 ;
        RECT 33.574 35.742 33.626 35.778 ;
        RECT 34.054 35.742 34.106 35.778 ;
        RECT 34.374 35.742 34.426 35.778 ;
        RECT 34.854 35.742 34.906 35.778 ;
        RECT 35.174 35.742 35.226 35.778 ;
        RECT 0.654 35.862 0.706 35.898 ;
        RECT 0.974 35.862 1.026 35.898 ;
        RECT 1.454 35.862 1.506 35.898 ;
        RECT 1.774 35.862 1.826 35.898 ;
        RECT 2.254 35.862 2.306 35.898 ;
        RECT 2.574 35.862 2.626 35.898 ;
        RECT 3.054 35.862 3.106 35.898 ;
        RECT 3.374 35.862 3.426 35.898 ;
        RECT 3.854 35.862 3.906 35.898 ;
        RECT 4.174 35.862 4.226 35.898 ;
        RECT 4.654 35.862 4.706 35.898 ;
        RECT 4.974 35.862 5.026 35.898 ;
        RECT 5.454 35.862 5.506 35.898 ;
        RECT 5.774 35.862 5.826 35.898 ;
        RECT 6.254 35.862 6.306 35.898 ;
        RECT 6.574 35.862 6.626 35.898 ;
        RECT 7.054 35.862 7.106 35.898 ;
        RECT 7.374 35.862 7.426 35.898 ;
        RECT 7.854 35.862 7.906 35.898 ;
        RECT 8.174 35.862 8.226 35.898 ;
        RECT 8.654 35.862 8.706 35.898 ;
        RECT 8.974 35.862 9.026 35.898 ;
        RECT 9.454 35.862 9.506 35.898 ;
        RECT 9.774 35.862 9.826 35.898 ;
        RECT 10.254 35.862 10.306 35.898 ;
        RECT 10.574 35.862 10.626 35.898 ;
        RECT 11.054 35.862 11.106 35.898 ;
        RECT 11.374 35.862 11.426 35.898 ;
        RECT 11.854 35.862 11.906 35.898 ;
        RECT 12.174 35.862 12.226 35.898 ;
        RECT 12.654 35.862 12.706 35.898 ;
        RECT 12.974 35.862 13.026 35.898 ;
        RECT 22.854 35.862 22.906 35.898 ;
        RECT 23.174 35.862 23.226 35.898 ;
        RECT 23.654 35.862 23.706 35.898 ;
        RECT 23.974 35.862 24.026 35.898 ;
        RECT 24.454 35.862 24.506 35.898 ;
        RECT 24.774 35.862 24.826 35.898 ;
        RECT 25.254 35.862 25.306 35.898 ;
        RECT 25.574 35.862 25.626 35.898 ;
        RECT 26.054 35.862 26.106 35.898 ;
        RECT 26.374 35.862 26.426 35.898 ;
        RECT 26.854 35.862 26.906 35.898 ;
        RECT 27.174 35.862 27.226 35.898 ;
        RECT 27.654 35.862 27.706 35.898 ;
        RECT 27.974 35.862 28.026 35.898 ;
        RECT 28.454 35.862 28.506 35.898 ;
        RECT 28.774 35.862 28.826 35.898 ;
        RECT 29.254 35.862 29.306 35.898 ;
        RECT 29.574 35.862 29.626 35.898 ;
        RECT 30.054 35.862 30.106 35.898 ;
        RECT 30.374 35.862 30.426 35.898 ;
        RECT 30.854 35.862 30.906 35.898 ;
        RECT 31.174 35.862 31.226 35.898 ;
        RECT 31.654 35.862 31.706 35.898 ;
        RECT 31.974 35.862 32.026 35.898 ;
        RECT 32.454 35.862 32.506 35.898 ;
        RECT 32.774 35.862 32.826 35.898 ;
        RECT 33.254 35.862 33.306 35.898 ;
        RECT 33.574 35.862 33.626 35.898 ;
        RECT 34.054 35.862 34.106 35.898 ;
        RECT 34.374 35.862 34.426 35.898 ;
        RECT 34.854 35.862 34.906 35.898 ;
        RECT 35.174 35.862 35.226 35.898 ;
        RECT 0.654 36.102 0.706 36.138 ;
        RECT 0.974 36.102 1.026 36.138 ;
        RECT 1.454 36.102 1.506 36.138 ;
        RECT 1.774 36.102 1.826 36.138 ;
        RECT 2.254 36.102 2.306 36.138 ;
        RECT 2.574 36.102 2.626 36.138 ;
        RECT 3.054 36.102 3.106 36.138 ;
        RECT 3.374 36.102 3.426 36.138 ;
        RECT 3.854 36.102 3.906 36.138 ;
        RECT 4.174 36.102 4.226 36.138 ;
        RECT 4.654 36.102 4.706 36.138 ;
        RECT 4.974 36.102 5.026 36.138 ;
        RECT 5.454 36.102 5.506 36.138 ;
        RECT 5.774 36.102 5.826 36.138 ;
        RECT 6.254 36.102 6.306 36.138 ;
        RECT 6.574 36.102 6.626 36.138 ;
        RECT 7.054 36.102 7.106 36.138 ;
        RECT 7.374 36.102 7.426 36.138 ;
        RECT 7.854 36.102 7.906 36.138 ;
        RECT 8.174 36.102 8.226 36.138 ;
        RECT 8.654 36.102 8.706 36.138 ;
        RECT 8.974 36.102 9.026 36.138 ;
        RECT 9.454 36.102 9.506 36.138 ;
        RECT 9.774 36.102 9.826 36.138 ;
        RECT 10.254 36.102 10.306 36.138 ;
        RECT 10.574 36.102 10.626 36.138 ;
        RECT 11.054 36.102 11.106 36.138 ;
        RECT 11.374 36.102 11.426 36.138 ;
        RECT 11.854 36.102 11.906 36.138 ;
        RECT 12.174 36.102 12.226 36.138 ;
        RECT 12.654 36.102 12.706 36.138 ;
        RECT 12.974 36.102 13.026 36.138 ;
        RECT 14.05 36.102 14.104 36.138 ;
        RECT 14.296 36.102 14.35 36.138 ;
        RECT 14.932 36.102 14.986 36.138 ;
        RECT 21.014 36.102 21.068 36.138 ;
        RECT 21.65 36.102 21.704 36.138 ;
        RECT 21.896 36.102 21.95 36.138 ;
        RECT 22.854 36.102 22.906 36.138 ;
        RECT 23.174 36.102 23.226 36.138 ;
        RECT 23.654 36.102 23.706 36.138 ;
        RECT 23.974 36.102 24.026 36.138 ;
        RECT 24.454 36.102 24.506 36.138 ;
        RECT 24.774 36.102 24.826 36.138 ;
        RECT 25.254 36.102 25.306 36.138 ;
        RECT 25.574 36.102 25.626 36.138 ;
        RECT 26.054 36.102 26.106 36.138 ;
        RECT 26.374 36.102 26.426 36.138 ;
        RECT 26.854 36.102 26.906 36.138 ;
        RECT 27.174 36.102 27.226 36.138 ;
        RECT 27.654 36.102 27.706 36.138 ;
        RECT 27.974 36.102 28.026 36.138 ;
        RECT 28.454 36.102 28.506 36.138 ;
        RECT 28.774 36.102 28.826 36.138 ;
        RECT 29.254 36.102 29.306 36.138 ;
        RECT 29.574 36.102 29.626 36.138 ;
        RECT 30.054 36.102 30.106 36.138 ;
        RECT 30.374 36.102 30.426 36.138 ;
        RECT 30.854 36.102 30.906 36.138 ;
        RECT 31.174 36.102 31.226 36.138 ;
        RECT 31.654 36.102 31.706 36.138 ;
        RECT 31.974 36.102 32.026 36.138 ;
        RECT 32.454 36.102 32.506 36.138 ;
        RECT 32.774 36.102 32.826 36.138 ;
        RECT 33.254 36.102 33.306 36.138 ;
        RECT 33.574 36.102 33.626 36.138 ;
        RECT 34.054 36.102 34.106 36.138 ;
        RECT 34.374 36.102 34.426 36.138 ;
        RECT 34.854 36.102 34.906 36.138 ;
        RECT 35.174 36.102 35.226 36.138 ;
        RECT 15.874 36.2275 15.926 36.2525 ;
        RECT 16.964 36.2275 17.036 36.2525 ;
        RECT 17.844 36.2275 17.916 36.2525 ;
        RECT 18.664 36.2275 18.736 36.2525 ;
        RECT 18.964 36.2275 19.036 36.2525 ;
        RECT 20.074 36.2275 20.126 36.2525 ;
        RECT 0.654 36.222 0.706 36.258 ;
        RECT 1.454 36.222 1.506 36.258 ;
        RECT 2.254 36.222 2.306 36.258 ;
        RECT 3.054 36.222 3.106 36.258 ;
        RECT 3.854 36.222 3.906 36.258 ;
        RECT 4.654 36.222 4.706 36.258 ;
        RECT 5.454 36.222 5.506 36.258 ;
        RECT 6.254 36.222 6.306 36.258 ;
        RECT 7.054 36.222 7.106 36.258 ;
        RECT 7.854 36.222 7.906 36.258 ;
        RECT 8.654 36.222 8.706 36.258 ;
        RECT 9.454 36.222 9.506 36.258 ;
        RECT 10.254 36.222 10.306 36.258 ;
        RECT 11.054 36.222 11.106 36.258 ;
        RECT 11.854 36.222 11.906 36.258 ;
        RECT 12.654 36.222 12.706 36.258 ;
        RECT 14.05 36.222 14.104 36.258 ;
        RECT 14.296 36.222 14.35 36.258 ;
        RECT 14.932 36.222 14.986 36.258 ;
        RECT 15.318 36.222 15.37 36.258 ;
        RECT 16.034 36.222 16.086 36.258 ;
        RECT 16.8 36.222 16.854 36.258 ;
        RECT 17.412 36.222 17.452 36.258 ;
        RECT 18.148 36.222 18.188 36.258 ;
        RECT 18.356 36.222 18.396 36.258 ;
        RECT 19.31 36.222 19.35 36.258 ;
        RECT 19.914 36.222 19.966 36.258 ;
        RECT 20.63 36.222 20.682 36.258 ;
        RECT 21.014 36.222 21.068 36.258 ;
        RECT 21.65 36.222 21.704 36.258 ;
        RECT 21.896 36.222 21.95 36.258 ;
        RECT 22.854 36.222 22.906 36.258 ;
        RECT 23.654 36.222 23.706 36.258 ;
        RECT 24.454 36.222 24.506 36.258 ;
        RECT 25.254 36.222 25.306 36.258 ;
        RECT 26.054 36.222 26.106 36.258 ;
        RECT 26.854 36.222 26.906 36.258 ;
        RECT 27.654 36.222 27.706 36.258 ;
        RECT 28.454 36.222 28.506 36.258 ;
        RECT 29.254 36.222 29.306 36.258 ;
        RECT 30.054 36.222 30.106 36.258 ;
        RECT 30.854 36.222 30.906 36.258 ;
        RECT 31.654 36.222 31.706 36.258 ;
        RECT 32.454 36.222 32.506 36.258 ;
        RECT 33.254 36.222 33.306 36.258 ;
        RECT 34.054 36.222 34.106 36.258 ;
        RECT 34.854 36.222 34.906 36.258 ;
        RECT 14.296 36.7075 14.35 36.7325 ;
        RECT 16.964 36.7075 17.036 36.7325 ;
        RECT 17.844 36.7075 17.916 36.7325 ;
        RECT 18.664 36.7075 18.736 36.7325 ;
        RECT 18.964 36.7075 19.036 36.7325 ;
        RECT 21.65 36.7075 21.704 36.7325 ;
        RECT 0.654 36.702 0.706 36.738 ;
        RECT 0.974 36.702 1.026 36.738 ;
        RECT 1.454 36.702 1.506 36.738 ;
        RECT 1.774 36.702 1.826 36.738 ;
        RECT 2.254 36.702 2.306 36.738 ;
        RECT 2.574 36.702 2.626 36.738 ;
        RECT 3.054 36.702 3.106 36.738 ;
        RECT 3.374 36.702 3.426 36.738 ;
        RECT 3.854 36.702 3.906 36.738 ;
        RECT 4.174 36.702 4.226 36.738 ;
        RECT 4.654 36.702 4.706 36.738 ;
        RECT 4.974 36.702 5.026 36.738 ;
        RECT 5.454 36.702 5.506 36.738 ;
        RECT 5.774 36.702 5.826 36.738 ;
        RECT 6.254 36.702 6.306 36.738 ;
        RECT 6.574 36.702 6.626 36.738 ;
        RECT 7.054 36.702 7.106 36.738 ;
        RECT 7.374 36.702 7.426 36.738 ;
        RECT 7.854 36.702 7.906 36.738 ;
        RECT 8.174 36.702 8.226 36.738 ;
        RECT 8.654 36.702 8.706 36.738 ;
        RECT 8.974 36.702 9.026 36.738 ;
        RECT 9.454 36.702 9.506 36.738 ;
        RECT 9.774 36.702 9.826 36.738 ;
        RECT 10.254 36.702 10.306 36.738 ;
        RECT 10.574 36.702 10.626 36.738 ;
        RECT 11.054 36.702 11.106 36.738 ;
        RECT 11.374 36.702 11.426 36.738 ;
        RECT 11.854 36.702 11.906 36.738 ;
        RECT 12.174 36.702 12.226 36.738 ;
        RECT 12.654 36.702 12.706 36.738 ;
        RECT 12.974 36.702 13.026 36.738 ;
        RECT 14.05 36.702 14.104 36.738 ;
        RECT 14.932 36.702 14.986 36.738 ;
        RECT 15.318 36.702 15.37 36.738 ;
        RECT 15.874 36.702 15.926 36.738 ;
        RECT 16.034 36.702 16.086 36.738 ;
        RECT 16.8 36.702 16.854 36.738 ;
        RECT 17.412 36.702 17.452 36.738 ;
        RECT 18.148 36.702 18.188 36.738 ;
        RECT 18.356 36.702 18.396 36.738 ;
        RECT 19.31 36.702 19.35 36.738 ;
        RECT 19.914 36.702 19.966 36.738 ;
        RECT 20.074 36.702 20.126 36.738 ;
        RECT 20.63 36.702 20.682 36.738 ;
        RECT 21.014 36.702 21.068 36.738 ;
        RECT 21.896 36.702 21.95 36.738 ;
        RECT 22.854 36.702 22.906 36.738 ;
        RECT 23.174 36.702 23.226 36.738 ;
        RECT 23.654 36.702 23.706 36.738 ;
        RECT 23.974 36.702 24.026 36.738 ;
        RECT 24.454 36.702 24.506 36.738 ;
        RECT 24.774 36.702 24.826 36.738 ;
        RECT 25.254 36.702 25.306 36.738 ;
        RECT 25.574 36.702 25.626 36.738 ;
        RECT 26.054 36.702 26.106 36.738 ;
        RECT 26.374 36.702 26.426 36.738 ;
        RECT 26.854 36.702 26.906 36.738 ;
        RECT 27.174 36.702 27.226 36.738 ;
        RECT 27.654 36.702 27.706 36.738 ;
        RECT 27.974 36.702 28.026 36.738 ;
        RECT 28.454 36.702 28.506 36.738 ;
        RECT 28.774 36.702 28.826 36.738 ;
        RECT 29.254 36.702 29.306 36.738 ;
        RECT 29.574 36.702 29.626 36.738 ;
        RECT 30.054 36.702 30.106 36.738 ;
        RECT 30.374 36.702 30.426 36.738 ;
        RECT 30.854 36.702 30.906 36.738 ;
        RECT 31.174 36.702 31.226 36.738 ;
        RECT 31.654 36.702 31.706 36.738 ;
        RECT 31.974 36.702 32.026 36.738 ;
        RECT 32.454 36.702 32.506 36.738 ;
        RECT 32.774 36.702 32.826 36.738 ;
        RECT 33.254 36.702 33.306 36.738 ;
        RECT 33.574 36.702 33.626 36.738 ;
        RECT 34.054 36.702 34.106 36.738 ;
        RECT 34.374 36.702 34.426 36.738 ;
        RECT 34.854 36.702 34.906 36.738 ;
        RECT 35.174 36.702 35.226 36.738 ;
        RECT 14.05 37.1875 14.104 37.2125 ;
        RECT 14.296 37.1875 14.35 37.2125 ;
        RECT 16.964 37.1875 17.036 37.2125 ;
        RECT 18.664 37.1875 18.736 37.2125 ;
        RECT 18.964 37.1875 19.036 37.2125 ;
        RECT 21.65 37.1875 21.704 37.2125 ;
        RECT 21.896 37.1875 21.95 37.2125 ;
        RECT 0.654 37.182 0.706 37.218 ;
        RECT 0.974 37.182 1.026 37.218 ;
        RECT 1.454 37.182 1.506 37.218 ;
        RECT 1.774 37.182 1.826 37.218 ;
        RECT 2.254 37.182 2.306 37.218 ;
        RECT 2.574 37.182 2.626 37.218 ;
        RECT 3.054 37.182 3.106 37.218 ;
        RECT 3.374 37.182 3.426 37.218 ;
        RECT 3.854 37.182 3.906 37.218 ;
        RECT 4.174 37.182 4.226 37.218 ;
        RECT 4.654 37.182 4.706 37.218 ;
        RECT 4.974 37.182 5.026 37.218 ;
        RECT 5.454 37.182 5.506 37.218 ;
        RECT 5.774 37.182 5.826 37.218 ;
        RECT 6.254 37.182 6.306 37.218 ;
        RECT 6.574 37.182 6.626 37.218 ;
        RECT 7.054 37.182 7.106 37.218 ;
        RECT 7.374 37.182 7.426 37.218 ;
        RECT 7.854 37.182 7.906 37.218 ;
        RECT 8.174 37.182 8.226 37.218 ;
        RECT 8.654 37.182 8.706 37.218 ;
        RECT 8.974 37.182 9.026 37.218 ;
        RECT 9.454 37.182 9.506 37.218 ;
        RECT 9.774 37.182 9.826 37.218 ;
        RECT 10.254 37.182 10.306 37.218 ;
        RECT 10.574 37.182 10.626 37.218 ;
        RECT 11.054 37.182 11.106 37.218 ;
        RECT 11.374 37.182 11.426 37.218 ;
        RECT 11.854 37.182 11.906 37.218 ;
        RECT 12.174 37.182 12.226 37.218 ;
        RECT 12.654 37.182 12.706 37.218 ;
        RECT 12.974 37.182 13.026 37.218 ;
        RECT 14.932 37.182 14.986 37.218 ;
        RECT 15.318 37.182 15.37 37.218 ;
        RECT 15.874 37.182 15.926 37.218 ;
        RECT 16.034 37.182 16.086 37.218 ;
        RECT 16.8 37.182 16.854 37.218 ;
        RECT 17.412 37.182 17.452 37.218 ;
        RECT 18.148 37.182 18.188 37.218 ;
        RECT 18.356 37.182 18.396 37.218 ;
        RECT 19.31 37.182 19.35 37.218 ;
        RECT 19.914 37.182 19.966 37.218 ;
        RECT 20.074 37.182 20.126 37.218 ;
        RECT 20.63 37.182 20.682 37.218 ;
        RECT 21.014 37.182 21.068 37.218 ;
        RECT 22.854 37.182 22.906 37.218 ;
        RECT 23.174 37.182 23.226 37.218 ;
        RECT 23.654 37.182 23.706 37.218 ;
        RECT 23.974 37.182 24.026 37.218 ;
        RECT 24.454 37.182 24.506 37.218 ;
        RECT 24.774 37.182 24.826 37.218 ;
        RECT 25.254 37.182 25.306 37.218 ;
        RECT 25.574 37.182 25.626 37.218 ;
        RECT 26.054 37.182 26.106 37.218 ;
        RECT 26.374 37.182 26.426 37.218 ;
        RECT 26.854 37.182 26.906 37.218 ;
        RECT 27.174 37.182 27.226 37.218 ;
        RECT 27.654 37.182 27.706 37.218 ;
        RECT 27.974 37.182 28.026 37.218 ;
        RECT 28.454 37.182 28.506 37.218 ;
        RECT 28.774 37.182 28.826 37.218 ;
        RECT 29.254 37.182 29.306 37.218 ;
        RECT 29.574 37.182 29.626 37.218 ;
        RECT 30.054 37.182 30.106 37.218 ;
        RECT 30.374 37.182 30.426 37.218 ;
        RECT 30.854 37.182 30.906 37.218 ;
        RECT 31.174 37.182 31.226 37.218 ;
        RECT 31.654 37.182 31.706 37.218 ;
        RECT 31.974 37.182 32.026 37.218 ;
        RECT 32.454 37.182 32.506 37.218 ;
        RECT 32.774 37.182 32.826 37.218 ;
        RECT 33.254 37.182 33.306 37.218 ;
        RECT 33.574 37.182 33.626 37.218 ;
        RECT 34.054 37.182 34.106 37.218 ;
        RECT 34.374 37.182 34.426 37.218 ;
        RECT 34.854 37.182 34.906 37.218 ;
        RECT 35.174 37.182 35.226 37.218 ;
        RECT 0.654 37.302 0.706 37.338 ;
        RECT 0.974 37.302 1.026 37.338 ;
        RECT 1.454 37.302 1.506 37.338 ;
        RECT 1.774 37.302 1.826 37.338 ;
        RECT 2.254 37.302 2.306 37.338 ;
        RECT 2.574 37.302 2.626 37.338 ;
        RECT 3.054 37.302 3.106 37.338 ;
        RECT 3.374 37.302 3.426 37.338 ;
        RECT 3.854 37.302 3.906 37.338 ;
        RECT 4.174 37.302 4.226 37.338 ;
        RECT 4.654 37.302 4.706 37.338 ;
        RECT 4.974 37.302 5.026 37.338 ;
        RECT 5.454 37.302 5.506 37.338 ;
        RECT 5.774 37.302 5.826 37.338 ;
        RECT 6.254 37.302 6.306 37.338 ;
        RECT 6.574 37.302 6.626 37.338 ;
        RECT 7.054 37.302 7.106 37.338 ;
        RECT 7.374 37.302 7.426 37.338 ;
        RECT 7.854 37.302 7.906 37.338 ;
        RECT 8.174 37.302 8.226 37.338 ;
        RECT 8.654 37.302 8.706 37.338 ;
        RECT 8.974 37.302 9.026 37.338 ;
        RECT 9.454 37.302 9.506 37.338 ;
        RECT 9.774 37.302 9.826 37.338 ;
        RECT 10.254 37.302 10.306 37.338 ;
        RECT 10.574 37.302 10.626 37.338 ;
        RECT 11.054 37.302 11.106 37.338 ;
        RECT 11.374 37.302 11.426 37.338 ;
        RECT 11.854 37.302 11.906 37.338 ;
        RECT 12.174 37.302 12.226 37.338 ;
        RECT 12.654 37.302 12.706 37.338 ;
        RECT 12.974 37.302 13.026 37.338 ;
        RECT 22.854 37.302 22.906 37.338 ;
        RECT 23.174 37.302 23.226 37.338 ;
        RECT 23.654 37.302 23.706 37.338 ;
        RECT 23.974 37.302 24.026 37.338 ;
        RECT 24.454 37.302 24.506 37.338 ;
        RECT 24.774 37.302 24.826 37.338 ;
        RECT 25.254 37.302 25.306 37.338 ;
        RECT 25.574 37.302 25.626 37.338 ;
        RECT 26.054 37.302 26.106 37.338 ;
        RECT 26.374 37.302 26.426 37.338 ;
        RECT 26.854 37.302 26.906 37.338 ;
        RECT 27.174 37.302 27.226 37.338 ;
        RECT 27.654 37.302 27.706 37.338 ;
        RECT 27.974 37.302 28.026 37.338 ;
        RECT 28.454 37.302 28.506 37.338 ;
        RECT 28.774 37.302 28.826 37.338 ;
        RECT 29.254 37.302 29.306 37.338 ;
        RECT 29.574 37.302 29.626 37.338 ;
        RECT 30.054 37.302 30.106 37.338 ;
        RECT 30.374 37.302 30.426 37.338 ;
        RECT 30.854 37.302 30.906 37.338 ;
        RECT 31.174 37.302 31.226 37.338 ;
        RECT 31.654 37.302 31.706 37.338 ;
        RECT 31.974 37.302 32.026 37.338 ;
        RECT 32.454 37.302 32.506 37.338 ;
        RECT 32.774 37.302 32.826 37.338 ;
        RECT 33.254 37.302 33.306 37.338 ;
        RECT 33.574 37.302 33.626 37.338 ;
        RECT 34.054 37.302 34.106 37.338 ;
        RECT 34.374 37.302 34.426 37.338 ;
        RECT 34.854 37.302 34.906 37.338 ;
        RECT 35.174 37.302 35.226 37.338 ;
        RECT 15.318 37.6675 15.37 37.6925 ;
        RECT 16.964 37.6675 17.036 37.6925 ;
        RECT 17.844 37.6675 17.916 37.6925 ;
        RECT 18.664 37.6675 18.736 37.6925 ;
        RECT 18.964 37.6675 19.036 37.6925 ;
        RECT 20.63 37.6675 20.682 37.6925 ;
        RECT 14.05 37.662 14.104 37.698 ;
        RECT 14.296 37.662 14.35 37.698 ;
        RECT 14.932 37.662 14.986 37.698 ;
        RECT 15.874 37.662 15.926 37.698 ;
        RECT 16.034 37.662 16.086 37.698 ;
        RECT 16.8 37.662 16.854 37.698 ;
        RECT 17.412 37.662 17.452 37.698 ;
        RECT 18.148 37.662 18.188 37.698 ;
        RECT 19.31 37.662 19.35 37.698 ;
        RECT 19.914 37.662 19.966 37.698 ;
        RECT 20.074 37.662 20.126 37.698 ;
        RECT 21.014 37.662 21.068 37.698 ;
        RECT 21.65 37.662 21.704 37.698 ;
        RECT 21.896 37.662 21.95 37.698 ;
        RECT 0.654 37.782 0.706 37.818 ;
        RECT 0.974 37.782 1.026 37.818 ;
        RECT 1.454 37.782 1.506 37.818 ;
        RECT 1.774 37.782 1.826 37.818 ;
        RECT 2.254 37.782 2.306 37.818 ;
        RECT 2.574 37.782 2.626 37.818 ;
        RECT 3.054 37.782 3.106 37.818 ;
        RECT 3.374 37.782 3.426 37.818 ;
        RECT 3.854 37.782 3.906 37.818 ;
        RECT 4.174 37.782 4.226 37.818 ;
        RECT 4.654 37.782 4.706 37.818 ;
        RECT 4.974 37.782 5.026 37.818 ;
        RECT 5.454 37.782 5.506 37.818 ;
        RECT 5.774 37.782 5.826 37.818 ;
        RECT 6.254 37.782 6.306 37.818 ;
        RECT 6.574 37.782 6.626 37.818 ;
        RECT 7.054 37.782 7.106 37.818 ;
        RECT 7.374 37.782 7.426 37.818 ;
        RECT 7.854 37.782 7.906 37.818 ;
        RECT 8.174 37.782 8.226 37.818 ;
        RECT 8.654 37.782 8.706 37.818 ;
        RECT 8.974 37.782 9.026 37.818 ;
        RECT 9.454 37.782 9.506 37.818 ;
        RECT 9.774 37.782 9.826 37.818 ;
        RECT 10.254 37.782 10.306 37.818 ;
        RECT 10.574 37.782 10.626 37.818 ;
        RECT 11.054 37.782 11.106 37.818 ;
        RECT 11.374 37.782 11.426 37.818 ;
        RECT 11.854 37.782 11.906 37.818 ;
        RECT 12.174 37.782 12.226 37.818 ;
        RECT 12.654 37.782 12.706 37.818 ;
        RECT 12.974 37.782 13.026 37.818 ;
        RECT 22.854 37.782 22.906 37.818 ;
        RECT 23.174 37.782 23.226 37.818 ;
        RECT 23.654 37.782 23.706 37.818 ;
        RECT 23.974 37.782 24.026 37.818 ;
        RECT 24.454 37.782 24.506 37.818 ;
        RECT 24.774 37.782 24.826 37.818 ;
        RECT 25.254 37.782 25.306 37.818 ;
        RECT 25.574 37.782 25.626 37.818 ;
        RECT 26.054 37.782 26.106 37.818 ;
        RECT 26.374 37.782 26.426 37.818 ;
        RECT 26.854 37.782 26.906 37.818 ;
        RECT 27.174 37.782 27.226 37.818 ;
        RECT 27.654 37.782 27.706 37.818 ;
        RECT 27.974 37.782 28.026 37.818 ;
        RECT 28.454 37.782 28.506 37.818 ;
        RECT 28.774 37.782 28.826 37.818 ;
        RECT 29.254 37.782 29.306 37.818 ;
        RECT 29.574 37.782 29.626 37.818 ;
        RECT 30.054 37.782 30.106 37.818 ;
        RECT 30.374 37.782 30.426 37.818 ;
        RECT 30.854 37.782 30.906 37.818 ;
        RECT 31.174 37.782 31.226 37.818 ;
        RECT 31.654 37.782 31.706 37.818 ;
        RECT 31.974 37.782 32.026 37.818 ;
        RECT 32.454 37.782 32.506 37.818 ;
        RECT 32.774 37.782 32.826 37.818 ;
        RECT 33.254 37.782 33.306 37.818 ;
        RECT 33.574 37.782 33.626 37.818 ;
        RECT 34.054 37.782 34.106 37.818 ;
        RECT 34.374 37.782 34.426 37.818 ;
        RECT 34.854 37.782 34.906 37.818 ;
        RECT 35.174 37.782 35.226 37.818 ;
        RECT 0.654 38.022 0.706 38.058 ;
        RECT 0.974 38.022 1.026 38.058 ;
        RECT 1.454 38.022 1.506 38.058 ;
        RECT 1.774 38.022 1.826 38.058 ;
        RECT 2.254 38.022 2.306 38.058 ;
        RECT 2.574 38.022 2.626 38.058 ;
        RECT 3.054 38.022 3.106 38.058 ;
        RECT 3.374 38.022 3.426 38.058 ;
        RECT 3.854 38.022 3.906 38.058 ;
        RECT 4.174 38.022 4.226 38.058 ;
        RECT 4.654 38.022 4.706 38.058 ;
        RECT 4.974 38.022 5.026 38.058 ;
        RECT 5.454 38.022 5.506 38.058 ;
        RECT 5.774 38.022 5.826 38.058 ;
        RECT 6.254 38.022 6.306 38.058 ;
        RECT 6.574 38.022 6.626 38.058 ;
        RECT 7.054 38.022 7.106 38.058 ;
        RECT 7.374 38.022 7.426 38.058 ;
        RECT 7.854 38.022 7.906 38.058 ;
        RECT 8.174 38.022 8.226 38.058 ;
        RECT 8.654 38.022 8.706 38.058 ;
        RECT 8.974 38.022 9.026 38.058 ;
        RECT 9.454 38.022 9.506 38.058 ;
        RECT 9.774 38.022 9.826 38.058 ;
        RECT 10.254 38.022 10.306 38.058 ;
        RECT 10.574 38.022 10.626 38.058 ;
        RECT 11.054 38.022 11.106 38.058 ;
        RECT 11.374 38.022 11.426 38.058 ;
        RECT 11.854 38.022 11.906 38.058 ;
        RECT 12.174 38.022 12.226 38.058 ;
        RECT 12.654 38.022 12.706 38.058 ;
        RECT 12.974 38.022 13.026 38.058 ;
        RECT 14.05 38.022 14.104 38.058 ;
        RECT 14.296 38.022 14.35 38.058 ;
        RECT 14.932 38.022 14.986 38.058 ;
        RECT 21.014 38.022 21.068 38.058 ;
        RECT 21.65 38.022 21.704 38.058 ;
        RECT 21.896 38.022 21.95 38.058 ;
        RECT 22.854 38.022 22.906 38.058 ;
        RECT 23.174 38.022 23.226 38.058 ;
        RECT 23.654 38.022 23.706 38.058 ;
        RECT 23.974 38.022 24.026 38.058 ;
        RECT 24.454 38.022 24.506 38.058 ;
        RECT 24.774 38.022 24.826 38.058 ;
        RECT 25.254 38.022 25.306 38.058 ;
        RECT 25.574 38.022 25.626 38.058 ;
        RECT 26.054 38.022 26.106 38.058 ;
        RECT 26.374 38.022 26.426 38.058 ;
        RECT 26.854 38.022 26.906 38.058 ;
        RECT 27.174 38.022 27.226 38.058 ;
        RECT 27.654 38.022 27.706 38.058 ;
        RECT 27.974 38.022 28.026 38.058 ;
        RECT 28.454 38.022 28.506 38.058 ;
        RECT 28.774 38.022 28.826 38.058 ;
        RECT 29.254 38.022 29.306 38.058 ;
        RECT 29.574 38.022 29.626 38.058 ;
        RECT 30.054 38.022 30.106 38.058 ;
        RECT 30.374 38.022 30.426 38.058 ;
        RECT 30.854 38.022 30.906 38.058 ;
        RECT 31.174 38.022 31.226 38.058 ;
        RECT 31.654 38.022 31.706 38.058 ;
        RECT 31.974 38.022 32.026 38.058 ;
        RECT 32.454 38.022 32.506 38.058 ;
        RECT 32.774 38.022 32.826 38.058 ;
        RECT 33.254 38.022 33.306 38.058 ;
        RECT 33.574 38.022 33.626 38.058 ;
        RECT 34.054 38.022 34.106 38.058 ;
        RECT 34.374 38.022 34.426 38.058 ;
        RECT 34.854 38.022 34.906 38.058 ;
        RECT 35.174 38.022 35.226 38.058 ;
        RECT 15.874 38.1475 15.926 38.1725 ;
        RECT 16.964 38.1475 17.036 38.1725 ;
        RECT 17.844 38.1475 17.916 38.1725 ;
        RECT 18.664 38.1475 18.736 38.1725 ;
        RECT 18.964 38.1475 19.036 38.1725 ;
        RECT 20.074 38.1475 20.126 38.1725 ;
        RECT 14.05 38.142 14.104 38.178 ;
        RECT 14.296 38.142 14.35 38.178 ;
        RECT 14.932 38.142 14.986 38.178 ;
        RECT 15.318 38.142 15.37 38.178 ;
        RECT 16.034 38.142 16.086 38.178 ;
        RECT 16.8 38.142 16.854 38.178 ;
        RECT 17.412 38.142 17.452 38.178 ;
        RECT 18.148 38.142 18.188 38.178 ;
        RECT 18.356 38.142 18.396 38.178 ;
        RECT 19.31 38.142 19.35 38.178 ;
        RECT 19.914 38.142 19.966 38.178 ;
        RECT 20.63 38.142 20.682 38.178 ;
        RECT 21.014 38.142 21.068 38.178 ;
        RECT 21.65 38.142 21.704 38.178 ;
        RECT 21.896 38.142 21.95 38.178 ;
        RECT 0.654 38.502 0.706 38.538 ;
        RECT 0.974 38.502 1.026 38.538 ;
        RECT 1.454 38.502 1.506 38.538 ;
        RECT 1.774 38.502 1.826 38.538 ;
        RECT 2.254 38.502 2.306 38.538 ;
        RECT 2.574 38.502 2.626 38.538 ;
        RECT 3.054 38.502 3.106 38.538 ;
        RECT 3.374 38.502 3.426 38.538 ;
        RECT 3.854 38.502 3.906 38.538 ;
        RECT 4.174 38.502 4.226 38.538 ;
        RECT 4.654 38.502 4.706 38.538 ;
        RECT 4.974 38.502 5.026 38.538 ;
        RECT 5.454 38.502 5.506 38.538 ;
        RECT 5.774 38.502 5.826 38.538 ;
        RECT 6.254 38.502 6.306 38.538 ;
        RECT 6.574 38.502 6.626 38.538 ;
        RECT 7.054 38.502 7.106 38.538 ;
        RECT 7.374 38.502 7.426 38.538 ;
        RECT 7.854 38.502 7.906 38.538 ;
        RECT 8.174 38.502 8.226 38.538 ;
        RECT 8.654 38.502 8.706 38.538 ;
        RECT 8.974 38.502 9.026 38.538 ;
        RECT 9.454 38.502 9.506 38.538 ;
        RECT 9.774 38.502 9.826 38.538 ;
        RECT 10.254 38.502 10.306 38.538 ;
        RECT 10.574 38.502 10.626 38.538 ;
        RECT 11.054 38.502 11.106 38.538 ;
        RECT 11.374 38.502 11.426 38.538 ;
        RECT 11.854 38.502 11.906 38.538 ;
        RECT 12.174 38.502 12.226 38.538 ;
        RECT 12.654 38.502 12.706 38.538 ;
        RECT 12.974 38.502 13.026 38.538 ;
        RECT 14.05 38.502 14.104 38.538 ;
        RECT 14.296 38.502 14.35 38.538 ;
        RECT 14.932 38.502 14.986 38.538 ;
        RECT 21.014 38.502 21.068 38.538 ;
        RECT 21.65 38.502 21.704 38.538 ;
        RECT 21.896 38.502 21.95 38.538 ;
        RECT 22.854 38.502 22.906 38.538 ;
        RECT 23.174 38.502 23.226 38.538 ;
        RECT 23.654 38.502 23.706 38.538 ;
        RECT 23.974 38.502 24.026 38.538 ;
        RECT 24.454 38.502 24.506 38.538 ;
        RECT 24.774 38.502 24.826 38.538 ;
        RECT 25.254 38.502 25.306 38.538 ;
        RECT 25.574 38.502 25.626 38.538 ;
        RECT 26.054 38.502 26.106 38.538 ;
        RECT 26.374 38.502 26.426 38.538 ;
        RECT 26.854 38.502 26.906 38.538 ;
        RECT 27.174 38.502 27.226 38.538 ;
        RECT 27.654 38.502 27.706 38.538 ;
        RECT 27.974 38.502 28.026 38.538 ;
        RECT 28.454 38.502 28.506 38.538 ;
        RECT 28.774 38.502 28.826 38.538 ;
        RECT 29.254 38.502 29.306 38.538 ;
        RECT 29.574 38.502 29.626 38.538 ;
        RECT 30.054 38.502 30.106 38.538 ;
        RECT 30.374 38.502 30.426 38.538 ;
        RECT 30.854 38.502 30.906 38.538 ;
        RECT 31.174 38.502 31.226 38.538 ;
        RECT 31.654 38.502 31.706 38.538 ;
        RECT 31.974 38.502 32.026 38.538 ;
        RECT 32.454 38.502 32.506 38.538 ;
        RECT 32.774 38.502 32.826 38.538 ;
        RECT 33.254 38.502 33.306 38.538 ;
        RECT 33.574 38.502 33.626 38.538 ;
        RECT 34.054 38.502 34.106 38.538 ;
        RECT 34.374 38.502 34.426 38.538 ;
        RECT 34.854 38.502 34.906 38.538 ;
        RECT 35.174 38.502 35.226 38.538 ;
        RECT 14.296 38.6275 14.35 38.6525 ;
        RECT 16.964 38.6275 17.036 38.6525 ;
        RECT 17.844 38.6275 17.916 38.6525 ;
        RECT 18.664 38.6275 18.736 38.6525 ;
        RECT 18.964 38.6275 19.036 38.6525 ;
        RECT 21.65 38.6275 21.704 38.6525 ;
        RECT 14.05 38.622 14.104 38.658 ;
        RECT 14.932 38.622 14.986 38.658 ;
        RECT 15.318 38.622 15.37 38.658 ;
        RECT 15.478 38.622 15.53 38.658 ;
        RECT 15.874 38.622 15.926 38.658 ;
        RECT 16.034 38.622 16.086 38.658 ;
        RECT 16.8 38.622 16.854 38.658 ;
        RECT 17.412 38.622 17.452 38.658 ;
        RECT 18.148 38.622 18.188 38.658 ;
        RECT 18.356 38.622 18.396 38.658 ;
        RECT 19.31 38.622 19.35 38.658 ;
        RECT 19.914 38.622 19.966 38.658 ;
        RECT 20.074 38.622 20.126 38.658 ;
        RECT 20.47 38.622 20.522 38.658 ;
        RECT 20.63 38.622 20.682 38.658 ;
        RECT 21.014 38.622 21.068 38.658 ;
        RECT 21.896 38.622 21.95 38.658 ;
        RECT 0.974 38.742 1.026 38.778 ;
        RECT 1.774 38.742 1.826 38.778 ;
        RECT 2.574 38.742 2.626 38.778 ;
        RECT 3.374 38.742 3.426 38.778 ;
        RECT 4.174 38.742 4.226 38.778 ;
        RECT 4.974 38.742 5.026 38.778 ;
        RECT 5.774 38.742 5.826 38.778 ;
        RECT 6.574 38.742 6.626 38.778 ;
        RECT 7.374 38.742 7.426 38.778 ;
        RECT 8.174 38.742 8.226 38.778 ;
        RECT 8.974 38.742 9.026 38.778 ;
        RECT 9.774 38.742 9.826 38.778 ;
        RECT 10.574 38.742 10.626 38.778 ;
        RECT 11.374 38.742 11.426 38.778 ;
        RECT 12.174 38.742 12.226 38.778 ;
        RECT 12.974 38.742 13.026 38.778 ;
        RECT 14.05 38.742 14.104 38.778 ;
        RECT 14.296 38.742 14.35 38.778 ;
        RECT 14.932 38.742 14.986 38.778 ;
        RECT 21.014 38.742 21.068 38.778 ;
        RECT 21.65 38.742 21.704 38.778 ;
        RECT 21.896 38.742 21.95 38.778 ;
        RECT 23.174 38.742 23.226 38.778 ;
        RECT 23.974 38.742 24.026 38.778 ;
        RECT 24.774 38.742 24.826 38.778 ;
        RECT 25.574 38.742 25.626 38.778 ;
        RECT 26.374 38.742 26.426 38.778 ;
        RECT 27.174 38.742 27.226 38.778 ;
        RECT 27.974 38.742 28.026 38.778 ;
        RECT 28.774 38.742 28.826 38.778 ;
        RECT 29.574 38.742 29.626 38.778 ;
        RECT 30.374 38.742 30.426 38.778 ;
        RECT 31.174 38.742 31.226 38.778 ;
        RECT 31.974 38.742 32.026 38.778 ;
        RECT 32.774 38.742 32.826 38.778 ;
        RECT 33.574 38.742 33.626 38.778 ;
        RECT 34.374 38.742 34.426 38.778 ;
        RECT 35.174 38.742 35.226 38.778 ;
        RECT 16.964 39.1075 17.036 39.1325 ;
        RECT 17.844 39.1075 17.916 39.1325 ;
        RECT 18.664 39.1075 18.736 39.1325 ;
        RECT 18.964 39.1075 19.036 39.1325 ;
        RECT 14.05 39.102 14.104 39.138 ;
        RECT 14.296 39.102 14.35 39.138 ;
        RECT 14.932 39.102 14.986 39.138 ;
        RECT 15.318 39.102 15.37 39.138 ;
        RECT 15.478 39.102 15.53 39.138 ;
        RECT 15.874 39.102 15.926 39.138 ;
        RECT 16.034 39.102 16.086 39.138 ;
        RECT 16.8 39.102 16.854 39.138 ;
        RECT 17.412 39.102 17.452 39.138 ;
        RECT 18.148 39.102 18.188 39.138 ;
        RECT 18.356 39.102 18.396 39.138 ;
        RECT 19.31 39.102 19.35 39.138 ;
        RECT 19.914 39.102 19.966 39.138 ;
        RECT 20.074 39.102 20.126 39.138 ;
        RECT 20.47 39.102 20.522 39.138 ;
        RECT 20.63 39.102 20.682 39.138 ;
        RECT 21.014 39.102 21.068 39.138 ;
        RECT 21.65 39.102 21.704 39.138 ;
        RECT 21.896 39.102 21.95 39.138 ;
        RECT 16.964 39.8545 17.036 39.8795 ;
        RECT 17.844 39.8545 17.916 39.8795 ;
        RECT 18.664 39.8545 18.736 39.8795 ;
        RECT 18.964 39.8545 19.036 39.8795 ;
        RECT 14.05 39.849 14.104 39.885 ;
        RECT 14.932 39.849 14.986 39.885 ;
        RECT 15.318 39.849 15.37 39.885 ;
        RECT 15.478 39.849 15.53 39.885 ;
        RECT 15.874 39.849 15.926 39.885 ;
        RECT 16.034 39.849 16.086 39.885 ;
        RECT 16.8 39.849 16.854 39.885 ;
        RECT 18.148 39.849 18.188 39.885 ;
        RECT 18.356 39.849 18.396 39.885 ;
        RECT 19.914 39.849 19.966 39.885 ;
        RECT 20.074 39.849 20.126 39.885 ;
        RECT 20.47 39.849 20.522 39.885 ;
        RECT 20.63 39.849 20.682 39.885 ;
        RECT 21.014 39.849 21.068 39.885 ;
        RECT 21.896 39.849 21.95 39.885 ;
        RECT 16.964 40.0835 17.036 40.1085 ;
        RECT 18.664 40.0835 18.736 40.1085 ;
        RECT 18.964 40.0835 19.036 40.1085 ;
        RECT 14.05 40.078 14.104 40.114 ;
        RECT 14.296 40.078 14.35 40.114 ;
        RECT 14.932 40.078 14.986 40.114 ;
        RECT 15.318 40.078 15.37 40.114 ;
        RECT 15.478 40.078 15.53 40.114 ;
        RECT 15.874 40.078 15.926 40.114 ;
        RECT 16.034 40.078 16.086 40.114 ;
        RECT 16.8 40.078 16.854 40.114 ;
        RECT 18.148 40.078 18.188 40.114 ;
        RECT 19.914 40.078 19.966 40.114 ;
        RECT 20.074 40.078 20.126 40.114 ;
        RECT 20.47 40.078 20.522 40.114 ;
        RECT 20.63 40.078 20.682 40.114 ;
        RECT 21.014 40.078 21.068 40.114 ;
        RECT 21.65 40.078 21.704 40.114 ;
        RECT 21.896 40.078 21.95 40.114 ;
        RECT 17.844 40.1605 17.916 40.1855 ;
        RECT 18.356 40.155 18.396 40.191 ;
        RECT 16.964 40.5315 17.036 40.5565 ;
        RECT 17.844 40.5315 17.916 40.5565 ;
        RECT 18.964 40.5315 19.036 40.5565 ;
        RECT 14.05 40.526 14.104 40.562 ;
        RECT 14.296 40.526 14.35 40.562 ;
        RECT 14.932 40.526 14.986 40.562 ;
        RECT 15.318 40.526 15.37 40.562 ;
        RECT 15.874 40.526 15.926 40.562 ;
        RECT 16.034 40.526 16.086 40.562 ;
        RECT 18.356 40.526 18.396 40.562 ;
        RECT 19.914 40.526 19.966 40.562 ;
        RECT 20.074 40.526 20.126 40.562 ;
        RECT 20.63 40.526 20.682 40.562 ;
        RECT 21.014 40.526 21.068 40.562 ;
        RECT 21.65 40.526 21.704 40.562 ;
        RECT 21.896 40.526 21.95 40.562 ;
        RECT 17.844 40.6835 17.916 40.7085 ;
        RECT 18.356 40.678 18.396 40.714 ;
        RECT 18.664 40.7605 18.736 40.7855 ;
        RECT 18.964 40.7605 19.036 40.7855 ;
        RECT 14.296 40.755 14.35 40.791 ;
        RECT 14.932 40.755 14.986 40.791 ;
        RECT 15.318 40.755 15.37 40.791 ;
        RECT 15.478 40.755 15.53 40.791 ;
        RECT 15.874 40.755 15.926 40.791 ;
        RECT 18.148 40.755 18.188 40.791 ;
        RECT 20.074 40.755 20.126 40.791 ;
        RECT 20.47 40.755 20.522 40.791 ;
        RECT 20.63 40.755 20.682 40.791 ;
        RECT 21.014 40.755 21.068 40.791 ;
        RECT 21.65 40.755 21.704 40.791 ;
        RECT 16.964 41.0545 17.036 41.0795 ;
        RECT 17.844 41.0545 17.916 41.0795 ;
        RECT 18.664 41.0545 18.736 41.0795 ;
        RECT 18.964 41.0545 19.036 41.0795 ;
        RECT 14.05 41.049 14.104 41.085 ;
        RECT 14.932 41.049 14.986 41.085 ;
        RECT 15.318 41.049 15.37 41.085 ;
        RECT 15.478 41.049 15.53 41.085 ;
        RECT 15.874 41.049 15.926 41.085 ;
        RECT 16.034 41.049 16.086 41.085 ;
        RECT 16.8 41.049 16.854 41.085 ;
        RECT 18.148 41.049 18.188 41.085 ;
        RECT 18.356 41.049 18.396 41.085 ;
        RECT 19.914 41.049 19.966 41.085 ;
        RECT 20.074 41.049 20.126 41.085 ;
        RECT 20.47 41.049 20.522 41.085 ;
        RECT 20.63 41.049 20.682 41.085 ;
        RECT 21.014 41.049 21.068 41.085 ;
        RECT 21.896 41.049 21.95 41.085 ;
        RECT 16.964 41.2835 17.036 41.3085 ;
        RECT 18.664 41.2835 18.736 41.3085 ;
        RECT 18.964 41.2835 19.036 41.3085 ;
        RECT 14.05 41.278 14.104 41.314 ;
        RECT 14.296 41.278 14.35 41.314 ;
        RECT 14.932 41.278 14.986 41.314 ;
        RECT 15.318 41.278 15.37 41.314 ;
        RECT 15.478 41.278 15.53 41.314 ;
        RECT 15.874 41.278 15.926 41.314 ;
        RECT 16.034 41.278 16.086 41.314 ;
        RECT 16.8 41.278 16.854 41.314 ;
        RECT 18.148 41.278 18.188 41.314 ;
        RECT 19.914 41.278 19.966 41.314 ;
        RECT 20.074 41.278 20.126 41.314 ;
        RECT 20.47 41.278 20.522 41.314 ;
        RECT 20.63 41.278 20.682 41.314 ;
        RECT 21.014 41.278 21.068 41.314 ;
        RECT 21.65 41.278 21.704 41.314 ;
        RECT 21.896 41.278 21.95 41.314 ;
        RECT 17.844 41.3605 17.916 41.3855 ;
        RECT 18.356 41.355 18.396 41.391 ;
        RECT 16.964 41.7315 17.036 41.7565 ;
        RECT 17.844 41.7315 17.916 41.7565 ;
        RECT 18.964 41.7315 19.036 41.7565 ;
        RECT 14.05 41.726 14.104 41.762 ;
        RECT 14.296 41.726 14.35 41.762 ;
        RECT 14.932 41.726 14.986 41.762 ;
        RECT 15.318 41.726 15.37 41.762 ;
        RECT 15.874 41.726 15.926 41.762 ;
        RECT 16.034 41.726 16.086 41.762 ;
        RECT 18.356 41.726 18.396 41.762 ;
        RECT 19.914 41.726 19.966 41.762 ;
        RECT 20.074 41.726 20.126 41.762 ;
        RECT 20.63 41.726 20.682 41.762 ;
        RECT 21.014 41.726 21.068 41.762 ;
        RECT 21.65 41.726 21.704 41.762 ;
        RECT 21.896 41.726 21.95 41.762 ;
        RECT 17.844 41.8835 17.916 41.9085 ;
        RECT 18.356 41.878 18.396 41.914 ;
        RECT 18.664 41.9605 18.736 41.9855 ;
        RECT 18.964 41.9605 19.036 41.9855 ;
        RECT 14.296 41.955 14.35 41.991 ;
        RECT 14.932 41.955 14.986 41.991 ;
        RECT 15.318 41.955 15.37 41.991 ;
        RECT 15.478 41.955 15.53 41.991 ;
        RECT 15.874 41.955 15.926 41.991 ;
        RECT 18.148 41.955 18.188 41.991 ;
        RECT 20.074 41.955 20.126 41.991 ;
        RECT 20.47 41.955 20.522 41.991 ;
        RECT 20.63 41.955 20.682 41.991 ;
        RECT 21.014 41.955 21.068 41.991 ;
        RECT 21.65 41.955 21.704 41.991 ;
        RECT 16.964 42.2545 17.036 42.2795 ;
        RECT 17.844 42.2545 17.916 42.2795 ;
        RECT 18.664 42.2545 18.736 42.2795 ;
        RECT 18.964 42.2545 19.036 42.2795 ;
        RECT 14.05 42.249 14.104 42.285 ;
        RECT 14.932 42.249 14.986 42.285 ;
        RECT 15.318 42.249 15.37 42.285 ;
        RECT 15.478 42.249 15.53 42.285 ;
        RECT 15.874 42.249 15.926 42.285 ;
        RECT 16.034 42.249 16.086 42.285 ;
        RECT 16.8 42.249 16.854 42.285 ;
        RECT 18.148 42.249 18.188 42.285 ;
        RECT 18.356 42.249 18.396 42.285 ;
        RECT 19.914 42.249 19.966 42.285 ;
        RECT 20.074 42.249 20.126 42.285 ;
        RECT 20.47 42.249 20.522 42.285 ;
        RECT 20.63 42.249 20.682 42.285 ;
        RECT 21.014 42.249 21.068 42.285 ;
        RECT 21.896 42.249 21.95 42.285 ;
        RECT 16.964 42.4835 17.036 42.5085 ;
        RECT 18.664 42.4835 18.736 42.5085 ;
        RECT 18.964 42.4835 19.036 42.5085 ;
        RECT 14.05 42.478 14.104 42.514 ;
        RECT 14.296 42.478 14.35 42.514 ;
        RECT 14.932 42.478 14.986 42.514 ;
        RECT 15.318 42.478 15.37 42.514 ;
        RECT 15.478 42.478 15.53 42.514 ;
        RECT 15.874 42.478 15.926 42.514 ;
        RECT 16.034 42.478 16.086 42.514 ;
        RECT 16.8 42.478 16.854 42.514 ;
        RECT 18.148 42.478 18.188 42.514 ;
        RECT 19.914 42.478 19.966 42.514 ;
        RECT 20.074 42.478 20.126 42.514 ;
        RECT 20.47 42.478 20.522 42.514 ;
        RECT 20.63 42.478 20.682 42.514 ;
        RECT 21.014 42.478 21.068 42.514 ;
        RECT 21.65 42.478 21.704 42.514 ;
        RECT 21.896 42.478 21.95 42.514 ;
        RECT 17.844 42.5605 17.916 42.5855 ;
        RECT 18.356 42.555 18.396 42.591 ;
        RECT 16.964 42.9315 17.036 42.9565 ;
        RECT 17.844 42.9315 17.916 42.9565 ;
        RECT 18.964 42.9315 19.036 42.9565 ;
        RECT 14.05 42.926 14.104 42.962 ;
        RECT 14.296 42.926 14.35 42.962 ;
        RECT 14.932 42.926 14.986 42.962 ;
        RECT 15.318 42.926 15.37 42.962 ;
        RECT 15.874 42.926 15.926 42.962 ;
        RECT 16.034 42.926 16.086 42.962 ;
        RECT 18.356 42.926 18.396 42.962 ;
        RECT 19.914 42.926 19.966 42.962 ;
        RECT 20.074 42.926 20.126 42.962 ;
        RECT 20.63 42.926 20.682 42.962 ;
        RECT 21.014 42.926 21.068 42.962 ;
        RECT 21.65 42.926 21.704 42.962 ;
        RECT 21.896 42.926 21.95 42.962 ;
        RECT 17.844 43.0835 17.916 43.1085 ;
        RECT 18.356 43.078 18.396 43.114 ;
        RECT 18.664 43.1605 18.736 43.1855 ;
        RECT 18.964 43.1605 19.036 43.1855 ;
        RECT 14.296 43.155 14.35 43.191 ;
        RECT 14.932 43.155 14.986 43.191 ;
        RECT 15.318 43.155 15.37 43.191 ;
        RECT 15.478 43.155 15.53 43.191 ;
        RECT 15.874 43.155 15.926 43.191 ;
        RECT 18.148 43.155 18.188 43.191 ;
        RECT 20.074 43.155 20.126 43.191 ;
        RECT 20.47 43.155 20.522 43.191 ;
        RECT 20.63 43.155 20.682 43.191 ;
        RECT 21.014 43.155 21.068 43.191 ;
        RECT 21.65 43.155 21.704 43.191 ;
        RECT 16.964 43.4545 17.036 43.4795 ;
        RECT 17.844 43.4545 17.916 43.4795 ;
        RECT 18.664 43.4545 18.736 43.4795 ;
        RECT 18.964 43.4545 19.036 43.4795 ;
        RECT 14.05 43.449 14.104 43.485 ;
        RECT 14.932 43.449 14.986 43.485 ;
        RECT 15.318 43.449 15.37 43.485 ;
        RECT 15.478 43.449 15.53 43.485 ;
        RECT 15.874 43.449 15.926 43.485 ;
        RECT 16.034 43.449 16.086 43.485 ;
        RECT 16.8 43.449 16.854 43.485 ;
        RECT 18.148 43.449 18.188 43.485 ;
        RECT 18.356 43.449 18.396 43.485 ;
        RECT 19.914 43.449 19.966 43.485 ;
        RECT 20.074 43.449 20.126 43.485 ;
        RECT 20.47 43.449 20.522 43.485 ;
        RECT 20.63 43.449 20.682 43.485 ;
        RECT 21.014 43.449 21.068 43.485 ;
        RECT 21.896 43.449 21.95 43.485 ;
        RECT 16.964 43.6835 17.036 43.7085 ;
        RECT 18.664 43.6835 18.736 43.7085 ;
        RECT 18.964 43.6835 19.036 43.7085 ;
        RECT 14.05 43.678 14.104 43.714 ;
        RECT 14.296 43.678 14.35 43.714 ;
        RECT 14.932 43.678 14.986 43.714 ;
        RECT 15.318 43.678 15.37 43.714 ;
        RECT 15.478 43.678 15.53 43.714 ;
        RECT 15.874 43.678 15.926 43.714 ;
        RECT 16.034 43.678 16.086 43.714 ;
        RECT 16.8 43.678 16.854 43.714 ;
        RECT 18.148 43.678 18.188 43.714 ;
        RECT 19.914 43.678 19.966 43.714 ;
        RECT 20.074 43.678 20.126 43.714 ;
        RECT 20.47 43.678 20.522 43.714 ;
        RECT 20.63 43.678 20.682 43.714 ;
        RECT 21.014 43.678 21.068 43.714 ;
        RECT 21.65 43.678 21.704 43.714 ;
        RECT 21.896 43.678 21.95 43.714 ;
        RECT 17.844 43.7605 17.916 43.7855 ;
        RECT 18.356 43.755 18.396 43.791 ;
        RECT 16.964 44.1315 17.036 44.1565 ;
        RECT 17.844 44.1315 17.916 44.1565 ;
        RECT 18.964 44.1315 19.036 44.1565 ;
        RECT 14.05 44.126 14.104 44.162 ;
        RECT 14.296 44.126 14.35 44.162 ;
        RECT 14.932 44.126 14.986 44.162 ;
        RECT 15.318 44.126 15.37 44.162 ;
        RECT 15.874 44.126 15.926 44.162 ;
        RECT 16.034 44.126 16.086 44.162 ;
        RECT 18.356 44.126 18.396 44.162 ;
        RECT 19.914 44.126 19.966 44.162 ;
        RECT 20.074 44.126 20.126 44.162 ;
        RECT 20.63 44.126 20.682 44.162 ;
        RECT 21.014 44.126 21.068 44.162 ;
        RECT 21.65 44.126 21.704 44.162 ;
        RECT 21.896 44.126 21.95 44.162 ;
        RECT 17.844 44.2835 17.916 44.3085 ;
        RECT 18.356 44.278 18.396 44.314 ;
        RECT 18.664 44.3605 18.736 44.3855 ;
        RECT 18.964 44.3605 19.036 44.3855 ;
        RECT 14.296 44.355 14.35 44.391 ;
        RECT 14.932 44.355 14.986 44.391 ;
        RECT 15.318 44.355 15.37 44.391 ;
        RECT 15.478 44.355 15.53 44.391 ;
        RECT 15.874 44.355 15.926 44.391 ;
        RECT 18.148 44.355 18.188 44.391 ;
        RECT 20.074 44.355 20.126 44.391 ;
        RECT 20.47 44.355 20.522 44.391 ;
        RECT 20.63 44.355 20.682 44.391 ;
        RECT 21.014 44.355 21.068 44.391 ;
        RECT 21.65 44.355 21.704 44.391 ;
        RECT 16.964 44.6545 17.036 44.6795 ;
        RECT 17.844 44.6545 17.916 44.6795 ;
        RECT 18.664 44.6545 18.736 44.6795 ;
        RECT 18.964 44.6545 19.036 44.6795 ;
        RECT 14.05 44.649 14.104 44.685 ;
        RECT 14.932 44.649 14.986 44.685 ;
        RECT 15.318 44.649 15.37 44.685 ;
        RECT 15.478 44.649 15.53 44.685 ;
        RECT 15.874 44.649 15.926 44.685 ;
        RECT 16.034 44.649 16.086 44.685 ;
        RECT 16.8 44.649 16.854 44.685 ;
        RECT 18.148 44.649 18.188 44.685 ;
        RECT 18.356 44.649 18.396 44.685 ;
        RECT 19.914 44.649 19.966 44.685 ;
        RECT 20.074 44.649 20.126 44.685 ;
        RECT 20.47 44.649 20.522 44.685 ;
        RECT 20.63 44.649 20.682 44.685 ;
        RECT 21.014 44.649 21.068 44.685 ;
        RECT 21.896 44.649 21.95 44.685 ;
        RECT 16.964 44.8835 17.036 44.9085 ;
        RECT 18.664 44.8835 18.736 44.9085 ;
        RECT 18.964 44.8835 19.036 44.9085 ;
        RECT 14.05 44.878 14.104 44.914 ;
        RECT 14.296 44.878 14.35 44.914 ;
        RECT 14.932 44.878 14.986 44.914 ;
        RECT 15.318 44.878 15.37 44.914 ;
        RECT 15.478 44.878 15.53 44.914 ;
        RECT 15.874 44.878 15.926 44.914 ;
        RECT 16.034 44.878 16.086 44.914 ;
        RECT 16.8 44.878 16.854 44.914 ;
        RECT 18.148 44.878 18.188 44.914 ;
        RECT 19.914 44.878 19.966 44.914 ;
        RECT 20.074 44.878 20.126 44.914 ;
        RECT 20.47 44.878 20.522 44.914 ;
        RECT 20.63 44.878 20.682 44.914 ;
        RECT 21.014 44.878 21.068 44.914 ;
        RECT 21.65 44.878 21.704 44.914 ;
        RECT 21.896 44.878 21.95 44.914 ;
        RECT 17.844 44.9605 17.916 44.9855 ;
        RECT 18.356 44.955 18.396 44.991 ;
        RECT 16.964 45.3315 17.036 45.3565 ;
        RECT 17.844 45.3315 17.916 45.3565 ;
        RECT 18.964 45.3315 19.036 45.3565 ;
        RECT 14.05 45.326 14.104 45.362 ;
        RECT 14.296 45.326 14.35 45.362 ;
        RECT 14.932 45.326 14.986 45.362 ;
        RECT 15.318 45.326 15.37 45.362 ;
        RECT 15.874 45.326 15.926 45.362 ;
        RECT 16.034 45.326 16.086 45.362 ;
        RECT 18.356 45.326 18.396 45.362 ;
        RECT 19.914 45.326 19.966 45.362 ;
        RECT 20.074 45.326 20.126 45.362 ;
        RECT 20.63 45.326 20.682 45.362 ;
        RECT 21.014 45.326 21.068 45.362 ;
        RECT 21.65 45.326 21.704 45.362 ;
        RECT 21.896 45.326 21.95 45.362 ;
        RECT 17.844 45.4835 17.916 45.5085 ;
        RECT 18.356 45.478 18.396 45.514 ;
        RECT 18.664 45.5605 18.736 45.5855 ;
        RECT 18.964 45.5605 19.036 45.5855 ;
        RECT 14.296 45.555 14.35 45.591 ;
        RECT 14.932 45.555 14.986 45.591 ;
        RECT 15.318 45.555 15.37 45.591 ;
        RECT 15.478 45.555 15.53 45.591 ;
        RECT 15.874 45.555 15.926 45.591 ;
        RECT 18.148 45.555 18.188 45.591 ;
        RECT 20.074 45.555 20.126 45.591 ;
        RECT 20.47 45.555 20.522 45.591 ;
        RECT 20.63 45.555 20.682 45.591 ;
        RECT 21.014 45.555 21.068 45.591 ;
        RECT 21.65 45.555 21.704 45.591 ;
        RECT 16.964 45.8545 17.036 45.8795 ;
        RECT 17.844 45.8545 17.916 45.8795 ;
        RECT 18.664 45.8545 18.736 45.8795 ;
        RECT 18.964 45.8545 19.036 45.8795 ;
        RECT 14.05 45.849 14.104 45.885 ;
        RECT 14.932 45.849 14.986 45.885 ;
        RECT 15.318 45.849 15.37 45.885 ;
        RECT 15.478 45.849 15.53 45.885 ;
        RECT 15.874 45.849 15.926 45.885 ;
        RECT 16.034 45.849 16.086 45.885 ;
        RECT 16.8 45.849 16.854 45.885 ;
        RECT 18.148 45.849 18.188 45.885 ;
        RECT 18.356 45.849 18.396 45.885 ;
        RECT 19.914 45.849 19.966 45.885 ;
        RECT 20.074 45.849 20.126 45.885 ;
        RECT 20.47 45.849 20.522 45.885 ;
        RECT 20.63 45.849 20.682 45.885 ;
        RECT 21.014 45.849 21.068 45.885 ;
        RECT 21.896 45.849 21.95 45.885 ;
        RECT 16.964 46.0835 17.036 46.1085 ;
        RECT 18.664 46.0835 18.736 46.1085 ;
        RECT 18.964 46.0835 19.036 46.1085 ;
        RECT 14.05 46.078 14.104 46.114 ;
        RECT 14.296 46.078 14.35 46.114 ;
        RECT 14.932 46.078 14.986 46.114 ;
        RECT 15.318 46.078 15.37 46.114 ;
        RECT 15.478 46.078 15.53 46.114 ;
        RECT 15.874 46.078 15.926 46.114 ;
        RECT 16.034 46.078 16.086 46.114 ;
        RECT 16.8 46.078 16.854 46.114 ;
        RECT 18.148 46.078 18.188 46.114 ;
        RECT 19.914 46.078 19.966 46.114 ;
        RECT 20.074 46.078 20.126 46.114 ;
        RECT 20.47 46.078 20.522 46.114 ;
        RECT 20.63 46.078 20.682 46.114 ;
        RECT 21.014 46.078 21.068 46.114 ;
        RECT 21.65 46.078 21.704 46.114 ;
        RECT 21.896 46.078 21.95 46.114 ;
        RECT 17.844 46.1605 17.916 46.1855 ;
        RECT 18.356 46.155 18.396 46.191 ;
        RECT 16.964 46.5315 17.036 46.5565 ;
        RECT 17.844 46.5315 17.916 46.5565 ;
        RECT 18.964 46.5315 19.036 46.5565 ;
        RECT 14.05 46.526 14.104 46.562 ;
        RECT 14.296 46.526 14.35 46.562 ;
        RECT 14.932 46.526 14.986 46.562 ;
        RECT 15.318 46.526 15.37 46.562 ;
        RECT 15.874 46.526 15.926 46.562 ;
        RECT 16.034 46.526 16.086 46.562 ;
        RECT 18.356 46.526 18.396 46.562 ;
        RECT 19.914 46.526 19.966 46.562 ;
        RECT 20.074 46.526 20.126 46.562 ;
        RECT 20.63 46.526 20.682 46.562 ;
        RECT 21.014 46.526 21.068 46.562 ;
        RECT 21.65 46.526 21.704 46.562 ;
        RECT 21.896 46.526 21.95 46.562 ;
        RECT 17.844 46.6835 17.916 46.7085 ;
        RECT 18.356 46.678 18.396 46.714 ;
        RECT 18.664 46.7605 18.736 46.7855 ;
        RECT 18.964 46.7605 19.036 46.7855 ;
        RECT 14.296 46.755 14.35 46.791 ;
        RECT 14.932 46.755 14.986 46.791 ;
        RECT 15.318 46.755 15.37 46.791 ;
        RECT 15.478 46.755 15.53 46.791 ;
        RECT 15.874 46.755 15.926 46.791 ;
        RECT 18.148 46.755 18.188 46.791 ;
        RECT 20.074 46.755 20.126 46.791 ;
        RECT 20.47 46.755 20.522 46.791 ;
        RECT 20.63 46.755 20.682 46.791 ;
        RECT 21.014 46.755 21.068 46.791 ;
        RECT 21.65 46.755 21.704 46.791 ;
        RECT 16.964 47.0545 17.036 47.0795 ;
        RECT 17.844 47.0545 17.916 47.0795 ;
        RECT 18.664 47.0545 18.736 47.0795 ;
        RECT 18.964 47.0545 19.036 47.0795 ;
        RECT 14.05 47.049 14.104 47.085 ;
        RECT 14.932 47.049 14.986 47.085 ;
        RECT 15.318 47.049 15.37 47.085 ;
        RECT 15.478 47.049 15.53 47.085 ;
        RECT 15.874 47.049 15.926 47.085 ;
        RECT 16.034 47.049 16.086 47.085 ;
        RECT 16.8 47.049 16.854 47.085 ;
        RECT 18.148 47.049 18.188 47.085 ;
        RECT 18.356 47.049 18.396 47.085 ;
        RECT 19.914 47.049 19.966 47.085 ;
        RECT 20.074 47.049 20.126 47.085 ;
        RECT 20.47 47.049 20.522 47.085 ;
        RECT 20.63 47.049 20.682 47.085 ;
        RECT 21.014 47.049 21.068 47.085 ;
        RECT 21.896 47.049 21.95 47.085 ;
        RECT 16.964 47.2835 17.036 47.3085 ;
        RECT 18.664 47.2835 18.736 47.3085 ;
        RECT 18.964 47.2835 19.036 47.3085 ;
        RECT 14.05 47.278 14.104 47.314 ;
        RECT 14.296 47.278 14.35 47.314 ;
        RECT 14.932 47.278 14.986 47.314 ;
        RECT 15.318 47.278 15.37 47.314 ;
        RECT 15.478 47.278 15.53 47.314 ;
        RECT 15.874 47.278 15.926 47.314 ;
        RECT 16.034 47.278 16.086 47.314 ;
        RECT 16.8 47.278 16.854 47.314 ;
        RECT 18.148 47.278 18.188 47.314 ;
        RECT 19.914 47.278 19.966 47.314 ;
        RECT 20.074 47.278 20.126 47.314 ;
        RECT 20.47 47.278 20.522 47.314 ;
        RECT 20.63 47.278 20.682 47.314 ;
        RECT 21.014 47.278 21.068 47.314 ;
        RECT 21.65 47.278 21.704 47.314 ;
        RECT 21.896 47.278 21.95 47.314 ;
        RECT 17.844 47.3605 17.916 47.3855 ;
        RECT 18.356 47.355 18.396 47.391 ;
        RECT 16.964 47.7315 17.036 47.7565 ;
        RECT 17.844 47.7315 17.916 47.7565 ;
        RECT 18.964 47.7315 19.036 47.7565 ;
        RECT 14.05 47.726 14.104 47.762 ;
        RECT 14.296 47.726 14.35 47.762 ;
        RECT 14.932 47.726 14.986 47.762 ;
        RECT 15.318 47.726 15.37 47.762 ;
        RECT 15.874 47.726 15.926 47.762 ;
        RECT 16.034 47.726 16.086 47.762 ;
        RECT 18.356 47.726 18.396 47.762 ;
        RECT 19.914 47.726 19.966 47.762 ;
        RECT 20.074 47.726 20.126 47.762 ;
        RECT 20.63 47.726 20.682 47.762 ;
        RECT 21.014 47.726 21.068 47.762 ;
        RECT 21.65 47.726 21.704 47.762 ;
        RECT 21.896 47.726 21.95 47.762 ;
        RECT 17.844 47.8835 17.916 47.9085 ;
        RECT 18.356 47.878 18.396 47.914 ;
        RECT 18.664 47.9605 18.736 47.9855 ;
        RECT 18.964 47.9605 19.036 47.9855 ;
        RECT 14.296 47.955 14.35 47.991 ;
        RECT 14.932 47.955 14.986 47.991 ;
        RECT 15.318 47.955 15.37 47.991 ;
        RECT 15.478 47.955 15.53 47.991 ;
        RECT 15.874 47.955 15.926 47.991 ;
        RECT 18.148 47.955 18.188 47.991 ;
        RECT 20.074 47.955 20.126 47.991 ;
        RECT 20.47 47.955 20.522 47.991 ;
        RECT 20.63 47.955 20.682 47.991 ;
        RECT 21.014 47.955 21.068 47.991 ;
        RECT 21.65 47.955 21.704 47.991 ;
        RECT 16.964 48.2545 17.036 48.2795 ;
        RECT 17.844 48.2545 17.916 48.2795 ;
        RECT 18.664 48.2545 18.736 48.2795 ;
        RECT 18.964 48.2545 19.036 48.2795 ;
        RECT 14.05 48.249 14.104 48.285 ;
        RECT 14.932 48.249 14.986 48.285 ;
        RECT 15.318 48.249 15.37 48.285 ;
        RECT 15.478 48.249 15.53 48.285 ;
        RECT 15.874 48.249 15.926 48.285 ;
        RECT 16.034 48.249 16.086 48.285 ;
        RECT 16.8 48.249 16.854 48.285 ;
        RECT 18.148 48.249 18.188 48.285 ;
        RECT 18.356 48.249 18.396 48.285 ;
        RECT 19.914 48.249 19.966 48.285 ;
        RECT 20.074 48.249 20.126 48.285 ;
        RECT 20.47 48.249 20.522 48.285 ;
        RECT 20.63 48.249 20.682 48.285 ;
        RECT 21.014 48.249 21.068 48.285 ;
        RECT 21.896 48.249 21.95 48.285 ;
        RECT 16.964 48.4835 17.036 48.5085 ;
        RECT 18.664 48.4835 18.736 48.5085 ;
        RECT 18.964 48.4835 19.036 48.5085 ;
        RECT 14.05 48.478 14.104 48.514 ;
        RECT 14.296 48.478 14.35 48.514 ;
        RECT 14.932 48.478 14.986 48.514 ;
        RECT 15.318 48.478 15.37 48.514 ;
        RECT 15.478 48.478 15.53 48.514 ;
        RECT 15.874 48.478 15.926 48.514 ;
        RECT 16.034 48.478 16.086 48.514 ;
        RECT 16.8 48.478 16.854 48.514 ;
        RECT 18.148 48.478 18.188 48.514 ;
        RECT 19.914 48.478 19.966 48.514 ;
        RECT 20.074 48.478 20.126 48.514 ;
        RECT 20.47 48.478 20.522 48.514 ;
        RECT 20.63 48.478 20.682 48.514 ;
        RECT 21.014 48.478 21.068 48.514 ;
        RECT 21.65 48.478 21.704 48.514 ;
        RECT 21.896 48.478 21.95 48.514 ;
        RECT 17.844 48.5605 17.916 48.5855 ;
        RECT 18.356 48.555 18.396 48.591 ;
        RECT 16.964 48.9315 17.036 48.9565 ;
        RECT 17.844 48.9315 17.916 48.9565 ;
        RECT 18.964 48.9315 19.036 48.9565 ;
        RECT 14.05 48.926 14.104 48.962 ;
        RECT 14.296 48.926 14.35 48.962 ;
        RECT 14.932 48.926 14.986 48.962 ;
        RECT 15.318 48.926 15.37 48.962 ;
        RECT 15.874 48.926 15.926 48.962 ;
        RECT 16.034 48.926 16.086 48.962 ;
        RECT 18.356 48.926 18.396 48.962 ;
        RECT 19.914 48.926 19.966 48.962 ;
        RECT 20.074 48.926 20.126 48.962 ;
        RECT 20.63 48.926 20.682 48.962 ;
        RECT 21.014 48.926 21.068 48.962 ;
        RECT 21.65 48.926 21.704 48.962 ;
        RECT 21.896 48.926 21.95 48.962 ;
        RECT 17.844 49.0835 17.916 49.1085 ;
        RECT 18.356 49.078 18.396 49.114 ;
        RECT 18.664 49.1605 18.736 49.1855 ;
        RECT 18.964 49.1605 19.036 49.1855 ;
        RECT 14.296 49.155 14.35 49.191 ;
        RECT 14.932 49.155 14.986 49.191 ;
        RECT 15.318 49.155 15.37 49.191 ;
        RECT 15.478 49.155 15.53 49.191 ;
        RECT 15.874 49.155 15.926 49.191 ;
        RECT 18.148 49.155 18.188 49.191 ;
        RECT 20.074 49.155 20.126 49.191 ;
        RECT 20.47 49.155 20.522 49.191 ;
        RECT 20.63 49.155 20.682 49.191 ;
        RECT 21.014 49.155 21.068 49.191 ;
        RECT 21.65 49.155 21.704 49.191 ;
        RECT 16.964 49.4545 17.036 49.4795 ;
        RECT 17.844 49.4545 17.916 49.4795 ;
        RECT 18.664 49.4545 18.736 49.4795 ;
        RECT 18.964 49.4545 19.036 49.4795 ;
        RECT 14.05 49.449 14.104 49.485 ;
        RECT 14.932 49.449 14.986 49.485 ;
        RECT 15.318 49.449 15.37 49.485 ;
        RECT 15.478 49.449 15.53 49.485 ;
        RECT 15.874 49.449 15.926 49.485 ;
        RECT 16.034 49.449 16.086 49.485 ;
        RECT 16.8 49.449 16.854 49.485 ;
        RECT 18.148 49.449 18.188 49.485 ;
        RECT 18.356 49.449 18.396 49.485 ;
        RECT 19.914 49.449 19.966 49.485 ;
        RECT 20.074 49.449 20.126 49.485 ;
        RECT 20.47 49.449 20.522 49.485 ;
        RECT 20.63 49.449 20.682 49.485 ;
        RECT 21.014 49.449 21.068 49.485 ;
        RECT 21.896 49.449 21.95 49.485 ;
        RECT 16.964 49.6835 17.036 49.7085 ;
        RECT 18.664 49.6835 18.736 49.7085 ;
        RECT 18.964 49.6835 19.036 49.7085 ;
        RECT 14.05 49.678 14.104 49.714 ;
        RECT 14.296 49.678 14.35 49.714 ;
        RECT 14.932 49.678 14.986 49.714 ;
        RECT 15.318 49.678 15.37 49.714 ;
        RECT 15.478 49.678 15.53 49.714 ;
        RECT 15.874 49.678 15.926 49.714 ;
        RECT 16.034 49.678 16.086 49.714 ;
        RECT 16.8 49.678 16.854 49.714 ;
        RECT 18.148 49.678 18.188 49.714 ;
        RECT 19.914 49.678 19.966 49.714 ;
        RECT 20.074 49.678 20.126 49.714 ;
        RECT 20.47 49.678 20.522 49.714 ;
        RECT 20.63 49.678 20.682 49.714 ;
        RECT 21.014 49.678 21.068 49.714 ;
        RECT 21.65 49.678 21.704 49.714 ;
        RECT 21.896 49.678 21.95 49.714 ;
        RECT 17.844 49.7605 17.916 49.7855 ;
        RECT 18.356 49.755 18.396 49.791 ;
        RECT 16.964 50.1315 17.036 50.1565 ;
        RECT 17.844 50.1315 17.916 50.1565 ;
        RECT 18.964 50.1315 19.036 50.1565 ;
        RECT 14.05 50.126 14.104 50.162 ;
        RECT 14.296 50.126 14.35 50.162 ;
        RECT 14.932 50.126 14.986 50.162 ;
        RECT 15.318 50.126 15.37 50.162 ;
        RECT 15.874 50.126 15.926 50.162 ;
        RECT 16.034 50.126 16.086 50.162 ;
        RECT 18.356 50.126 18.396 50.162 ;
        RECT 19.914 50.126 19.966 50.162 ;
        RECT 20.074 50.126 20.126 50.162 ;
        RECT 20.63 50.126 20.682 50.162 ;
        RECT 21.014 50.126 21.068 50.162 ;
        RECT 21.65 50.126 21.704 50.162 ;
        RECT 21.896 50.126 21.95 50.162 ;
        RECT 17.844 50.2835 17.916 50.3085 ;
        RECT 18.356 50.278 18.396 50.314 ;
        RECT 18.664 50.3605 18.736 50.3855 ;
        RECT 18.964 50.3605 19.036 50.3855 ;
        RECT 14.296 50.355 14.35 50.391 ;
        RECT 14.932 50.355 14.986 50.391 ;
        RECT 15.318 50.355 15.37 50.391 ;
        RECT 15.478 50.355 15.53 50.391 ;
        RECT 15.874 50.355 15.926 50.391 ;
        RECT 18.148 50.355 18.188 50.391 ;
        RECT 20.074 50.355 20.126 50.391 ;
        RECT 20.47 50.355 20.522 50.391 ;
        RECT 20.63 50.355 20.682 50.391 ;
        RECT 21.014 50.355 21.068 50.391 ;
        RECT 21.65 50.355 21.704 50.391 ;
        RECT 16.964 50.6545 17.036 50.6795 ;
        RECT 17.844 50.6545 17.916 50.6795 ;
        RECT 18.664 50.6545 18.736 50.6795 ;
        RECT 18.964 50.6545 19.036 50.6795 ;
        RECT 14.05 50.649 14.104 50.685 ;
        RECT 14.932 50.649 14.986 50.685 ;
        RECT 15.318 50.649 15.37 50.685 ;
        RECT 15.478 50.649 15.53 50.685 ;
        RECT 15.874 50.649 15.926 50.685 ;
        RECT 16.034 50.649 16.086 50.685 ;
        RECT 16.8 50.649 16.854 50.685 ;
        RECT 18.148 50.649 18.188 50.685 ;
        RECT 18.356 50.649 18.396 50.685 ;
        RECT 19.914 50.649 19.966 50.685 ;
        RECT 20.074 50.649 20.126 50.685 ;
        RECT 20.47 50.649 20.522 50.685 ;
        RECT 20.63 50.649 20.682 50.685 ;
        RECT 21.014 50.649 21.068 50.685 ;
        RECT 21.896 50.649 21.95 50.685 ;
        RECT 16.964 50.8835 17.036 50.9085 ;
        RECT 18.664 50.8835 18.736 50.9085 ;
        RECT 18.964 50.8835 19.036 50.9085 ;
        RECT 14.05 50.878 14.104 50.914 ;
        RECT 14.296 50.878 14.35 50.914 ;
        RECT 14.932 50.878 14.986 50.914 ;
        RECT 15.318 50.878 15.37 50.914 ;
        RECT 15.478 50.878 15.53 50.914 ;
        RECT 15.874 50.878 15.926 50.914 ;
        RECT 16.034 50.878 16.086 50.914 ;
        RECT 16.8 50.878 16.854 50.914 ;
        RECT 18.148 50.878 18.188 50.914 ;
        RECT 19.914 50.878 19.966 50.914 ;
        RECT 20.074 50.878 20.126 50.914 ;
        RECT 20.47 50.878 20.522 50.914 ;
        RECT 20.63 50.878 20.682 50.914 ;
        RECT 21.014 50.878 21.068 50.914 ;
        RECT 21.65 50.878 21.704 50.914 ;
        RECT 21.896 50.878 21.95 50.914 ;
        RECT 17.844 50.9605 17.916 50.9855 ;
        RECT 18.356 50.955 18.396 50.991 ;
        RECT 16.964 51.3315 17.036 51.3565 ;
        RECT 17.844 51.3315 17.916 51.3565 ;
        RECT 18.964 51.3315 19.036 51.3565 ;
        RECT 14.05 51.326 14.104 51.362 ;
        RECT 14.296 51.326 14.35 51.362 ;
        RECT 14.932 51.326 14.986 51.362 ;
        RECT 15.318 51.326 15.37 51.362 ;
        RECT 15.874 51.326 15.926 51.362 ;
        RECT 16.034 51.326 16.086 51.362 ;
        RECT 18.356 51.326 18.396 51.362 ;
        RECT 19.914 51.326 19.966 51.362 ;
        RECT 20.074 51.326 20.126 51.362 ;
        RECT 20.63 51.326 20.682 51.362 ;
        RECT 21.014 51.326 21.068 51.362 ;
        RECT 21.65 51.326 21.704 51.362 ;
        RECT 21.896 51.326 21.95 51.362 ;
        RECT 17.844 51.4835 17.916 51.5085 ;
        RECT 18.356 51.478 18.396 51.514 ;
        RECT 18.664 51.5605 18.736 51.5855 ;
        RECT 18.964 51.5605 19.036 51.5855 ;
        RECT 14.296 51.555 14.35 51.591 ;
        RECT 14.932 51.555 14.986 51.591 ;
        RECT 15.318 51.555 15.37 51.591 ;
        RECT 15.478 51.555 15.53 51.591 ;
        RECT 15.874 51.555 15.926 51.591 ;
        RECT 18.148 51.555 18.188 51.591 ;
        RECT 20.074 51.555 20.126 51.591 ;
        RECT 20.47 51.555 20.522 51.591 ;
        RECT 20.63 51.555 20.682 51.591 ;
        RECT 21.014 51.555 21.068 51.591 ;
        RECT 21.65 51.555 21.704 51.591 ;
        RECT 16.964 51.8545 17.036 51.8795 ;
        RECT 17.844 51.8545 17.916 51.8795 ;
        RECT 18.664 51.8545 18.736 51.8795 ;
        RECT 18.964 51.8545 19.036 51.8795 ;
        RECT 14.05 51.849 14.104 51.885 ;
        RECT 14.932 51.849 14.986 51.885 ;
        RECT 15.318 51.849 15.37 51.885 ;
        RECT 15.478 51.849 15.53 51.885 ;
        RECT 15.874 51.849 15.926 51.885 ;
        RECT 16.034 51.849 16.086 51.885 ;
        RECT 16.8 51.849 16.854 51.885 ;
        RECT 18.148 51.849 18.188 51.885 ;
        RECT 18.356 51.849 18.396 51.885 ;
        RECT 19.914 51.849 19.966 51.885 ;
        RECT 20.074 51.849 20.126 51.885 ;
        RECT 20.47 51.849 20.522 51.885 ;
        RECT 20.63 51.849 20.682 51.885 ;
        RECT 21.014 51.849 21.068 51.885 ;
        RECT 21.896 51.849 21.95 51.885 ;
        RECT 16.964 52.0835 17.036 52.1085 ;
        RECT 18.664 52.0835 18.736 52.1085 ;
        RECT 18.964 52.0835 19.036 52.1085 ;
        RECT 14.05 52.078 14.104 52.114 ;
        RECT 14.296 52.078 14.35 52.114 ;
        RECT 14.932 52.078 14.986 52.114 ;
        RECT 15.318 52.078 15.37 52.114 ;
        RECT 15.478 52.078 15.53 52.114 ;
        RECT 15.874 52.078 15.926 52.114 ;
        RECT 16.034 52.078 16.086 52.114 ;
        RECT 16.8 52.078 16.854 52.114 ;
        RECT 18.148 52.078 18.188 52.114 ;
        RECT 19.914 52.078 19.966 52.114 ;
        RECT 20.074 52.078 20.126 52.114 ;
        RECT 20.47 52.078 20.522 52.114 ;
        RECT 20.63 52.078 20.682 52.114 ;
        RECT 21.014 52.078 21.068 52.114 ;
        RECT 21.65 52.078 21.704 52.114 ;
        RECT 21.896 52.078 21.95 52.114 ;
        RECT 17.844 52.1605 17.916 52.1855 ;
        RECT 18.356 52.155 18.396 52.191 ;
        RECT 16.964 52.5315 17.036 52.5565 ;
        RECT 17.844 52.5315 17.916 52.5565 ;
        RECT 18.964 52.5315 19.036 52.5565 ;
        RECT 14.05 52.526 14.104 52.562 ;
        RECT 14.296 52.526 14.35 52.562 ;
        RECT 14.932 52.526 14.986 52.562 ;
        RECT 15.318 52.526 15.37 52.562 ;
        RECT 15.874 52.526 15.926 52.562 ;
        RECT 16.034 52.526 16.086 52.562 ;
        RECT 18.356 52.526 18.396 52.562 ;
        RECT 19.914 52.526 19.966 52.562 ;
        RECT 20.074 52.526 20.126 52.562 ;
        RECT 20.63 52.526 20.682 52.562 ;
        RECT 21.014 52.526 21.068 52.562 ;
        RECT 21.65 52.526 21.704 52.562 ;
        RECT 21.896 52.526 21.95 52.562 ;
        RECT 17.844 52.6835 17.916 52.7085 ;
        RECT 18.356 52.678 18.396 52.714 ;
        RECT 18.664 52.7605 18.736 52.7855 ;
        RECT 18.964 52.7605 19.036 52.7855 ;
        RECT 14.296 52.755 14.35 52.791 ;
        RECT 14.932 52.755 14.986 52.791 ;
        RECT 15.318 52.755 15.37 52.791 ;
        RECT 15.478 52.755 15.53 52.791 ;
        RECT 15.874 52.755 15.926 52.791 ;
        RECT 18.148 52.755 18.188 52.791 ;
        RECT 20.074 52.755 20.126 52.791 ;
        RECT 20.47 52.755 20.522 52.791 ;
        RECT 20.63 52.755 20.682 52.791 ;
        RECT 21.014 52.755 21.068 52.791 ;
        RECT 21.65 52.755 21.704 52.791 ;
        RECT 16.964 53.0545 17.036 53.0795 ;
        RECT 17.844 53.0545 17.916 53.0795 ;
        RECT 18.664 53.0545 18.736 53.0795 ;
        RECT 18.964 53.0545 19.036 53.0795 ;
        RECT 14.05 53.049 14.104 53.085 ;
        RECT 14.932 53.049 14.986 53.085 ;
        RECT 15.318 53.049 15.37 53.085 ;
        RECT 15.478 53.049 15.53 53.085 ;
        RECT 15.874 53.049 15.926 53.085 ;
        RECT 16.034 53.049 16.086 53.085 ;
        RECT 16.8 53.049 16.854 53.085 ;
        RECT 18.148 53.049 18.188 53.085 ;
        RECT 18.356 53.049 18.396 53.085 ;
        RECT 19.914 53.049 19.966 53.085 ;
        RECT 20.074 53.049 20.126 53.085 ;
        RECT 20.47 53.049 20.522 53.085 ;
        RECT 20.63 53.049 20.682 53.085 ;
        RECT 21.014 53.049 21.068 53.085 ;
        RECT 21.896 53.049 21.95 53.085 ;
        RECT 16.964 53.2835 17.036 53.3085 ;
        RECT 18.664 53.2835 18.736 53.3085 ;
        RECT 18.964 53.2835 19.036 53.3085 ;
        RECT 14.05 53.278 14.104 53.314 ;
        RECT 14.296 53.278 14.35 53.314 ;
        RECT 14.932 53.278 14.986 53.314 ;
        RECT 15.318 53.278 15.37 53.314 ;
        RECT 15.478 53.278 15.53 53.314 ;
        RECT 15.874 53.278 15.926 53.314 ;
        RECT 16.034 53.278 16.086 53.314 ;
        RECT 16.8 53.278 16.854 53.314 ;
        RECT 18.148 53.278 18.188 53.314 ;
        RECT 19.914 53.278 19.966 53.314 ;
        RECT 20.074 53.278 20.126 53.314 ;
        RECT 20.47 53.278 20.522 53.314 ;
        RECT 20.63 53.278 20.682 53.314 ;
        RECT 21.014 53.278 21.068 53.314 ;
        RECT 21.65 53.278 21.704 53.314 ;
        RECT 21.896 53.278 21.95 53.314 ;
        RECT 17.844 53.3605 17.916 53.3855 ;
        RECT 18.356 53.355 18.396 53.391 ;
        RECT 16.964 53.7315 17.036 53.7565 ;
        RECT 17.844 53.7315 17.916 53.7565 ;
        RECT 18.964 53.7315 19.036 53.7565 ;
        RECT 14.05 53.726 14.104 53.762 ;
        RECT 14.296 53.726 14.35 53.762 ;
        RECT 14.932 53.726 14.986 53.762 ;
        RECT 15.318 53.726 15.37 53.762 ;
        RECT 15.874 53.726 15.926 53.762 ;
        RECT 16.034 53.726 16.086 53.762 ;
        RECT 18.356 53.726 18.396 53.762 ;
        RECT 19.914 53.726 19.966 53.762 ;
        RECT 20.074 53.726 20.126 53.762 ;
        RECT 20.63 53.726 20.682 53.762 ;
        RECT 21.014 53.726 21.068 53.762 ;
        RECT 21.65 53.726 21.704 53.762 ;
        RECT 21.896 53.726 21.95 53.762 ;
        RECT 17.844 53.8835 17.916 53.9085 ;
        RECT 18.356 53.878 18.396 53.914 ;
        RECT 18.664 53.9605 18.736 53.9855 ;
        RECT 18.964 53.9605 19.036 53.9855 ;
        RECT 14.296 53.955 14.35 53.991 ;
        RECT 14.932 53.955 14.986 53.991 ;
        RECT 15.318 53.955 15.37 53.991 ;
        RECT 15.478 53.955 15.53 53.991 ;
        RECT 15.874 53.955 15.926 53.991 ;
        RECT 18.148 53.955 18.188 53.991 ;
        RECT 20.074 53.955 20.126 53.991 ;
        RECT 20.47 53.955 20.522 53.991 ;
        RECT 20.63 53.955 20.682 53.991 ;
        RECT 21.014 53.955 21.068 53.991 ;
        RECT 21.65 53.955 21.704 53.991 ;
        RECT 16.964 54.2545 17.036 54.2795 ;
        RECT 17.844 54.2545 17.916 54.2795 ;
        RECT 18.664 54.2545 18.736 54.2795 ;
        RECT 18.964 54.2545 19.036 54.2795 ;
        RECT 14.05 54.249 14.104 54.285 ;
        RECT 14.932 54.249 14.986 54.285 ;
        RECT 15.318 54.249 15.37 54.285 ;
        RECT 15.478 54.249 15.53 54.285 ;
        RECT 15.874 54.249 15.926 54.285 ;
        RECT 16.034 54.249 16.086 54.285 ;
        RECT 16.8 54.249 16.854 54.285 ;
        RECT 18.148 54.249 18.188 54.285 ;
        RECT 18.356 54.249 18.396 54.285 ;
        RECT 19.914 54.249 19.966 54.285 ;
        RECT 20.074 54.249 20.126 54.285 ;
        RECT 20.47 54.249 20.522 54.285 ;
        RECT 20.63 54.249 20.682 54.285 ;
        RECT 21.014 54.249 21.068 54.285 ;
        RECT 21.896 54.249 21.95 54.285 ;
        RECT 16.964 54.4835 17.036 54.5085 ;
        RECT 18.664 54.4835 18.736 54.5085 ;
        RECT 18.964 54.4835 19.036 54.5085 ;
        RECT 14.05 54.478 14.104 54.514 ;
        RECT 14.296 54.478 14.35 54.514 ;
        RECT 14.932 54.478 14.986 54.514 ;
        RECT 15.318 54.478 15.37 54.514 ;
        RECT 15.478 54.478 15.53 54.514 ;
        RECT 15.874 54.478 15.926 54.514 ;
        RECT 16.034 54.478 16.086 54.514 ;
        RECT 16.8 54.478 16.854 54.514 ;
        RECT 18.148 54.478 18.188 54.514 ;
        RECT 19.914 54.478 19.966 54.514 ;
        RECT 20.074 54.478 20.126 54.514 ;
        RECT 20.47 54.478 20.522 54.514 ;
        RECT 20.63 54.478 20.682 54.514 ;
        RECT 21.014 54.478 21.068 54.514 ;
        RECT 21.65 54.478 21.704 54.514 ;
        RECT 21.896 54.478 21.95 54.514 ;
        RECT 17.844 54.5605 17.916 54.5855 ;
        RECT 18.356 54.555 18.396 54.591 ;
        RECT 16.964 54.9315 17.036 54.9565 ;
        RECT 17.844 54.9315 17.916 54.9565 ;
        RECT 18.964 54.9315 19.036 54.9565 ;
        RECT 14.05 54.926 14.104 54.962 ;
        RECT 14.296 54.926 14.35 54.962 ;
        RECT 14.932 54.926 14.986 54.962 ;
        RECT 15.318 54.926 15.37 54.962 ;
        RECT 15.874 54.926 15.926 54.962 ;
        RECT 16.034 54.926 16.086 54.962 ;
        RECT 18.356 54.926 18.396 54.962 ;
        RECT 19.914 54.926 19.966 54.962 ;
        RECT 20.074 54.926 20.126 54.962 ;
        RECT 20.63 54.926 20.682 54.962 ;
        RECT 21.014 54.926 21.068 54.962 ;
        RECT 21.65 54.926 21.704 54.962 ;
        RECT 21.896 54.926 21.95 54.962 ;
        RECT 17.844 55.0835 17.916 55.1085 ;
        RECT 18.356 55.078 18.396 55.114 ;
        RECT 18.664 55.1605 18.736 55.1855 ;
        RECT 18.964 55.1605 19.036 55.1855 ;
        RECT 14.296 55.155 14.35 55.191 ;
        RECT 14.932 55.155 14.986 55.191 ;
        RECT 15.318 55.155 15.37 55.191 ;
        RECT 15.478 55.155 15.53 55.191 ;
        RECT 15.874 55.155 15.926 55.191 ;
        RECT 18.148 55.155 18.188 55.191 ;
        RECT 20.074 55.155 20.126 55.191 ;
        RECT 20.47 55.155 20.522 55.191 ;
        RECT 20.63 55.155 20.682 55.191 ;
        RECT 21.014 55.155 21.068 55.191 ;
        RECT 21.65 55.155 21.704 55.191 ;
        RECT 16.964 55.4545 17.036 55.4795 ;
        RECT 17.844 55.4545 17.916 55.4795 ;
        RECT 18.664 55.4545 18.736 55.4795 ;
        RECT 18.964 55.4545 19.036 55.4795 ;
        RECT 14.05 55.449 14.104 55.485 ;
        RECT 14.932 55.449 14.986 55.485 ;
        RECT 15.318 55.449 15.37 55.485 ;
        RECT 15.478 55.449 15.53 55.485 ;
        RECT 15.874 55.449 15.926 55.485 ;
        RECT 16.034 55.449 16.086 55.485 ;
        RECT 16.8 55.449 16.854 55.485 ;
        RECT 18.148 55.449 18.188 55.485 ;
        RECT 18.356 55.449 18.396 55.485 ;
        RECT 19.914 55.449 19.966 55.485 ;
        RECT 20.074 55.449 20.126 55.485 ;
        RECT 20.47 55.449 20.522 55.485 ;
        RECT 20.63 55.449 20.682 55.485 ;
        RECT 21.014 55.449 21.068 55.485 ;
        RECT 21.896 55.449 21.95 55.485 ;
        RECT 16.964 55.6835 17.036 55.7085 ;
        RECT 18.664 55.6835 18.736 55.7085 ;
        RECT 18.964 55.6835 19.036 55.7085 ;
        RECT 14.05 55.678 14.104 55.714 ;
        RECT 14.296 55.678 14.35 55.714 ;
        RECT 14.932 55.678 14.986 55.714 ;
        RECT 15.318 55.678 15.37 55.714 ;
        RECT 15.478 55.678 15.53 55.714 ;
        RECT 15.874 55.678 15.926 55.714 ;
        RECT 16.034 55.678 16.086 55.714 ;
        RECT 16.8 55.678 16.854 55.714 ;
        RECT 18.148 55.678 18.188 55.714 ;
        RECT 19.914 55.678 19.966 55.714 ;
        RECT 20.074 55.678 20.126 55.714 ;
        RECT 20.47 55.678 20.522 55.714 ;
        RECT 20.63 55.678 20.682 55.714 ;
        RECT 21.014 55.678 21.068 55.714 ;
        RECT 21.65 55.678 21.704 55.714 ;
        RECT 21.896 55.678 21.95 55.714 ;
        RECT 17.844 55.7605 17.916 55.7855 ;
        RECT 18.356 55.755 18.396 55.791 ;
        RECT 16.964 56.1315 17.036 56.1565 ;
        RECT 17.844 56.1315 17.916 56.1565 ;
        RECT 18.964 56.1315 19.036 56.1565 ;
        RECT 14.05 56.126 14.104 56.162 ;
        RECT 14.296 56.126 14.35 56.162 ;
        RECT 14.932 56.126 14.986 56.162 ;
        RECT 15.318 56.126 15.37 56.162 ;
        RECT 15.874 56.126 15.926 56.162 ;
        RECT 16.034 56.126 16.086 56.162 ;
        RECT 18.356 56.126 18.396 56.162 ;
        RECT 19.914 56.126 19.966 56.162 ;
        RECT 20.074 56.126 20.126 56.162 ;
        RECT 20.63 56.126 20.682 56.162 ;
        RECT 21.014 56.126 21.068 56.162 ;
        RECT 21.65 56.126 21.704 56.162 ;
        RECT 21.896 56.126 21.95 56.162 ;
        RECT 17.844 56.2835 17.916 56.3085 ;
        RECT 18.356 56.278 18.396 56.314 ;
        RECT 18.664 56.3605 18.736 56.3855 ;
        RECT 18.964 56.3605 19.036 56.3855 ;
        RECT 14.296 56.355 14.35 56.391 ;
        RECT 14.932 56.355 14.986 56.391 ;
        RECT 15.318 56.355 15.37 56.391 ;
        RECT 15.478 56.355 15.53 56.391 ;
        RECT 15.874 56.355 15.926 56.391 ;
        RECT 18.148 56.355 18.188 56.391 ;
        RECT 20.074 56.355 20.126 56.391 ;
        RECT 20.47 56.355 20.522 56.391 ;
        RECT 20.63 56.355 20.682 56.391 ;
        RECT 21.014 56.355 21.068 56.391 ;
        RECT 21.65 56.355 21.704 56.391 ;
        RECT 16.964 56.6545 17.036 56.6795 ;
        RECT 17.844 56.6545 17.916 56.6795 ;
        RECT 18.664 56.6545 18.736 56.6795 ;
        RECT 18.964 56.6545 19.036 56.6795 ;
        RECT 14.05 56.649 14.104 56.685 ;
        RECT 14.932 56.649 14.986 56.685 ;
        RECT 15.318 56.649 15.37 56.685 ;
        RECT 15.478 56.649 15.53 56.685 ;
        RECT 15.874 56.649 15.926 56.685 ;
        RECT 16.034 56.649 16.086 56.685 ;
        RECT 16.8 56.649 16.854 56.685 ;
        RECT 18.148 56.649 18.188 56.685 ;
        RECT 18.356 56.649 18.396 56.685 ;
        RECT 19.914 56.649 19.966 56.685 ;
        RECT 20.074 56.649 20.126 56.685 ;
        RECT 20.47 56.649 20.522 56.685 ;
        RECT 20.63 56.649 20.682 56.685 ;
        RECT 21.014 56.649 21.068 56.685 ;
        RECT 21.896 56.649 21.95 56.685 ;
        RECT 16.964 56.8835 17.036 56.9085 ;
        RECT 18.664 56.8835 18.736 56.9085 ;
        RECT 18.964 56.8835 19.036 56.9085 ;
        RECT 14.05 56.878 14.104 56.914 ;
        RECT 14.296 56.878 14.35 56.914 ;
        RECT 14.932 56.878 14.986 56.914 ;
        RECT 15.318 56.878 15.37 56.914 ;
        RECT 15.478 56.878 15.53 56.914 ;
        RECT 15.874 56.878 15.926 56.914 ;
        RECT 16.034 56.878 16.086 56.914 ;
        RECT 16.8 56.878 16.854 56.914 ;
        RECT 18.148 56.878 18.188 56.914 ;
        RECT 19.914 56.878 19.966 56.914 ;
        RECT 20.074 56.878 20.126 56.914 ;
        RECT 20.47 56.878 20.522 56.914 ;
        RECT 20.63 56.878 20.682 56.914 ;
        RECT 21.014 56.878 21.068 56.914 ;
        RECT 21.65 56.878 21.704 56.914 ;
        RECT 21.896 56.878 21.95 56.914 ;
        RECT 17.844 56.9605 17.916 56.9855 ;
        RECT 18.356 56.955 18.396 56.991 ;
        RECT 16.964 57.3315 17.036 57.3565 ;
        RECT 17.844 57.3315 17.916 57.3565 ;
        RECT 18.964 57.3315 19.036 57.3565 ;
        RECT 14.05 57.326 14.104 57.362 ;
        RECT 14.296 57.326 14.35 57.362 ;
        RECT 14.932 57.326 14.986 57.362 ;
        RECT 15.318 57.326 15.37 57.362 ;
        RECT 15.874 57.326 15.926 57.362 ;
        RECT 16.034 57.326 16.086 57.362 ;
        RECT 18.356 57.326 18.396 57.362 ;
        RECT 19.914 57.326 19.966 57.362 ;
        RECT 20.074 57.326 20.126 57.362 ;
        RECT 20.63 57.326 20.682 57.362 ;
        RECT 21.014 57.326 21.068 57.362 ;
        RECT 21.65 57.326 21.704 57.362 ;
        RECT 21.896 57.326 21.95 57.362 ;
        RECT 17.844 57.4835 17.916 57.5085 ;
        RECT 18.356 57.478 18.396 57.514 ;
        RECT 18.664 57.5605 18.736 57.5855 ;
        RECT 18.964 57.5605 19.036 57.5855 ;
        RECT 14.296 57.555 14.35 57.591 ;
        RECT 14.932 57.555 14.986 57.591 ;
        RECT 15.318 57.555 15.37 57.591 ;
        RECT 15.478 57.555 15.53 57.591 ;
        RECT 15.874 57.555 15.926 57.591 ;
        RECT 18.148 57.555 18.188 57.591 ;
        RECT 20.074 57.555 20.126 57.591 ;
        RECT 20.47 57.555 20.522 57.591 ;
        RECT 20.63 57.555 20.682 57.591 ;
        RECT 21.014 57.555 21.068 57.591 ;
        RECT 21.65 57.555 21.704 57.591 ;
        RECT 16.964 57.8545 17.036 57.8795 ;
        RECT 17.844 57.8545 17.916 57.8795 ;
        RECT 18.664 57.8545 18.736 57.8795 ;
        RECT 18.964 57.8545 19.036 57.8795 ;
        RECT 14.05 57.849 14.104 57.885 ;
        RECT 14.932 57.849 14.986 57.885 ;
        RECT 15.318 57.849 15.37 57.885 ;
        RECT 15.478 57.849 15.53 57.885 ;
        RECT 15.874 57.849 15.926 57.885 ;
        RECT 16.034 57.849 16.086 57.885 ;
        RECT 16.8 57.849 16.854 57.885 ;
        RECT 18.148 57.849 18.188 57.885 ;
        RECT 18.356 57.849 18.396 57.885 ;
        RECT 19.914 57.849 19.966 57.885 ;
        RECT 20.074 57.849 20.126 57.885 ;
        RECT 20.47 57.849 20.522 57.885 ;
        RECT 20.63 57.849 20.682 57.885 ;
        RECT 21.014 57.849 21.068 57.885 ;
        RECT 21.896 57.849 21.95 57.885 ;
        RECT 16.964 58.0835 17.036 58.1085 ;
        RECT 18.664 58.0835 18.736 58.1085 ;
        RECT 18.964 58.0835 19.036 58.1085 ;
        RECT 14.05 58.078 14.104 58.114 ;
        RECT 14.296 58.078 14.35 58.114 ;
        RECT 14.932 58.078 14.986 58.114 ;
        RECT 15.318 58.078 15.37 58.114 ;
        RECT 15.478 58.078 15.53 58.114 ;
        RECT 15.874 58.078 15.926 58.114 ;
        RECT 16.034 58.078 16.086 58.114 ;
        RECT 16.8 58.078 16.854 58.114 ;
        RECT 18.148 58.078 18.188 58.114 ;
        RECT 19.914 58.078 19.966 58.114 ;
        RECT 20.074 58.078 20.126 58.114 ;
        RECT 20.47 58.078 20.522 58.114 ;
        RECT 20.63 58.078 20.682 58.114 ;
        RECT 21.014 58.078 21.068 58.114 ;
        RECT 21.65 58.078 21.704 58.114 ;
        RECT 21.896 58.078 21.95 58.114 ;
        RECT 17.844 58.1605 17.916 58.1855 ;
        RECT 18.356 58.155 18.396 58.191 ;
        RECT 16.964 58.5315 17.036 58.5565 ;
        RECT 17.844 58.5315 17.916 58.5565 ;
        RECT 18.964 58.5315 19.036 58.5565 ;
        RECT 14.05 58.526 14.104 58.562 ;
        RECT 14.296 58.526 14.35 58.562 ;
        RECT 14.932 58.526 14.986 58.562 ;
        RECT 15.318 58.526 15.37 58.562 ;
        RECT 15.874 58.526 15.926 58.562 ;
        RECT 16.034 58.526 16.086 58.562 ;
        RECT 18.356 58.526 18.396 58.562 ;
        RECT 19.914 58.526 19.966 58.562 ;
        RECT 20.074 58.526 20.126 58.562 ;
        RECT 20.63 58.526 20.682 58.562 ;
        RECT 21.014 58.526 21.068 58.562 ;
        RECT 21.65 58.526 21.704 58.562 ;
        RECT 21.896 58.526 21.95 58.562 ;
        RECT 17.844 58.6835 17.916 58.7085 ;
        RECT 18.356 58.678 18.396 58.714 ;
        RECT 18.664 58.7605 18.736 58.7855 ;
        RECT 18.964 58.7605 19.036 58.7855 ;
        RECT 14.296 58.755 14.35 58.791 ;
        RECT 14.932 58.755 14.986 58.791 ;
        RECT 15.318 58.755 15.37 58.791 ;
        RECT 15.478 58.755 15.53 58.791 ;
        RECT 15.874 58.755 15.926 58.791 ;
        RECT 18.148 58.755 18.188 58.791 ;
        RECT 20.074 58.755 20.126 58.791 ;
        RECT 20.47 58.755 20.522 58.791 ;
        RECT 20.63 58.755 20.682 58.791 ;
        RECT 21.014 58.755 21.068 58.791 ;
        RECT 21.65 58.755 21.704 58.791 ;
        RECT 16.964 59.0545 17.036 59.0795 ;
        RECT 17.844 59.0545 17.916 59.0795 ;
        RECT 18.664 59.0545 18.736 59.0795 ;
        RECT 18.964 59.0545 19.036 59.0795 ;
        RECT 14.05 59.049 14.104 59.085 ;
        RECT 14.932 59.049 14.986 59.085 ;
        RECT 15.318 59.049 15.37 59.085 ;
        RECT 15.478 59.049 15.53 59.085 ;
        RECT 15.874 59.049 15.926 59.085 ;
        RECT 16.034 59.049 16.086 59.085 ;
        RECT 16.8 59.049 16.854 59.085 ;
        RECT 18.148 59.049 18.188 59.085 ;
        RECT 18.356 59.049 18.396 59.085 ;
        RECT 19.914 59.049 19.966 59.085 ;
        RECT 20.074 59.049 20.126 59.085 ;
        RECT 20.47 59.049 20.522 59.085 ;
        RECT 20.63 59.049 20.682 59.085 ;
        RECT 21.014 59.049 21.068 59.085 ;
        RECT 21.896 59.049 21.95 59.085 ;
        RECT 16.964 59.2835 17.036 59.3085 ;
        RECT 18.664 59.2835 18.736 59.3085 ;
        RECT 18.964 59.2835 19.036 59.3085 ;
        RECT 14.05 59.278 14.104 59.314 ;
        RECT 14.296 59.278 14.35 59.314 ;
        RECT 14.932 59.278 14.986 59.314 ;
        RECT 15.318 59.278 15.37 59.314 ;
        RECT 15.478 59.278 15.53 59.314 ;
        RECT 15.874 59.278 15.926 59.314 ;
        RECT 16.034 59.278 16.086 59.314 ;
        RECT 16.8 59.278 16.854 59.314 ;
        RECT 18.148 59.278 18.188 59.314 ;
        RECT 19.914 59.278 19.966 59.314 ;
        RECT 20.074 59.278 20.126 59.314 ;
        RECT 20.47 59.278 20.522 59.314 ;
        RECT 20.63 59.278 20.682 59.314 ;
        RECT 21.014 59.278 21.068 59.314 ;
        RECT 21.65 59.278 21.704 59.314 ;
        RECT 21.896 59.278 21.95 59.314 ;
        RECT 17.844 59.3605 17.916 59.3855 ;
        RECT 18.356 59.355 18.396 59.391 ;
        RECT 16.964 59.7315 17.036 59.7565 ;
        RECT 17.844 59.7315 17.916 59.7565 ;
        RECT 18.964 59.7315 19.036 59.7565 ;
        RECT 14.05 59.726 14.104 59.762 ;
        RECT 14.296 59.726 14.35 59.762 ;
        RECT 14.932 59.726 14.986 59.762 ;
        RECT 15.318 59.726 15.37 59.762 ;
        RECT 15.874 59.726 15.926 59.762 ;
        RECT 16.034 59.726 16.086 59.762 ;
        RECT 18.356 59.726 18.396 59.762 ;
        RECT 19.914 59.726 19.966 59.762 ;
        RECT 20.074 59.726 20.126 59.762 ;
        RECT 20.63 59.726 20.682 59.762 ;
        RECT 21.014 59.726 21.068 59.762 ;
        RECT 21.65 59.726 21.704 59.762 ;
        RECT 21.896 59.726 21.95 59.762 ;
        RECT 17.844 59.8835 17.916 59.9085 ;
        RECT 18.356 59.878 18.396 59.914 ;
        RECT 18.664 59.9605 18.736 59.9855 ;
        RECT 18.964 59.9605 19.036 59.9855 ;
        RECT 14.296 59.955 14.35 59.991 ;
        RECT 14.932 59.955 14.986 59.991 ;
        RECT 15.318 59.955 15.37 59.991 ;
        RECT 15.478 59.955 15.53 59.991 ;
        RECT 15.874 59.955 15.926 59.991 ;
        RECT 18.148 59.955 18.188 59.991 ;
        RECT 20.074 59.955 20.126 59.991 ;
        RECT 20.47 59.955 20.522 59.991 ;
        RECT 20.63 59.955 20.682 59.991 ;
        RECT 21.014 59.955 21.068 59.991 ;
        RECT 21.65 59.955 21.704 59.991 ;
        RECT 16.964 60.2545 17.036 60.2795 ;
        RECT 17.844 60.2545 17.916 60.2795 ;
        RECT 18.664 60.2545 18.736 60.2795 ;
        RECT 18.964 60.2545 19.036 60.2795 ;
        RECT 14.05 60.249 14.104 60.285 ;
        RECT 14.932 60.249 14.986 60.285 ;
        RECT 15.318 60.249 15.37 60.285 ;
        RECT 15.478 60.249 15.53 60.285 ;
        RECT 15.874 60.249 15.926 60.285 ;
        RECT 16.034 60.249 16.086 60.285 ;
        RECT 16.8 60.249 16.854 60.285 ;
        RECT 18.148 60.249 18.188 60.285 ;
        RECT 18.356 60.249 18.396 60.285 ;
        RECT 19.914 60.249 19.966 60.285 ;
        RECT 20.074 60.249 20.126 60.285 ;
        RECT 20.47 60.249 20.522 60.285 ;
        RECT 20.63 60.249 20.682 60.285 ;
        RECT 21.014 60.249 21.068 60.285 ;
        RECT 21.896 60.249 21.95 60.285 ;
        RECT 16.964 60.4835 17.036 60.5085 ;
        RECT 18.664 60.4835 18.736 60.5085 ;
        RECT 18.964 60.4835 19.036 60.5085 ;
        RECT 14.05 60.478 14.104 60.514 ;
        RECT 14.296 60.478 14.35 60.514 ;
        RECT 14.932 60.478 14.986 60.514 ;
        RECT 15.318 60.478 15.37 60.514 ;
        RECT 15.478 60.478 15.53 60.514 ;
        RECT 15.874 60.478 15.926 60.514 ;
        RECT 16.034 60.478 16.086 60.514 ;
        RECT 16.8 60.478 16.854 60.514 ;
        RECT 18.148 60.478 18.188 60.514 ;
        RECT 19.914 60.478 19.966 60.514 ;
        RECT 20.074 60.478 20.126 60.514 ;
        RECT 20.47 60.478 20.522 60.514 ;
        RECT 20.63 60.478 20.682 60.514 ;
        RECT 21.014 60.478 21.068 60.514 ;
        RECT 21.65 60.478 21.704 60.514 ;
        RECT 21.896 60.478 21.95 60.514 ;
        RECT 17.844 60.5605 17.916 60.5855 ;
        RECT 18.356 60.555 18.396 60.591 ;
        RECT 16.964 60.9315 17.036 60.9565 ;
        RECT 17.844 60.9315 17.916 60.9565 ;
        RECT 18.964 60.9315 19.036 60.9565 ;
        RECT 14.05 60.926 14.104 60.962 ;
        RECT 14.296 60.926 14.35 60.962 ;
        RECT 14.932 60.926 14.986 60.962 ;
        RECT 15.318 60.926 15.37 60.962 ;
        RECT 15.874 60.926 15.926 60.962 ;
        RECT 16.034 60.926 16.086 60.962 ;
        RECT 18.356 60.926 18.396 60.962 ;
        RECT 19.914 60.926 19.966 60.962 ;
        RECT 20.074 60.926 20.126 60.962 ;
        RECT 20.63 60.926 20.682 60.962 ;
        RECT 21.014 60.926 21.068 60.962 ;
        RECT 21.65 60.926 21.704 60.962 ;
        RECT 21.896 60.926 21.95 60.962 ;
        RECT 17.844 61.0835 17.916 61.1085 ;
        RECT 18.356 61.078 18.396 61.114 ;
        RECT 18.664 61.1605 18.736 61.1855 ;
        RECT 18.964 61.1605 19.036 61.1855 ;
        RECT 14.296 61.155 14.35 61.191 ;
        RECT 14.932 61.155 14.986 61.191 ;
        RECT 15.318 61.155 15.37 61.191 ;
        RECT 15.478 61.155 15.53 61.191 ;
        RECT 15.874 61.155 15.926 61.191 ;
        RECT 18.148 61.155 18.188 61.191 ;
        RECT 20.074 61.155 20.126 61.191 ;
        RECT 20.47 61.155 20.522 61.191 ;
        RECT 20.63 61.155 20.682 61.191 ;
        RECT 21.014 61.155 21.068 61.191 ;
        RECT 21.65 61.155 21.704 61.191 ;
        RECT 16.964 61.4545 17.036 61.4795 ;
        RECT 17.844 61.4545 17.916 61.4795 ;
        RECT 18.664 61.4545 18.736 61.4795 ;
        RECT 18.964 61.4545 19.036 61.4795 ;
        RECT 14.05 61.449 14.104 61.485 ;
        RECT 14.932 61.449 14.986 61.485 ;
        RECT 15.318 61.449 15.37 61.485 ;
        RECT 15.478 61.449 15.53 61.485 ;
        RECT 15.874 61.449 15.926 61.485 ;
        RECT 16.034 61.449 16.086 61.485 ;
        RECT 16.8 61.449 16.854 61.485 ;
        RECT 18.148 61.449 18.188 61.485 ;
        RECT 18.356 61.449 18.396 61.485 ;
        RECT 19.914 61.449 19.966 61.485 ;
        RECT 20.074 61.449 20.126 61.485 ;
        RECT 20.47 61.449 20.522 61.485 ;
        RECT 20.63 61.449 20.682 61.485 ;
        RECT 21.014 61.449 21.068 61.485 ;
        RECT 21.896 61.449 21.95 61.485 ;
        RECT 16.964 61.6835 17.036 61.7085 ;
        RECT 18.664 61.6835 18.736 61.7085 ;
        RECT 18.964 61.6835 19.036 61.7085 ;
        RECT 14.05 61.678 14.104 61.714 ;
        RECT 14.296 61.678 14.35 61.714 ;
        RECT 14.932 61.678 14.986 61.714 ;
        RECT 15.318 61.678 15.37 61.714 ;
        RECT 15.478 61.678 15.53 61.714 ;
        RECT 15.874 61.678 15.926 61.714 ;
        RECT 16.034 61.678 16.086 61.714 ;
        RECT 16.8 61.678 16.854 61.714 ;
        RECT 18.148 61.678 18.188 61.714 ;
        RECT 19.914 61.678 19.966 61.714 ;
        RECT 20.074 61.678 20.126 61.714 ;
        RECT 20.47 61.678 20.522 61.714 ;
        RECT 20.63 61.678 20.682 61.714 ;
        RECT 21.014 61.678 21.068 61.714 ;
        RECT 21.65 61.678 21.704 61.714 ;
        RECT 21.896 61.678 21.95 61.714 ;
        RECT 17.844 61.7605 17.916 61.7855 ;
        RECT 18.356 61.755 18.396 61.791 ;
        RECT 16.964 62.1315 17.036 62.1565 ;
        RECT 17.844 62.1315 17.916 62.1565 ;
        RECT 18.964 62.1315 19.036 62.1565 ;
        RECT 14.05 62.126 14.104 62.162 ;
        RECT 14.296 62.126 14.35 62.162 ;
        RECT 14.932 62.126 14.986 62.162 ;
        RECT 15.318 62.126 15.37 62.162 ;
        RECT 15.874 62.126 15.926 62.162 ;
        RECT 16.034 62.126 16.086 62.162 ;
        RECT 18.356 62.126 18.396 62.162 ;
        RECT 19.914 62.126 19.966 62.162 ;
        RECT 20.074 62.126 20.126 62.162 ;
        RECT 20.63 62.126 20.682 62.162 ;
        RECT 21.014 62.126 21.068 62.162 ;
        RECT 21.65 62.126 21.704 62.162 ;
        RECT 21.896 62.126 21.95 62.162 ;
        RECT 17.844 62.2835 17.916 62.3085 ;
        RECT 18.356 62.278 18.396 62.314 ;
        RECT 18.664 62.3605 18.736 62.3855 ;
        RECT 18.964 62.3605 19.036 62.3855 ;
        RECT 14.296 62.355 14.35 62.391 ;
        RECT 14.932 62.355 14.986 62.391 ;
        RECT 15.318 62.355 15.37 62.391 ;
        RECT 15.478 62.355 15.53 62.391 ;
        RECT 15.874 62.355 15.926 62.391 ;
        RECT 18.148 62.355 18.188 62.391 ;
        RECT 20.074 62.355 20.126 62.391 ;
        RECT 20.47 62.355 20.522 62.391 ;
        RECT 20.63 62.355 20.682 62.391 ;
        RECT 21.014 62.355 21.068 62.391 ;
        RECT 21.65 62.355 21.704 62.391 ;
        RECT 16.964 62.6545 17.036 62.6795 ;
        RECT 17.844 62.6545 17.916 62.6795 ;
        RECT 18.664 62.6545 18.736 62.6795 ;
        RECT 18.964 62.6545 19.036 62.6795 ;
        RECT 14.05 62.649 14.104 62.685 ;
        RECT 14.932 62.649 14.986 62.685 ;
        RECT 15.318 62.649 15.37 62.685 ;
        RECT 15.478 62.649 15.53 62.685 ;
        RECT 15.874 62.649 15.926 62.685 ;
        RECT 16.034 62.649 16.086 62.685 ;
        RECT 16.8 62.649 16.854 62.685 ;
        RECT 18.148 62.649 18.188 62.685 ;
        RECT 18.356 62.649 18.396 62.685 ;
        RECT 19.914 62.649 19.966 62.685 ;
        RECT 20.074 62.649 20.126 62.685 ;
        RECT 20.47 62.649 20.522 62.685 ;
        RECT 20.63 62.649 20.682 62.685 ;
        RECT 21.014 62.649 21.068 62.685 ;
        RECT 21.896 62.649 21.95 62.685 ;
        RECT 16.964 62.8835 17.036 62.9085 ;
        RECT 18.664 62.8835 18.736 62.9085 ;
        RECT 18.964 62.8835 19.036 62.9085 ;
        RECT 14.05 62.878 14.104 62.914 ;
        RECT 14.296 62.878 14.35 62.914 ;
        RECT 14.932 62.878 14.986 62.914 ;
        RECT 15.318 62.878 15.37 62.914 ;
        RECT 15.478 62.878 15.53 62.914 ;
        RECT 15.874 62.878 15.926 62.914 ;
        RECT 16.034 62.878 16.086 62.914 ;
        RECT 16.8 62.878 16.854 62.914 ;
        RECT 18.148 62.878 18.188 62.914 ;
        RECT 19.914 62.878 19.966 62.914 ;
        RECT 20.074 62.878 20.126 62.914 ;
        RECT 20.47 62.878 20.522 62.914 ;
        RECT 20.63 62.878 20.682 62.914 ;
        RECT 21.014 62.878 21.068 62.914 ;
        RECT 21.65 62.878 21.704 62.914 ;
        RECT 21.896 62.878 21.95 62.914 ;
        RECT 17.844 62.9605 17.916 62.9855 ;
        RECT 18.356 62.955 18.396 62.991 ;
        RECT 16.964 63.3315 17.036 63.3565 ;
        RECT 17.844 63.3315 17.916 63.3565 ;
        RECT 18.964 63.3315 19.036 63.3565 ;
        RECT 14.05 63.326 14.104 63.362 ;
        RECT 14.296 63.326 14.35 63.362 ;
        RECT 14.932 63.326 14.986 63.362 ;
        RECT 15.318 63.326 15.37 63.362 ;
        RECT 15.874 63.326 15.926 63.362 ;
        RECT 16.034 63.326 16.086 63.362 ;
        RECT 18.356 63.326 18.396 63.362 ;
        RECT 19.914 63.326 19.966 63.362 ;
        RECT 20.074 63.326 20.126 63.362 ;
        RECT 20.63 63.326 20.682 63.362 ;
        RECT 21.014 63.326 21.068 63.362 ;
        RECT 21.65 63.326 21.704 63.362 ;
        RECT 21.896 63.326 21.95 63.362 ;
        RECT 17.844 63.4835 17.916 63.5085 ;
        RECT 18.356 63.478 18.396 63.514 ;
        RECT 18.664 63.5605 18.736 63.5855 ;
        RECT 18.964 63.5605 19.036 63.5855 ;
        RECT 14.296 63.555 14.35 63.591 ;
        RECT 14.932 63.555 14.986 63.591 ;
        RECT 15.318 63.555 15.37 63.591 ;
        RECT 15.478 63.555 15.53 63.591 ;
        RECT 15.874 63.555 15.926 63.591 ;
        RECT 18.148 63.555 18.188 63.591 ;
        RECT 20.074 63.555 20.126 63.591 ;
        RECT 20.47 63.555 20.522 63.591 ;
        RECT 20.63 63.555 20.682 63.591 ;
        RECT 21.014 63.555 21.068 63.591 ;
        RECT 21.65 63.555 21.704 63.591 ;
        RECT 16.964 63.8545 17.036 63.8795 ;
        RECT 17.844 63.8545 17.916 63.8795 ;
        RECT 18.664 63.8545 18.736 63.8795 ;
        RECT 18.964 63.8545 19.036 63.8795 ;
        RECT 14.05 63.849 14.104 63.885 ;
        RECT 14.932 63.849 14.986 63.885 ;
        RECT 15.318 63.849 15.37 63.885 ;
        RECT 15.478 63.849 15.53 63.885 ;
        RECT 15.874 63.849 15.926 63.885 ;
        RECT 16.034 63.849 16.086 63.885 ;
        RECT 16.8 63.849 16.854 63.885 ;
        RECT 18.148 63.849 18.188 63.885 ;
        RECT 18.356 63.849 18.396 63.885 ;
        RECT 19.914 63.849 19.966 63.885 ;
        RECT 20.074 63.849 20.126 63.885 ;
        RECT 20.47 63.849 20.522 63.885 ;
        RECT 20.63 63.849 20.682 63.885 ;
        RECT 21.014 63.849 21.068 63.885 ;
        RECT 21.896 63.849 21.95 63.885 ;
        RECT 16.964 64.0835 17.036 64.1085 ;
        RECT 18.664 64.0835 18.736 64.1085 ;
        RECT 18.964 64.0835 19.036 64.1085 ;
        RECT 14.05 64.078 14.104 64.114 ;
        RECT 14.296 64.078 14.35 64.114 ;
        RECT 14.932 64.078 14.986 64.114 ;
        RECT 15.318 64.078 15.37 64.114 ;
        RECT 15.478 64.078 15.53 64.114 ;
        RECT 15.874 64.078 15.926 64.114 ;
        RECT 16.034 64.078 16.086 64.114 ;
        RECT 16.8 64.078 16.854 64.114 ;
        RECT 18.148 64.078 18.188 64.114 ;
        RECT 19.914 64.078 19.966 64.114 ;
        RECT 20.074 64.078 20.126 64.114 ;
        RECT 20.47 64.078 20.522 64.114 ;
        RECT 20.63 64.078 20.682 64.114 ;
        RECT 21.014 64.078 21.068 64.114 ;
        RECT 21.65 64.078 21.704 64.114 ;
        RECT 21.896 64.078 21.95 64.114 ;
        RECT 17.844 64.1605 17.916 64.1855 ;
        RECT 18.356 64.155 18.396 64.191 ;
        RECT 16.964 64.5315 17.036 64.5565 ;
        RECT 17.844 64.5315 17.916 64.5565 ;
        RECT 18.964 64.5315 19.036 64.5565 ;
        RECT 14.05 64.526 14.104 64.562 ;
        RECT 14.296 64.526 14.35 64.562 ;
        RECT 14.932 64.526 14.986 64.562 ;
        RECT 15.318 64.526 15.37 64.562 ;
        RECT 15.874 64.526 15.926 64.562 ;
        RECT 16.034 64.526 16.086 64.562 ;
        RECT 18.356 64.526 18.396 64.562 ;
        RECT 19.914 64.526 19.966 64.562 ;
        RECT 20.074 64.526 20.126 64.562 ;
        RECT 20.63 64.526 20.682 64.562 ;
        RECT 21.014 64.526 21.068 64.562 ;
        RECT 21.65 64.526 21.704 64.562 ;
        RECT 21.896 64.526 21.95 64.562 ;
        RECT 17.844 64.6835 17.916 64.7085 ;
        RECT 18.356 64.678 18.396 64.714 ;
        RECT 18.664 64.7605 18.736 64.7855 ;
        RECT 18.964 64.7605 19.036 64.7855 ;
        RECT 14.296 64.755 14.35 64.791 ;
        RECT 14.932 64.755 14.986 64.791 ;
        RECT 15.318 64.755 15.37 64.791 ;
        RECT 15.478 64.755 15.53 64.791 ;
        RECT 15.874 64.755 15.926 64.791 ;
        RECT 18.148 64.755 18.188 64.791 ;
        RECT 20.074 64.755 20.126 64.791 ;
        RECT 20.47 64.755 20.522 64.791 ;
        RECT 20.63 64.755 20.682 64.791 ;
        RECT 21.014 64.755 21.068 64.791 ;
        RECT 21.65 64.755 21.704 64.791 ;
        RECT 16.964 65.0545 17.036 65.0795 ;
        RECT 17.844 65.0545 17.916 65.0795 ;
        RECT 18.664 65.0545 18.736 65.0795 ;
        RECT 18.964 65.0545 19.036 65.0795 ;
        RECT 14.05 65.049 14.104 65.085 ;
        RECT 14.932 65.049 14.986 65.085 ;
        RECT 15.318 65.049 15.37 65.085 ;
        RECT 15.478 65.049 15.53 65.085 ;
        RECT 15.874 65.049 15.926 65.085 ;
        RECT 16.034 65.049 16.086 65.085 ;
        RECT 16.8 65.049 16.854 65.085 ;
        RECT 18.148 65.049 18.188 65.085 ;
        RECT 18.356 65.049 18.396 65.085 ;
        RECT 19.914 65.049 19.966 65.085 ;
        RECT 20.074 65.049 20.126 65.085 ;
        RECT 20.47 65.049 20.522 65.085 ;
        RECT 20.63 65.049 20.682 65.085 ;
        RECT 21.014 65.049 21.068 65.085 ;
        RECT 21.896 65.049 21.95 65.085 ;
        RECT 16.964 65.2835 17.036 65.3085 ;
        RECT 18.664 65.2835 18.736 65.3085 ;
        RECT 18.964 65.2835 19.036 65.3085 ;
        RECT 14.05 65.278 14.104 65.314 ;
        RECT 14.296 65.278 14.35 65.314 ;
        RECT 14.932 65.278 14.986 65.314 ;
        RECT 15.318 65.278 15.37 65.314 ;
        RECT 15.478 65.278 15.53 65.314 ;
        RECT 15.874 65.278 15.926 65.314 ;
        RECT 16.034 65.278 16.086 65.314 ;
        RECT 16.8 65.278 16.854 65.314 ;
        RECT 18.148 65.278 18.188 65.314 ;
        RECT 19.914 65.278 19.966 65.314 ;
        RECT 20.074 65.278 20.126 65.314 ;
        RECT 20.47 65.278 20.522 65.314 ;
        RECT 20.63 65.278 20.682 65.314 ;
        RECT 21.014 65.278 21.068 65.314 ;
        RECT 21.65 65.278 21.704 65.314 ;
        RECT 21.896 65.278 21.95 65.314 ;
        RECT 17.844 65.3605 17.916 65.3855 ;
        RECT 18.356 65.355 18.396 65.391 ;
        RECT 16.964 65.7315 17.036 65.7565 ;
        RECT 17.844 65.7315 17.916 65.7565 ;
        RECT 18.964 65.7315 19.036 65.7565 ;
        RECT 14.05 65.726 14.104 65.762 ;
        RECT 14.296 65.726 14.35 65.762 ;
        RECT 14.932 65.726 14.986 65.762 ;
        RECT 15.318 65.726 15.37 65.762 ;
        RECT 15.874 65.726 15.926 65.762 ;
        RECT 16.034 65.726 16.086 65.762 ;
        RECT 18.356 65.726 18.396 65.762 ;
        RECT 19.914 65.726 19.966 65.762 ;
        RECT 20.074 65.726 20.126 65.762 ;
        RECT 20.63 65.726 20.682 65.762 ;
        RECT 21.014 65.726 21.068 65.762 ;
        RECT 21.65 65.726 21.704 65.762 ;
        RECT 21.896 65.726 21.95 65.762 ;
        RECT 17.844 65.8835 17.916 65.9085 ;
        RECT 18.356 65.878 18.396 65.914 ;
        RECT 18.664 65.9605 18.736 65.9855 ;
        RECT 18.964 65.9605 19.036 65.9855 ;
        RECT 14.296 65.955 14.35 65.991 ;
        RECT 14.932 65.955 14.986 65.991 ;
        RECT 15.318 65.955 15.37 65.991 ;
        RECT 15.478 65.955 15.53 65.991 ;
        RECT 15.874 65.955 15.926 65.991 ;
        RECT 18.148 65.955 18.188 65.991 ;
        RECT 20.074 65.955 20.126 65.991 ;
        RECT 20.47 65.955 20.522 65.991 ;
        RECT 20.63 65.955 20.682 65.991 ;
        RECT 21.014 65.955 21.068 65.991 ;
        RECT 21.65 65.955 21.704 65.991 ;
        RECT 16.964 66.2545 17.036 66.2795 ;
        RECT 17.844 66.2545 17.916 66.2795 ;
        RECT 18.664 66.2545 18.736 66.2795 ;
        RECT 18.964 66.2545 19.036 66.2795 ;
        RECT 14.05 66.249 14.104 66.285 ;
        RECT 14.932 66.249 14.986 66.285 ;
        RECT 15.318 66.249 15.37 66.285 ;
        RECT 15.478 66.249 15.53 66.285 ;
        RECT 15.874 66.249 15.926 66.285 ;
        RECT 16.034 66.249 16.086 66.285 ;
        RECT 16.8 66.249 16.854 66.285 ;
        RECT 18.148 66.249 18.188 66.285 ;
        RECT 18.356 66.249 18.396 66.285 ;
        RECT 19.914 66.249 19.966 66.285 ;
        RECT 20.074 66.249 20.126 66.285 ;
        RECT 20.47 66.249 20.522 66.285 ;
        RECT 20.63 66.249 20.682 66.285 ;
        RECT 21.014 66.249 21.068 66.285 ;
        RECT 21.896 66.249 21.95 66.285 ;
        RECT 16.964 66.4835 17.036 66.5085 ;
        RECT 18.664 66.4835 18.736 66.5085 ;
        RECT 18.964 66.4835 19.036 66.5085 ;
        RECT 14.05 66.478 14.104 66.514 ;
        RECT 14.296 66.478 14.35 66.514 ;
        RECT 14.932 66.478 14.986 66.514 ;
        RECT 15.318 66.478 15.37 66.514 ;
        RECT 15.478 66.478 15.53 66.514 ;
        RECT 15.874 66.478 15.926 66.514 ;
        RECT 16.034 66.478 16.086 66.514 ;
        RECT 16.8 66.478 16.854 66.514 ;
        RECT 18.148 66.478 18.188 66.514 ;
        RECT 19.914 66.478 19.966 66.514 ;
        RECT 20.074 66.478 20.126 66.514 ;
        RECT 20.47 66.478 20.522 66.514 ;
        RECT 20.63 66.478 20.682 66.514 ;
        RECT 21.014 66.478 21.068 66.514 ;
        RECT 21.65 66.478 21.704 66.514 ;
        RECT 21.896 66.478 21.95 66.514 ;
        RECT 17.844 66.5605 17.916 66.5855 ;
        RECT 18.356 66.555 18.396 66.591 ;
        RECT 16.964 66.9315 17.036 66.9565 ;
        RECT 17.844 66.9315 17.916 66.9565 ;
        RECT 18.964 66.9315 19.036 66.9565 ;
        RECT 14.05 66.926 14.104 66.962 ;
        RECT 14.296 66.926 14.35 66.962 ;
        RECT 14.932 66.926 14.986 66.962 ;
        RECT 15.318 66.926 15.37 66.962 ;
        RECT 15.874 66.926 15.926 66.962 ;
        RECT 16.034 66.926 16.086 66.962 ;
        RECT 18.356 66.926 18.396 66.962 ;
        RECT 19.914 66.926 19.966 66.962 ;
        RECT 20.074 66.926 20.126 66.962 ;
        RECT 20.63 66.926 20.682 66.962 ;
        RECT 21.014 66.926 21.068 66.962 ;
        RECT 21.65 66.926 21.704 66.962 ;
        RECT 21.896 66.926 21.95 66.962 ;
        RECT 17.844 67.0835 17.916 67.1085 ;
        RECT 18.356 67.078 18.396 67.114 ;
        RECT 18.664 67.1605 18.736 67.1855 ;
        RECT 18.964 67.1605 19.036 67.1855 ;
        RECT 14.296 67.155 14.35 67.191 ;
        RECT 14.932 67.155 14.986 67.191 ;
        RECT 15.318 67.155 15.37 67.191 ;
        RECT 15.478 67.155 15.53 67.191 ;
        RECT 15.874 67.155 15.926 67.191 ;
        RECT 18.148 67.155 18.188 67.191 ;
        RECT 20.074 67.155 20.126 67.191 ;
        RECT 20.47 67.155 20.522 67.191 ;
        RECT 20.63 67.155 20.682 67.191 ;
        RECT 21.014 67.155 21.068 67.191 ;
        RECT 21.65 67.155 21.704 67.191 ;
        RECT 16.964 67.4545 17.036 67.4795 ;
        RECT 17.844 67.4545 17.916 67.4795 ;
        RECT 18.664 67.4545 18.736 67.4795 ;
        RECT 18.964 67.4545 19.036 67.4795 ;
        RECT 14.05 67.449 14.104 67.485 ;
        RECT 14.932 67.449 14.986 67.485 ;
        RECT 15.318 67.449 15.37 67.485 ;
        RECT 15.478 67.449 15.53 67.485 ;
        RECT 15.874 67.449 15.926 67.485 ;
        RECT 16.034 67.449 16.086 67.485 ;
        RECT 16.8 67.449 16.854 67.485 ;
        RECT 18.148 67.449 18.188 67.485 ;
        RECT 18.356 67.449 18.396 67.485 ;
        RECT 19.914 67.449 19.966 67.485 ;
        RECT 20.074 67.449 20.126 67.485 ;
        RECT 20.47 67.449 20.522 67.485 ;
        RECT 20.63 67.449 20.682 67.485 ;
        RECT 21.014 67.449 21.068 67.485 ;
        RECT 21.896 67.449 21.95 67.485 ;
        RECT 16.964 67.6835 17.036 67.7085 ;
        RECT 18.664 67.6835 18.736 67.7085 ;
        RECT 18.964 67.6835 19.036 67.7085 ;
        RECT 14.05 67.678 14.104 67.714 ;
        RECT 14.296 67.678 14.35 67.714 ;
        RECT 14.932 67.678 14.986 67.714 ;
        RECT 15.318 67.678 15.37 67.714 ;
        RECT 15.478 67.678 15.53 67.714 ;
        RECT 15.874 67.678 15.926 67.714 ;
        RECT 16.034 67.678 16.086 67.714 ;
        RECT 16.8 67.678 16.854 67.714 ;
        RECT 18.148 67.678 18.188 67.714 ;
        RECT 19.914 67.678 19.966 67.714 ;
        RECT 20.074 67.678 20.126 67.714 ;
        RECT 20.47 67.678 20.522 67.714 ;
        RECT 20.63 67.678 20.682 67.714 ;
        RECT 21.014 67.678 21.068 67.714 ;
        RECT 21.65 67.678 21.704 67.714 ;
        RECT 21.896 67.678 21.95 67.714 ;
        RECT 17.844 67.7605 17.916 67.7855 ;
        RECT 18.356 67.755 18.396 67.791 ;
        RECT 16.964 68.1315 17.036 68.1565 ;
        RECT 17.844 68.1315 17.916 68.1565 ;
        RECT 18.964 68.1315 19.036 68.1565 ;
        RECT 14.05 68.126 14.104 68.162 ;
        RECT 14.296 68.126 14.35 68.162 ;
        RECT 14.932 68.126 14.986 68.162 ;
        RECT 15.318 68.126 15.37 68.162 ;
        RECT 15.874 68.126 15.926 68.162 ;
        RECT 16.034 68.126 16.086 68.162 ;
        RECT 18.356 68.126 18.396 68.162 ;
        RECT 19.914 68.126 19.966 68.162 ;
        RECT 20.074 68.126 20.126 68.162 ;
        RECT 20.63 68.126 20.682 68.162 ;
        RECT 21.014 68.126 21.068 68.162 ;
        RECT 21.65 68.126 21.704 68.162 ;
        RECT 21.896 68.126 21.95 68.162 ;
        RECT 17.844 68.2835 17.916 68.3085 ;
        RECT 18.356 68.278 18.396 68.314 ;
        RECT 18.664 68.3605 18.736 68.3855 ;
        RECT 18.964 68.3605 19.036 68.3855 ;
        RECT 14.296 68.355 14.35 68.391 ;
        RECT 14.932 68.355 14.986 68.391 ;
        RECT 15.318 68.355 15.37 68.391 ;
        RECT 15.478 68.355 15.53 68.391 ;
        RECT 15.874 68.355 15.926 68.391 ;
        RECT 18.148 68.355 18.188 68.391 ;
        RECT 20.074 68.355 20.126 68.391 ;
        RECT 20.47 68.355 20.522 68.391 ;
        RECT 20.63 68.355 20.682 68.391 ;
        RECT 21.014 68.355 21.068 68.391 ;
        RECT 21.65 68.355 21.704 68.391 ;
        RECT 16.964 68.6545 17.036 68.6795 ;
        RECT 17.844 68.6545 17.916 68.6795 ;
        RECT 18.664 68.6545 18.736 68.6795 ;
        RECT 18.964 68.6545 19.036 68.6795 ;
        RECT 14.05 68.649 14.104 68.685 ;
        RECT 14.932 68.649 14.986 68.685 ;
        RECT 15.318 68.649 15.37 68.685 ;
        RECT 15.478 68.649 15.53 68.685 ;
        RECT 15.874 68.649 15.926 68.685 ;
        RECT 16.034 68.649 16.086 68.685 ;
        RECT 16.8 68.649 16.854 68.685 ;
        RECT 18.148 68.649 18.188 68.685 ;
        RECT 18.356 68.649 18.396 68.685 ;
        RECT 19.914 68.649 19.966 68.685 ;
        RECT 20.074 68.649 20.126 68.685 ;
        RECT 20.47 68.649 20.522 68.685 ;
        RECT 20.63 68.649 20.682 68.685 ;
        RECT 21.014 68.649 21.068 68.685 ;
        RECT 21.896 68.649 21.95 68.685 ;
        RECT 16.964 68.8835 17.036 68.9085 ;
        RECT 18.664 68.8835 18.736 68.9085 ;
        RECT 18.964 68.8835 19.036 68.9085 ;
        RECT 14.05 68.878 14.104 68.914 ;
        RECT 14.296 68.878 14.35 68.914 ;
        RECT 14.932 68.878 14.986 68.914 ;
        RECT 15.318 68.878 15.37 68.914 ;
        RECT 15.478 68.878 15.53 68.914 ;
        RECT 15.874 68.878 15.926 68.914 ;
        RECT 16.034 68.878 16.086 68.914 ;
        RECT 16.8 68.878 16.854 68.914 ;
        RECT 18.148 68.878 18.188 68.914 ;
        RECT 19.914 68.878 19.966 68.914 ;
        RECT 20.074 68.878 20.126 68.914 ;
        RECT 20.47 68.878 20.522 68.914 ;
        RECT 20.63 68.878 20.682 68.914 ;
        RECT 21.014 68.878 21.068 68.914 ;
        RECT 21.65 68.878 21.704 68.914 ;
        RECT 21.896 68.878 21.95 68.914 ;
        RECT 17.844 68.9605 17.916 68.9855 ;
        RECT 18.356 68.955 18.396 68.991 ;
        RECT 16.964 69.3315 17.036 69.3565 ;
        RECT 17.844 69.3315 17.916 69.3565 ;
        RECT 18.964 69.3315 19.036 69.3565 ;
        RECT 14.05 69.326 14.104 69.362 ;
        RECT 14.296 69.326 14.35 69.362 ;
        RECT 14.932 69.326 14.986 69.362 ;
        RECT 15.318 69.326 15.37 69.362 ;
        RECT 15.874 69.326 15.926 69.362 ;
        RECT 16.034 69.326 16.086 69.362 ;
        RECT 18.356 69.326 18.396 69.362 ;
        RECT 19.914 69.326 19.966 69.362 ;
        RECT 20.074 69.326 20.126 69.362 ;
        RECT 20.63 69.326 20.682 69.362 ;
        RECT 21.014 69.326 21.068 69.362 ;
        RECT 21.65 69.326 21.704 69.362 ;
        RECT 21.896 69.326 21.95 69.362 ;
        RECT 17.844 69.4835 17.916 69.5085 ;
        RECT 18.356 69.478 18.396 69.514 ;
        RECT 18.664 69.5605 18.736 69.5855 ;
        RECT 18.964 69.5605 19.036 69.5855 ;
        RECT 14.296 69.555 14.35 69.591 ;
        RECT 14.932 69.555 14.986 69.591 ;
        RECT 15.318 69.555 15.37 69.591 ;
        RECT 15.478 69.555 15.53 69.591 ;
        RECT 15.874 69.555 15.926 69.591 ;
        RECT 18.148 69.555 18.188 69.591 ;
        RECT 20.074 69.555 20.126 69.591 ;
        RECT 20.47 69.555 20.522 69.591 ;
        RECT 20.63 69.555 20.682 69.591 ;
        RECT 21.014 69.555 21.068 69.591 ;
        RECT 21.65 69.555 21.704 69.591 ;
        RECT 16.964 69.8545 17.036 69.8795 ;
        RECT 17.844 69.8545 17.916 69.8795 ;
        RECT 18.664 69.8545 18.736 69.8795 ;
        RECT 18.964 69.8545 19.036 69.8795 ;
        RECT 14.05 69.849 14.104 69.885 ;
        RECT 14.932 69.849 14.986 69.885 ;
        RECT 15.318 69.849 15.37 69.885 ;
        RECT 15.478 69.849 15.53 69.885 ;
        RECT 15.874 69.849 15.926 69.885 ;
        RECT 16.034 69.849 16.086 69.885 ;
        RECT 16.8 69.849 16.854 69.885 ;
        RECT 18.148 69.849 18.188 69.885 ;
        RECT 18.356 69.849 18.396 69.885 ;
        RECT 19.914 69.849 19.966 69.885 ;
        RECT 20.074 69.849 20.126 69.885 ;
        RECT 20.47 69.849 20.522 69.885 ;
        RECT 20.63 69.849 20.682 69.885 ;
        RECT 21.014 69.849 21.068 69.885 ;
        RECT 21.896 69.849 21.95 69.885 ;
        RECT 16.964 70.0835 17.036 70.1085 ;
        RECT 18.664 70.0835 18.736 70.1085 ;
        RECT 18.964 70.0835 19.036 70.1085 ;
        RECT 14.05 70.078 14.104 70.114 ;
        RECT 14.296 70.078 14.35 70.114 ;
        RECT 14.932 70.078 14.986 70.114 ;
        RECT 15.318 70.078 15.37 70.114 ;
        RECT 15.478 70.078 15.53 70.114 ;
        RECT 15.874 70.078 15.926 70.114 ;
        RECT 16.034 70.078 16.086 70.114 ;
        RECT 16.8 70.078 16.854 70.114 ;
        RECT 18.148 70.078 18.188 70.114 ;
        RECT 19.914 70.078 19.966 70.114 ;
        RECT 20.074 70.078 20.126 70.114 ;
        RECT 20.47 70.078 20.522 70.114 ;
        RECT 20.63 70.078 20.682 70.114 ;
        RECT 21.014 70.078 21.068 70.114 ;
        RECT 21.65 70.078 21.704 70.114 ;
        RECT 21.896 70.078 21.95 70.114 ;
        RECT 17.844 70.1605 17.916 70.1855 ;
        RECT 18.356 70.155 18.396 70.191 ;
        RECT 16.964 70.5315 17.036 70.5565 ;
        RECT 17.844 70.5315 17.916 70.5565 ;
        RECT 18.964 70.5315 19.036 70.5565 ;
        RECT 14.05 70.526 14.104 70.562 ;
        RECT 14.296 70.526 14.35 70.562 ;
        RECT 14.932 70.526 14.986 70.562 ;
        RECT 15.318 70.526 15.37 70.562 ;
        RECT 15.874 70.526 15.926 70.562 ;
        RECT 16.034 70.526 16.086 70.562 ;
        RECT 18.356 70.526 18.396 70.562 ;
        RECT 19.914 70.526 19.966 70.562 ;
        RECT 20.074 70.526 20.126 70.562 ;
        RECT 20.63 70.526 20.682 70.562 ;
        RECT 21.014 70.526 21.068 70.562 ;
        RECT 21.65 70.526 21.704 70.562 ;
        RECT 21.896 70.526 21.95 70.562 ;
        RECT 17.844 70.6835 17.916 70.7085 ;
        RECT 18.356 70.678 18.396 70.714 ;
        RECT 18.664 70.7605 18.736 70.7855 ;
        RECT 18.964 70.7605 19.036 70.7855 ;
        RECT 14.296 70.755 14.35 70.791 ;
        RECT 14.932 70.755 14.986 70.791 ;
        RECT 15.318 70.755 15.37 70.791 ;
        RECT 15.478 70.755 15.53 70.791 ;
        RECT 15.874 70.755 15.926 70.791 ;
        RECT 18.148 70.755 18.188 70.791 ;
        RECT 20.074 70.755 20.126 70.791 ;
        RECT 20.47 70.755 20.522 70.791 ;
        RECT 20.63 70.755 20.682 70.791 ;
        RECT 21.014 70.755 21.068 70.791 ;
        RECT 21.65 70.755 21.704 70.791 ;
        RECT 16.964 71.0545 17.036 71.0795 ;
        RECT 17.844 71.0545 17.916 71.0795 ;
        RECT 18.664 71.0545 18.736 71.0795 ;
        RECT 18.964 71.0545 19.036 71.0795 ;
        RECT 14.05 71.049 14.104 71.085 ;
        RECT 14.932 71.049 14.986 71.085 ;
        RECT 15.318 71.049 15.37 71.085 ;
        RECT 15.478 71.049 15.53 71.085 ;
        RECT 15.874 71.049 15.926 71.085 ;
        RECT 16.034 71.049 16.086 71.085 ;
        RECT 16.8 71.049 16.854 71.085 ;
        RECT 18.148 71.049 18.188 71.085 ;
        RECT 18.356 71.049 18.396 71.085 ;
        RECT 19.914 71.049 19.966 71.085 ;
        RECT 20.074 71.049 20.126 71.085 ;
        RECT 20.47 71.049 20.522 71.085 ;
        RECT 20.63 71.049 20.682 71.085 ;
        RECT 21.014 71.049 21.068 71.085 ;
        RECT 21.896 71.049 21.95 71.085 ;
        RECT 16.964 71.2835 17.036 71.3085 ;
        RECT 18.664 71.2835 18.736 71.3085 ;
        RECT 18.964 71.2835 19.036 71.3085 ;
        RECT 14.05 71.278 14.104 71.314 ;
        RECT 14.296 71.278 14.35 71.314 ;
        RECT 14.932 71.278 14.986 71.314 ;
        RECT 15.318 71.278 15.37 71.314 ;
        RECT 15.478 71.278 15.53 71.314 ;
        RECT 15.874 71.278 15.926 71.314 ;
        RECT 16.034 71.278 16.086 71.314 ;
        RECT 16.8 71.278 16.854 71.314 ;
        RECT 18.148 71.278 18.188 71.314 ;
        RECT 19.914 71.278 19.966 71.314 ;
        RECT 20.074 71.278 20.126 71.314 ;
        RECT 20.47 71.278 20.522 71.314 ;
        RECT 20.63 71.278 20.682 71.314 ;
        RECT 21.014 71.278 21.068 71.314 ;
        RECT 21.65 71.278 21.704 71.314 ;
        RECT 21.896 71.278 21.95 71.314 ;
        RECT 17.844 71.3605 17.916 71.3855 ;
        RECT 18.356 71.355 18.396 71.391 ;
        RECT 16.964 71.7315 17.036 71.7565 ;
        RECT 17.844 71.7315 17.916 71.7565 ;
        RECT 18.964 71.7315 19.036 71.7565 ;
        RECT 14.05 71.726 14.104 71.762 ;
        RECT 14.296 71.726 14.35 71.762 ;
        RECT 14.932 71.726 14.986 71.762 ;
        RECT 15.318 71.726 15.37 71.762 ;
        RECT 15.874 71.726 15.926 71.762 ;
        RECT 16.034 71.726 16.086 71.762 ;
        RECT 18.356 71.726 18.396 71.762 ;
        RECT 19.914 71.726 19.966 71.762 ;
        RECT 20.074 71.726 20.126 71.762 ;
        RECT 20.63 71.726 20.682 71.762 ;
        RECT 21.014 71.726 21.068 71.762 ;
        RECT 21.65 71.726 21.704 71.762 ;
        RECT 21.896 71.726 21.95 71.762 ;
        RECT 17.844 71.8835 17.916 71.9085 ;
        RECT 18.356 71.878 18.396 71.914 ;
        RECT 18.664 71.9605 18.736 71.9855 ;
        RECT 18.964 71.9605 19.036 71.9855 ;
        RECT 14.296 71.955 14.35 71.991 ;
        RECT 14.932 71.955 14.986 71.991 ;
        RECT 15.318 71.955 15.37 71.991 ;
        RECT 15.478 71.955 15.53 71.991 ;
        RECT 15.874 71.955 15.926 71.991 ;
        RECT 18.148 71.955 18.188 71.991 ;
        RECT 20.074 71.955 20.126 71.991 ;
        RECT 20.47 71.955 20.522 71.991 ;
        RECT 20.63 71.955 20.682 71.991 ;
        RECT 21.014 71.955 21.068 71.991 ;
        RECT 21.65 71.955 21.704 71.991 ;
      LAYER m5 ;
        RECT 15.478 0.5695 15.53 32.8595 ;
        RECT 20.47 0.5695 20.522 32.8595 ;
        RECT 0.654 32.9505 0.706 38.5695 ;
        RECT 1.454 32.9505 1.506 38.5695 ;
        RECT 2.254 32.9505 2.306 38.5695 ;
        RECT 3.054 32.9505 3.106 38.5695 ;
        RECT 3.854 32.9505 3.906 38.5695 ;
        RECT 4.654 32.9505 4.706 38.5695 ;
        RECT 5.454 32.9505 5.506 38.5695 ;
        RECT 6.254 32.9505 6.306 38.5695 ;
        RECT 7.054 32.9505 7.106 38.5695 ;
        RECT 7.854 32.9505 7.906 38.5695 ;
        RECT 8.654 32.9505 8.706 38.5695 ;
        RECT 9.454 32.9505 9.506 38.5695 ;
        RECT 10.254 32.9505 10.306 38.5695 ;
        RECT 11.054 32.9505 11.106 38.5695 ;
        RECT 11.854 32.9505 11.906 38.5695 ;
        RECT 12.654 32.9505 12.706 38.5695 ;
        RECT 22.854 32.9505 22.906 38.5695 ;
        RECT 23.654 32.9505 23.706 38.5695 ;
        RECT 24.454 32.9505 24.506 38.5695 ;
        RECT 25.254 32.9505 25.306 38.5695 ;
        RECT 26.054 32.9505 26.106 38.5695 ;
        RECT 26.854 32.9505 26.906 38.5695 ;
        RECT 27.654 32.9505 27.706 38.5695 ;
        RECT 28.454 32.9505 28.506 38.5695 ;
        RECT 29.254 32.9505 29.306 38.5695 ;
        RECT 30.054 32.9505 30.106 38.5695 ;
        RECT 30.854 32.9505 30.906 38.5695 ;
        RECT 31.654 32.9505 31.706 38.5695 ;
        RECT 32.454 32.9505 32.506 38.5695 ;
        RECT 33.254 32.9505 33.306 38.5695 ;
        RECT 34.054 32.9505 34.106 38.5695 ;
        RECT 34.854 32.9505 34.906 38.5695 ;
        RECT 17.412 32.18 17.452 39.34 ;
        RECT 19.31 31.8 19.35 39.72 ;
        RECT 0.974 0.6 1.026 72.12 ;
        RECT 1.774 0.6 1.826 72.12 ;
        RECT 2.574 0.6 2.626 72.12 ;
        RECT 3.374 0.6 3.426 72.12 ;
        RECT 4.174 0.6 4.226 72.12 ;
        RECT 4.974 0.6 5.026 72.12 ;
        RECT 5.774 0.6 5.826 72.12 ;
        RECT 6.574 0.6 6.626 72.12 ;
        RECT 7.374 0.6 7.426 72.12 ;
        RECT 8.174 0.6 8.226 72.12 ;
        RECT 8.974 0.6 9.026 72.12 ;
        RECT 9.774 0.6 9.826 72.12 ;
        RECT 10.574 0.6 10.626 72.12 ;
        RECT 11.374 0.6 11.426 72.12 ;
        RECT 12.174 0.6 12.226 72.12 ;
        RECT 12.974 0.6 13.026 72.12 ;
        RECT 15.874 0.6 15.926 72.12 ;
        RECT 20.074 0.6 20.126 72.12 ;
        RECT 23.174 0.6 23.226 72.12 ;
        RECT 23.974 0.6 24.026 72.12 ;
        RECT 24.774 0.6 24.826 72.12 ;
        RECT 25.574 0.6 25.626 72.12 ;
        RECT 26.374 0.6 26.426 72.12 ;
        RECT 27.174 0.6 27.226 72.12 ;
        RECT 27.974 0.6 28.026 72.12 ;
        RECT 28.774 0.6 28.826 72.12 ;
        RECT 29.574 0.6 29.626 72.12 ;
        RECT 30.374 0.6 30.426 72.12 ;
        RECT 31.174 0.6 31.226 72.12 ;
        RECT 31.974 0.6 32.026 72.12 ;
        RECT 32.774 0.6 32.826 72.12 ;
        RECT 33.574 0.6 33.626 72.12 ;
        RECT 34.374 0.6 34.426 72.12 ;
        RECT 35.174 0.6 35.226 72.12 ;
        RECT 14.05 0.5695 14.104 72.1505 ;
        RECT 14.296 0.5695 14.35 72.1505 ;
        RECT 14.932 0.5695 14.986 72.1505 ;
        RECT 15.318 0.5695 15.37 72.1505 ;
        RECT 15.478 38.199 15.53 72.1505 ;
        RECT 16.034 0.5695 16.086 72.1505 ;
        RECT 16.8 0.5695 16.854 72.1505 ;
        RECT 16.964 0.5695 17.036 72.1505 ;
        RECT 17.844 0.5695 17.916 72.1505 ;
        RECT 18.148 0.5695 18.188 72.1505 ;
        RECT 18.356 0.5695 18.396 72.1505 ;
        RECT 18.664 0.5695 18.736 72.1505 ;
        RECT 18.964 0.5695 19.036 72.1505 ;
        RECT 19.914 0.5695 19.966 72.1505 ;
        RECT 20.47 38.199 20.522 72.1505 ;
        RECT 20.63 0.5695 20.682 72.1505 ;
        RECT 21.014 0.5695 21.068 72.1505 ;
        RECT 21.65 0.5695 21.704 72.1505 ;
        RECT 21.896 0.5695 21.95 72.1505 ;
    END
  END vddp
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER v4 ;
        RECT 18.564 0.5875 18.636 0.6125 ;
        RECT 18.864 0.5875 18.936 0.6125 ;
        RECT 0.574 0.582 0.626 0.618 ;
        RECT 1.374 0.582 1.426 0.618 ;
        RECT 2.174 0.582 2.226 0.618 ;
        RECT 2.974 0.582 3.026 0.618 ;
        RECT 3.774 0.582 3.826 0.618 ;
        RECT 4.574 0.582 4.626 0.618 ;
        RECT 5.374 0.582 5.426 0.618 ;
        RECT 6.174 0.582 6.226 0.618 ;
        RECT 6.974 0.582 7.026 0.618 ;
        RECT 7.774 0.582 7.826 0.618 ;
        RECT 8.574 0.582 8.626 0.618 ;
        RECT 9.374 0.582 9.426 0.618 ;
        RECT 10.174 0.582 10.226 0.618 ;
        RECT 10.974 0.582 11.026 0.618 ;
        RECT 11.774 0.582 11.826 0.618 ;
        RECT 12.574 0.582 12.626 0.618 ;
        RECT 13.374 0.582 13.426 0.618 ;
        RECT 14.45 0.582 14.504 0.618 ;
        RECT 15.658 0.582 15.71 0.618 ;
        RECT 15.954 0.582 16.006 0.618 ;
        RECT 16.266 0.582 16.318 0.618 ;
        RECT 16.498 0.582 16.55 0.618 ;
        RECT 17.344 0.582 17.384 0.618 ;
        RECT 17.684 0.582 17.736 0.618 ;
        RECT 19.45 0.582 19.502 0.618 ;
        RECT 19.682 0.582 19.734 0.618 ;
        RECT 19.994 0.582 20.046 0.618 ;
        RECT 20.29 0.582 20.342 0.618 ;
        RECT 21.496 0.582 21.55 0.618 ;
        RECT 22.774 0.582 22.826 0.618 ;
        RECT 23.574 0.582 23.626 0.618 ;
        RECT 24.374 0.582 24.426 0.618 ;
        RECT 25.174 0.582 25.226 0.618 ;
        RECT 25.974 0.582 26.026 0.618 ;
        RECT 26.774 0.582 26.826 0.618 ;
        RECT 27.574 0.582 27.626 0.618 ;
        RECT 28.374 0.582 28.426 0.618 ;
        RECT 29.174 0.582 29.226 0.618 ;
        RECT 29.974 0.582 30.026 0.618 ;
        RECT 30.774 0.582 30.826 0.618 ;
        RECT 31.574 0.582 31.626 0.618 ;
        RECT 32.374 0.582 32.426 0.618 ;
        RECT 33.174 0.582 33.226 0.618 ;
        RECT 33.974 0.582 34.026 0.618 ;
        RECT 34.774 0.582 34.826 0.618 ;
        RECT 35.574 0.582 35.626 0.618 ;
        RECT 18.564 1.1875 18.636 1.2125 ;
        RECT 18.864 1.1875 18.936 1.2125 ;
        RECT 0.574 1.182 0.626 1.218 ;
        RECT 1.374 1.182 1.426 1.218 ;
        RECT 2.174 1.182 2.226 1.218 ;
        RECT 2.974 1.182 3.026 1.218 ;
        RECT 3.774 1.182 3.826 1.218 ;
        RECT 4.574 1.182 4.626 1.218 ;
        RECT 5.374 1.182 5.426 1.218 ;
        RECT 6.174 1.182 6.226 1.218 ;
        RECT 6.974 1.182 7.026 1.218 ;
        RECT 7.774 1.182 7.826 1.218 ;
        RECT 8.574 1.182 8.626 1.218 ;
        RECT 9.374 1.182 9.426 1.218 ;
        RECT 10.174 1.182 10.226 1.218 ;
        RECT 10.974 1.182 11.026 1.218 ;
        RECT 11.774 1.182 11.826 1.218 ;
        RECT 12.574 1.182 12.626 1.218 ;
        RECT 13.374 1.182 13.426 1.218 ;
        RECT 14.45 1.182 14.504 1.218 ;
        RECT 15.658 1.182 15.71 1.218 ;
        RECT 15.954 1.182 16.006 1.218 ;
        RECT 16.266 1.182 16.318 1.218 ;
        RECT 16.498 1.182 16.55 1.218 ;
        RECT 17.344 1.182 17.384 1.218 ;
        RECT 17.684 1.182 17.736 1.218 ;
        RECT 19.45 1.182 19.502 1.218 ;
        RECT 19.682 1.182 19.734 1.218 ;
        RECT 19.994 1.182 20.046 1.218 ;
        RECT 20.29 1.182 20.342 1.218 ;
        RECT 21.496 1.182 21.55 1.218 ;
        RECT 22.774 1.182 22.826 1.218 ;
        RECT 23.574 1.182 23.626 1.218 ;
        RECT 24.374 1.182 24.426 1.218 ;
        RECT 25.174 1.182 25.226 1.218 ;
        RECT 25.974 1.182 26.026 1.218 ;
        RECT 26.774 1.182 26.826 1.218 ;
        RECT 27.574 1.182 27.626 1.218 ;
        RECT 28.374 1.182 28.426 1.218 ;
        RECT 29.174 1.182 29.226 1.218 ;
        RECT 29.974 1.182 30.026 1.218 ;
        RECT 30.774 1.182 30.826 1.218 ;
        RECT 31.574 1.182 31.626 1.218 ;
        RECT 32.374 1.182 32.426 1.218 ;
        RECT 33.174 1.182 33.226 1.218 ;
        RECT 33.974 1.182 34.026 1.218 ;
        RECT 34.774 1.182 34.826 1.218 ;
        RECT 35.574 1.182 35.626 1.218 ;
        RECT 18.564 1.7875 18.636 1.8125 ;
        RECT 18.864 1.7875 18.936 1.8125 ;
        RECT 0.574 1.782 0.626 1.818 ;
        RECT 1.374 1.782 1.426 1.818 ;
        RECT 2.174 1.782 2.226 1.818 ;
        RECT 2.974 1.782 3.026 1.818 ;
        RECT 3.774 1.782 3.826 1.818 ;
        RECT 4.574 1.782 4.626 1.818 ;
        RECT 5.374 1.782 5.426 1.818 ;
        RECT 6.174 1.782 6.226 1.818 ;
        RECT 6.974 1.782 7.026 1.818 ;
        RECT 7.774 1.782 7.826 1.818 ;
        RECT 8.574 1.782 8.626 1.818 ;
        RECT 9.374 1.782 9.426 1.818 ;
        RECT 10.174 1.782 10.226 1.818 ;
        RECT 10.974 1.782 11.026 1.818 ;
        RECT 11.774 1.782 11.826 1.818 ;
        RECT 12.574 1.782 12.626 1.818 ;
        RECT 13.374 1.782 13.426 1.818 ;
        RECT 14.45 1.782 14.504 1.818 ;
        RECT 15.658 1.782 15.71 1.818 ;
        RECT 15.954 1.782 16.006 1.818 ;
        RECT 16.266 1.782 16.318 1.818 ;
        RECT 16.498 1.782 16.55 1.818 ;
        RECT 17.344 1.782 17.384 1.818 ;
        RECT 17.684 1.782 17.736 1.818 ;
        RECT 19.45 1.782 19.502 1.818 ;
        RECT 19.682 1.782 19.734 1.818 ;
        RECT 19.994 1.782 20.046 1.818 ;
        RECT 20.29 1.782 20.342 1.818 ;
        RECT 21.496 1.782 21.55 1.818 ;
        RECT 22.774 1.782 22.826 1.818 ;
        RECT 23.574 1.782 23.626 1.818 ;
        RECT 24.374 1.782 24.426 1.818 ;
        RECT 25.174 1.782 25.226 1.818 ;
        RECT 25.974 1.782 26.026 1.818 ;
        RECT 26.774 1.782 26.826 1.818 ;
        RECT 27.574 1.782 27.626 1.818 ;
        RECT 28.374 1.782 28.426 1.818 ;
        RECT 29.174 1.782 29.226 1.818 ;
        RECT 29.974 1.782 30.026 1.818 ;
        RECT 30.774 1.782 30.826 1.818 ;
        RECT 31.574 1.782 31.626 1.818 ;
        RECT 32.374 1.782 32.426 1.818 ;
        RECT 33.174 1.782 33.226 1.818 ;
        RECT 33.974 1.782 34.026 1.818 ;
        RECT 34.774 1.782 34.826 1.818 ;
        RECT 35.574 1.782 35.626 1.818 ;
        RECT 18.564 2.3875 18.636 2.4125 ;
        RECT 18.864 2.3875 18.936 2.4125 ;
        RECT 0.574 2.382 0.626 2.418 ;
        RECT 1.374 2.382 1.426 2.418 ;
        RECT 2.174 2.382 2.226 2.418 ;
        RECT 2.974 2.382 3.026 2.418 ;
        RECT 3.774 2.382 3.826 2.418 ;
        RECT 4.574 2.382 4.626 2.418 ;
        RECT 5.374 2.382 5.426 2.418 ;
        RECT 6.174 2.382 6.226 2.418 ;
        RECT 6.974 2.382 7.026 2.418 ;
        RECT 7.774 2.382 7.826 2.418 ;
        RECT 8.574 2.382 8.626 2.418 ;
        RECT 9.374 2.382 9.426 2.418 ;
        RECT 10.174 2.382 10.226 2.418 ;
        RECT 10.974 2.382 11.026 2.418 ;
        RECT 11.774 2.382 11.826 2.418 ;
        RECT 12.574 2.382 12.626 2.418 ;
        RECT 13.374 2.382 13.426 2.418 ;
        RECT 14.45 2.382 14.504 2.418 ;
        RECT 15.658 2.382 15.71 2.418 ;
        RECT 15.954 2.382 16.006 2.418 ;
        RECT 16.266 2.382 16.318 2.418 ;
        RECT 16.498 2.382 16.55 2.418 ;
        RECT 17.344 2.382 17.384 2.418 ;
        RECT 17.684 2.382 17.736 2.418 ;
        RECT 19.45 2.382 19.502 2.418 ;
        RECT 19.682 2.382 19.734 2.418 ;
        RECT 19.994 2.382 20.046 2.418 ;
        RECT 20.29 2.382 20.342 2.418 ;
        RECT 21.496 2.382 21.55 2.418 ;
        RECT 22.774 2.382 22.826 2.418 ;
        RECT 23.574 2.382 23.626 2.418 ;
        RECT 24.374 2.382 24.426 2.418 ;
        RECT 25.174 2.382 25.226 2.418 ;
        RECT 25.974 2.382 26.026 2.418 ;
        RECT 26.774 2.382 26.826 2.418 ;
        RECT 27.574 2.382 27.626 2.418 ;
        RECT 28.374 2.382 28.426 2.418 ;
        RECT 29.174 2.382 29.226 2.418 ;
        RECT 29.974 2.382 30.026 2.418 ;
        RECT 30.774 2.382 30.826 2.418 ;
        RECT 31.574 2.382 31.626 2.418 ;
        RECT 32.374 2.382 32.426 2.418 ;
        RECT 33.174 2.382 33.226 2.418 ;
        RECT 33.974 2.382 34.026 2.418 ;
        RECT 34.774 2.382 34.826 2.418 ;
        RECT 35.574 2.382 35.626 2.418 ;
        RECT 18.564 2.9875 18.636 3.0125 ;
        RECT 18.864 2.9875 18.936 3.0125 ;
        RECT 0.574 2.982 0.626 3.018 ;
        RECT 1.374 2.982 1.426 3.018 ;
        RECT 2.174 2.982 2.226 3.018 ;
        RECT 2.974 2.982 3.026 3.018 ;
        RECT 3.774 2.982 3.826 3.018 ;
        RECT 4.574 2.982 4.626 3.018 ;
        RECT 5.374 2.982 5.426 3.018 ;
        RECT 6.174 2.982 6.226 3.018 ;
        RECT 6.974 2.982 7.026 3.018 ;
        RECT 7.774 2.982 7.826 3.018 ;
        RECT 8.574 2.982 8.626 3.018 ;
        RECT 9.374 2.982 9.426 3.018 ;
        RECT 10.174 2.982 10.226 3.018 ;
        RECT 10.974 2.982 11.026 3.018 ;
        RECT 11.774 2.982 11.826 3.018 ;
        RECT 12.574 2.982 12.626 3.018 ;
        RECT 13.374 2.982 13.426 3.018 ;
        RECT 14.45 2.982 14.504 3.018 ;
        RECT 15.658 2.982 15.71 3.018 ;
        RECT 15.954 2.982 16.006 3.018 ;
        RECT 16.266 2.982 16.318 3.018 ;
        RECT 16.498 2.982 16.55 3.018 ;
        RECT 17.344 2.982 17.384 3.018 ;
        RECT 17.684 2.982 17.736 3.018 ;
        RECT 19.45 2.982 19.502 3.018 ;
        RECT 19.682 2.982 19.734 3.018 ;
        RECT 19.994 2.982 20.046 3.018 ;
        RECT 20.29 2.982 20.342 3.018 ;
        RECT 21.496 2.982 21.55 3.018 ;
        RECT 22.774 2.982 22.826 3.018 ;
        RECT 23.574 2.982 23.626 3.018 ;
        RECT 24.374 2.982 24.426 3.018 ;
        RECT 25.174 2.982 25.226 3.018 ;
        RECT 25.974 2.982 26.026 3.018 ;
        RECT 26.774 2.982 26.826 3.018 ;
        RECT 27.574 2.982 27.626 3.018 ;
        RECT 28.374 2.982 28.426 3.018 ;
        RECT 29.174 2.982 29.226 3.018 ;
        RECT 29.974 2.982 30.026 3.018 ;
        RECT 30.774 2.982 30.826 3.018 ;
        RECT 31.574 2.982 31.626 3.018 ;
        RECT 32.374 2.982 32.426 3.018 ;
        RECT 33.174 2.982 33.226 3.018 ;
        RECT 33.974 2.982 34.026 3.018 ;
        RECT 34.774 2.982 34.826 3.018 ;
        RECT 35.574 2.982 35.626 3.018 ;
        RECT 18.564 3.5875 18.636 3.6125 ;
        RECT 18.864 3.5875 18.936 3.6125 ;
        RECT 0.574 3.582 0.626 3.618 ;
        RECT 1.374 3.582 1.426 3.618 ;
        RECT 2.174 3.582 2.226 3.618 ;
        RECT 2.974 3.582 3.026 3.618 ;
        RECT 3.774 3.582 3.826 3.618 ;
        RECT 4.574 3.582 4.626 3.618 ;
        RECT 5.374 3.582 5.426 3.618 ;
        RECT 6.174 3.582 6.226 3.618 ;
        RECT 6.974 3.582 7.026 3.618 ;
        RECT 7.774 3.582 7.826 3.618 ;
        RECT 8.574 3.582 8.626 3.618 ;
        RECT 9.374 3.582 9.426 3.618 ;
        RECT 10.174 3.582 10.226 3.618 ;
        RECT 10.974 3.582 11.026 3.618 ;
        RECT 11.774 3.582 11.826 3.618 ;
        RECT 12.574 3.582 12.626 3.618 ;
        RECT 13.374 3.582 13.426 3.618 ;
        RECT 14.45 3.582 14.504 3.618 ;
        RECT 15.658 3.582 15.71 3.618 ;
        RECT 15.954 3.582 16.006 3.618 ;
        RECT 16.266 3.582 16.318 3.618 ;
        RECT 16.498 3.582 16.55 3.618 ;
        RECT 17.344 3.582 17.384 3.618 ;
        RECT 17.684 3.582 17.736 3.618 ;
        RECT 19.45 3.582 19.502 3.618 ;
        RECT 19.682 3.582 19.734 3.618 ;
        RECT 19.994 3.582 20.046 3.618 ;
        RECT 20.29 3.582 20.342 3.618 ;
        RECT 21.496 3.582 21.55 3.618 ;
        RECT 22.774 3.582 22.826 3.618 ;
        RECT 23.574 3.582 23.626 3.618 ;
        RECT 24.374 3.582 24.426 3.618 ;
        RECT 25.174 3.582 25.226 3.618 ;
        RECT 25.974 3.582 26.026 3.618 ;
        RECT 26.774 3.582 26.826 3.618 ;
        RECT 27.574 3.582 27.626 3.618 ;
        RECT 28.374 3.582 28.426 3.618 ;
        RECT 29.174 3.582 29.226 3.618 ;
        RECT 29.974 3.582 30.026 3.618 ;
        RECT 30.774 3.582 30.826 3.618 ;
        RECT 31.574 3.582 31.626 3.618 ;
        RECT 32.374 3.582 32.426 3.618 ;
        RECT 33.174 3.582 33.226 3.618 ;
        RECT 33.974 3.582 34.026 3.618 ;
        RECT 34.774 3.582 34.826 3.618 ;
        RECT 35.574 3.582 35.626 3.618 ;
        RECT 18.564 4.1875 18.636 4.2125 ;
        RECT 18.864 4.1875 18.936 4.2125 ;
        RECT 0.574 4.182 0.626 4.218 ;
        RECT 1.374 4.182 1.426 4.218 ;
        RECT 2.174 4.182 2.226 4.218 ;
        RECT 2.974 4.182 3.026 4.218 ;
        RECT 3.774 4.182 3.826 4.218 ;
        RECT 4.574 4.182 4.626 4.218 ;
        RECT 5.374 4.182 5.426 4.218 ;
        RECT 6.174 4.182 6.226 4.218 ;
        RECT 6.974 4.182 7.026 4.218 ;
        RECT 7.774 4.182 7.826 4.218 ;
        RECT 8.574 4.182 8.626 4.218 ;
        RECT 9.374 4.182 9.426 4.218 ;
        RECT 10.174 4.182 10.226 4.218 ;
        RECT 10.974 4.182 11.026 4.218 ;
        RECT 11.774 4.182 11.826 4.218 ;
        RECT 12.574 4.182 12.626 4.218 ;
        RECT 13.374 4.182 13.426 4.218 ;
        RECT 14.45 4.182 14.504 4.218 ;
        RECT 15.658 4.182 15.71 4.218 ;
        RECT 15.954 4.182 16.006 4.218 ;
        RECT 16.266 4.182 16.318 4.218 ;
        RECT 16.498 4.182 16.55 4.218 ;
        RECT 17.344 4.182 17.384 4.218 ;
        RECT 17.684 4.182 17.736 4.218 ;
        RECT 19.45 4.182 19.502 4.218 ;
        RECT 19.682 4.182 19.734 4.218 ;
        RECT 19.994 4.182 20.046 4.218 ;
        RECT 20.29 4.182 20.342 4.218 ;
        RECT 21.496 4.182 21.55 4.218 ;
        RECT 22.774 4.182 22.826 4.218 ;
        RECT 23.574 4.182 23.626 4.218 ;
        RECT 24.374 4.182 24.426 4.218 ;
        RECT 25.174 4.182 25.226 4.218 ;
        RECT 25.974 4.182 26.026 4.218 ;
        RECT 26.774 4.182 26.826 4.218 ;
        RECT 27.574 4.182 27.626 4.218 ;
        RECT 28.374 4.182 28.426 4.218 ;
        RECT 29.174 4.182 29.226 4.218 ;
        RECT 29.974 4.182 30.026 4.218 ;
        RECT 30.774 4.182 30.826 4.218 ;
        RECT 31.574 4.182 31.626 4.218 ;
        RECT 32.374 4.182 32.426 4.218 ;
        RECT 33.174 4.182 33.226 4.218 ;
        RECT 33.974 4.182 34.026 4.218 ;
        RECT 34.774 4.182 34.826 4.218 ;
        RECT 35.574 4.182 35.626 4.218 ;
        RECT 18.564 4.7875 18.636 4.8125 ;
        RECT 18.864 4.7875 18.936 4.8125 ;
        RECT 0.574 4.782 0.626 4.818 ;
        RECT 1.374 4.782 1.426 4.818 ;
        RECT 2.174 4.782 2.226 4.818 ;
        RECT 2.974 4.782 3.026 4.818 ;
        RECT 3.774 4.782 3.826 4.818 ;
        RECT 4.574 4.782 4.626 4.818 ;
        RECT 5.374 4.782 5.426 4.818 ;
        RECT 6.174 4.782 6.226 4.818 ;
        RECT 6.974 4.782 7.026 4.818 ;
        RECT 7.774 4.782 7.826 4.818 ;
        RECT 8.574 4.782 8.626 4.818 ;
        RECT 9.374 4.782 9.426 4.818 ;
        RECT 10.174 4.782 10.226 4.818 ;
        RECT 10.974 4.782 11.026 4.818 ;
        RECT 11.774 4.782 11.826 4.818 ;
        RECT 12.574 4.782 12.626 4.818 ;
        RECT 13.374 4.782 13.426 4.818 ;
        RECT 14.45 4.782 14.504 4.818 ;
        RECT 15.658 4.782 15.71 4.818 ;
        RECT 15.954 4.782 16.006 4.818 ;
        RECT 16.266 4.782 16.318 4.818 ;
        RECT 16.498 4.782 16.55 4.818 ;
        RECT 17.344 4.782 17.384 4.818 ;
        RECT 17.684 4.782 17.736 4.818 ;
        RECT 19.45 4.782 19.502 4.818 ;
        RECT 19.682 4.782 19.734 4.818 ;
        RECT 19.994 4.782 20.046 4.818 ;
        RECT 20.29 4.782 20.342 4.818 ;
        RECT 21.496 4.782 21.55 4.818 ;
        RECT 22.774 4.782 22.826 4.818 ;
        RECT 23.574 4.782 23.626 4.818 ;
        RECT 24.374 4.782 24.426 4.818 ;
        RECT 25.174 4.782 25.226 4.818 ;
        RECT 25.974 4.782 26.026 4.818 ;
        RECT 26.774 4.782 26.826 4.818 ;
        RECT 27.574 4.782 27.626 4.818 ;
        RECT 28.374 4.782 28.426 4.818 ;
        RECT 29.174 4.782 29.226 4.818 ;
        RECT 29.974 4.782 30.026 4.818 ;
        RECT 30.774 4.782 30.826 4.818 ;
        RECT 31.574 4.782 31.626 4.818 ;
        RECT 32.374 4.782 32.426 4.818 ;
        RECT 33.174 4.782 33.226 4.818 ;
        RECT 33.974 4.782 34.026 4.818 ;
        RECT 34.774 4.782 34.826 4.818 ;
        RECT 35.574 4.782 35.626 4.818 ;
        RECT 18.564 5.3875 18.636 5.4125 ;
        RECT 18.864 5.3875 18.936 5.4125 ;
        RECT 0.574 5.382 0.626 5.418 ;
        RECT 1.374 5.382 1.426 5.418 ;
        RECT 2.174 5.382 2.226 5.418 ;
        RECT 2.974 5.382 3.026 5.418 ;
        RECT 3.774 5.382 3.826 5.418 ;
        RECT 4.574 5.382 4.626 5.418 ;
        RECT 5.374 5.382 5.426 5.418 ;
        RECT 6.174 5.382 6.226 5.418 ;
        RECT 6.974 5.382 7.026 5.418 ;
        RECT 7.774 5.382 7.826 5.418 ;
        RECT 8.574 5.382 8.626 5.418 ;
        RECT 9.374 5.382 9.426 5.418 ;
        RECT 10.174 5.382 10.226 5.418 ;
        RECT 10.974 5.382 11.026 5.418 ;
        RECT 11.774 5.382 11.826 5.418 ;
        RECT 12.574 5.382 12.626 5.418 ;
        RECT 13.374 5.382 13.426 5.418 ;
        RECT 14.45 5.382 14.504 5.418 ;
        RECT 15.658 5.382 15.71 5.418 ;
        RECT 15.954 5.382 16.006 5.418 ;
        RECT 16.266 5.382 16.318 5.418 ;
        RECT 16.498 5.382 16.55 5.418 ;
        RECT 17.344 5.382 17.384 5.418 ;
        RECT 17.684 5.382 17.736 5.418 ;
        RECT 19.45 5.382 19.502 5.418 ;
        RECT 19.682 5.382 19.734 5.418 ;
        RECT 19.994 5.382 20.046 5.418 ;
        RECT 20.29 5.382 20.342 5.418 ;
        RECT 21.496 5.382 21.55 5.418 ;
        RECT 22.774 5.382 22.826 5.418 ;
        RECT 23.574 5.382 23.626 5.418 ;
        RECT 24.374 5.382 24.426 5.418 ;
        RECT 25.174 5.382 25.226 5.418 ;
        RECT 25.974 5.382 26.026 5.418 ;
        RECT 26.774 5.382 26.826 5.418 ;
        RECT 27.574 5.382 27.626 5.418 ;
        RECT 28.374 5.382 28.426 5.418 ;
        RECT 29.174 5.382 29.226 5.418 ;
        RECT 29.974 5.382 30.026 5.418 ;
        RECT 30.774 5.382 30.826 5.418 ;
        RECT 31.574 5.382 31.626 5.418 ;
        RECT 32.374 5.382 32.426 5.418 ;
        RECT 33.174 5.382 33.226 5.418 ;
        RECT 33.974 5.382 34.026 5.418 ;
        RECT 34.774 5.382 34.826 5.418 ;
        RECT 35.574 5.382 35.626 5.418 ;
        RECT 18.564 5.9875 18.636 6.0125 ;
        RECT 18.864 5.9875 18.936 6.0125 ;
        RECT 0.574 5.982 0.626 6.018 ;
        RECT 1.374 5.982 1.426 6.018 ;
        RECT 2.174 5.982 2.226 6.018 ;
        RECT 2.974 5.982 3.026 6.018 ;
        RECT 3.774 5.982 3.826 6.018 ;
        RECT 4.574 5.982 4.626 6.018 ;
        RECT 5.374 5.982 5.426 6.018 ;
        RECT 6.174 5.982 6.226 6.018 ;
        RECT 6.974 5.982 7.026 6.018 ;
        RECT 7.774 5.982 7.826 6.018 ;
        RECT 8.574 5.982 8.626 6.018 ;
        RECT 9.374 5.982 9.426 6.018 ;
        RECT 10.174 5.982 10.226 6.018 ;
        RECT 10.974 5.982 11.026 6.018 ;
        RECT 11.774 5.982 11.826 6.018 ;
        RECT 12.574 5.982 12.626 6.018 ;
        RECT 13.374 5.982 13.426 6.018 ;
        RECT 14.45 5.982 14.504 6.018 ;
        RECT 15.658 5.982 15.71 6.018 ;
        RECT 15.954 5.982 16.006 6.018 ;
        RECT 16.266 5.982 16.318 6.018 ;
        RECT 16.498 5.982 16.55 6.018 ;
        RECT 17.344 5.982 17.384 6.018 ;
        RECT 17.684 5.982 17.736 6.018 ;
        RECT 19.45 5.982 19.502 6.018 ;
        RECT 19.682 5.982 19.734 6.018 ;
        RECT 19.994 5.982 20.046 6.018 ;
        RECT 20.29 5.982 20.342 6.018 ;
        RECT 21.496 5.982 21.55 6.018 ;
        RECT 22.774 5.982 22.826 6.018 ;
        RECT 23.574 5.982 23.626 6.018 ;
        RECT 24.374 5.982 24.426 6.018 ;
        RECT 25.174 5.982 25.226 6.018 ;
        RECT 25.974 5.982 26.026 6.018 ;
        RECT 26.774 5.982 26.826 6.018 ;
        RECT 27.574 5.982 27.626 6.018 ;
        RECT 28.374 5.982 28.426 6.018 ;
        RECT 29.174 5.982 29.226 6.018 ;
        RECT 29.974 5.982 30.026 6.018 ;
        RECT 30.774 5.982 30.826 6.018 ;
        RECT 31.574 5.982 31.626 6.018 ;
        RECT 32.374 5.982 32.426 6.018 ;
        RECT 33.174 5.982 33.226 6.018 ;
        RECT 33.974 5.982 34.026 6.018 ;
        RECT 34.774 5.982 34.826 6.018 ;
        RECT 35.574 5.982 35.626 6.018 ;
        RECT 18.564 6.5875 18.636 6.6125 ;
        RECT 18.864 6.5875 18.936 6.6125 ;
        RECT 0.574 6.582 0.626 6.618 ;
        RECT 1.374 6.582 1.426 6.618 ;
        RECT 2.174 6.582 2.226 6.618 ;
        RECT 2.974 6.582 3.026 6.618 ;
        RECT 3.774 6.582 3.826 6.618 ;
        RECT 4.574 6.582 4.626 6.618 ;
        RECT 5.374 6.582 5.426 6.618 ;
        RECT 6.174 6.582 6.226 6.618 ;
        RECT 6.974 6.582 7.026 6.618 ;
        RECT 7.774 6.582 7.826 6.618 ;
        RECT 8.574 6.582 8.626 6.618 ;
        RECT 9.374 6.582 9.426 6.618 ;
        RECT 10.174 6.582 10.226 6.618 ;
        RECT 10.974 6.582 11.026 6.618 ;
        RECT 11.774 6.582 11.826 6.618 ;
        RECT 12.574 6.582 12.626 6.618 ;
        RECT 13.374 6.582 13.426 6.618 ;
        RECT 14.45 6.582 14.504 6.618 ;
        RECT 15.658 6.582 15.71 6.618 ;
        RECT 15.954 6.582 16.006 6.618 ;
        RECT 16.266 6.582 16.318 6.618 ;
        RECT 16.498 6.582 16.55 6.618 ;
        RECT 17.344 6.582 17.384 6.618 ;
        RECT 17.684 6.582 17.736 6.618 ;
        RECT 19.45 6.582 19.502 6.618 ;
        RECT 19.682 6.582 19.734 6.618 ;
        RECT 19.994 6.582 20.046 6.618 ;
        RECT 20.29 6.582 20.342 6.618 ;
        RECT 21.496 6.582 21.55 6.618 ;
        RECT 22.774 6.582 22.826 6.618 ;
        RECT 23.574 6.582 23.626 6.618 ;
        RECT 24.374 6.582 24.426 6.618 ;
        RECT 25.174 6.582 25.226 6.618 ;
        RECT 25.974 6.582 26.026 6.618 ;
        RECT 26.774 6.582 26.826 6.618 ;
        RECT 27.574 6.582 27.626 6.618 ;
        RECT 28.374 6.582 28.426 6.618 ;
        RECT 29.174 6.582 29.226 6.618 ;
        RECT 29.974 6.582 30.026 6.618 ;
        RECT 30.774 6.582 30.826 6.618 ;
        RECT 31.574 6.582 31.626 6.618 ;
        RECT 32.374 6.582 32.426 6.618 ;
        RECT 33.174 6.582 33.226 6.618 ;
        RECT 33.974 6.582 34.026 6.618 ;
        RECT 34.774 6.582 34.826 6.618 ;
        RECT 35.574 6.582 35.626 6.618 ;
        RECT 18.564 7.1875 18.636 7.2125 ;
        RECT 18.864 7.1875 18.936 7.2125 ;
        RECT 0.574 7.182 0.626 7.218 ;
        RECT 1.374 7.182 1.426 7.218 ;
        RECT 2.174 7.182 2.226 7.218 ;
        RECT 2.974 7.182 3.026 7.218 ;
        RECT 3.774 7.182 3.826 7.218 ;
        RECT 4.574 7.182 4.626 7.218 ;
        RECT 5.374 7.182 5.426 7.218 ;
        RECT 6.174 7.182 6.226 7.218 ;
        RECT 6.974 7.182 7.026 7.218 ;
        RECT 7.774 7.182 7.826 7.218 ;
        RECT 8.574 7.182 8.626 7.218 ;
        RECT 9.374 7.182 9.426 7.218 ;
        RECT 10.174 7.182 10.226 7.218 ;
        RECT 10.974 7.182 11.026 7.218 ;
        RECT 11.774 7.182 11.826 7.218 ;
        RECT 12.574 7.182 12.626 7.218 ;
        RECT 13.374 7.182 13.426 7.218 ;
        RECT 14.45 7.182 14.504 7.218 ;
        RECT 15.658 7.182 15.71 7.218 ;
        RECT 15.954 7.182 16.006 7.218 ;
        RECT 16.266 7.182 16.318 7.218 ;
        RECT 16.498 7.182 16.55 7.218 ;
        RECT 17.344 7.182 17.384 7.218 ;
        RECT 17.684 7.182 17.736 7.218 ;
        RECT 19.45 7.182 19.502 7.218 ;
        RECT 19.682 7.182 19.734 7.218 ;
        RECT 19.994 7.182 20.046 7.218 ;
        RECT 20.29 7.182 20.342 7.218 ;
        RECT 21.496 7.182 21.55 7.218 ;
        RECT 22.774 7.182 22.826 7.218 ;
        RECT 23.574 7.182 23.626 7.218 ;
        RECT 24.374 7.182 24.426 7.218 ;
        RECT 25.174 7.182 25.226 7.218 ;
        RECT 25.974 7.182 26.026 7.218 ;
        RECT 26.774 7.182 26.826 7.218 ;
        RECT 27.574 7.182 27.626 7.218 ;
        RECT 28.374 7.182 28.426 7.218 ;
        RECT 29.174 7.182 29.226 7.218 ;
        RECT 29.974 7.182 30.026 7.218 ;
        RECT 30.774 7.182 30.826 7.218 ;
        RECT 31.574 7.182 31.626 7.218 ;
        RECT 32.374 7.182 32.426 7.218 ;
        RECT 33.174 7.182 33.226 7.218 ;
        RECT 33.974 7.182 34.026 7.218 ;
        RECT 34.774 7.182 34.826 7.218 ;
        RECT 35.574 7.182 35.626 7.218 ;
        RECT 18.564 7.7875 18.636 7.8125 ;
        RECT 18.864 7.7875 18.936 7.8125 ;
        RECT 0.574 7.782 0.626 7.818 ;
        RECT 1.374 7.782 1.426 7.818 ;
        RECT 2.174 7.782 2.226 7.818 ;
        RECT 2.974 7.782 3.026 7.818 ;
        RECT 3.774 7.782 3.826 7.818 ;
        RECT 4.574 7.782 4.626 7.818 ;
        RECT 5.374 7.782 5.426 7.818 ;
        RECT 6.174 7.782 6.226 7.818 ;
        RECT 6.974 7.782 7.026 7.818 ;
        RECT 7.774 7.782 7.826 7.818 ;
        RECT 8.574 7.782 8.626 7.818 ;
        RECT 9.374 7.782 9.426 7.818 ;
        RECT 10.174 7.782 10.226 7.818 ;
        RECT 10.974 7.782 11.026 7.818 ;
        RECT 11.774 7.782 11.826 7.818 ;
        RECT 12.574 7.782 12.626 7.818 ;
        RECT 13.374 7.782 13.426 7.818 ;
        RECT 14.45 7.782 14.504 7.818 ;
        RECT 15.658 7.782 15.71 7.818 ;
        RECT 15.954 7.782 16.006 7.818 ;
        RECT 16.266 7.782 16.318 7.818 ;
        RECT 16.498 7.782 16.55 7.818 ;
        RECT 17.344 7.782 17.384 7.818 ;
        RECT 17.684 7.782 17.736 7.818 ;
        RECT 19.45 7.782 19.502 7.818 ;
        RECT 19.682 7.782 19.734 7.818 ;
        RECT 19.994 7.782 20.046 7.818 ;
        RECT 20.29 7.782 20.342 7.818 ;
        RECT 21.496 7.782 21.55 7.818 ;
        RECT 22.774 7.782 22.826 7.818 ;
        RECT 23.574 7.782 23.626 7.818 ;
        RECT 24.374 7.782 24.426 7.818 ;
        RECT 25.174 7.782 25.226 7.818 ;
        RECT 25.974 7.782 26.026 7.818 ;
        RECT 26.774 7.782 26.826 7.818 ;
        RECT 27.574 7.782 27.626 7.818 ;
        RECT 28.374 7.782 28.426 7.818 ;
        RECT 29.174 7.782 29.226 7.818 ;
        RECT 29.974 7.782 30.026 7.818 ;
        RECT 30.774 7.782 30.826 7.818 ;
        RECT 31.574 7.782 31.626 7.818 ;
        RECT 32.374 7.782 32.426 7.818 ;
        RECT 33.174 7.782 33.226 7.818 ;
        RECT 33.974 7.782 34.026 7.818 ;
        RECT 34.774 7.782 34.826 7.818 ;
        RECT 35.574 7.782 35.626 7.818 ;
        RECT 18.564 8.3875 18.636 8.4125 ;
        RECT 18.864 8.3875 18.936 8.4125 ;
        RECT 0.574 8.382 0.626 8.418 ;
        RECT 1.374 8.382 1.426 8.418 ;
        RECT 2.174 8.382 2.226 8.418 ;
        RECT 2.974 8.382 3.026 8.418 ;
        RECT 3.774 8.382 3.826 8.418 ;
        RECT 4.574 8.382 4.626 8.418 ;
        RECT 5.374 8.382 5.426 8.418 ;
        RECT 6.174 8.382 6.226 8.418 ;
        RECT 6.974 8.382 7.026 8.418 ;
        RECT 7.774 8.382 7.826 8.418 ;
        RECT 8.574 8.382 8.626 8.418 ;
        RECT 9.374 8.382 9.426 8.418 ;
        RECT 10.174 8.382 10.226 8.418 ;
        RECT 10.974 8.382 11.026 8.418 ;
        RECT 11.774 8.382 11.826 8.418 ;
        RECT 12.574 8.382 12.626 8.418 ;
        RECT 13.374 8.382 13.426 8.418 ;
        RECT 14.45 8.382 14.504 8.418 ;
        RECT 15.658 8.382 15.71 8.418 ;
        RECT 15.954 8.382 16.006 8.418 ;
        RECT 16.266 8.382 16.318 8.418 ;
        RECT 16.498 8.382 16.55 8.418 ;
        RECT 17.344 8.382 17.384 8.418 ;
        RECT 17.684 8.382 17.736 8.418 ;
        RECT 19.45 8.382 19.502 8.418 ;
        RECT 19.682 8.382 19.734 8.418 ;
        RECT 19.994 8.382 20.046 8.418 ;
        RECT 20.29 8.382 20.342 8.418 ;
        RECT 21.496 8.382 21.55 8.418 ;
        RECT 22.774 8.382 22.826 8.418 ;
        RECT 23.574 8.382 23.626 8.418 ;
        RECT 24.374 8.382 24.426 8.418 ;
        RECT 25.174 8.382 25.226 8.418 ;
        RECT 25.974 8.382 26.026 8.418 ;
        RECT 26.774 8.382 26.826 8.418 ;
        RECT 27.574 8.382 27.626 8.418 ;
        RECT 28.374 8.382 28.426 8.418 ;
        RECT 29.174 8.382 29.226 8.418 ;
        RECT 29.974 8.382 30.026 8.418 ;
        RECT 30.774 8.382 30.826 8.418 ;
        RECT 31.574 8.382 31.626 8.418 ;
        RECT 32.374 8.382 32.426 8.418 ;
        RECT 33.174 8.382 33.226 8.418 ;
        RECT 33.974 8.382 34.026 8.418 ;
        RECT 34.774 8.382 34.826 8.418 ;
        RECT 35.574 8.382 35.626 8.418 ;
        RECT 18.564 8.9875 18.636 9.0125 ;
        RECT 18.864 8.9875 18.936 9.0125 ;
        RECT 0.574 8.982 0.626 9.018 ;
        RECT 1.374 8.982 1.426 9.018 ;
        RECT 2.174 8.982 2.226 9.018 ;
        RECT 2.974 8.982 3.026 9.018 ;
        RECT 3.774 8.982 3.826 9.018 ;
        RECT 4.574 8.982 4.626 9.018 ;
        RECT 5.374 8.982 5.426 9.018 ;
        RECT 6.174 8.982 6.226 9.018 ;
        RECT 6.974 8.982 7.026 9.018 ;
        RECT 7.774 8.982 7.826 9.018 ;
        RECT 8.574 8.982 8.626 9.018 ;
        RECT 9.374 8.982 9.426 9.018 ;
        RECT 10.174 8.982 10.226 9.018 ;
        RECT 10.974 8.982 11.026 9.018 ;
        RECT 11.774 8.982 11.826 9.018 ;
        RECT 12.574 8.982 12.626 9.018 ;
        RECT 13.374 8.982 13.426 9.018 ;
        RECT 14.45 8.982 14.504 9.018 ;
        RECT 15.658 8.982 15.71 9.018 ;
        RECT 15.954 8.982 16.006 9.018 ;
        RECT 16.266 8.982 16.318 9.018 ;
        RECT 16.498 8.982 16.55 9.018 ;
        RECT 17.344 8.982 17.384 9.018 ;
        RECT 17.684 8.982 17.736 9.018 ;
        RECT 19.45 8.982 19.502 9.018 ;
        RECT 19.682 8.982 19.734 9.018 ;
        RECT 19.994 8.982 20.046 9.018 ;
        RECT 20.29 8.982 20.342 9.018 ;
        RECT 21.496 8.982 21.55 9.018 ;
        RECT 22.774 8.982 22.826 9.018 ;
        RECT 23.574 8.982 23.626 9.018 ;
        RECT 24.374 8.982 24.426 9.018 ;
        RECT 25.174 8.982 25.226 9.018 ;
        RECT 25.974 8.982 26.026 9.018 ;
        RECT 26.774 8.982 26.826 9.018 ;
        RECT 27.574 8.982 27.626 9.018 ;
        RECT 28.374 8.982 28.426 9.018 ;
        RECT 29.174 8.982 29.226 9.018 ;
        RECT 29.974 8.982 30.026 9.018 ;
        RECT 30.774 8.982 30.826 9.018 ;
        RECT 31.574 8.982 31.626 9.018 ;
        RECT 32.374 8.982 32.426 9.018 ;
        RECT 33.174 8.982 33.226 9.018 ;
        RECT 33.974 8.982 34.026 9.018 ;
        RECT 34.774 8.982 34.826 9.018 ;
        RECT 35.574 8.982 35.626 9.018 ;
        RECT 18.564 9.5875 18.636 9.6125 ;
        RECT 18.864 9.5875 18.936 9.6125 ;
        RECT 0.574 9.582 0.626 9.618 ;
        RECT 1.374 9.582 1.426 9.618 ;
        RECT 2.174 9.582 2.226 9.618 ;
        RECT 2.974 9.582 3.026 9.618 ;
        RECT 3.774 9.582 3.826 9.618 ;
        RECT 4.574 9.582 4.626 9.618 ;
        RECT 5.374 9.582 5.426 9.618 ;
        RECT 6.174 9.582 6.226 9.618 ;
        RECT 6.974 9.582 7.026 9.618 ;
        RECT 7.774 9.582 7.826 9.618 ;
        RECT 8.574 9.582 8.626 9.618 ;
        RECT 9.374 9.582 9.426 9.618 ;
        RECT 10.174 9.582 10.226 9.618 ;
        RECT 10.974 9.582 11.026 9.618 ;
        RECT 11.774 9.582 11.826 9.618 ;
        RECT 12.574 9.582 12.626 9.618 ;
        RECT 13.374 9.582 13.426 9.618 ;
        RECT 14.45 9.582 14.504 9.618 ;
        RECT 15.658 9.582 15.71 9.618 ;
        RECT 15.954 9.582 16.006 9.618 ;
        RECT 16.266 9.582 16.318 9.618 ;
        RECT 16.498 9.582 16.55 9.618 ;
        RECT 17.344 9.582 17.384 9.618 ;
        RECT 17.684 9.582 17.736 9.618 ;
        RECT 19.45 9.582 19.502 9.618 ;
        RECT 19.682 9.582 19.734 9.618 ;
        RECT 19.994 9.582 20.046 9.618 ;
        RECT 20.29 9.582 20.342 9.618 ;
        RECT 21.496 9.582 21.55 9.618 ;
        RECT 22.774 9.582 22.826 9.618 ;
        RECT 23.574 9.582 23.626 9.618 ;
        RECT 24.374 9.582 24.426 9.618 ;
        RECT 25.174 9.582 25.226 9.618 ;
        RECT 25.974 9.582 26.026 9.618 ;
        RECT 26.774 9.582 26.826 9.618 ;
        RECT 27.574 9.582 27.626 9.618 ;
        RECT 28.374 9.582 28.426 9.618 ;
        RECT 29.174 9.582 29.226 9.618 ;
        RECT 29.974 9.582 30.026 9.618 ;
        RECT 30.774 9.582 30.826 9.618 ;
        RECT 31.574 9.582 31.626 9.618 ;
        RECT 32.374 9.582 32.426 9.618 ;
        RECT 33.174 9.582 33.226 9.618 ;
        RECT 33.974 9.582 34.026 9.618 ;
        RECT 34.774 9.582 34.826 9.618 ;
        RECT 35.574 9.582 35.626 9.618 ;
        RECT 18.564 10.1875 18.636 10.2125 ;
        RECT 18.864 10.1875 18.936 10.2125 ;
        RECT 0.574 10.182 0.626 10.218 ;
        RECT 1.374 10.182 1.426 10.218 ;
        RECT 2.174 10.182 2.226 10.218 ;
        RECT 2.974 10.182 3.026 10.218 ;
        RECT 3.774 10.182 3.826 10.218 ;
        RECT 4.574 10.182 4.626 10.218 ;
        RECT 5.374 10.182 5.426 10.218 ;
        RECT 6.174 10.182 6.226 10.218 ;
        RECT 6.974 10.182 7.026 10.218 ;
        RECT 7.774 10.182 7.826 10.218 ;
        RECT 8.574 10.182 8.626 10.218 ;
        RECT 9.374 10.182 9.426 10.218 ;
        RECT 10.174 10.182 10.226 10.218 ;
        RECT 10.974 10.182 11.026 10.218 ;
        RECT 11.774 10.182 11.826 10.218 ;
        RECT 12.574 10.182 12.626 10.218 ;
        RECT 13.374 10.182 13.426 10.218 ;
        RECT 14.45 10.182 14.504 10.218 ;
        RECT 15.658 10.182 15.71 10.218 ;
        RECT 15.954 10.182 16.006 10.218 ;
        RECT 16.266 10.182 16.318 10.218 ;
        RECT 16.498 10.182 16.55 10.218 ;
        RECT 17.344 10.182 17.384 10.218 ;
        RECT 17.684 10.182 17.736 10.218 ;
        RECT 19.45 10.182 19.502 10.218 ;
        RECT 19.682 10.182 19.734 10.218 ;
        RECT 19.994 10.182 20.046 10.218 ;
        RECT 20.29 10.182 20.342 10.218 ;
        RECT 21.496 10.182 21.55 10.218 ;
        RECT 22.774 10.182 22.826 10.218 ;
        RECT 23.574 10.182 23.626 10.218 ;
        RECT 24.374 10.182 24.426 10.218 ;
        RECT 25.174 10.182 25.226 10.218 ;
        RECT 25.974 10.182 26.026 10.218 ;
        RECT 26.774 10.182 26.826 10.218 ;
        RECT 27.574 10.182 27.626 10.218 ;
        RECT 28.374 10.182 28.426 10.218 ;
        RECT 29.174 10.182 29.226 10.218 ;
        RECT 29.974 10.182 30.026 10.218 ;
        RECT 30.774 10.182 30.826 10.218 ;
        RECT 31.574 10.182 31.626 10.218 ;
        RECT 32.374 10.182 32.426 10.218 ;
        RECT 33.174 10.182 33.226 10.218 ;
        RECT 33.974 10.182 34.026 10.218 ;
        RECT 34.774 10.182 34.826 10.218 ;
        RECT 35.574 10.182 35.626 10.218 ;
        RECT 18.564 10.7875 18.636 10.8125 ;
        RECT 18.864 10.7875 18.936 10.8125 ;
        RECT 0.574 10.782 0.626 10.818 ;
        RECT 1.374 10.782 1.426 10.818 ;
        RECT 2.174 10.782 2.226 10.818 ;
        RECT 2.974 10.782 3.026 10.818 ;
        RECT 3.774 10.782 3.826 10.818 ;
        RECT 4.574 10.782 4.626 10.818 ;
        RECT 5.374 10.782 5.426 10.818 ;
        RECT 6.174 10.782 6.226 10.818 ;
        RECT 6.974 10.782 7.026 10.818 ;
        RECT 7.774 10.782 7.826 10.818 ;
        RECT 8.574 10.782 8.626 10.818 ;
        RECT 9.374 10.782 9.426 10.818 ;
        RECT 10.174 10.782 10.226 10.818 ;
        RECT 10.974 10.782 11.026 10.818 ;
        RECT 11.774 10.782 11.826 10.818 ;
        RECT 12.574 10.782 12.626 10.818 ;
        RECT 13.374 10.782 13.426 10.818 ;
        RECT 14.45 10.782 14.504 10.818 ;
        RECT 15.658 10.782 15.71 10.818 ;
        RECT 15.954 10.782 16.006 10.818 ;
        RECT 16.266 10.782 16.318 10.818 ;
        RECT 16.498 10.782 16.55 10.818 ;
        RECT 17.344 10.782 17.384 10.818 ;
        RECT 17.684 10.782 17.736 10.818 ;
        RECT 19.45 10.782 19.502 10.818 ;
        RECT 19.682 10.782 19.734 10.818 ;
        RECT 19.994 10.782 20.046 10.818 ;
        RECT 20.29 10.782 20.342 10.818 ;
        RECT 21.496 10.782 21.55 10.818 ;
        RECT 22.774 10.782 22.826 10.818 ;
        RECT 23.574 10.782 23.626 10.818 ;
        RECT 24.374 10.782 24.426 10.818 ;
        RECT 25.174 10.782 25.226 10.818 ;
        RECT 25.974 10.782 26.026 10.818 ;
        RECT 26.774 10.782 26.826 10.818 ;
        RECT 27.574 10.782 27.626 10.818 ;
        RECT 28.374 10.782 28.426 10.818 ;
        RECT 29.174 10.782 29.226 10.818 ;
        RECT 29.974 10.782 30.026 10.818 ;
        RECT 30.774 10.782 30.826 10.818 ;
        RECT 31.574 10.782 31.626 10.818 ;
        RECT 32.374 10.782 32.426 10.818 ;
        RECT 33.174 10.782 33.226 10.818 ;
        RECT 33.974 10.782 34.026 10.818 ;
        RECT 34.774 10.782 34.826 10.818 ;
        RECT 35.574 10.782 35.626 10.818 ;
        RECT 18.564 11.3875 18.636 11.4125 ;
        RECT 18.864 11.3875 18.936 11.4125 ;
        RECT 0.574 11.382 0.626 11.418 ;
        RECT 1.374 11.382 1.426 11.418 ;
        RECT 2.174 11.382 2.226 11.418 ;
        RECT 2.974 11.382 3.026 11.418 ;
        RECT 3.774 11.382 3.826 11.418 ;
        RECT 4.574 11.382 4.626 11.418 ;
        RECT 5.374 11.382 5.426 11.418 ;
        RECT 6.174 11.382 6.226 11.418 ;
        RECT 6.974 11.382 7.026 11.418 ;
        RECT 7.774 11.382 7.826 11.418 ;
        RECT 8.574 11.382 8.626 11.418 ;
        RECT 9.374 11.382 9.426 11.418 ;
        RECT 10.174 11.382 10.226 11.418 ;
        RECT 10.974 11.382 11.026 11.418 ;
        RECT 11.774 11.382 11.826 11.418 ;
        RECT 12.574 11.382 12.626 11.418 ;
        RECT 13.374 11.382 13.426 11.418 ;
        RECT 14.45 11.382 14.504 11.418 ;
        RECT 15.658 11.382 15.71 11.418 ;
        RECT 15.954 11.382 16.006 11.418 ;
        RECT 16.266 11.382 16.318 11.418 ;
        RECT 16.498 11.382 16.55 11.418 ;
        RECT 17.344 11.382 17.384 11.418 ;
        RECT 17.684 11.382 17.736 11.418 ;
        RECT 19.45 11.382 19.502 11.418 ;
        RECT 19.682 11.382 19.734 11.418 ;
        RECT 19.994 11.382 20.046 11.418 ;
        RECT 20.29 11.382 20.342 11.418 ;
        RECT 21.496 11.382 21.55 11.418 ;
        RECT 22.774 11.382 22.826 11.418 ;
        RECT 23.574 11.382 23.626 11.418 ;
        RECT 24.374 11.382 24.426 11.418 ;
        RECT 25.174 11.382 25.226 11.418 ;
        RECT 25.974 11.382 26.026 11.418 ;
        RECT 26.774 11.382 26.826 11.418 ;
        RECT 27.574 11.382 27.626 11.418 ;
        RECT 28.374 11.382 28.426 11.418 ;
        RECT 29.174 11.382 29.226 11.418 ;
        RECT 29.974 11.382 30.026 11.418 ;
        RECT 30.774 11.382 30.826 11.418 ;
        RECT 31.574 11.382 31.626 11.418 ;
        RECT 32.374 11.382 32.426 11.418 ;
        RECT 33.174 11.382 33.226 11.418 ;
        RECT 33.974 11.382 34.026 11.418 ;
        RECT 34.774 11.382 34.826 11.418 ;
        RECT 35.574 11.382 35.626 11.418 ;
        RECT 18.564 11.9875 18.636 12.0125 ;
        RECT 18.864 11.9875 18.936 12.0125 ;
        RECT 0.574 11.982 0.626 12.018 ;
        RECT 1.374 11.982 1.426 12.018 ;
        RECT 2.174 11.982 2.226 12.018 ;
        RECT 2.974 11.982 3.026 12.018 ;
        RECT 3.774 11.982 3.826 12.018 ;
        RECT 4.574 11.982 4.626 12.018 ;
        RECT 5.374 11.982 5.426 12.018 ;
        RECT 6.174 11.982 6.226 12.018 ;
        RECT 6.974 11.982 7.026 12.018 ;
        RECT 7.774 11.982 7.826 12.018 ;
        RECT 8.574 11.982 8.626 12.018 ;
        RECT 9.374 11.982 9.426 12.018 ;
        RECT 10.174 11.982 10.226 12.018 ;
        RECT 10.974 11.982 11.026 12.018 ;
        RECT 11.774 11.982 11.826 12.018 ;
        RECT 12.574 11.982 12.626 12.018 ;
        RECT 13.374 11.982 13.426 12.018 ;
        RECT 14.45 11.982 14.504 12.018 ;
        RECT 15.658 11.982 15.71 12.018 ;
        RECT 15.954 11.982 16.006 12.018 ;
        RECT 16.266 11.982 16.318 12.018 ;
        RECT 16.498 11.982 16.55 12.018 ;
        RECT 17.344 11.982 17.384 12.018 ;
        RECT 17.684 11.982 17.736 12.018 ;
        RECT 19.45 11.982 19.502 12.018 ;
        RECT 19.682 11.982 19.734 12.018 ;
        RECT 19.994 11.982 20.046 12.018 ;
        RECT 20.29 11.982 20.342 12.018 ;
        RECT 21.496 11.982 21.55 12.018 ;
        RECT 22.774 11.982 22.826 12.018 ;
        RECT 23.574 11.982 23.626 12.018 ;
        RECT 24.374 11.982 24.426 12.018 ;
        RECT 25.174 11.982 25.226 12.018 ;
        RECT 25.974 11.982 26.026 12.018 ;
        RECT 26.774 11.982 26.826 12.018 ;
        RECT 27.574 11.982 27.626 12.018 ;
        RECT 28.374 11.982 28.426 12.018 ;
        RECT 29.174 11.982 29.226 12.018 ;
        RECT 29.974 11.982 30.026 12.018 ;
        RECT 30.774 11.982 30.826 12.018 ;
        RECT 31.574 11.982 31.626 12.018 ;
        RECT 32.374 11.982 32.426 12.018 ;
        RECT 33.174 11.982 33.226 12.018 ;
        RECT 33.974 11.982 34.026 12.018 ;
        RECT 34.774 11.982 34.826 12.018 ;
        RECT 35.574 11.982 35.626 12.018 ;
        RECT 18.564 12.5875 18.636 12.6125 ;
        RECT 18.864 12.5875 18.936 12.6125 ;
        RECT 0.574 12.582 0.626 12.618 ;
        RECT 1.374 12.582 1.426 12.618 ;
        RECT 2.174 12.582 2.226 12.618 ;
        RECT 2.974 12.582 3.026 12.618 ;
        RECT 3.774 12.582 3.826 12.618 ;
        RECT 4.574 12.582 4.626 12.618 ;
        RECT 5.374 12.582 5.426 12.618 ;
        RECT 6.174 12.582 6.226 12.618 ;
        RECT 6.974 12.582 7.026 12.618 ;
        RECT 7.774 12.582 7.826 12.618 ;
        RECT 8.574 12.582 8.626 12.618 ;
        RECT 9.374 12.582 9.426 12.618 ;
        RECT 10.174 12.582 10.226 12.618 ;
        RECT 10.974 12.582 11.026 12.618 ;
        RECT 11.774 12.582 11.826 12.618 ;
        RECT 12.574 12.582 12.626 12.618 ;
        RECT 13.374 12.582 13.426 12.618 ;
        RECT 14.45 12.582 14.504 12.618 ;
        RECT 15.658 12.582 15.71 12.618 ;
        RECT 15.954 12.582 16.006 12.618 ;
        RECT 16.266 12.582 16.318 12.618 ;
        RECT 16.498 12.582 16.55 12.618 ;
        RECT 17.344 12.582 17.384 12.618 ;
        RECT 17.684 12.582 17.736 12.618 ;
        RECT 19.45 12.582 19.502 12.618 ;
        RECT 19.682 12.582 19.734 12.618 ;
        RECT 19.994 12.582 20.046 12.618 ;
        RECT 20.29 12.582 20.342 12.618 ;
        RECT 21.496 12.582 21.55 12.618 ;
        RECT 22.774 12.582 22.826 12.618 ;
        RECT 23.574 12.582 23.626 12.618 ;
        RECT 24.374 12.582 24.426 12.618 ;
        RECT 25.174 12.582 25.226 12.618 ;
        RECT 25.974 12.582 26.026 12.618 ;
        RECT 26.774 12.582 26.826 12.618 ;
        RECT 27.574 12.582 27.626 12.618 ;
        RECT 28.374 12.582 28.426 12.618 ;
        RECT 29.174 12.582 29.226 12.618 ;
        RECT 29.974 12.582 30.026 12.618 ;
        RECT 30.774 12.582 30.826 12.618 ;
        RECT 31.574 12.582 31.626 12.618 ;
        RECT 32.374 12.582 32.426 12.618 ;
        RECT 33.174 12.582 33.226 12.618 ;
        RECT 33.974 12.582 34.026 12.618 ;
        RECT 34.774 12.582 34.826 12.618 ;
        RECT 35.574 12.582 35.626 12.618 ;
        RECT 18.564 13.1875 18.636 13.2125 ;
        RECT 18.864 13.1875 18.936 13.2125 ;
        RECT 0.574 13.182 0.626 13.218 ;
        RECT 1.374 13.182 1.426 13.218 ;
        RECT 2.174 13.182 2.226 13.218 ;
        RECT 2.974 13.182 3.026 13.218 ;
        RECT 3.774 13.182 3.826 13.218 ;
        RECT 4.574 13.182 4.626 13.218 ;
        RECT 5.374 13.182 5.426 13.218 ;
        RECT 6.174 13.182 6.226 13.218 ;
        RECT 6.974 13.182 7.026 13.218 ;
        RECT 7.774 13.182 7.826 13.218 ;
        RECT 8.574 13.182 8.626 13.218 ;
        RECT 9.374 13.182 9.426 13.218 ;
        RECT 10.174 13.182 10.226 13.218 ;
        RECT 10.974 13.182 11.026 13.218 ;
        RECT 11.774 13.182 11.826 13.218 ;
        RECT 12.574 13.182 12.626 13.218 ;
        RECT 13.374 13.182 13.426 13.218 ;
        RECT 14.45 13.182 14.504 13.218 ;
        RECT 15.658 13.182 15.71 13.218 ;
        RECT 15.954 13.182 16.006 13.218 ;
        RECT 16.266 13.182 16.318 13.218 ;
        RECT 16.498 13.182 16.55 13.218 ;
        RECT 17.344 13.182 17.384 13.218 ;
        RECT 17.684 13.182 17.736 13.218 ;
        RECT 19.45 13.182 19.502 13.218 ;
        RECT 19.682 13.182 19.734 13.218 ;
        RECT 19.994 13.182 20.046 13.218 ;
        RECT 20.29 13.182 20.342 13.218 ;
        RECT 21.496 13.182 21.55 13.218 ;
        RECT 22.774 13.182 22.826 13.218 ;
        RECT 23.574 13.182 23.626 13.218 ;
        RECT 24.374 13.182 24.426 13.218 ;
        RECT 25.174 13.182 25.226 13.218 ;
        RECT 25.974 13.182 26.026 13.218 ;
        RECT 26.774 13.182 26.826 13.218 ;
        RECT 27.574 13.182 27.626 13.218 ;
        RECT 28.374 13.182 28.426 13.218 ;
        RECT 29.174 13.182 29.226 13.218 ;
        RECT 29.974 13.182 30.026 13.218 ;
        RECT 30.774 13.182 30.826 13.218 ;
        RECT 31.574 13.182 31.626 13.218 ;
        RECT 32.374 13.182 32.426 13.218 ;
        RECT 33.174 13.182 33.226 13.218 ;
        RECT 33.974 13.182 34.026 13.218 ;
        RECT 34.774 13.182 34.826 13.218 ;
        RECT 35.574 13.182 35.626 13.218 ;
        RECT 18.564 13.7875 18.636 13.8125 ;
        RECT 18.864 13.7875 18.936 13.8125 ;
        RECT 0.574 13.782 0.626 13.818 ;
        RECT 1.374 13.782 1.426 13.818 ;
        RECT 2.174 13.782 2.226 13.818 ;
        RECT 2.974 13.782 3.026 13.818 ;
        RECT 3.774 13.782 3.826 13.818 ;
        RECT 4.574 13.782 4.626 13.818 ;
        RECT 5.374 13.782 5.426 13.818 ;
        RECT 6.174 13.782 6.226 13.818 ;
        RECT 6.974 13.782 7.026 13.818 ;
        RECT 7.774 13.782 7.826 13.818 ;
        RECT 8.574 13.782 8.626 13.818 ;
        RECT 9.374 13.782 9.426 13.818 ;
        RECT 10.174 13.782 10.226 13.818 ;
        RECT 10.974 13.782 11.026 13.818 ;
        RECT 11.774 13.782 11.826 13.818 ;
        RECT 12.574 13.782 12.626 13.818 ;
        RECT 13.374 13.782 13.426 13.818 ;
        RECT 14.45 13.782 14.504 13.818 ;
        RECT 15.658 13.782 15.71 13.818 ;
        RECT 15.954 13.782 16.006 13.818 ;
        RECT 16.266 13.782 16.318 13.818 ;
        RECT 16.498 13.782 16.55 13.818 ;
        RECT 17.344 13.782 17.384 13.818 ;
        RECT 17.684 13.782 17.736 13.818 ;
        RECT 19.45 13.782 19.502 13.818 ;
        RECT 19.682 13.782 19.734 13.818 ;
        RECT 19.994 13.782 20.046 13.818 ;
        RECT 20.29 13.782 20.342 13.818 ;
        RECT 21.496 13.782 21.55 13.818 ;
        RECT 22.774 13.782 22.826 13.818 ;
        RECT 23.574 13.782 23.626 13.818 ;
        RECT 24.374 13.782 24.426 13.818 ;
        RECT 25.174 13.782 25.226 13.818 ;
        RECT 25.974 13.782 26.026 13.818 ;
        RECT 26.774 13.782 26.826 13.818 ;
        RECT 27.574 13.782 27.626 13.818 ;
        RECT 28.374 13.782 28.426 13.818 ;
        RECT 29.174 13.782 29.226 13.818 ;
        RECT 29.974 13.782 30.026 13.818 ;
        RECT 30.774 13.782 30.826 13.818 ;
        RECT 31.574 13.782 31.626 13.818 ;
        RECT 32.374 13.782 32.426 13.818 ;
        RECT 33.174 13.782 33.226 13.818 ;
        RECT 33.974 13.782 34.026 13.818 ;
        RECT 34.774 13.782 34.826 13.818 ;
        RECT 35.574 13.782 35.626 13.818 ;
        RECT 18.564 14.3875 18.636 14.4125 ;
        RECT 18.864 14.3875 18.936 14.4125 ;
        RECT 0.574 14.382 0.626 14.418 ;
        RECT 1.374 14.382 1.426 14.418 ;
        RECT 2.174 14.382 2.226 14.418 ;
        RECT 2.974 14.382 3.026 14.418 ;
        RECT 3.774 14.382 3.826 14.418 ;
        RECT 4.574 14.382 4.626 14.418 ;
        RECT 5.374 14.382 5.426 14.418 ;
        RECT 6.174 14.382 6.226 14.418 ;
        RECT 6.974 14.382 7.026 14.418 ;
        RECT 7.774 14.382 7.826 14.418 ;
        RECT 8.574 14.382 8.626 14.418 ;
        RECT 9.374 14.382 9.426 14.418 ;
        RECT 10.174 14.382 10.226 14.418 ;
        RECT 10.974 14.382 11.026 14.418 ;
        RECT 11.774 14.382 11.826 14.418 ;
        RECT 12.574 14.382 12.626 14.418 ;
        RECT 13.374 14.382 13.426 14.418 ;
        RECT 14.45 14.382 14.504 14.418 ;
        RECT 15.658 14.382 15.71 14.418 ;
        RECT 15.954 14.382 16.006 14.418 ;
        RECT 16.266 14.382 16.318 14.418 ;
        RECT 16.498 14.382 16.55 14.418 ;
        RECT 17.344 14.382 17.384 14.418 ;
        RECT 17.684 14.382 17.736 14.418 ;
        RECT 19.45 14.382 19.502 14.418 ;
        RECT 19.682 14.382 19.734 14.418 ;
        RECT 19.994 14.382 20.046 14.418 ;
        RECT 20.29 14.382 20.342 14.418 ;
        RECT 21.496 14.382 21.55 14.418 ;
        RECT 22.774 14.382 22.826 14.418 ;
        RECT 23.574 14.382 23.626 14.418 ;
        RECT 24.374 14.382 24.426 14.418 ;
        RECT 25.174 14.382 25.226 14.418 ;
        RECT 25.974 14.382 26.026 14.418 ;
        RECT 26.774 14.382 26.826 14.418 ;
        RECT 27.574 14.382 27.626 14.418 ;
        RECT 28.374 14.382 28.426 14.418 ;
        RECT 29.174 14.382 29.226 14.418 ;
        RECT 29.974 14.382 30.026 14.418 ;
        RECT 30.774 14.382 30.826 14.418 ;
        RECT 31.574 14.382 31.626 14.418 ;
        RECT 32.374 14.382 32.426 14.418 ;
        RECT 33.174 14.382 33.226 14.418 ;
        RECT 33.974 14.382 34.026 14.418 ;
        RECT 34.774 14.382 34.826 14.418 ;
        RECT 35.574 14.382 35.626 14.418 ;
        RECT 18.564 14.9875 18.636 15.0125 ;
        RECT 18.864 14.9875 18.936 15.0125 ;
        RECT 0.574 14.982 0.626 15.018 ;
        RECT 1.374 14.982 1.426 15.018 ;
        RECT 2.174 14.982 2.226 15.018 ;
        RECT 2.974 14.982 3.026 15.018 ;
        RECT 3.774 14.982 3.826 15.018 ;
        RECT 4.574 14.982 4.626 15.018 ;
        RECT 5.374 14.982 5.426 15.018 ;
        RECT 6.174 14.982 6.226 15.018 ;
        RECT 6.974 14.982 7.026 15.018 ;
        RECT 7.774 14.982 7.826 15.018 ;
        RECT 8.574 14.982 8.626 15.018 ;
        RECT 9.374 14.982 9.426 15.018 ;
        RECT 10.174 14.982 10.226 15.018 ;
        RECT 10.974 14.982 11.026 15.018 ;
        RECT 11.774 14.982 11.826 15.018 ;
        RECT 12.574 14.982 12.626 15.018 ;
        RECT 13.374 14.982 13.426 15.018 ;
        RECT 14.45 14.982 14.504 15.018 ;
        RECT 15.658 14.982 15.71 15.018 ;
        RECT 15.954 14.982 16.006 15.018 ;
        RECT 16.266 14.982 16.318 15.018 ;
        RECT 16.498 14.982 16.55 15.018 ;
        RECT 17.344 14.982 17.384 15.018 ;
        RECT 17.684 14.982 17.736 15.018 ;
        RECT 19.45 14.982 19.502 15.018 ;
        RECT 19.682 14.982 19.734 15.018 ;
        RECT 19.994 14.982 20.046 15.018 ;
        RECT 20.29 14.982 20.342 15.018 ;
        RECT 21.496 14.982 21.55 15.018 ;
        RECT 22.774 14.982 22.826 15.018 ;
        RECT 23.574 14.982 23.626 15.018 ;
        RECT 24.374 14.982 24.426 15.018 ;
        RECT 25.174 14.982 25.226 15.018 ;
        RECT 25.974 14.982 26.026 15.018 ;
        RECT 26.774 14.982 26.826 15.018 ;
        RECT 27.574 14.982 27.626 15.018 ;
        RECT 28.374 14.982 28.426 15.018 ;
        RECT 29.174 14.982 29.226 15.018 ;
        RECT 29.974 14.982 30.026 15.018 ;
        RECT 30.774 14.982 30.826 15.018 ;
        RECT 31.574 14.982 31.626 15.018 ;
        RECT 32.374 14.982 32.426 15.018 ;
        RECT 33.174 14.982 33.226 15.018 ;
        RECT 33.974 14.982 34.026 15.018 ;
        RECT 34.774 14.982 34.826 15.018 ;
        RECT 35.574 14.982 35.626 15.018 ;
        RECT 18.564 15.5875 18.636 15.6125 ;
        RECT 18.864 15.5875 18.936 15.6125 ;
        RECT 0.574 15.582 0.626 15.618 ;
        RECT 1.374 15.582 1.426 15.618 ;
        RECT 2.174 15.582 2.226 15.618 ;
        RECT 2.974 15.582 3.026 15.618 ;
        RECT 3.774 15.582 3.826 15.618 ;
        RECT 4.574 15.582 4.626 15.618 ;
        RECT 5.374 15.582 5.426 15.618 ;
        RECT 6.174 15.582 6.226 15.618 ;
        RECT 6.974 15.582 7.026 15.618 ;
        RECT 7.774 15.582 7.826 15.618 ;
        RECT 8.574 15.582 8.626 15.618 ;
        RECT 9.374 15.582 9.426 15.618 ;
        RECT 10.174 15.582 10.226 15.618 ;
        RECT 10.974 15.582 11.026 15.618 ;
        RECT 11.774 15.582 11.826 15.618 ;
        RECT 12.574 15.582 12.626 15.618 ;
        RECT 13.374 15.582 13.426 15.618 ;
        RECT 14.45 15.582 14.504 15.618 ;
        RECT 15.658 15.582 15.71 15.618 ;
        RECT 15.954 15.582 16.006 15.618 ;
        RECT 16.266 15.582 16.318 15.618 ;
        RECT 16.498 15.582 16.55 15.618 ;
        RECT 17.344 15.582 17.384 15.618 ;
        RECT 17.684 15.582 17.736 15.618 ;
        RECT 19.45 15.582 19.502 15.618 ;
        RECT 19.682 15.582 19.734 15.618 ;
        RECT 19.994 15.582 20.046 15.618 ;
        RECT 20.29 15.582 20.342 15.618 ;
        RECT 21.496 15.582 21.55 15.618 ;
        RECT 22.774 15.582 22.826 15.618 ;
        RECT 23.574 15.582 23.626 15.618 ;
        RECT 24.374 15.582 24.426 15.618 ;
        RECT 25.174 15.582 25.226 15.618 ;
        RECT 25.974 15.582 26.026 15.618 ;
        RECT 26.774 15.582 26.826 15.618 ;
        RECT 27.574 15.582 27.626 15.618 ;
        RECT 28.374 15.582 28.426 15.618 ;
        RECT 29.174 15.582 29.226 15.618 ;
        RECT 29.974 15.582 30.026 15.618 ;
        RECT 30.774 15.582 30.826 15.618 ;
        RECT 31.574 15.582 31.626 15.618 ;
        RECT 32.374 15.582 32.426 15.618 ;
        RECT 33.174 15.582 33.226 15.618 ;
        RECT 33.974 15.582 34.026 15.618 ;
        RECT 34.774 15.582 34.826 15.618 ;
        RECT 35.574 15.582 35.626 15.618 ;
        RECT 18.564 16.1875 18.636 16.2125 ;
        RECT 18.864 16.1875 18.936 16.2125 ;
        RECT 0.574 16.182 0.626 16.218 ;
        RECT 1.374 16.182 1.426 16.218 ;
        RECT 2.174 16.182 2.226 16.218 ;
        RECT 2.974 16.182 3.026 16.218 ;
        RECT 3.774 16.182 3.826 16.218 ;
        RECT 4.574 16.182 4.626 16.218 ;
        RECT 5.374 16.182 5.426 16.218 ;
        RECT 6.174 16.182 6.226 16.218 ;
        RECT 6.974 16.182 7.026 16.218 ;
        RECT 7.774 16.182 7.826 16.218 ;
        RECT 8.574 16.182 8.626 16.218 ;
        RECT 9.374 16.182 9.426 16.218 ;
        RECT 10.174 16.182 10.226 16.218 ;
        RECT 10.974 16.182 11.026 16.218 ;
        RECT 11.774 16.182 11.826 16.218 ;
        RECT 12.574 16.182 12.626 16.218 ;
        RECT 13.374 16.182 13.426 16.218 ;
        RECT 14.45 16.182 14.504 16.218 ;
        RECT 15.658 16.182 15.71 16.218 ;
        RECT 15.954 16.182 16.006 16.218 ;
        RECT 16.266 16.182 16.318 16.218 ;
        RECT 16.498 16.182 16.55 16.218 ;
        RECT 17.344 16.182 17.384 16.218 ;
        RECT 17.684 16.182 17.736 16.218 ;
        RECT 19.45 16.182 19.502 16.218 ;
        RECT 19.682 16.182 19.734 16.218 ;
        RECT 19.994 16.182 20.046 16.218 ;
        RECT 20.29 16.182 20.342 16.218 ;
        RECT 21.496 16.182 21.55 16.218 ;
        RECT 22.774 16.182 22.826 16.218 ;
        RECT 23.574 16.182 23.626 16.218 ;
        RECT 24.374 16.182 24.426 16.218 ;
        RECT 25.174 16.182 25.226 16.218 ;
        RECT 25.974 16.182 26.026 16.218 ;
        RECT 26.774 16.182 26.826 16.218 ;
        RECT 27.574 16.182 27.626 16.218 ;
        RECT 28.374 16.182 28.426 16.218 ;
        RECT 29.174 16.182 29.226 16.218 ;
        RECT 29.974 16.182 30.026 16.218 ;
        RECT 30.774 16.182 30.826 16.218 ;
        RECT 31.574 16.182 31.626 16.218 ;
        RECT 32.374 16.182 32.426 16.218 ;
        RECT 33.174 16.182 33.226 16.218 ;
        RECT 33.974 16.182 34.026 16.218 ;
        RECT 34.774 16.182 34.826 16.218 ;
        RECT 35.574 16.182 35.626 16.218 ;
        RECT 18.564 16.7875 18.636 16.8125 ;
        RECT 18.864 16.7875 18.936 16.8125 ;
        RECT 0.574 16.782 0.626 16.818 ;
        RECT 1.374 16.782 1.426 16.818 ;
        RECT 2.174 16.782 2.226 16.818 ;
        RECT 2.974 16.782 3.026 16.818 ;
        RECT 3.774 16.782 3.826 16.818 ;
        RECT 4.574 16.782 4.626 16.818 ;
        RECT 5.374 16.782 5.426 16.818 ;
        RECT 6.174 16.782 6.226 16.818 ;
        RECT 6.974 16.782 7.026 16.818 ;
        RECT 7.774 16.782 7.826 16.818 ;
        RECT 8.574 16.782 8.626 16.818 ;
        RECT 9.374 16.782 9.426 16.818 ;
        RECT 10.174 16.782 10.226 16.818 ;
        RECT 10.974 16.782 11.026 16.818 ;
        RECT 11.774 16.782 11.826 16.818 ;
        RECT 12.574 16.782 12.626 16.818 ;
        RECT 13.374 16.782 13.426 16.818 ;
        RECT 14.45 16.782 14.504 16.818 ;
        RECT 15.658 16.782 15.71 16.818 ;
        RECT 15.954 16.782 16.006 16.818 ;
        RECT 16.266 16.782 16.318 16.818 ;
        RECT 16.498 16.782 16.55 16.818 ;
        RECT 17.344 16.782 17.384 16.818 ;
        RECT 17.684 16.782 17.736 16.818 ;
        RECT 19.45 16.782 19.502 16.818 ;
        RECT 19.682 16.782 19.734 16.818 ;
        RECT 19.994 16.782 20.046 16.818 ;
        RECT 20.29 16.782 20.342 16.818 ;
        RECT 21.496 16.782 21.55 16.818 ;
        RECT 22.774 16.782 22.826 16.818 ;
        RECT 23.574 16.782 23.626 16.818 ;
        RECT 24.374 16.782 24.426 16.818 ;
        RECT 25.174 16.782 25.226 16.818 ;
        RECT 25.974 16.782 26.026 16.818 ;
        RECT 26.774 16.782 26.826 16.818 ;
        RECT 27.574 16.782 27.626 16.818 ;
        RECT 28.374 16.782 28.426 16.818 ;
        RECT 29.174 16.782 29.226 16.818 ;
        RECT 29.974 16.782 30.026 16.818 ;
        RECT 30.774 16.782 30.826 16.818 ;
        RECT 31.574 16.782 31.626 16.818 ;
        RECT 32.374 16.782 32.426 16.818 ;
        RECT 33.174 16.782 33.226 16.818 ;
        RECT 33.974 16.782 34.026 16.818 ;
        RECT 34.774 16.782 34.826 16.818 ;
        RECT 35.574 16.782 35.626 16.818 ;
        RECT 18.564 17.3875 18.636 17.4125 ;
        RECT 18.864 17.3875 18.936 17.4125 ;
        RECT 0.574 17.382 0.626 17.418 ;
        RECT 1.374 17.382 1.426 17.418 ;
        RECT 2.174 17.382 2.226 17.418 ;
        RECT 2.974 17.382 3.026 17.418 ;
        RECT 3.774 17.382 3.826 17.418 ;
        RECT 4.574 17.382 4.626 17.418 ;
        RECT 5.374 17.382 5.426 17.418 ;
        RECT 6.174 17.382 6.226 17.418 ;
        RECT 6.974 17.382 7.026 17.418 ;
        RECT 7.774 17.382 7.826 17.418 ;
        RECT 8.574 17.382 8.626 17.418 ;
        RECT 9.374 17.382 9.426 17.418 ;
        RECT 10.174 17.382 10.226 17.418 ;
        RECT 10.974 17.382 11.026 17.418 ;
        RECT 11.774 17.382 11.826 17.418 ;
        RECT 12.574 17.382 12.626 17.418 ;
        RECT 13.374 17.382 13.426 17.418 ;
        RECT 14.45 17.382 14.504 17.418 ;
        RECT 15.658 17.382 15.71 17.418 ;
        RECT 15.954 17.382 16.006 17.418 ;
        RECT 16.266 17.382 16.318 17.418 ;
        RECT 16.498 17.382 16.55 17.418 ;
        RECT 17.344 17.382 17.384 17.418 ;
        RECT 17.684 17.382 17.736 17.418 ;
        RECT 19.45 17.382 19.502 17.418 ;
        RECT 19.682 17.382 19.734 17.418 ;
        RECT 19.994 17.382 20.046 17.418 ;
        RECT 20.29 17.382 20.342 17.418 ;
        RECT 21.496 17.382 21.55 17.418 ;
        RECT 22.774 17.382 22.826 17.418 ;
        RECT 23.574 17.382 23.626 17.418 ;
        RECT 24.374 17.382 24.426 17.418 ;
        RECT 25.174 17.382 25.226 17.418 ;
        RECT 25.974 17.382 26.026 17.418 ;
        RECT 26.774 17.382 26.826 17.418 ;
        RECT 27.574 17.382 27.626 17.418 ;
        RECT 28.374 17.382 28.426 17.418 ;
        RECT 29.174 17.382 29.226 17.418 ;
        RECT 29.974 17.382 30.026 17.418 ;
        RECT 30.774 17.382 30.826 17.418 ;
        RECT 31.574 17.382 31.626 17.418 ;
        RECT 32.374 17.382 32.426 17.418 ;
        RECT 33.174 17.382 33.226 17.418 ;
        RECT 33.974 17.382 34.026 17.418 ;
        RECT 34.774 17.382 34.826 17.418 ;
        RECT 35.574 17.382 35.626 17.418 ;
        RECT 18.564 17.9875 18.636 18.0125 ;
        RECT 18.864 17.9875 18.936 18.0125 ;
        RECT 0.574 17.982 0.626 18.018 ;
        RECT 1.374 17.982 1.426 18.018 ;
        RECT 2.174 17.982 2.226 18.018 ;
        RECT 2.974 17.982 3.026 18.018 ;
        RECT 3.774 17.982 3.826 18.018 ;
        RECT 4.574 17.982 4.626 18.018 ;
        RECT 5.374 17.982 5.426 18.018 ;
        RECT 6.174 17.982 6.226 18.018 ;
        RECT 6.974 17.982 7.026 18.018 ;
        RECT 7.774 17.982 7.826 18.018 ;
        RECT 8.574 17.982 8.626 18.018 ;
        RECT 9.374 17.982 9.426 18.018 ;
        RECT 10.174 17.982 10.226 18.018 ;
        RECT 10.974 17.982 11.026 18.018 ;
        RECT 11.774 17.982 11.826 18.018 ;
        RECT 12.574 17.982 12.626 18.018 ;
        RECT 13.374 17.982 13.426 18.018 ;
        RECT 14.45 17.982 14.504 18.018 ;
        RECT 15.658 17.982 15.71 18.018 ;
        RECT 15.954 17.982 16.006 18.018 ;
        RECT 16.266 17.982 16.318 18.018 ;
        RECT 16.498 17.982 16.55 18.018 ;
        RECT 17.344 17.982 17.384 18.018 ;
        RECT 17.684 17.982 17.736 18.018 ;
        RECT 19.45 17.982 19.502 18.018 ;
        RECT 19.682 17.982 19.734 18.018 ;
        RECT 19.994 17.982 20.046 18.018 ;
        RECT 20.29 17.982 20.342 18.018 ;
        RECT 21.496 17.982 21.55 18.018 ;
        RECT 22.774 17.982 22.826 18.018 ;
        RECT 23.574 17.982 23.626 18.018 ;
        RECT 24.374 17.982 24.426 18.018 ;
        RECT 25.174 17.982 25.226 18.018 ;
        RECT 25.974 17.982 26.026 18.018 ;
        RECT 26.774 17.982 26.826 18.018 ;
        RECT 27.574 17.982 27.626 18.018 ;
        RECT 28.374 17.982 28.426 18.018 ;
        RECT 29.174 17.982 29.226 18.018 ;
        RECT 29.974 17.982 30.026 18.018 ;
        RECT 30.774 17.982 30.826 18.018 ;
        RECT 31.574 17.982 31.626 18.018 ;
        RECT 32.374 17.982 32.426 18.018 ;
        RECT 33.174 17.982 33.226 18.018 ;
        RECT 33.974 17.982 34.026 18.018 ;
        RECT 34.774 17.982 34.826 18.018 ;
        RECT 35.574 17.982 35.626 18.018 ;
        RECT 18.564 18.5875 18.636 18.6125 ;
        RECT 18.864 18.5875 18.936 18.6125 ;
        RECT 0.574 18.582 0.626 18.618 ;
        RECT 1.374 18.582 1.426 18.618 ;
        RECT 2.174 18.582 2.226 18.618 ;
        RECT 2.974 18.582 3.026 18.618 ;
        RECT 3.774 18.582 3.826 18.618 ;
        RECT 4.574 18.582 4.626 18.618 ;
        RECT 5.374 18.582 5.426 18.618 ;
        RECT 6.174 18.582 6.226 18.618 ;
        RECT 6.974 18.582 7.026 18.618 ;
        RECT 7.774 18.582 7.826 18.618 ;
        RECT 8.574 18.582 8.626 18.618 ;
        RECT 9.374 18.582 9.426 18.618 ;
        RECT 10.174 18.582 10.226 18.618 ;
        RECT 10.974 18.582 11.026 18.618 ;
        RECT 11.774 18.582 11.826 18.618 ;
        RECT 12.574 18.582 12.626 18.618 ;
        RECT 13.374 18.582 13.426 18.618 ;
        RECT 14.45 18.582 14.504 18.618 ;
        RECT 15.658 18.582 15.71 18.618 ;
        RECT 15.954 18.582 16.006 18.618 ;
        RECT 16.266 18.582 16.318 18.618 ;
        RECT 16.498 18.582 16.55 18.618 ;
        RECT 17.344 18.582 17.384 18.618 ;
        RECT 17.684 18.582 17.736 18.618 ;
        RECT 19.45 18.582 19.502 18.618 ;
        RECT 19.682 18.582 19.734 18.618 ;
        RECT 19.994 18.582 20.046 18.618 ;
        RECT 20.29 18.582 20.342 18.618 ;
        RECT 21.496 18.582 21.55 18.618 ;
        RECT 22.774 18.582 22.826 18.618 ;
        RECT 23.574 18.582 23.626 18.618 ;
        RECT 24.374 18.582 24.426 18.618 ;
        RECT 25.174 18.582 25.226 18.618 ;
        RECT 25.974 18.582 26.026 18.618 ;
        RECT 26.774 18.582 26.826 18.618 ;
        RECT 27.574 18.582 27.626 18.618 ;
        RECT 28.374 18.582 28.426 18.618 ;
        RECT 29.174 18.582 29.226 18.618 ;
        RECT 29.974 18.582 30.026 18.618 ;
        RECT 30.774 18.582 30.826 18.618 ;
        RECT 31.574 18.582 31.626 18.618 ;
        RECT 32.374 18.582 32.426 18.618 ;
        RECT 33.174 18.582 33.226 18.618 ;
        RECT 33.974 18.582 34.026 18.618 ;
        RECT 34.774 18.582 34.826 18.618 ;
        RECT 35.574 18.582 35.626 18.618 ;
        RECT 18.564 19.1875 18.636 19.2125 ;
        RECT 18.864 19.1875 18.936 19.2125 ;
        RECT 0.574 19.182 0.626 19.218 ;
        RECT 1.374 19.182 1.426 19.218 ;
        RECT 2.174 19.182 2.226 19.218 ;
        RECT 2.974 19.182 3.026 19.218 ;
        RECT 3.774 19.182 3.826 19.218 ;
        RECT 4.574 19.182 4.626 19.218 ;
        RECT 5.374 19.182 5.426 19.218 ;
        RECT 6.174 19.182 6.226 19.218 ;
        RECT 6.974 19.182 7.026 19.218 ;
        RECT 7.774 19.182 7.826 19.218 ;
        RECT 8.574 19.182 8.626 19.218 ;
        RECT 9.374 19.182 9.426 19.218 ;
        RECT 10.174 19.182 10.226 19.218 ;
        RECT 10.974 19.182 11.026 19.218 ;
        RECT 11.774 19.182 11.826 19.218 ;
        RECT 12.574 19.182 12.626 19.218 ;
        RECT 13.374 19.182 13.426 19.218 ;
        RECT 14.45 19.182 14.504 19.218 ;
        RECT 15.658 19.182 15.71 19.218 ;
        RECT 15.954 19.182 16.006 19.218 ;
        RECT 16.266 19.182 16.318 19.218 ;
        RECT 16.498 19.182 16.55 19.218 ;
        RECT 17.344 19.182 17.384 19.218 ;
        RECT 17.684 19.182 17.736 19.218 ;
        RECT 19.45 19.182 19.502 19.218 ;
        RECT 19.682 19.182 19.734 19.218 ;
        RECT 19.994 19.182 20.046 19.218 ;
        RECT 20.29 19.182 20.342 19.218 ;
        RECT 21.496 19.182 21.55 19.218 ;
        RECT 22.774 19.182 22.826 19.218 ;
        RECT 23.574 19.182 23.626 19.218 ;
        RECT 24.374 19.182 24.426 19.218 ;
        RECT 25.174 19.182 25.226 19.218 ;
        RECT 25.974 19.182 26.026 19.218 ;
        RECT 26.774 19.182 26.826 19.218 ;
        RECT 27.574 19.182 27.626 19.218 ;
        RECT 28.374 19.182 28.426 19.218 ;
        RECT 29.174 19.182 29.226 19.218 ;
        RECT 29.974 19.182 30.026 19.218 ;
        RECT 30.774 19.182 30.826 19.218 ;
        RECT 31.574 19.182 31.626 19.218 ;
        RECT 32.374 19.182 32.426 19.218 ;
        RECT 33.174 19.182 33.226 19.218 ;
        RECT 33.974 19.182 34.026 19.218 ;
        RECT 34.774 19.182 34.826 19.218 ;
        RECT 35.574 19.182 35.626 19.218 ;
        RECT 18.564 19.7875 18.636 19.8125 ;
        RECT 18.864 19.7875 18.936 19.8125 ;
        RECT 0.574 19.782 0.626 19.818 ;
        RECT 1.374 19.782 1.426 19.818 ;
        RECT 2.174 19.782 2.226 19.818 ;
        RECT 2.974 19.782 3.026 19.818 ;
        RECT 3.774 19.782 3.826 19.818 ;
        RECT 4.574 19.782 4.626 19.818 ;
        RECT 5.374 19.782 5.426 19.818 ;
        RECT 6.174 19.782 6.226 19.818 ;
        RECT 6.974 19.782 7.026 19.818 ;
        RECT 7.774 19.782 7.826 19.818 ;
        RECT 8.574 19.782 8.626 19.818 ;
        RECT 9.374 19.782 9.426 19.818 ;
        RECT 10.174 19.782 10.226 19.818 ;
        RECT 10.974 19.782 11.026 19.818 ;
        RECT 11.774 19.782 11.826 19.818 ;
        RECT 12.574 19.782 12.626 19.818 ;
        RECT 13.374 19.782 13.426 19.818 ;
        RECT 14.45 19.782 14.504 19.818 ;
        RECT 15.658 19.782 15.71 19.818 ;
        RECT 15.954 19.782 16.006 19.818 ;
        RECT 16.266 19.782 16.318 19.818 ;
        RECT 16.498 19.782 16.55 19.818 ;
        RECT 17.344 19.782 17.384 19.818 ;
        RECT 17.684 19.782 17.736 19.818 ;
        RECT 19.45 19.782 19.502 19.818 ;
        RECT 19.682 19.782 19.734 19.818 ;
        RECT 19.994 19.782 20.046 19.818 ;
        RECT 20.29 19.782 20.342 19.818 ;
        RECT 21.496 19.782 21.55 19.818 ;
        RECT 22.774 19.782 22.826 19.818 ;
        RECT 23.574 19.782 23.626 19.818 ;
        RECT 24.374 19.782 24.426 19.818 ;
        RECT 25.174 19.782 25.226 19.818 ;
        RECT 25.974 19.782 26.026 19.818 ;
        RECT 26.774 19.782 26.826 19.818 ;
        RECT 27.574 19.782 27.626 19.818 ;
        RECT 28.374 19.782 28.426 19.818 ;
        RECT 29.174 19.782 29.226 19.818 ;
        RECT 29.974 19.782 30.026 19.818 ;
        RECT 30.774 19.782 30.826 19.818 ;
        RECT 31.574 19.782 31.626 19.818 ;
        RECT 32.374 19.782 32.426 19.818 ;
        RECT 33.174 19.782 33.226 19.818 ;
        RECT 33.974 19.782 34.026 19.818 ;
        RECT 34.774 19.782 34.826 19.818 ;
        RECT 35.574 19.782 35.626 19.818 ;
        RECT 18.564 20.3875 18.636 20.4125 ;
        RECT 18.864 20.3875 18.936 20.4125 ;
        RECT 0.574 20.382 0.626 20.418 ;
        RECT 1.374 20.382 1.426 20.418 ;
        RECT 2.174 20.382 2.226 20.418 ;
        RECT 2.974 20.382 3.026 20.418 ;
        RECT 3.774 20.382 3.826 20.418 ;
        RECT 4.574 20.382 4.626 20.418 ;
        RECT 5.374 20.382 5.426 20.418 ;
        RECT 6.174 20.382 6.226 20.418 ;
        RECT 6.974 20.382 7.026 20.418 ;
        RECT 7.774 20.382 7.826 20.418 ;
        RECT 8.574 20.382 8.626 20.418 ;
        RECT 9.374 20.382 9.426 20.418 ;
        RECT 10.174 20.382 10.226 20.418 ;
        RECT 10.974 20.382 11.026 20.418 ;
        RECT 11.774 20.382 11.826 20.418 ;
        RECT 12.574 20.382 12.626 20.418 ;
        RECT 13.374 20.382 13.426 20.418 ;
        RECT 14.45 20.382 14.504 20.418 ;
        RECT 15.658 20.382 15.71 20.418 ;
        RECT 15.954 20.382 16.006 20.418 ;
        RECT 16.266 20.382 16.318 20.418 ;
        RECT 16.498 20.382 16.55 20.418 ;
        RECT 17.344 20.382 17.384 20.418 ;
        RECT 17.684 20.382 17.736 20.418 ;
        RECT 19.45 20.382 19.502 20.418 ;
        RECT 19.682 20.382 19.734 20.418 ;
        RECT 19.994 20.382 20.046 20.418 ;
        RECT 20.29 20.382 20.342 20.418 ;
        RECT 21.496 20.382 21.55 20.418 ;
        RECT 22.774 20.382 22.826 20.418 ;
        RECT 23.574 20.382 23.626 20.418 ;
        RECT 24.374 20.382 24.426 20.418 ;
        RECT 25.174 20.382 25.226 20.418 ;
        RECT 25.974 20.382 26.026 20.418 ;
        RECT 26.774 20.382 26.826 20.418 ;
        RECT 27.574 20.382 27.626 20.418 ;
        RECT 28.374 20.382 28.426 20.418 ;
        RECT 29.174 20.382 29.226 20.418 ;
        RECT 29.974 20.382 30.026 20.418 ;
        RECT 30.774 20.382 30.826 20.418 ;
        RECT 31.574 20.382 31.626 20.418 ;
        RECT 32.374 20.382 32.426 20.418 ;
        RECT 33.174 20.382 33.226 20.418 ;
        RECT 33.974 20.382 34.026 20.418 ;
        RECT 34.774 20.382 34.826 20.418 ;
        RECT 35.574 20.382 35.626 20.418 ;
        RECT 18.564 20.9875 18.636 21.0125 ;
        RECT 18.864 20.9875 18.936 21.0125 ;
        RECT 0.574 20.982 0.626 21.018 ;
        RECT 1.374 20.982 1.426 21.018 ;
        RECT 2.174 20.982 2.226 21.018 ;
        RECT 2.974 20.982 3.026 21.018 ;
        RECT 3.774 20.982 3.826 21.018 ;
        RECT 4.574 20.982 4.626 21.018 ;
        RECT 5.374 20.982 5.426 21.018 ;
        RECT 6.174 20.982 6.226 21.018 ;
        RECT 6.974 20.982 7.026 21.018 ;
        RECT 7.774 20.982 7.826 21.018 ;
        RECT 8.574 20.982 8.626 21.018 ;
        RECT 9.374 20.982 9.426 21.018 ;
        RECT 10.174 20.982 10.226 21.018 ;
        RECT 10.974 20.982 11.026 21.018 ;
        RECT 11.774 20.982 11.826 21.018 ;
        RECT 12.574 20.982 12.626 21.018 ;
        RECT 13.374 20.982 13.426 21.018 ;
        RECT 14.45 20.982 14.504 21.018 ;
        RECT 15.658 20.982 15.71 21.018 ;
        RECT 15.954 20.982 16.006 21.018 ;
        RECT 16.266 20.982 16.318 21.018 ;
        RECT 16.498 20.982 16.55 21.018 ;
        RECT 17.344 20.982 17.384 21.018 ;
        RECT 17.684 20.982 17.736 21.018 ;
        RECT 19.45 20.982 19.502 21.018 ;
        RECT 19.682 20.982 19.734 21.018 ;
        RECT 19.994 20.982 20.046 21.018 ;
        RECT 20.29 20.982 20.342 21.018 ;
        RECT 21.496 20.982 21.55 21.018 ;
        RECT 22.774 20.982 22.826 21.018 ;
        RECT 23.574 20.982 23.626 21.018 ;
        RECT 24.374 20.982 24.426 21.018 ;
        RECT 25.174 20.982 25.226 21.018 ;
        RECT 25.974 20.982 26.026 21.018 ;
        RECT 26.774 20.982 26.826 21.018 ;
        RECT 27.574 20.982 27.626 21.018 ;
        RECT 28.374 20.982 28.426 21.018 ;
        RECT 29.174 20.982 29.226 21.018 ;
        RECT 29.974 20.982 30.026 21.018 ;
        RECT 30.774 20.982 30.826 21.018 ;
        RECT 31.574 20.982 31.626 21.018 ;
        RECT 32.374 20.982 32.426 21.018 ;
        RECT 33.174 20.982 33.226 21.018 ;
        RECT 33.974 20.982 34.026 21.018 ;
        RECT 34.774 20.982 34.826 21.018 ;
        RECT 35.574 20.982 35.626 21.018 ;
        RECT 18.564 21.5875 18.636 21.6125 ;
        RECT 18.864 21.5875 18.936 21.6125 ;
        RECT 0.574 21.582 0.626 21.618 ;
        RECT 1.374 21.582 1.426 21.618 ;
        RECT 2.174 21.582 2.226 21.618 ;
        RECT 2.974 21.582 3.026 21.618 ;
        RECT 3.774 21.582 3.826 21.618 ;
        RECT 4.574 21.582 4.626 21.618 ;
        RECT 5.374 21.582 5.426 21.618 ;
        RECT 6.174 21.582 6.226 21.618 ;
        RECT 6.974 21.582 7.026 21.618 ;
        RECT 7.774 21.582 7.826 21.618 ;
        RECT 8.574 21.582 8.626 21.618 ;
        RECT 9.374 21.582 9.426 21.618 ;
        RECT 10.174 21.582 10.226 21.618 ;
        RECT 10.974 21.582 11.026 21.618 ;
        RECT 11.774 21.582 11.826 21.618 ;
        RECT 12.574 21.582 12.626 21.618 ;
        RECT 13.374 21.582 13.426 21.618 ;
        RECT 14.45 21.582 14.504 21.618 ;
        RECT 15.658 21.582 15.71 21.618 ;
        RECT 15.954 21.582 16.006 21.618 ;
        RECT 16.266 21.582 16.318 21.618 ;
        RECT 16.498 21.582 16.55 21.618 ;
        RECT 17.344 21.582 17.384 21.618 ;
        RECT 17.684 21.582 17.736 21.618 ;
        RECT 19.45 21.582 19.502 21.618 ;
        RECT 19.682 21.582 19.734 21.618 ;
        RECT 19.994 21.582 20.046 21.618 ;
        RECT 20.29 21.582 20.342 21.618 ;
        RECT 21.496 21.582 21.55 21.618 ;
        RECT 22.774 21.582 22.826 21.618 ;
        RECT 23.574 21.582 23.626 21.618 ;
        RECT 24.374 21.582 24.426 21.618 ;
        RECT 25.174 21.582 25.226 21.618 ;
        RECT 25.974 21.582 26.026 21.618 ;
        RECT 26.774 21.582 26.826 21.618 ;
        RECT 27.574 21.582 27.626 21.618 ;
        RECT 28.374 21.582 28.426 21.618 ;
        RECT 29.174 21.582 29.226 21.618 ;
        RECT 29.974 21.582 30.026 21.618 ;
        RECT 30.774 21.582 30.826 21.618 ;
        RECT 31.574 21.582 31.626 21.618 ;
        RECT 32.374 21.582 32.426 21.618 ;
        RECT 33.174 21.582 33.226 21.618 ;
        RECT 33.974 21.582 34.026 21.618 ;
        RECT 34.774 21.582 34.826 21.618 ;
        RECT 35.574 21.582 35.626 21.618 ;
        RECT 18.564 22.1875 18.636 22.2125 ;
        RECT 18.864 22.1875 18.936 22.2125 ;
        RECT 0.574 22.182 0.626 22.218 ;
        RECT 1.374 22.182 1.426 22.218 ;
        RECT 2.174 22.182 2.226 22.218 ;
        RECT 2.974 22.182 3.026 22.218 ;
        RECT 3.774 22.182 3.826 22.218 ;
        RECT 4.574 22.182 4.626 22.218 ;
        RECT 5.374 22.182 5.426 22.218 ;
        RECT 6.174 22.182 6.226 22.218 ;
        RECT 6.974 22.182 7.026 22.218 ;
        RECT 7.774 22.182 7.826 22.218 ;
        RECT 8.574 22.182 8.626 22.218 ;
        RECT 9.374 22.182 9.426 22.218 ;
        RECT 10.174 22.182 10.226 22.218 ;
        RECT 10.974 22.182 11.026 22.218 ;
        RECT 11.774 22.182 11.826 22.218 ;
        RECT 12.574 22.182 12.626 22.218 ;
        RECT 13.374 22.182 13.426 22.218 ;
        RECT 14.45 22.182 14.504 22.218 ;
        RECT 15.658 22.182 15.71 22.218 ;
        RECT 15.954 22.182 16.006 22.218 ;
        RECT 16.266 22.182 16.318 22.218 ;
        RECT 16.498 22.182 16.55 22.218 ;
        RECT 17.344 22.182 17.384 22.218 ;
        RECT 17.684 22.182 17.736 22.218 ;
        RECT 19.45 22.182 19.502 22.218 ;
        RECT 19.682 22.182 19.734 22.218 ;
        RECT 19.994 22.182 20.046 22.218 ;
        RECT 20.29 22.182 20.342 22.218 ;
        RECT 21.496 22.182 21.55 22.218 ;
        RECT 22.774 22.182 22.826 22.218 ;
        RECT 23.574 22.182 23.626 22.218 ;
        RECT 24.374 22.182 24.426 22.218 ;
        RECT 25.174 22.182 25.226 22.218 ;
        RECT 25.974 22.182 26.026 22.218 ;
        RECT 26.774 22.182 26.826 22.218 ;
        RECT 27.574 22.182 27.626 22.218 ;
        RECT 28.374 22.182 28.426 22.218 ;
        RECT 29.174 22.182 29.226 22.218 ;
        RECT 29.974 22.182 30.026 22.218 ;
        RECT 30.774 22.182 30.826 22.218 ;
        RECT 31.574 22.182 31.626 22.218 ;
        RECT 32.374 22.182 32.426 22.218 ;
        RECT 33.174 22.182 33.226 22.218 ;
        RECT 33.974 22.182 34.026 22.218 ;
        RECT 34.774 22.182 34.826 22.218 ;
        RECT 35.574 22.182 35.626 22.218 ;
        RECT 18.564 22.7875 18.636 22.8125 ;
        RECT 18.864 22.7875 18.936 22.8125 ;
        RECT 0.574 22.782 0.626 22.818 ;
        RECT 1.374 22.782 1.426 22.818 ;
        RECT 2.174 22.782 2.226 22.818 ;
        RECT 2.974 22.782 3.026 22.818 ;
        RECT 3.774 22.782 3.826 22.818 ;
        RECT 4.574 22.782 4.626 22.818 ;
        RECT 5.374 22.782 5.426 22.818 ;
        RECT 6.174 22.782 6.226 22.818 ;
        RECT 6.974 22.782 7.026 22.818 ;
        RECT 7.774 22.782 7.826 22.818 ;
        RECT 8.574 22.782 8.626 22.818 ;
        RECT 9.374 22.782 9.426 22.818 ;
        RECT 10.174 22.782 10.226 22.818 ;
        RECT 10.974 22.782 11.026 22.818 ;
        RECT 11.774 22.782 11.826 22.818 ;
        RECT 12.574 22.782 12.626 22.818 ;
        RECT 13.374 22.782 13.426 22.818 ;
        RECT 14.45 22.782 14.504 22.818 ;
        RECT 15.658 22.782 15.71 22.818 ;
        RECT 15.954 22.782 16.006 22.818 ;
        RECT 16.266 22.782 16.318 22.818 ;
        RECT 16.498 22.782 16.55 22.818 ;
        RECT 17.344 22.782 17.384 22.818 ;
        RECT 17.684 22.782 17.736 22.818 ;
        RECT 19.45 22.782 19.502 22.818 ;
        RECT 19.682 22.782 19.734 22.818 ;
        RECT 19.994 22.782 20.046 22.818 ;
        RECT 20.29 22.782 20.342 22.818 ;
        RECT 21.496 22.782 21.55 22.818 ;
        RECT 22.774 22.782 22.826 22.818 ;
        RECT 23.574 22.782 23.626 22.818 ;
        RECT 24.374 22.782 24.426 22.818 ;
        RECT 25.174 22.782 25.226 22.818 ;
        RECT 25.974 22.782 26.026 22.818 ;
        RECT 26.774 22.782 26.826 22.818 ;
        RECT 27.574 22.782 27.626 22.818 ;
        RECT 28.374 22.782 28.426 22.818 ;
        RECT 29.174 22.782 29.226 22.818 ;
        RECT 29.974 22.782 30.026 22.818 ;
        RECT 30.774 22.782 30.826 22.818 ;
        RECT 31.574 22.782 31.626 22.818 ;
        RECT 32.374 22.782 32.426 22.818 ;
        RECT 33.174 22.782 33.226 22.818 ;
        RECT 33.974 22.782 34.026 22.818 ;
        RECT 34.774 22.782 34.826 22.818 ;
        RECT 35.574 22.782 35.626 22.818 ;
        RECT 18.564 23.3875 18.636 23.4125 ;
        RECT 18.864 23.3875 18.936 23.4125 ;
        RECT 0.574 23.382 0.626 23.418 ;
        RECT 1.374 23.382 1.426 23.418 ;
        RECT 2.174 23.382 2.226 23.418 ;
        RECT 2.974 23.382 3.026 23.418 ;
        RECT 3.774 23.382 3.826 23.418 ;
        RECT 4.574 23.382 4.626 23.418 ;
        RECT 5.374 23.382 5.426 23.418 ;
        RECT 6.174 23.382 6.226 23.418 ;
        RECT 6.974 23.382 7.026 23.418 ;
        RECT 7.774 23.382 7.826 23.418 ;
        RECT 8.574 23.382 8.626 23.418 ;
        RECT 9.374 23.382 9.426 23.418 ;
        RECT 10.174 23.382 10.226 23.418 ;
        RECT 10.974 23.382 11.026 23.418 ;
        RECT 11.774 23.382 11.826 23.418 ;
        RECT 12.574 23.382 12.626 23.418 ;
        RECT 13.374 23.382 13.426 23.418 ;
        RECT 14.45 23.382 14.504 23.418 ;
        RECT 15.658 23.382 15.71 23.418 ;
        RECT 15.954 23.382 16.006 23.418 ;
        RECT 16.266 23.382 16.318 23.418 ;
        RECT 16.498 23.382 16.55 23.418 ;
        RECT 17.344 23.382 17.384 23.418 ;
        RECT 17.684 23.382 17.736 23.418 ;
        RECT 19.45 23.382 19.502 23.418 ;
        RECT 19.682 23.382 19.734 23.418 ;
        RECT 19.994 23.382 20.046 23.418 ;
        RECT 20.29 23.382 20.342 23.418 ;
        RECT 21.496 23.382 21.55 23.418 ;
        RECT 22.774 23.382 22.826 23.418 ;
        RECT 23.574 23.382 23.626 23.418 ;
        RECT 24.374 23.382 24.426 23.418 ;
        RECT 25.174 23.382 25.226 23.418 ;
        RECT 25.974 23.382 26.026 23.418 ;
        RECT 26.774 23.382 26.826 23.418 ;
        RECT 27.574 23.382 27.626 23.418 ;
        RECT 28.374 23.382 28.426 23.418 ;
        RECT 29.174 23.382 29.226 23.418 ;
        RECT 29.974 23.382 30.026 23.418 ;
        RECT 30.774 23.382 30.826 23.418 ;
        RECT 31.574 23.382 31.626 23.418 ;
        RECT 32.374 23.382 32.426 23.418 ;
        RECT 33.174 23.382 33.226 23.418 ;
        RECT 33.974 23.382 34.026 23.418 ;
        RECT 34.774 23.382 34.826 23.418 ;
        RECT 35.574 23.382 35.626 23.418 ;
        RECT 18.564 23.9875 18.636 24.0125 ;
        RECT 18.864 23.9875 18.936 24.0125 ;
        RECT 0.574 23.982 0.626 24.018 ;
        RECT 1.374 23.982 1.426 24.018 ;
        RECT 2.174 23.982 2.226 24.018 ;
        RECT 2.974 23.982 3.026 24.018 ;
        RECT 3.774 23.982 3.826 24.018 ;
        RECT 4.574 23.982 4.626 24.018 ;
        RECT 5.374 23.982 5.426 24.018 ;
        RECT 6.174 23.982 6.226 24.018 ;
        RECT 6.974 23.982 7.026 24.018 ;
        RECT 7.774 23.982 7.826 24.018 ;
        RECT 8.574 23.982 8.626 24.018 ;
        RECT 9.374 23.982 9.426 24.018 ;
        RECT 10.174 23.982 10.226 24.018 ;
        RECT 10.974 23.982 11.026 24.018 ;
        RECT 11.774 23.982 11.826 24.018 ;
        RECT 12.574 23.982 12.626 24.018 ;
        RECT 13.374 23.982 13.426 24.018 ;
        RECT 14.45 23.982 14.504 24.018 ;
        RECT 15.658 23.982 15.71 24.018 ;
        RECT 15.954 23.982 16.006 24.018 ;
        RECT 16.266 23.982 16.318 24.018 ;
        RECT 16.498 23.982 16.55 24.018 ;
        RECT 17.344 23.982 17.384 24.018 ;
        RECT 17.684 23.982 17.736 24.018 ;
        RECT 19.45 23.982 19.502 24.018 ;
        RECT 19.682 23.982 19.734 24.018 ;
        RECT 19.994 23.982 20.046 24.018 ;
        RECT 20.29 23.982 20.342 24.018 ;
        RECT 21.496 23.982 21.55 24.018 ;
        RECT 22.774 23.982 22.826 24.018 ;
        RECT 23.574 23.982 23.626 24.018 ;
        RECT 24.374 23.982 24.426 24.018 ;
        RECT 25.174 23.982 25.226 24.018 ;
        RECT 25.974 23.982 26.026 24.018 ;
        RECT 26.774 23.982 26.826 24.018 ;
        RECT 27.574 23.982 27.626 24.018 ;
        RECT 28.374 23.982 28.426 24.018 ;
        RECT 29.174 23.982 29.226 24.018 ;
        RECT 29.974 23.982 30.026 24.018 ;
        RECT 30.774 23.982 30.826 24.018 ;
        RECT 31.574 23.982 31.626 24.018 ;
        RECT 32.374 23.982 32.426 24.018 ;
        RECT 33.174 23.982 33.226 24.018 ;
        RECT 33.974 23.982 34.026 24.018 ;
        RECT 34.774 23.982 34.826 24.018 ;
        RECT 35.574 23.982 35.626 24.018 ;
        RECT 18.564 24.5875 18.636 24.6125 ;
        RECT 18.864 24.5875 18.936 24.6125 ;
        RECT 0.574 24.582 0.626 24.618 ;
        RECT 1.374 24.582 1.426 24.618 ;
        RECT 2.174 24.582 2.226 24.618 ;
        RECT 2.974 24.582 3.026 24.618 ;
        RECT 3.774 24.582 3.826 24.618 ;
        RECT 4.574 24.582 4.626 24.618 ;
        RECT 5.374 24.582 5.426 24.618 ;
        RECT 6.174 24.582 6.226 24.618 ;
        RECT 6.974 24.582 7.026 24.618 ;
        RECT 7.774 24.582 7.826 24.618 ;
        RECT 8.574 24.582 8.626 24.618 ;
        RECT 9.374 24.582 9.426 24.618 ;
        RECT 10.174 24.582 10.226 24.618 ;
        RECT 10.974 24.582 11.026 24.618 ;
        RECT 11.774 24.582 11.826 24.618 ;
        RECT 12.574 24.582 12.626 24.618 ;
        RECT 13.374 24.582 13.426 24.618 ;
        RECT 14.45 24.582 14.504 24.618 ;
        RECT 15.658 24.582 15.71 24.618 ;
        RECT 15.954 24.582 16.006 24.618 ;
        RECT 16.266 24.582 16.318 24.618 ;
        RECT 16.498 24.582 16.55 24.618 ;
        RECT 17.344 24.582 17.384 24.618 ;
        RECT 17.684 24.582 17.736 24.618 ;
        RECT 19.45 24.582 19.502 24.618 ;
        RECT 19.682 24.582 19.734 24.618 ;
        RECT 19.994 24.582 20.046 24.618 ;
        RECT 20.29 24.582 20.342 24.618 ;
        RECT 21.496 24.582 21.55 24.618 ;
        RECT 22.774 24.582 22.826 24.618 ;
        RECT 23.574 24.582 23.626 24.618 ;
        RECT 24.374 24.582 24.426 24.618 ;
        RECT 25.174 24.582 25.226 24.618 ;
        RECT 25.974 24.582 26.026 24.618 ;
        RECT 26.774 24.582 26.826 24.618 ;
        RECT 27.574 24.582 27.626 24.618 ;
        RECT 28.374 24.582 28.426 24.618 ;
        RECT 29.174 24.582 29.226 24.618 ;
        RECT 29.974 24.582 30.026 24.618 ;
        RECT 30.774 24.582 30.826 24.618 ;
        RECT 31.574 24.582 31.626 24.618 ;
        RECT 32.374 24.582 32.426 24.618 ;
        RECT 33.174 24.582 33.226 24.618 ;
        RECT 33.974 24.582 34.026 24.618 ;
        RECT 34.774 24.582 34.826 24.618 ;
        RECT 35.574 24.582 35.626 24.618 ;
        RECT 18.564 25.1875 18.636 25.2125 ;
        RECT 18.864 25.1875 18.936 25.2125 ;
        RECT 0.574 25.182 0.626 25.218 ;
        RECT 1.374 25.182 1.426 25.218 ;
        RECT 2.174 25.182 2.226 25.218 ;
        RECT 2.974 25.182 3.026 25.218 ;
        RECT 3.774 25.182 3.826 25.218 ;
        RECT 4.574 25.182 4.626 25.218 ;
        RECT 5.374 25.182 5.426 25.218 ;
        RECT 6.174 25.182 6.226 25.218 ;
        RECT 6.974 25.182 7.026 25.218 ;
        RECT 7.774 25.182 7.826 25.218 ;
        RECT 8.574 25.182 8.626 25.218 ;
        RECT 9.374 25.182 9.426 25.218 ;
        RECT 10.174 25.182 10.226 25.218 ;
        RECT 10.974 25.182 11.026 25.218 ;
        RECT 11.774 25.182 11.826 25.218 ;
        RECT 12.574 25.182 12.626 25.218 ;
        RECT 13.374 25.182 13.426 25.218 ;
        RECT 14.45 25.182 14.504 25.218 ;
        RECT 15.658 25.182 15.71 25.218 ;
        RECT 15.954 25.182 16.006 25.218 ;
        RECT 16.266 25.182 16.318 25.218 ;
        RECT 16.498 25.182 16.55 25.218 ;
        RECT 17.344 25.182 17.384 25.218 ;
        RECT 17.684 25.182 17.736 25.218 ;
        RECT 19.45 25.182 19.502 25.218 ;
        RECT 19.682 25.182 19.734 25.218 ;
        RECT 19.994 25.182 20.046 25.218 ;
        RECT 20.29 25.182 20.342 25.218 ;
        RECT 21.496 25.182 21.55 25.218 ;
        RECT 22.774 25.182 22.826 25.218 ;
        RECT 23.574 25.182 23.626 25.218 ;
        RECT 24.374 25.182 24.426 25.218 ;
        RECT 25.174 25.182 25.226 25.218 ;
        RECT 25.974 25.182 26.026 25.218 ;
        RECT 26.774 25.182 26.826 25.218 ;
        RECT 27.574 25.182 27.626 25.218 ;
        RECT 28.374 25.182 28.426 25.218 ;
        RECT 29.174 25.182 29.226 25.218 ;
        RECT 29.974 25.182 30.026 25.218 ;
        RECT 30.774 25.182 30.826 25.218 ;
        RECT 31.574 25.182 31.626 25.218 ;
        RECT 32.374 25.182 32.426 25.218 ;
        RECT 33.174 25.182 33.226 25.218 ;
        RECT 33.974 25.182 34.026 25.218 ;
        RECT 34.774 25.182 34.826 25.218 ;
        RECT 35.574 25.182 35.626 25.218 ;
        RECT 18.564 25.7875 18.636 25.8125 ;
        RECT 18.864 25.7875 18.936 25.8125 ;
        RECT 0.574 25.782 0.626 25.818 ;
        RECT 1.374 25.782 1.426 25.818 ;
        RECT 2.174 25.782 2.226 25.818 ;
        RECT 2.974 25.782 3.026 25.818 ;
        RECT 3.774 25.782 3.826 25.818 ;
        RECT 4.574 25.782 4.626 25.818 ;
        RECT 5.374 25.782 5.426 25.818 ;
        RECT 6.174 25.782 6.226 25.818 ;
        RECT 6.974 25.782 7.026 25.818 ;
        RECT 7.774 25.782 7.826 25.818 ;
        RECT 8.574 25.782 8.626 25.818 ;
        RECT 9.374 25.782 9.426 25.818 ;
        RECT 10.174 25.782 10.226 25.818 ;
        RECT 10.974 25.782 11.026 25.818 ;
        RECT 11.774 25.782 11.826 25.818 ;
        RECT 12.574 25.782 12.626 25.818 ;
        RECT 13.374 25.782 13.426 25.818 ;
        RECT 14.45 25.782 14.504 25.818 ;
        RECT 15.658 25.782 15.71 25.818 ;
        RECT 15.954 25.782 16.006 25.818 ;
        RECT 16.266 25.782 16.318 25.818 ;
        RECT 16.498 25.782 16.55 25.818 ;
        RECT 17.344 25.782 17.384 25.818 ;
        RECT 17.684 25.782 17.736 25.818 ;
        RECT 19.45 25.782 19.502 25.818 ;
        RECT 19.682 25.782 19.734 25.818 ;
        RECT 19.994 25.782 20.046 25.818 ;
        RECT 20.29 25.782 20.342 25.818 ;
        RECT 21.496 25.782 21.55 25.818 ;
        RECT 22.774 25.782 22.826 25.818 ;
        RECT 23.574 25.782 23.626 25.818 ;
        RECT 24.374 25.782 24.426 25.818 ;
        RECT 25.174 25.782 25.226 25.818 ;
        RECT 25.974 25.782 26.026 25.818 ;
        RECT 26.774 25.782 26.826 25.818 ;
        RECT 27.574 25.782 27.626 25.818 ;
        RECT 28.374 25.782 28.426 25.818 ;
        RECT 29.174 25.782 29.226 25.818 ;
        RECT 29.974 25.782 30.026 25.818 ;
        RECT 30.774 25.782 30.826 25.818 ;
        RECT 31.574 25.782 31.626 25.818 ;
        RECT 32.374 25.782 32.426 25.818 ;
        RECT 33.174 25.782 33.226 25.818 ;
        RECT 33.974 25.782 34.026 25.818 ;
        RECT 34.774 25.782 34.826 25.818 ;
        RECT 35.574 25.782 35.626 25.818 ;
        RECT 18.564 26.3875 18.636 26.4125 ;
        RECT 18.864 26.3875 18.936 26.4125 ;
        RECT 0.574 26.382 0.626 26.418 ;
        RECT 1.374 26.382 1.426 26.418 ;
        RECT 2.174 26.382 2.226 26.418 ;
        RECT 2.974 26.382 3.026 26.418 ;
        RECT 3.774 26.382 3.826 26.418 ;
        RECT 4.574 26.382 4.626 26.418 ;
        RECT 5.374 26.382 5.426 26.418 ;
        RECT 6.174 26.382 6.226 26.418 ;
        RECT 6.974 26.382 7.026 26.418 ;
        RECT 7.774 26.382 7.826 26.418 ;
        RECT 8.574 26.382 8.626 26.418 ;
        RECT 9.374 26.382 9.426 26.418 ;
        RECT 10.174 26.382 10.226 26.418 ;
        RECT 10.974 26.382 11.026 26.418 ;
        RECT 11.774 26.382 11.826 26.418 ;
        RECT 12.574 26.382 12.626 26.418 ;
        RECT 13.374 26.382 13.426 26.418 ;
        RECT 14.45 26.382 14.504 26.418 ;
        RECT 15.658 26.382 15.71 26.418 ;
        RECT 15.954 26.382 16.006 26.418 ;
        RECT 16.266 26.382 16.318 26.418 ;
        RECT 16.498 26.382 16.55 26.418 ;
        RECT 17.344 26.382 17.384 26.418 ;
        RECT 17.684 26.382 17.736 26.418 ;
        RECT 19.45 26.382 19.502 26.418 ;
        RECT 19.682 26.382 19.734 26.418 ;
        RECT 19.994 26.382 20.046 26.418 ;
        RECT 20.29 26.382 20.342 26.418 ;
        RECT 21.496 26.382 21.55 26.418 ;
        RECT 22.774 26.382 22.826 26.418 ;
        RECT 23.574 26.382 23.626 26.418 ;
        RECT 24.374 26.382 24.426 26.418 ;
        RECT 25.174 26.382 25.226 26.418 ;
        RECT 25.974 26.382 26.026 26.418 ;
        RECT 26.774 26.382 26.826 26.418 ;
        RECT 27.574 26.382 27.626 26.418 ;
        RECT 28.374 26.382 28.426 26.418 ;
        RECT 29.174 26.382 29.226 26.418 ;
        RECT 29.974 26.382 30.026 26.418 ;
        RECT 30.774 26.382 30.826 26.418 ;
        RECT 31.574 26.382 31.626 26.418 ;
        RECT 32.374 26.382 32.426 26.418 ;
        RECT 33.174 26.382 33.226 26.418 ;
        RECT 33.974 26.382 34.026 26.418 ;
        RECT 34.774 26.382 34.826 26.418 ;
        RECT 35.574 26.382 35.626 26.418 ;
        RECT 18.564 26.9875 18.636 27.0125 ;
        RECT 18.864 26.9875 18.936 27.0125 ;
        RECT 0.574 26.982 0.626 27.018 ;
        RECT 1.374 26.982 1.426 27.018 ;
        RECT 2.174 26.982 2.226 27.018 ;
        RECT 2.974 26.982 3.026 27.018 ;
        RECT 3.774 26.982 3.826 27.018 ;
        RECT 4.574 26.982 4.626 27.018 ;
        RECT 5.374 26.982 5.426 27.018 ;
        RECT 6.174 26.982 6.226 27.018 ;
        RECT 6.974 26.982 7.026 27.018 ;
        RECT 7.774 26.982 7.826 27.018 ;
        RECT 8.574 26.982 8.626 27.018 ;
        RECT 9.374 26.982 9.426 27.018 ;
        RECT 10.174 26.982 10.226 27.018 ;
        RECT 10.974 26.982 11.026 27.018 ;
        RECT 11.774 26.982 11.826 27.018 ;
        RECT 12.574 26.982 12.626 27.018 ;
        RECT 13.374 26.982 13.426 27.018 ;
        RECT 14.45 26.982 14.504 27.018 ;
        RECT 15.658 26.982 15.71 27.018 ;
        RECT 15.954 26.982 16.006 27.018 ;
        RECT 16.266 26.982 16.318 27.018 ;
        RECT 16.498 26.982 16.55 27.018 ;
        RECT 17.344 26.982 17.384 27.018 ;
        RECT 17.684 26.982 17.736 27.018 ;
        RECT 19.45 26.982 19.502 27.018 ;
        RECT 19.682 26.982 19.734 27.018 ;
        RECT 19.994 26.982 20.046 27.018 ;
        RECT 20.29 26.982 20.342 27.018 ;
        RECT 21.496 26.982 21.55 27.018 ;
        RECT 22.774 26.982 22.826 27.018 ;
        RECT 23.574 26.982 23.626 27.018 ;
        RECT 24.374 26.982 24.426 27.018 ;
        RECT 25.174 26.982 25.226 27.018 ;
        RECT 25.974 26.982 26.026 27.018 ;
        RECT 26.774 26.982 26.826 27.018 ;
        RECT 27.574 26.982 27.626 27.018 ;
        RECT 28.374 26.982 28.426 27.018 ;
        RECT 29.174 26.982 29.226 27.018 ;
        RECT 29.974 26.982 30.026 27.018 ;
        RECT 30.774 26.982 30.826 27.018 ;
        RECT 31.574 26.982 31.626 27.018 ;
        RECT 32.374 26.982 32.426 27.018 ;
        RECT 33.174 26.982 33.226 27.018 ;
        RECT 33.974 26.982 34.026 27.018 ;
        RECT 34.774 26.982 34.826 27.018 ;
        RECT 35.574 26.982 35.626 27.018 ;
        RECT 18.564 27.5875 18.636 27.6125 ;
        RECT 18.864 27.5875 18.936 27.6125 ;
        RECT 0.574 27.582 0.626 27.618 ;
        RECT 1.374 27.582 1.426 27.618 ;
        RECT 2.174 27.582 2.226 27.618 ;
        RECT 2.974 27.582 3.026 27.618 ;
        RECT 3.774 27.582 3.826 27.618 ;
        RECT 4.574 27.582 4.626 27.618 ;
        RECT 5.374 27.582 5.426 27.618 ;
        RECT 6.174 27.582 6.226 27.618 ;
        RECT 6.974 27.582 7.026 27.618 ;
        RECT 7.774 27.582 7.826 27.618 ;
        RECT 8.574 27.582 8.626 27.618 ;
        RECT 9.374 27.582 9.426 27.618 ;
        RECT 10.174 27.582 10.226 27.618 ;
        RECT 10.974 27.582 11.026 27.618 ;
        RECT 11.774 27.582 11.826 27.618 ;
        RECT 12.574 27.582 12.626 27.618 ;
        RECT 13.374 27.582 13.426 27.618 ;
        RECT 14.45 27.582 14.504 27.618 ;
        RECT 15.658 27.582 15.71 27.618 ;
        RECT 15.954 27.582 16.006 27.618 ;
        RECT 16.266 27.582 16.318 27.618 ;
        RECT 16.498 27.582 16.55 27.618 ;
        RECT 17.344 27.582 17.384 27.618 ;
        RECT 17.684 27.582 17.736 27.618 ;
        RECT 19.45 27.582 19.502 27.618 ;
        RECT 19.682 27.582 19.734 27.618 ;
        RECT 19.994 27.582 20.046 27.618 ;
        RECT 20.29 27.582 20.342 27.618 ;
        RECT 21.496 27.582 21.55 27.618 ;
        RECT 22.774 27.582 22.826 27.618 ;
        RECT 23.574 27.582 23.626 27.618 ;
        RECT 24.374 27.582 24.426 27.618 ;
        RECT 25.174 27.582 25.226 27.618 ;
        RECT 25.974 27.582 26.026 27.618 ;
        RECT 26.774 27.582 26.826 27.618 ;
        RECT 27.574 27.582 27.626 27.618 ;
        RECT 28.374 27.582 28.426 27.618 ;
        RECT 29.174 27.582 29.226 27.618 ;
        RECT 29.974 27.582 30.026 27.618 ;
        RECT 30.774 27.582 30.826 27.618 ;
        RECT 31.574 27.582 31.626 27.618 ;
        RECT 32.374 27.582 32.426 27.618 ;
        RECT 33.174 27.582 33.226 27.618 ;
        RECT 33.974 27.582 34.026 27.618 ;
        RECT 34.774 27.582 34.826 27.618 ;
        RECT 35.574 27.582 35.626 27.618 ;
        RECT 18.564 28.1875 18.636 28.2125 ;
        RECT 18.864 28.1875 18.936 28.2125 ;
        RECT 0.574 28.182 0.626 28.218 ;
        RECT 1.374 28.182 1.426 28.218 ;
        RECT 2.174 28.182 2.226 28.218 ;
        RECT 2.974 28.182 3.026 28.218 ;
        RECT 3.774 28.182 3.826 28.218 ;
        RECT 4.574 28.182 4.626 28.218 ;
        RECT 5.374 28.182 5.426 28.218 ;
        RECT 6.174 28.182 6.226 28.218 ;
        RECT 6.974 28.182 7.026 28.218 ;
        RECT 7.774 28.182 7.826 28.218 ;
        RECT 8.574 28.182 8.626 28.218 ;
        RECT 9.374 28.182 9.426 28.218 ;
        RECT 10.174 28.182 10.226 28.218 ;
        RECT 10.974 28.182 11.026 28.218 ;
        RECT 11.774 28.182 11.826 28.218 ;
        RECT 12.574 28.182 12.626 28.218 ;
        RECT 13.374 28.182 13.426 28.218 ;
        RECT 14.45 28.182 14.504 28.218 ;
        RECT 15.658 28.182 15.71 28.218 ;
        RECT 15.954 28.182 16.006 28.218 ;
        RECT 16.266 28.182 16.318 28.218 ;
        RECT 16.498 28.182 16.55 28.218 ;
        RECT 17.344 28.182 17.384 28.218 ;
        RECT 17.684 28.182 17.736 28.218 ;
        RECT 19.45 28.182 19.502 28.218 ;
        RECT 19.682 28.182 19.734 28.218 ;
        RECT 19.994 28.182 20.046 28.218 ;
        RECT 20.29 28.182 20.342 28.218 ;
        RECT 21.496 28.182 21.55 28.218 ;
        RECT 22.774 28.182 22.826 28.218 ;
        RECT 23.574 28.182 23.626 28.218 ;
        RECT 24.374 28.182 24.426 28.218 ;
        RECT 25.174 28.182 25.226 28.218 ;
        RECT 25.974 28.182 26.026 28.218 ;
        RECT 26.774 28.182 26.826 28.218 ;
        RECT 27.574 28.182 27.626 28.218 ;
        RECT 28.374 28.182 28.426 28.218 ;
        RECT 29.174 28.182 29.226 28.218 ;
        RECT 29.974 28.182 30.026 28.218 ;
        RECT 30.774 28.182 30.826 28.218 ;
        RECT 31.574 28.182 31.626 28.218 ;
        RECT 32.374 28.182 32.426 28.218 ;
        RECT 33.174 28.182 33.226 28.218 ;
        RECT 33.974 28.182 34.026 28.218 ;
        RECT 34.774 28.182 34.826 28.218 ;
        RECT 35.574 28.182 35.626 28.218 ;
        RECT 18.564 28.7875 18.636 28.8125 ;
        RECT 18.864 28.7875 18.936 28.8125 ;
        RECT 0.574 28.782 0.626 28.818 ;
        RECT 1.374 28.782 1.426 28.818 ;
        RECT 2.174 28.782 2.226 28.818 ;
        RECT 2.974 28.782 3.026 28.818 ;
        RECT 3.774 28.782 3.826 28.818 ;
        RECT 4.574 28.782 4.626 28.818 ;
        RECT 5.374 28.782 5.426 28.818 ;
        RECT 6.174 28.782 6.226 28.818 ;
        RECT 6.974 28.782 7.026 28.818 ;
        RECT 7.774 28.782 7.826 28.818 ;
        RECT 8.574 28.782 8.626 28.818 ;
        RECT 9.374 28.782 9.426 28.818 ;
        RECT 10.174 28.782 10.226 28.818 ;
        RECT 10.974 28.782 11.026 28.818 ;
        RECT 11.774 28.782 11.826 28.818 ;
        RECT 12.574 28.782 12.626 28.818 ;
        RECT 13.374 28.782 13.426 28.818 ;
        RECT 14.45 28.782 14.504 28.818 ;
        RECT 15.658 28.782 15.71 28.818 ;
        RECT 15.954 28.782 16.006 28.818 ;
        RECT 16.266 28.782 16.318 28.818 ;
        RECT 16.498 28.782 16.55 28.818 ;
        RECT 17.344 28.782 17.384 28.818 ;
        RECT 17.684 28.782 17.736 28.818 ;
        RECT 19.45 28.782 19.502 28.818 ;
        RECT 19.682 28.782 19.734 28.818 ;
        RECT 19.994 28.782 20.046 28.818 ;
        RECT 20.29 28.782 20.342 28.818 ;
        RECT 21.496 28.782 21.55 28.818 ;
        RECT 22.774 28.782 22.826 28.818 ;
        RECT 23.574 28.782 23.626 28.818 ;
        RECT 24.374 28.782 24.426 28.818 ;
        RECT 25.174 28.782 25.226 28.818 ;
        RECT 25.974 28.782 26.026 28.818 ;
        RECT 26.774 28.782 26.826 28.818 ;
        RECT 27.574 28.782 27.626 28.818 ;
        RECT 28.374 28.782 28.426 28.818 ;
        RECT 29.174 28.782 29.226 28.818 ;
        RECT 29.974 28.782 30.026 28.818 ;
        RECT 30.774 28.782 30.826 28.818 ;
        RECT 31.574 28.782 31.626 28.818 ;
        RECT 32.374 28.782 32.426 28.818 ;
        RECT 33.174 28.782 33.226 28.818 ;
        RECT 33.974 28.782 34.026 28.818 ;
        RECT 34.774 28.782 34.826 28.818 ;
        RECT 35.574 28.782 35.626 28.818 ;
        RECT 18.564 29.3875 18.636 29.4125 ;
        RECT 18.864 29.3875 18.936 29.4125 ;
        RECT 0.574 29.382 0.626 29.418 ;
        RECT 1.374 29.382 1.426 29.418 ;
        RECT 2.174 29.382 2.226 29.418 ;
        RECT 2.974 29.382 3.026 29.418 ;
        RECT 3.774 29.382 3.826 29.418 ;
        RECT 4.574 29.382 4.626 29.418 ;
        RECT 5.374 29.382 5.426 29.418 ;
        RECT 6.174 29.382 6.226 29.418 ;
        RECT 6.974 29.382 7.026 29.418 ;
        RECT 7.774 29.382 7.826 29.418 ;
        RECT 8.574 29.382 8.626 29.418 ;
        RECT 9.374 29.382 9.426 29.418 ;
        RECT 10.174 29.382 10.226 29.418 ;
        RECT 10.974 29.382 11.026 29.418 ;
        RECT 11.774 29.382 11.826 29.418 ;
        RECT 12.574 29.382 12.626 29.418 ;
        RECT 13.374 29.382 13.426 29.418 ;
        RECT 14.45 29.382 14.504 29.418 ;
        RECT 15.658 29.382 15.71 29.418 ;
        RECT 15.954 29.382 16.006 29.418 ;
        RECT 16.266 29.382 16.318 29.418 ;
        RECT 16.498 29.382 16.55 29.418 ;
        RECT 17.344 29.382 17.384 29.418 ;
        RECT 17.684 29.382 17.736 29.418 ;
        RECT 19.45 29.382 19.502 29.418 ;
        RECT 19.682 29.382 19.734 29.418 ;
        RECT 19.994 29.382 20.046 29.418 ;
        RECT 20.29 29.382 20.342 29.418 ;
        RECT 21.496 29.382 21.55 29.418 ;
        RECT 22.774 29.382 22.826 29.418 ;
        RECT 23.574 29.382 23.626 29.418 ;
        RECT 24.374 29.382 24.426 29.418 ;
        RECT 25.174 29.382 25.226 29.418 ;
        RECT 25.974 29.382 26.026 29.418 ;
        RECT 26.774 29.382 26.826 29.418 ;
        RECT 27.574 29.382 27.626 29.418 ;
        RECT 28.374 29.382 28.426 29.418 ;
        RECT 29.174 29.382 29.226 29.418 ;
        RECT 29.974 29.382 30.026 29.418 ;
        RECT 30.774 29.382 30.826 29.418 ;
        RECT 31.574 29.382 31.626 29.418 ;
        RECT 32.374 29.382 32.426 29.418 ;
        RECT 33.174 29.382 33.226 29.418 ;
        RECT 33.974 29.382 34.026 29.418 ;
        RECT 34.774 29.382 34.826 29.418 ;
        RECT 35.574 29.382 35.626 29.418 ;
        RECT 18.564 29.9875 18.636 30.0125 ;
        RECT 18.864 29.9875 18.936 30.0125 ;
        RECT 0.574 29.982 0.626 30.018 ;
        RECT 1.374 29.982 1.426 30.018 ;
        RECT 2.174 29.982 2.226 30.018 ;
        RECT 2.974 29.982 3.026 30.018 ;
        RECT 3.774 29.982 3.826 30.018 ;
        RECT 4.574 29.982 4.626 30.018 ;
        RECT 5.374 29.982 5.426 30.018 ;
        RECT 6.174 29.982 6.226 30.018 ;
        RECT 6.974 29.982 7.026 30.018 ;
        RECT 7.774 29.982 7.826 30.018 ;
        RECT 8.574 29.982 8.626 30.018 ;
        RECT 9.374 29.982 9.426 30.018 ;
        RECT 10.174 29.982 10.226 30.018 ;
        RECT 10.974 29.982 11.026 30.018 ;
        RECT 11.774 29.982 11.826 30.018 ;
        RECT 12.574 29.982 12.626 30.018 ;
        RECT 13.374 29.982 13.426 30.018 ;
        RECT 14.45 29.982 14.504 30.018 ;
        RECT 15.658 29.982 15.71 30.018 ;
        RECT 15.954 29.982 16.006 30.018 ;
        RECT 16.266 29.982 16.318 30.018 ;
        RECT 16.498 29.982 16.55 30.018 ;
        RECT 17.344 29.982 17.384 30.018 ;
        RECT 17.684 29.982 17.736 30.018 ;
        RECT 19.45 29.982 19.502 30.018 ;
        RECT 19.682 29.982 19.734 30.018 ;
        RECT 19.994 29.982 20.046 30.018 ;
        RECT 20.29 29.982 20.342 30.018 ;
        RECT 21.496 29.982 21.55 30.018 ;
        RECT 22.774 29.982 22.826 30.018 ;
        RECT 23.574 29.982 23.626 30.018 ;
        RECT 24.374 29.982 24.426 30.018 ;
        RECT 25.174 29.982 25.226 30.018 ;
        RECT 25.974 29.982 26.026 30.018 ;
        RECT 26.774 29.982 26.826 30.018 ;
        RECT 27.574 29.982 27.626 30.018 ;
        RECT 28.374 29.982 28.426 30.018 ;
        RECT 29.174 29.982 29.226 30.018 ;
        RECT 29.974 29.982 30.026 30.018 ;
        RECT 30.774 29.982 30.826 30.018 ;
        RECT 31.574 29.982 31.626 30.018 ;
        RECT 32.374 29.982 32.426 30.018 ;
        RECT 33.174 29.982 33.226 30.018 ;
        RECT 33.974 29.982 34.026 30.018 ;
        RECT 34.774 29.982 34.826 30.018 ;
        RECT 35.574 29.982 35.626 30.018 ;
        RECT 18.564 30.5875 18.636 30.6125 ;
        RECT 18.864 30.5875 18.936 30.6125 ;
        RECT 0.574 30.582 0.626 30.618 ;
        RECT 1.374 30.582 1.426 30.618 ;
        RECT 2.174 30.582 2.226 30.618 ;
        RECT 2.974 30.582 3.026 30.618 ;
        RECT 3.774 30.582 3.826 30.618 ;
        RECT 4.574 30.582 4.626 30.618 ;
        RECT 5.374 30.582 5.426 30.618 ;
        RECT 6.174 30.582 6.226 30.618 ;
        RECT 6.974 30.582 7.026 30.618 ;
        RECT 7.774 30.582 7.826 30.618 ;
        RECT 8.574 30.582 8.626 30.618 ;
        RECT 9.374 30.582 9.426 30.618 ;
        RECT 10.174 30.582 10.226 30.618 ;
        RECT 10.974 30.582 11.026 30.618 ;
        RECT 11.774 30.582 11.826 30.618 ;
        RECT 12.574 30.582 12.626 30.618 ;
        RECT 13.374 30.582 13.426 30.618 ;
        RECT 14.45 30.582 14.504 30.618 ;
        RECT 15.658 30.582 15.71 30.618 ;
        RECT 15.954 30.582 16.006 30.618 ;
        RECT 16.266 30.582 16.318 30.618 ;
        RECT 16.498 30.582 16.55 30.618 ;
        RECT 17.344 30.582 17.384 30.618 ;
        RECT 17.684 30.582 17.736 30.618 ;
        RECT 19.45 30.582 19.502 30.618 ;
        RECT 19.682 30.582 19.734 30.618 ;
        RECT 19.994 30.582 20.046 30.618 ;
        RECT 20.29 30.582 20.342 30.618 ;
        RECT 21.496 30.582 21.55 30.618 ;
        RECT 22.774 30.582 22.826 30.618 ;
        RECT 23.574 30.582 23.626 30.618 ;
        RECT 24.374 30.582 24.426 30.618 ;
        RECT 25.174 30.582 25.226 30.618 ;
        RECT 25.974 30.582 26.026 30.618 ;
        RECT 26.774 30.582 26.826 30.618 ;
        RECT 27.574 30.582 27.626 30.618 ;
        RECT 28.374 30.582 28.426 30.618 ;
        RECT 29.174 30.582 29.226 30.618 ;
        RECT 29.974 30.582 30.026 30.618 ;
        RECT 30.774 30.582 30.826 30.618 ;
        RECT 31.574 30.582 31.626 30.618 ;
        RECT 32.374 30.582 32.426 30.618 ;
        RECT 33.174 30.582 33.226 30.618 ;
        RECT 33.974 30.582 34.026 30.618 ;
        RECT 34.774 30.582 34.826 30.618 ;
        RECT 35.574 30.582 35.626 30.618 ;
        RECT 18.564 31.1875 18.636 31.2125 ;
        RECT 18.864 31.1875 18.936 31.2125 ;
        RECT 0.574 31.182 0.626 31.218 ;
        RECT 1.374 31.182 1.426 31.218 ;
        RECT 2.174 31.182 2.226 31.218 ;
        RECT 2.974 31.182 3.026 31.218 ;
        RECT 3.774 31.182 3.826 31.218 ;
        RECT 4.574 31.182 4.626 31.218 ;
        RECT 5.374 31.182 5.426 31.218 ;
        RECT 6.174 31.182 6.226 31.218 ;
        RECT 6.974 31.182 7.026 31.218 ;
        RECT 7.774 31.182 7.826 31.218 ;
        RECT 8.574 31.182 8.626 31.218 ;
        RECT 9.374 31.182 9.426 31.218 ;
        RECT 10.174 31.182 10.226 31.218 ;
        RECT 10.974 31.182 11.026 31.218 ;
        RECT 11.774 31.182 11.826 31.218 ;
        RECT 12.574 31.182 12.626 31.218 ;
        RECT 13.374 31.182 13.426 31.218 ;
        RECT 14.45 31.182 14.504 31.218 ;
        RECT 15.658 31.182 15.71 31.218 ;
        RECT 15.954 31.182 16.006 31.218 ;
        RECT 16.266 31.182 16.318 31.218 ;
        RECT 16.498 31.182 16.55 31.218 ;
        RECT 17.344 31.182 17.384 31.218 ;
        RECT 17.684 31.182 17.736 31.218 ;
        RECT 19.45 31.182 19.502 31.218 ;
        RECT 19.682 31.182 19.734 31.218 ;
        RECT 19.994 31.182 20.046 31.218 ;
        RECT 20.29 31.182 20.342 31.218 ;
        RECT 21.496 31.182 21.55 31.218 ;
        RECT 22.774 31.182 22.826 31.218 ;
        RECT 23.574 31.182 23.626 31.218 ;
        RECT 24.374 31.182 24.426 31.218 ;
        RECT 25.174 31.182 25.226 31.218 ;
        RECT 25.974 31.182 26.026 31.218 ;
        RECT 26.774 31.182 26.826 31.218 ;
        RECT 27.574 31.182 27.626 31.218 ;
        RECT 28.374 31.182 28.426 31.218 ;
        RECT 29.174 31.182 29.226 31.218 ;
        RECT 29.974 31.182 30.026 31.218 ;
        RECT 30.774 31.182 30.826 31.218 ;
        RECT 31.574 31.182 31.626 31.218 ;
        RECT 32.374 31.182 32.426 31.218 ;
        RECT 33.174 31.182 33.226 31.218 ;
        RECT 33.974 31.182 34.026 31.218 ;
        RECT 34.774 31.182 34.826 31.218 ;
        RECT 35.574 31.182 35.626 31.218 ;
        RECT 18.564 31.7875 18.636 31.8125 ;
        RECT 18.864 31.7875 18.936 31.8125 ;
        RECT 0.574 31.782 0.626 31.818 ;
        RECT 1.374 31.782 1.426 31.818 ;
        RECT 2.174 31.782 2.226 31.818 ;
        RECT 2.974 31.782 3.026 31.818 ;
        RECT 3.774 31.782 3.826 31.818 ;
        RECT 4.574 31.782 4.626 31.818 ;
        RECT 5.374 31.782 5.426 31.818 ;
        RECT 6.174 31.782 6.226 31.818 ;
        RECT 6.974 31.782 7.026 31.818 ;
        RECT 7.774 31.782 7.826 31.818 ;
        RECT 8.574 31.782 8.626 31.818 ;
        RECT 9.374 31.782 9.426 31.818 ;
        RECT 10.174 31.782 10.226 31.818 ;
        RECT 10.974 31.782 11.026 31.818 ;
        RECT 11.774 31.782 11.826 31.818 ;
        RECT 12.574 31.782 12.626 31.818 ;
        RECT 13.374 31.782 13.426 31.818 ;
        RECT 14.45 31.782 14.504 31.818 ;
        RECT 15.658 31.782 15.71 31.818 ;
        RECT 15.954 31.782 16.006 31.818 ;
        RECT 16.266 31.782 16.318 31.818 ;
        RECT 16.498 31.782 16.55 31.818 ;
        RECT 17.344 31.782 17.384 31.818 ;
        RECT 17.684 31.782 17.736 31.818 ;
        RECT 19.45 31.782 19.502 31.818 ;
        RECT 19.682 31.782 19.734 31.818 ;
        RECT 19.994 31.782 20.046 31.818 ;
        RECT 20.29 31.782 20.342 31.818 ;
        RECT 21.496 31.782 21.55 31.818 ;
        RECT 22.774 31.782 22.826 31.818 ;
        RECT 23.574 31.782 23.626 31.818 ;
        RECT 24.374 31.782 24.426 31.818 ;
        RECT 25.174 31.782 25.226 31.818 ;
        RECT 25.974 31.782 26.026 31.818 ;
        RECT 26.774 31.782 26.826 31.818 ;
        RECT 27.574 31.782 27.626 31.818 ;
        RECT 28.374 31.782 28.426 31.818 ;
        RECT 29.174 31.782 29.226 31.818 ;
        RECT 29.974 31.782 30.026 31.818 ;
        RECT 30.774 31.782 30.826 31.818 ;
        RECT 31.574 31.782 31.626 31.818 ;
        RECT 32.374 31.782 32.426 31.818 ;
        RECT 33.174 31.782 33.226 31.818 ;
        RECT 33.974 31.782 34.026 31.818 ;
        RECT 34.774 31.782 34.826 31.818 ;
        RECT 35.574 31.782 35.626 31.818 ;
        RECT 13.374 32.1475 13.426 32.1725 ;
        RECT 18.564 32.1475 18.636 32.1725 ;
        RECT 18.864 32.1475 18.936 32.1725 ;
        RECT 35.574 32.1475 35.626 32.1725 ;
        RECT 0.574 32.142 0.626 32.178 ;
        RECT 1.374 32.142 1.426 32.178 ;
        RECT 2.174 32.142 2.226 32.178 ;
        RECT 2.974 32.142 3.026 32.178 ;
        RECT 3.774 32.142 3.826 32.178 ;
        RECT 4.574 32.142 4.626 32.178 ;
        RECT 5.374 32.142 5.426 32.178 ;
        RECT 6.174 32.142 6.226 32.178 ;
        RECT 6.974 32.142 7.026 32.178 ;
        RECT 7.774 32.142 7.826 32.178 ;
        RECT 8.574 32.142 8.626 32.178 ;
        RECT 9.374 32.142 9.426 32.178 ;
        RECT 10.174 32.142 10.226 32.178 ;
        RECT 10.974 32.142 11.026 32.178 ;
        RECT 11.774 32.142 11.826 32.178 ;
        RECT 12.574 32.142 12.626 32.178 ;
        RECT 14.45 32.142 14.504 32.178 ;
        RECT 15.658 32.142 15.71 32.178 ;
        RECT 15.954 32.142 16.006 32.178 ;
        RECT 16.266 32.142 16.318 32.178 ;
        RECT 16.498 32.142 16.55 32.178 ;
        RECT 17.204 32.142 17.244 32.178 ;
        RECT 17.684 32.142 17.736 32.178 ;
        RECT 18.216 32.142 18.256 32.178 ;
        RECT 19.228 32.142 19.282 32.178 ;
        RECT 19.45 32.142 19.502 32.178 ;
        RECT 19.682 32.142 19.734 32.178 ;
        RECT 19.994 32.142 20.046 32.178 ;
        RECT 20.29 32.142 20.342 32.178 ;
        RECT 21.496 32.142 21.55 32.178 ;
        RECT 22.774 32.142 22.826 32.178 ;
        RECT 23.574 32.142 23.626 32.178 ;
        RECT 24.374 32.142 24.426 32.178 ;
        RECT 25.174 32.142 25.226 32.178 ;
        RECT 25.974 32.142 26.026 32.178 ;
        RECT 26.774 32.142 26.826 32.178 ;
        RECT 27.574 32.142 27.626 32.178 ;
        RECT 28.374 32.142 28.426 32.178 ;
        RECT 29.174 32.142 29.226 32.178 ;
        RECT 29.974 32.142 30.026 32.178 ;
        RECT 30.774 32.142 30.826 32.178 ;
        RECT 31.574 32.142 31.626 32.178 ;
        RECT 32.374 32.142 32.426 32.178 ;
        RECT 33.174 32.142 33.226 32.178 ;
        RECT 33.974 32.142 34.026 32.178 ;
        RECT 34.774 32.142 34.826 32.178 ;
        RECT 0.574 32.382 0.626 32.418 ;
        RECT 1.374 32.382 1.426 32.418 ;
        RECT 2.174 32.382 2.226 32.418 ;
        RECT 2.974 32.382 3.026 32.418 ;
        RECT 3.774 32.382 3.826 32.418 ;
        RECT 4.574 32.382 4.626 32.418 ;
        RECT 5.374 32.382 5.426 32.418 ;
        RECT 6.174 32.382 6.226 32.418 ;
        RECT 6.974 32.382 7.026 32.418 ;
        RECT 7.774 32.382 7.826 32.418 ;
        RECT 8.574 32.382 8.626 32.418 ;
        RECT 9.374 32.382 9.426 32.418 ;
        RECT 10.174 32.382 10.226 32.418 ;
        RECT 10.974 32.382 11.026 32.418 ;
        RECT 11.774 32.382 11.826 32.418 ;
        RECT 12.574 32.382 12.626 32.418 ;
        RECT 13.374 32.382 13.426 32.418 ;
        RECT 22.774 32.382 22.826 32.418 ;
        RECT 23.574 32.382 23.626 32.418 ;
        RECT 24.374 32.382 24.426 32.418 ;
        RECT 25.174 32.382 25.226 32.418 ;
        RECT 25.974 32.382 26.026 32.418 ;
        RECT 26.774 32.382 26.826 32.418 ;
        RECT 27.574 32.382 27.626 32.418 ;
        RECT 28.374 32.382 28.426 32.418 ;
        RECT 29.174 32.382 29.226 32.418 ;
        RECT 29.974 32.382 30.026 32.418 ;
        RECT 30.774 32.382 30.826 32.418 ;
        RECT 31.574 32.382 31.626 32.418 ;
        RECT 32.374 32.382 32.426 32.418 ;
        RECT 33.174 32.382 33.226 32.418 ;
        RECT 33.974 32.382 34.026 32.418 ;
        RECT 34.774 32.382 34.826 32.418 ;
        RECT 35.574 32.382 35.626 32.418 ;
        RECT 18.564 32.6275 18.636 32.6525 ;
        RECT 18.864 32.6275 18.936 32.6525 ;
        RECT 14.45 32.622 14.504 32.658 ;
        RECT 15.658 32.622 15.71 32.658 ;
        RECT 15.954 32.622 16.006 32.658 ;
        RECT 16.498 32.622 16.55 32.658 ;
        RECT 16.882 32.622 16.936 32.658 ;
        RECT 17.204 32.622 17.244 32.658 ;
        RECT 17.684 32.622 17.736 32.658 ;
        RECT 18.216 32.622 18.256 32.658 ;
        RECT 19.228 32.622 19.282 32.658 ;
        RECT 19.45 32.622 19.502 32.658 ;
        RECT 19.682 32.622 19.734 32.658 ;
        RECT 19.994 32.622 20.046 32.658 ;
        RECT 20.29 32.622 20.342 32.658 ;
        RECT 21.496 32.622 21.55 32.658 ;
        RECT 17.204 32.9205 17.244 32.9565 ;
        RECT 17.684 32.9205 17.736 32.9565 ;
        RECT 19.45 32.9205 19.502 32.9565 ;
        RECT 19.682 32.9205 19.734 32.9565 ;
        RECT 20.29 32.9205 20.342 32.9565 ;
        RECT 18.864 33.1075 18.936 33.1325 ;
        RECT 0.574 33.102 0.626 33.138 ;
        RECT 1.374 33.102 1.426 33.138 ;
        RECT 2.174 33.102 2.226 33.138 ;
        RECT 2.974 33.102 3.026 33.138 ;
        RECT 3.774 33.102 3.826 33.138 ;
        RECT 4.574 33.102 4.626 33.138 ;
        RECT 5.374 33.102 5.426 33.138 ;
        RECT 6.174 33.102 6.226 33.138 ;
        RECT 6.974 33.102 7.026 33.138 ;
        RECT 7.774 33.102 7.826 33.138 ;
        RECT 8.574 33.102 8.626 33.138 ;
        RECT 9.374 33.102 9.426 33.138 ;
        RECT 10.174 33.102 10.226 33.138 ;
        RECT 10.974 33.102 11.026 33.138 ;
        RECT 11.774 33.102 11.826 33.138 ;
        RECT 12.574 33.102 12.626 33.138 ;
        RECT 13.374 33.102 13.426 33.138 ;
        RECT 14.45 33.102 14.504 33.138 ;
        RECT 15.658 33.102 15.71 33.138 ;
        RECT 15.954 33.102 16.006 33.138 ;
        RECT 16.266 33.102 16.318 33.138 ;
        RECT 16.498 33.102 16.55 33.138 ;
        RECT 17.204 33.102 17.244 33.138 ;
        RECT 17.684 33.102 17.736 33.138 ;
        RECT 18.216 33.102 18.256 33.138 ;
        RECT 19.228 33.102 19.282 33.138 ;
        RECT 19.45 33.102 19.502 33.138 ;
        RECT 19.682 33.102 19.734 33.138 ;
        RECT 19.994 33.102 20.046 33.138 ;
        RECT 20.29 33.102 20.342 33.138 ;
        RECT 21.496 33.102 21.55 33.138 ;
        RECT 22.774 33.102 22.826 33.138 ;
        RECT 23.574 33.102 23.626 33.138 ;
        RECT 24.374 33.102 24.426 33.138 ;
        RECT 25.174 33.102 25.226 33.138 ;
        RECT 25.974 33.102 26.026 33.138 ;
        RECT 26.774 33.102 26.826 33.138 ;
        RECT 27.574 33.102 27.626 33.138 ;
        RECT 28.374 33.102 28.426 33.138 ;
        RECT 29.174 33.102 29.226 33.138 ;
        RECT 29.974 33.102 30.026 33.138 ;
        RECT 30.774 33.102 30.826 33.138 ;
        RECT 31.574 33.102 31.626 33.138 ;
        RECT 32.374 33.102 32.426 33.138 ;
        RECT 33.174 33.102 33.226 33.138 ;
        RECT 33.974 33.102 34.026 33.138 ;
        RECT 34.774 33.102 34.826 33.138 ;
        RECT 35.574 33.102 35.626 33.138 ;
        RECT 14.45 33.2835 14.504 33.3195 ;
        RECT 21.496 33.2835 21.55 33.3195 ;
        RECT 16.882 33.5875 16.936 33.6125 ;
        RECT 18.564 33.5875 18.636 33.6125 ;
        RECT 18.864 33.5875 18.936 33.6125 ;
        RECT 14.45 33.582 14.504 33.618 ;
        RECT 15.658 33.582 15.71 33.618 ;
        RECT 15.954 33.582 16.006 33.618 ;
        RECT 16.266 33.582 16.318 33.618 ;
        RECT 16.498 33.582 16.55 33.618 ;
        RECT 17.204 33.582 17.244 33.618 ;
        RECT 17.684 33.582 17.736 33.618 ;
        RECT 18.216 33.582 18.256 33.618 ;
        RECT 19.228 33.582 19.282 33.618 ;
        RECT 19.45 33.582 19.502 33.618 ;
        RECT 19.682 33.582 19.734 33.618 ;
        RECT 19.994 33.582 20.046 33.618 ;
        RECT 20.29 33.582 20.342 33.618 ;
        RECT 21.496 33.582 21.55 33.618 ;
        RECT 0.574 33.822 0.626 33.858 ;
        RECT 1.374 33.822 1.426 33.858 ;
        RECT 2.174 33.822 2.226 33.858 ;
        RECT 2.974 33.822 3.026 33.858 ;
        RECT 3.774 33.822 3.826 33.858 ;
        RECT 4.574 33.822 4.626 33.858 ;
        RECT 5.374 33.822 5.426 33.858 ;
        RECT 6.174 33.822 6.226 33.858 ;
        RECT 6.974 33.822 7.026 33.858 ;
        RECT 7.774 33.822 7.826 33.858 ;
        RECT 8.574 33.822 8.626 33.858 ;
        RECT 9.374 33.822 9.426 33.858 ;
        RECT 10.174 33.822 10.226 33.858 ;
        RECT 10.974 33.822 11.026 33.858 ;
        RECT 11.774 33.822 11.826 33.858 ;
        RECT 12.574 33.822 12.626 33.858 ;
        RECT 13.374 33.822 13.426 33.858 ;
        RECT 22.774 33.822 22.826 33.858 ;
        RECT 23.574 33.822 23.626 33.858 ;
        RECT 24.374 33.822 24.426 33.858 ;
        RECT 25.174 33.822 25.226 33.858 ;
        RECT 25.974 33.822 26.026 33.858 ;
        RECT 26.774 33.822 26.826 33.858 ;
        RECT 27.574 33.822 27.626 33.858 ;
        RECT 28.374 33.822 28.426 33.858 ;
        RECT 29.174 33.822 29.226 33.858 ;
        RECT 29.974 33.822 30.026 33.858 ;
        RECT 30.774 33.822 30.826 33.858 ;
        RECT 31.574 33.822 31.626 33.858 ;
        RECT 32.374 33.822 32.426 33.858 ;
        RECT 33.174 33.822 33.226 33.858 ;
        RECT 33.974 33.822 34.026 33.858 ;
        RECT 34.774 33.822 34.826 33.858 ;
        RECT 35.574 33.822 35.626 33.858 ;
        RECT 18.564 34.0675 18.636 34.0925 ;
        RECT 18.864 34.0675 18.936 34.0925 ;
        RECT 0.574 34.062 0.626 34.098 ;
        RECT 1.374 34.062 1.426 34.098 ;
        RECT 2.174 34.062 2.226 34.098 ;
        RECT 2.974 34.062 3.026 34.098 ;
        RECT 3.774 34.062 3.826 34.098 ;
        RECT 4.574 34.062 4.626 34.098 ;
        RECT 5.374 34.062 5.426 34.098 ;
        RECT 6.174 34.062 6.226 34.098 ;
        RECT 6.974 34.062 7.026 34.098 ;
        RECT 7.774 34.062 7.826 34.098 ;
        RECT 8.574 34.062 8.626 34.098 ;
        RECT 9.374 34.062 9.426 34.098 ;
        RECT 10.174 34.062 10.226 34.098 ;
        RECT 10.974 34.062 11.026 34.098 ;
        RECT 11.774 34.062 11.826 34.098 ;
        RECT 12.574 34.062 12.626 34.098 ;
        RECT 13.374 34.062 13.426 34.098 ;
        RECT 14.45 34.062 14.504 34.098 ;
        RECT 15.658 34.062 15.71 34.098 ;
        RECT 15.954 34.062 16.006 34.098 ;
        RECT 16.266 34.062 16.318 34.098 ;
        RECT 16.498 34.062 16.55 34.098 ;
        RECT 16.882 34.062 16.936 34.098 ;
        RECT 17.204 34.062 17.244 34.098 ;
        RECT 17.684 34.062 17.736 34.098 ;
        RECT 18.216 34.062 18.256 34.098 ;
        RECT 19.228 34.062 19.282 34.098 ;
        RECT 19.45 34.062 19.502 34.098 ;
        RECT 19.682 34.062 19.734 34.098 ;
        RECT 19.994 34.062 20.046 34.098 ;
        RECT 20.29 34.062 20.342 34.098 ;
        RECT 21.496 34.062 21.55 34.098 ;
        RECT 22.774 34.062 22.826 34.098 ;
        RECT 23.574 34.062 23.626 34.098 ;
        RECT 24.374 34.062 24.426 34.098 ;
        RECT 25.174 34.062 25.226 34.098 ;
        RECT 25.974 34.062 26.026 34.098 ;
        RECT 26.774 34.062 26.826 34.098 ;
        RECT 27.574 34.062 27.626 34.098 ;
        RECT 28.374 34.062 28.426 34.098 ;
        RECT 29.174 34.062 29.226 34.098 ;
        RECT 29.974 34.062 30.026 34.098 ;
        RECT 30.774 34.062 30.826 34.098 ;
        RECT 31.574 34.062 31.626 34.098 ;
        RECT 32.374 34.062 32.426 34.098 ;
        RECT 33.174 34.062 33.226 34.098 ;
        RECT 33.974 34.062 34.026 34.098 ;
        RECT 34.774 34.062 34.826 34.098 ;
        RECT 35.574 34.062 35.626 34.098 ;
        RECT 16.882 34.5475 16.936 34.5725 ;
        RECT 18.564 34.5475 18.636 34.5725 ;
        RECT 18.864 34.5475 18.936 34.5725 ;
        RECT 0.574 34.542 0.626 34.578 ;
        RECT 1.374 34.542 1.426 34.578 ;
        RECT 2.174 34.542 2.226 34.578 ;
        RECT 2.974 34.542 3.026 34.578 ;
        RECT 3.774 34.542 3.826 34.578 ;
        RECT 4.574 34.542 4.626 34.578 ;
        RECT 5.374 34.542 5.426 34.578 ;
        RECT 6.174 34.542 6.226 34.578 ;
        RECT 6.974 34.542 7.026 34.578 ;
        RECT 7.774 34.542 7.826 34.578 ;
        RECT 8.574 34.542 8.626 34.578 ;
        RECT 9.374 34.542 9.426 34.578 ;
        RECT 10.174 34.542 10.226 34.578 ;
        RECT 10.974 34.542 11.026 34.578 ;
        RECT 11.774 34.542 11.826 34.578 ;
        RECT 12.574 34.542 12.626 34.578 ;
        RECT 13.374 34.542 13.426 34.578 ;
        RECT 14.45 34.542 14.504 34.578 ;
        RECT 15.658 34.542 15.71 34.578 ;
        RECT 15.954 34.542 16.006 34.578 ;
        RECT 16.266 34.542 16.318 34.578 ;
        RECT 16.498 34.542 16.55 34.578 ;
        RECT 17.204 34.542 17.244 34.578 ;
        RECT 17.684 34.542 17.736 34.578 ;
        RECT 18.216 34.542 18.256 34.578 ;
        RECT 19.228 34.542 19.282 34.578 ;
        RECT 19.45 34.542 19.502 34.578 ;
        RECT 19.682 34.542 19.734 34.578 ;
        RECT 19.994 34.542 20.046 34.578 ;
        RECT 20.29 34.542 20.342 34.578 ;
        RECT 21.496 34.542 21.55 34.578 ;
        RECT 22.774 34.542 22.826 34.578 ;
        RECT 23.574 34.542 23.626 34.578 ;
        RECT 24.374 34.542 24.426 34.578 ;
        RECT 25.174 34.542 25.226 34.578 ;
        RECT 25.974 34.542 26.026 34.578 ;
        RECT 26.774 34.542 26.826 34.578 ;
        RECT 27.574 34.542 27.626 34.578 ;
        RECT 28.374 34.542 28.426 34.578 ;
        RECT 29.174 34.542 29.226 34.578 ;
        RECT 29.974 34.542 30.026 34.578 ;
        RECT 30.774 34.542 30.826 34.578 ;
        RECT 31.574 34.542 31.626 34.578 ;
        RECT 32.374 34.542 32.426 34.578 ;
        RECT 33.174 34.542 33.226 34.578 ;
        RECT 33.974 34.542 34.026 34.578 ;
        RECT 34.774 34.542 34.826 34.578 ;
        RECT 35.574 34.542 35.626 34.578 ;
        RECT 18.564 35.0275 18.636 35.0525 ;
        RECT 18.864 35.0275 18.936 35.0525 ;
        RECT 0.574 35.022 0.626 35.058 ;
        RECT 1.374 35.022 1.426 35.058 ;
        RECT 2.174 35.022 2.226 35.058 ;
        RECT 2.974 35.022 3.026 35.058 ;
        RECT 3.774 35.022 3.826 35.058 ;
        RECT 4.574 35.022 4.626 35.058 ;
        RECT 5.374 35.022 5.426 35.058 ;
        RECT 6.174 35.022 6.226 35.058 ;
        RECT 6.974 35.022 7.026 35.058 ;
        RECT 7.774 35.022 7.826 35.058 ;
        RECT 8.574 35.022 8.626 35.058 ;
        RECT 9.374 35.022 9.426 35.058 ;
        RECT 10.174 35.022 10.226 35.058 ;
        RECT 10.974 35.022 11.026 35.058 ;
        RECT 11.774 35.022 11.826 35.058 ;
        RECT 12.574 35.022 12.626 35.058 ;
        RECT 13.374 35.022 13.426 35.058 ;
        RECT 14.45 35.022 14.504 35.058 ;
        RECT 15.658 35.022 15.71 35.058 ;
        RECT 15.954 35.022 16.006 35.058 ;
        RECT 16.266 35.022 16.318 35.058 ;
        RECT 16.498 35.022 16.55 35.058 ;
        RECT 16.882 35.022 16.936 35.058 ;
        RECT 17.204 35.022 17.244 35.058 ;
        RECT 17.684 35.022 17.736 35.058 ;
        RECT 18.216 35.022 18.256 35.058 ;
        RECT 19.228 35.022 19.282 35.058 ;
        RECT 19.45 35.022 19.502 35.058 ;
        RECT 19.682 35.022 19.734 35.058 ;
        RECT 19.994 35.022 20.046 35.058 ;
        RECT 20.29 35.022 20.342 35.058 ;
        RECT 21.496 35.022 21.55 35.058 ;
        RECT 22.774 35.022 22.826 35.058 ;
        RECT 23.574 35.022 23.626 35.058 ;
        RECT 24.374 35.022 24.426 35.058 ;
        RECT 25.174 35.022 25.226 35.058 ;
        RECT 25.974 35.022 26.026 35.058 ;
        RECT 26.774 35.022 26.826 35.058 ;
        RECT 27.574 35.022 27.626 35.058 ;
        RECT 28.374 35.022 28.426 35.058 ;
        RECT 29.174 35.022 29.226 35.058 ;
        RECT 29.974 35.022 30.026 35.058 ;
        RECT 30.774 35.022 30.826 35.058 ;
        RECT 31.574 35.022 31.626 35.058 ;
        RECT 32.374 35.022 32.426 35.058 ;
        RECT 33.174 35.022 33.226 35.058 ;
        RECT 33.974 35.022 34.026 35.058 ;
        RECT 34.774 35.022 34.826 35.058 ;
        RECT 35.574 35.022 35.626 35.058 ;
        RECT 16.882 35.5075 16.936 35.5325 ;
        RECT 18.564 35.5075 18.636 35.5325 ;
        RECT 18.864 35.5075 18.936 35.5325 ;
        RECT 0.574 35.502 0.626 35.538 ;
        RECT 1.374 35.502 1.426 35.538 ;
        RECT 2.174 35.502 2.226 35.538 ;
        RECT 2.974 35.502 3.026 35.538 ;
        RECT 3.774 35.502 3.826 35.538 ;
        RECT 4.574 35.502 4.626 35.538 ;
        RECT 5.374 35.502 5.426 35.538 ;
        RECT 6.174 35.502 6.226 35.538 ;
        RECT 6.974 35.502 7.026 35.538 ;
        RECT 7.774 35.502 7.826 35.538 ;
        RECT 8.574 35.502 8.626 35.538 ;
        RECT 9.374 35.502 9.426 35.538 ;
        RECT 10.174 35.502 10.226 35.538 ;
        RECT 10.974 35.502 11.026 35.538 ;
        RECT 11.774 35.502 11.826 35.538 ;
        RECT 12.574 35.502 12.626 35.538 ;
        RECT 13.374 35.502 13.426 35.538 ;
        RECT 14.45 35.502 14.504 35.538 ;
        RECT 15.658 35.502 15.71 35.538 ;
        RECT 15.954 35.502 16.006 35.538 ;
        RECT 16.266 35.502 16.318 35.538 ;
        RECT 16.498 35.502 16.55 35.538 ;
        RECT 17.204 35.502 17.244 35.538 ;
        RECT 17.684 35.502 17.736 35.538 ;
        RECT 18.216 35.502 18.256 35.538 ;
        RECT 19.228 35.502 19.282 35.538 ;
        RECT 19.45 35.502 19.502 35.538 ;
        RECT 19.682 35.502 19.734 35.538 ;
        RECT 19.994 35.502 20.046 35.538 ;
        RECT 20.29 35.502 20.342 35.538 ;
        RECT 21.496 35.502 21.55 35.538 ;
        RECT 22.774 35.502 22.826 35.538 ;
        RECT 23.574 35.502 23.626 35.538 ;
        RECT 24.374 35.502 24.426 35.538 ;
        RECT 25.174 35.502 25.226 35.538 ;
        RECT 25.974 35.502 26.026 35.538 ;
        RECT 26.774 35.502 26.826 35.538 ;
        RECT 27.574 35.502 27.626 35.538 ;
        RECT 28.374 35.502 28.426 35.538 ;
        RECT 29.174 35.502 29.226 35.538 ;
        RECT 29.974 35.502 30.026 35.538 ;
        RECT 30.774 35.502 30.826 35.538 ;
        RECT 31.574 35.502 31.626 35.538 ;
        RECT 32.374 35.502 32.426 35.538 ;
        RECT 33.174 35.502 33.226 35.538 ;
        RECT 33.974 35.502 34.026 35.538 ;
        RECT 34.774 35.502 34.826 35.538 ;
        RECT 35.574 35.502 35.626 35.538 ;
        RECT 18.564 35.8675 18.636 35.8925 ;
        RECT 18.864 35.8675 18.936 35.8925 ;
        RECT 14.45 35.862 14.504 35.898 ;
        RECT 15.658 35.862 15.71 35.898 ;
        RECT 15.954 35.862 16.006 35.898 ;
        RECT 16.266 35.862 16.318 35.898 ;
        RECT 16.498 35.862 16.55 35.898 ;
        RECT 16.882 35.862 16.936 35.898 ;
        RECT 17.204 35.862 17.244 35.898 ;
        RECT 18.216 35.862 18.256 35.898 ;
        RECT 19.228 35.862 19.282 35.898 ;
        RECT 19.45 35.862 19.502 35.898 ;
        RECT 19.994 35.862 20.046 35.898 ;
        RECT 20.29 35.862 20.342 35.898 ;
        RECT 21.496 35.862 21.55 35.898 ;
        RECT 18.564 35.9875 18.636 36.0125 ;
        RECT 18.864 35.9875 18.936 36.0125 ;
        RECT 0.574 35.982 0.626 36.018 ;
        RECT 1.374 35.982 1.426 36.018 ;
        RECT 2.174 35.982 2.226 36.018 ;
        RECT 2.974 35.982 3.026 36.018 ;
        RECT 3.774 35.982 3.826 36.018 ;
        RECT 4.574 35.982 4.626 36.018 ;
        RECT 5.374 35.982 5.426 36.018 ;
        RECT 6.174 35.982 6.226 36.018 ;
        RECT 6.974 35.982 7.026 36.018 ;
        RECT 7.774 35.982 7.826 36.018 ;
        RECT 8.574 35.982 8.626 36.018 ;
        RECT 9.374 35.982 9.426 36.018 ;
        RECT 10.174 35.982 10.226 36.018 ;
        RECT 10.974 35.982 11.026 36.018 ;
        RECT 11.774 35.982 11.826 36.018 ;
        RECT 12.574 35.982 12.626 36.018 ;
        RECT 13.374 35.982 13.426 36.018 ;
        RECT 14.45 35.982 14.504 36.018 ;
        RECT 15.658 35.982 15.71 36.018 ;
        RECT 15.954 35.982 16.006 36.018 ;
        RECT 16.266 35.982 16.318 36.018 ;
        RECT 16.498 35.982 16.55 36.018 ;
        RECT 16.882 35.982 16.936 36.018 ;
        RECT 17.204 35.982 17.244 36.018 ;
        RECT 17.684 35.982 17.736 36.018 ;
        RECT 18.216 35.982 18.256 36.018 ;
        RECT 19.228 35.982 19.282 36.018 ;
        RECT 19.45 35.982 19.502 36.018 ;
        RECT 19.682 35.982 19.734 36.018 ;
        RECT 19.994 35.982 20.046 36.018 ;
        RECT 20.29 35.982 20.342 36.018 ;
        RECT 21.496 35.982 21.55 36.018 ;
        RECT 22.774 35.982 22.826 36.018 ;
        RECT 23.574 35.982 23.626 36.018 ;
        RECT 24.374 35.982 24.426 36.018 ;
        RECT 25.174 35.982 25.226 36.018 ;
        RECT 25.974 35.982 26.026 36.018 ;
        RECT 26.774 35.982 26.826 36.018 ;
        RECT 27.574 35.982 27.626 36.018 ;
        RECT 28.374 35.982 28.426 36.018 ;
        RECT 29.174 35.982 29.226 36.018 ;
        RECT 29.974 35.982 30.026 36.018 ;
        RECT 30.774 35.982 30.826 36.018 ;
        RECT 31.574 35.982 31.626 36.018 ;
        RECT 32.374 35.982 32.426 36.018 ;
        RECT 33.174 35.982 33.226 36.018 ;
        RECT 33.974 35.982 34.026 36.018 ;
        RECT 34.774 35.982 34.826 36.018 ;
        RECT 35.574 35.982 35.626 36.018 ;
        RECT 15.954 36.4675 16.006 36.4925 ;
        RECT 18.564 36.4675 18.636 36.4925 ;
        RECT 18.864 36.4675 18.936 36.4925 ;
        RECT 19.994 36.4675 20.046 36.4925 ;
        RECT 0.574 36.462 0.626 36.498 ;
        RECT 1.374 36.462 1.426 36.498 ;
        RECT 2.174 36.462 2.226 36.498 ;
        RECT 2.974 36.462 3.026 36.498 ;
        RECT 3.774 36.462 3.826 36.498 ;
        RECT 4.574 36.462 4.626 36.498 ;
        RECT 5.374 36.462 5.426 36.498 ;
        RECT 6.174 36.462 6.226 36.498 ;
        RECT 6.974 36.462 7.026 36.498 ;
        RECT 7.774 36.462 7.826 36.498 ;
        RECT 8.574 36.462 8.626 36.498 ;
        RECT 9.374 36.462 9.426 36.498 ;
        RECT 10.174 36.462 10.226 36.498 ;
        RECT 10.974 36.462 11.026 36.498 ;
        RECT 11.774 36.462 11.826 36.498 ;
        RECT 12.574 36.462 12.626 36.498 ;
        RECT 13.374 36.462 13.426 36.498 ;
        RECT 14.45 36.462 14.504 36.498 ;
        RECT 15.658 36.462 15.71 36.498 ;
        RECT 16.266 36.462 16.318 36.498 ;
        RECT 16.498 36.462 16.55 36.498 ;
        RECT 16.882 36.462 16.936 36.498 ;
        RECT 17.204 36.462 17.244 36.498 ;
        RECT 17.684 36.462 17.736 36.498 ;
        RECT 18.216 36.462 18.256 36.498 ;
        RECT 19.228 36.462 19.282 36.498 ;
        RECT 19.45 36.462 19.502 36.498 ;
        RECT 19.682 36.462 19.734 36.498 ;
        RECT 20.29 36.462 20.342 36.498 ;
        RECT 21.496 36.462 21.55 36.498 ;
        RECT 22.774 36.462 22.826 36.498 ;
        RECT 23.574 36.462 23.626 36.498 ;
        RECT 24.374 36.462 24.426 36.498 ;
        RECT 25.174 36.462 25.226 36.498 ;
        RECT 25.974 36.462 26.026 36.498 ;
        RECT 26.774 36.462 26.826 36.498 ;
        RECT 27.574 36.462 27.626 36.498 ;
        RECT 28.374 36.462 28.426 36.498 ;
        RECT 29.174 36.462 29.226 36.498 ;
        RECT 29.974 36.462 30.026 36.498 ;
        RECT 30.774 36.462 30.826 36.498 ;
        RECT 31.574 36.462 31.626 36.498 ;
        RECT 32.374 36.462 32.426 36.498 ;
        RECT 33.174 36.462 33.226 36.498 ;
        RECT 33.974 36.462 34.026 36.498 ;
        RECT 34.774 36.462 34.826 36.498 ;
        RECT 35.574 36.462 35.626 36.498 ;
        RECT 16.882 36.9475 16.936 36.9725 ;
        RECT 18.564 36.9475 18.636 36.9725 ;
        RECT 18.864 36.9475 18.936 36.9725 ;
        RECT 0.574 36.942 0.626 36.978 ;
        RECT 1.374 36.942 1.426 36.978 ;
        RECT 2.174 36.942 2.226 36.978 ;
        RECT 2.974 36.942 3.026 36.978 ;
        RECT 3.774 36.942 3.826 36.978 ;
        RECT 4.574 36.942 4.626 36.978 ;
        RECT 5.374 36.942 5.426 36.978 ;
        RECT 6.174 36.942 6.226 36.978 ;
        RECT 6.974 36.942 7.026 36.978 ;
        RECT 7.774 36.942 7.826 36.978 ;
        RECT 8.574 36.942 8.626 36.978 ;
        RECT 9.374 36.942 9.426 36.978 ;
        RECT 10.174 36.942 10.226 36.978 ;
        RECT 10.974 36.942 11.026 36.978 ;
        RECT 11.774 36.942 11.826 36.978 ;
        RECT 12.574 36.942 12.626 36.978 ;
        RECT 13.374 36.942 13.426 36.978 ;
        RECT 14.45 36.942 14.504 36.978 ;
        RECT 15.658 36.942 15.71 36.978 ;
        RECT 15.954 36.942 16.006 36.978 ;
        RECT 16.266 36.942 16.318 36.978 ;
        RECT 16.498 36.942 16.55 36.978 ;
        RECT 17.204 36.942 17.244 36.978 ;
        RECT 17.684 36.942 17.736 36.978 ;
        RECT 19.228 36.942 19.282 36.978 ;
        RECT 19.45 36.942 19.502 36.978 ;
        RECT 19.682 36.942 19.734 36.978 ;
        RECT 19.994 36.942 20.046 36.978 ;
        RECT 20.29 36.942 20.342 36.978 ;
        RECT 21.496 36.942 21.55 36.978 ;
        RECT 22.774 36.942 22.826 36.978 ;
        RECT 23.574 36.942 23.626 36.978 ;
        RECT 24.374 36.942 24.426 36.978 ;
        RECT 25.174 36.942 25.226 36.978 ;
        RECT 25.974 36.942 26.026 36.978 ;
        RECT 26.774 36.942 26.826 36.978 ;
        RECT 27.574 36.942 27.626 36.978 ;
        RECT 28.374 36.942 28.426 36.978 ;
        RECT 29.174 36.942 29.226 36.978 ;
        RECT 29.974 36.942 30.026 36.978 ;
        RECT 30.774 36.942 30.826 36.978 ;
        RECT 31.574 36.942 31.626 36.978 ;
        RECT 32.374 36.942 32.426 36.978 ;
        RECT 33.174 36.942 33.226 36.978 ;
        RECT 33.974 36.942 34.026 36.978 ;
        RECT 34.774 36.942 34.826 36.978 ;
        RECT 35.574 36.942 35.626 36.978 ;
        RECT 15.658 37.4275 15.71 37.4525 ;
        RECT 16.882 37.4275 16.936 37.4525 ;
        RECT 18.564 37.4275 18.636 37.4525 ;
        RECT 18.864 37.4275 18.936 37.4525 ;
        RECT 20.29 37.4275 20.342 37.4525 ;
        RECT 0.574 37.422 0.626 37.458 ;
        RECT 1.374 37.422 1.426 37.458 ;
        RECT 2.174 37.422 2.226 37.458 ;
        RECT 2.974 37.422 3.026 37.458 ;
        RECT 3.774 37.422 3.826 37.458 ;
        RECT 4.574 37.422 4.626 37.458 ;
        RECT 5.374 37.422 5.426 37.458 ;
        RECT 6.174 37.422 6.226 37.458 ;
        RECT 6.974 37.422 7.026 37.458 ;
        RECT 7.774 37.422 7.826 37.458 ;
        RECT 8.574 37.422 8.626 37.458 ;
        RECT 9.374 37.422 9.426 37.458 ;
        RECT 10.174 37.422 10.226 37.458 ;
        RECT 10.974 37.422 11.026 37.458 ;
        RECT 11.774 37.422 11.826 37.458 ;
        RECT 12.574 37.422 12.626 37.458 ;
        RECT 13.374 37.422 13.426 37.458 ;
        RECT 14.45 37.422 14.504 37.458 ;
        RECT 15.954 37.422 16.006 37.458 ;
        RECT 16.266 37.422 16.318 37.458 ;
        RECT 16.498 37.422 16.55 37.458 ;
        RECT 17.204 37.422 17.244 37.458 ;
        RECT 17.684 37.422 17.736 37.458 ;
        RECT 18.216 37.422 18.256 37.458 ;
        RECT 19.228 37.422 19.282 37.458 ;
        RECT 19.45 37.422 19.502 37.458 ;
        RECT 19.682 37.422 19.734 37.458 ;
        RECT 19.994 37.422 20.046 37.458 ;
        RECT 21.496 37.422 21.55 37.458 ;
        RECT 22.774 37.422 22.826 37.458 ;
        RECT 23.574 37.422 23.626 37.458 ;
        RECT 24.374 37.422 24.426 37.458 ;
        RECT 25.174 37.422 25.226 37.458 ;
        RECT 25.974 37.422 26.026 37.458 ;
        RECT 26.774 37.422 26.826 37.458 ;
        RECT 27.574 37.422 27.626 37.458 ;
        RECT 28.374 37.422 28.426 37.458 ;
        RECT 29.174 37.422 29.226 37.458 ;
        RECT 29.974 37.422 30.026 37.458 ;
        RECT 30.774 37.422 30.826 37.458 ;
        RECT 31.574 37.422 31.626 37.458 ;
        RECT 32.374 37.422 32.426 37.458 ;
        RECT 33.174 37.422 33.226 37.458 ;
        RECT 33.974 37.422 34.026 37.458 ;
        RECT 34.774 37.422 34.826 37.458 ;
        RECT 35.574 37.422 35.626 37.458 ;
        RECT 0.574 37.662 0.626 37.698 ;
        RECT 1.374 37.662 1.426 37.698 ;
        RECT 2.174 37.662 2.226 37.698 ;
        RECT 2.974 37.662 3.026 37.698 ;
        RECT 3.774 37.662 3.826 37.698 ;
        RECT 4.574 37.662 4.626 37.698 ;
        RECT 5.374 37.662 5.426 37.698 ;
        RECT 6.174 37.662 6.226 37.698 ;
        RECT 6.974 37.662 7.026 37.698 ;
        RECT 7.774 37.662 7.826 37.698 ;
        RECT 8.574 37.662 8.626 37.698 ;
        RECT 9.374 37.662 9.426 37.698 ;
        RECT 10.174 37.662 10.226 37.698 ;
        RECT 10.974 37.662 11.026 37.698 ;
        RECT 11.774 37.662 11.826 37.698 ;
        RECT 12.574 37.662 12.626 37.698 ;
        RECT 13.374 37.662 13.426 37.698 ;
        RECT 22.774 37.662 22.826 37.698 ;
        RECT 23.574 37.662 23.626 37.698 ;
        RECT 24.374 37.662 24.426 37.698 ;
        RECT 25.174 37.662 25.226 37.698 ;
        RECT 25.974 37.662 26.026 37.698 ;
        RECT 26.774 37.662 26.826 37.698 ;
        RECT 27.574 37.662 27.626 37.698 ;
        RECT 28.374 37.662 28.426 37.698 ;
        RECT 29.174 37.662 29.226 37.698 ;
        RECT 29.974 37.662 30.026 37.698 ;
        RECT 30.774 37.662 30.826 37.698 ;
        RECT 31.574 37.662 31.626 37.698 ;
        RECT 32.374 37.662 32.426 37.698 ;
        RECT 33.174 37.662 33.226 37.698 ;
        RECT 33.974 37.662 34.026 37.698 ;
        RECT 34.774 37.662 34.826 37.698 ;
        RECT 35.574 37.662 35.626 37.698 ;
        RECT 16.882 37.9075 16.936 37.9325 ;
        RECT 18.564 37.9075 18.636 37.9325 ;
        RECT 18.864 37.9075 18.936 37.9325 ;
        RECT 14.45 37.902 14.504 37.938 ;
        RECT 15.658 37.902 15.71 37.938 ;
        RECT 15.954 37.902 16.006 37.938 ;
        RECT 16.266 37.902 16.318 37.938 ;
        RECT 16.498 37.902 16.55 37.938 ;
        RECT 17.204 37.902 17.244 37.938 ;
        RECT 17.684 37.902 17.736 37.938 ;
        RECT 18.216 37.902 18.256 37.938 ;
        RECT 19.228 37.902 19.282 37.938 ;
        RECT 19.45 37.902 19.502 37.938 ;
        RECT 19.682 37.902 19.734 37.938 ;
        RECT 19.994 37.902 20.046 37.938 ;
        RECT 20.29 37.902 20.342 37.938 ;
        RECT 21.496 37.902 21.55 37.938 ;
        RECT 18.564 38.3875 18.636 38.4125 ;
        RECT 18.864 38.3875 18.936 38.4125 ;
        RECT 0.574 38.382 0.626 38.418 ;
        RECT 1.374 38.382 1.426 38.418 ;
        RECT 2.174 38.382 2.226 38.418 ;
        RECT 2.974 38.382 3.026 38.418 ;
        RECT 3.774 38.382 3.826 38.418 ;
        RECT 4.574 38.382 4.626 38.418 ;
        RECT 5.374 38.382 5.426 38.418 ;
        RECT 6.174 38.382 6.226 38.418 ;
        RECT 6.974 38.382 7.026 38.418 ;
        RECT 7.774 38.382 7.826 38.418 ;
        RECT 8.574 38.382 8.626 38.418 ;
        RECT 9.374 38.382 9.426 38.418 ;
        RECT 10.174 38.382 10.226 38.418 ;
        RECT 10.974 38.382 11.026 38.418 ;
        RECT 11.774 38.382 11.826 38.418 ;
        RECT 12.574 38.382 12.626 38.418 ;
        RECT 13.374 38.382 13.426 38.418 ;
        RECT 14.45 38.382 14.504 38.418 ;
        RECT 15.658 38.382 15.71 38.418 ;
        RECT 15.954 38.382 16.006 38.418 ;
        RECT 16.498 38.382 16.55 38.418 ;
        RECT 16.882 38.382 16.936 38.418 ;
        RECT 17.204 38.382 17.244 38.418 ;
        RECT 17.684 38.382 17.736 38.418 ;
        RECT 18.216 38.382 18.256 38.418 ;
        RECT 19.228 38.382 19.282 38.418 ;
        RECT 19.45 38.382 19.502 38.418 ;
        RECT 19.994 38.382 20.046 38.418 ;
        RECT 20.29 38.382 20.342 38.418 ;
        RECT 21.496 38.382 21.55 38.418 ;
        RECT 22.774 38.382 22.826 38.418 ;
        RECT 23.574 38.382 23.626 38.418 ;
        RECT 24.374 38.382 24.426 38.418 ;
        RECT 25.174 38.382 25.226 38.418 ;
        RECT 25.974 38.382 26.026 38.418 ;
        RECT 26.774 38.382 26.826 38.418 ;
        RECT 27.574 38.382 27.626 38.418 ;
        RECT 28.374 38.382 28.426 38.418 ;
        RECT 29.174 38.382 29.226 38.418 ;
        RECT 29.974 38.382 30.026 38.418 ;
        RECT 30.774 38.382 30.826 38.418 ;
        RECT 31.574 38.382 31.626 38.418 ;
        RECT 32.374 38.382 32.426 38.418 ;
        RECT 33.174 38.382 33.226 38.418 ;
        RECT 33.974 38.382 34.026 38.418 ;
        RECT 34.774 38.382 34.826 38.418 ;
        RECT 35.574 38.382 35.626 38.418 ;
        RECT 15.658 38.8675 15.71 38.8925 ;
        RECT 18.564 38.8675 18.636 38.8925 ;
        RECT 18.864 38.8675 18.936 38.8925 ;
        RECT 20.29 38.8675 20.342 38.8925 ;
        RECT 14.45 38.862 14.504 38.898 ;
        RECT 15.954 38.862 16.006 38.898 ;
        RECT 16.266 38.862 16.318 38.898 ;
        RECT 16.498 38.862 16.55 38.898 ;
        RECT 16.882 38.862 16.936 38.898 ;
        RECT 17.204 38.862 17.244 38.898 ;
        RECT 17.684 38.862 17.736 38.898 ;
        RECT 18.216 38.862 18.256 38.898 ;
        RECT 19.228 38.862 19.282 38.898 ;
        RECT 19.45 38.862 19.502 38.898 ;
        RECT 19.682 38.862 19.734 38.898 ;
        RECT 19.994 38.862 20.046 38.898 ;
        RECT 21.496 38.862 21.55 38.898 ;
        RECT 0.574 39.102 0.626 39.138 ;
        RECT 1.374 39.102 1.426 39.138 ;
        RECT 2.174 39.102 2.226 39.138 ;
        RECT 2.974 39.102 3.026 39.138 ;
        RECT 3.774 39.102 3.826 39.138 ;
        RECT 4.574 39.102 4.626 39.138 ;
        RECT 5.374 39.102 5.426 39.138 ;
        RECT 6.174 39.102 6.226 39.138 ;
        RECT 6.974 39.102 7.026 39.138 ;
        RECT 7.774 39.102 7.826 39.138 ;
        RECT 8.574 39.102 8.626 39.138 ;
        RECT 9.374 39.102 9.426 39.138 ;
        RECT 10.174 39.102 10.226 39.138 ;
        RECT 10.974 39.102 11.026 39.138 ;
        RECT 11.774 39.102 11.826 39.138 ;
        RECT 12.574 39.102 12.626 39.138 ;
        RECT 13.374 39.102 13.426 39.138 ;
        RECT 22.774 39.102 22.826 39.138 ;
        RECT 23.574 39.102 23.626 39.138 ;
        RECT 24.374 39.102 24.426 39.138 ;
        RECT 25.174 39.102 25.226 39.138 ;
        RECT 25.974 39.102 26.026 39.138 ;
        RECT 26.774 39.102 26.826 39.138 ;
        RECT 27.574 39.102 27.626 39.138 ;
        RECT 28.374 39.102 28.426 39.138 ;
        RECT 29.174 39.102 29.226 39.138 ;
        RECT 29.974 39.102 30.026 39.138 ;
        RECT 30.774 39.102 30.826 39.138 ;
        RECT 31.574 39.102 31.626 39.138 ;
        RECT 32.374 39.102 32.426 39.138 ;
        RECT 33.174 39.102 33.226 39.138 ;
        RECT 33.974 39.102 34.026 39.138 ;
        RECT 34.774 39.102 34.826 39.138 ;
        RECT 35.574 39.102 35.626 39.138 ;
        RECT 13.374 39.3475 13.426 39.3725 ;
        RECT 18.216 39.3475 18.256 39.3725 ;
        RECT 18.564 39.3475 18.636 39.3725 ;
        RECT 18.864 39.3475 18.936 39.3725 ;
        RECT 35.574 39.3475 35.626 39.3725 ;
        RECT 0.574 39.342 0.626 39.378 ;
        RECT 1.374 39.342 1.426 39.378 ;
        RECT 2.174 39.342 2.226 39.378 ;
        RECT 2.974 39.342 3.026 39.378 ;
        RECT 3.774 39.342 3.826 39.378 ;
        RECT 4.574 39.342 4.626 39.378 ;
        RECT 5.374 39.342 5.426 39.378 ;
        RECT 6.174 39.342 6.226 39.378 ;
        RECT 6.974 39.342 7.026 39.378 ;
        RECT 7.774 39.342 7.826 39.378 ;
        RECT 8.574 39.342 8.626 39.378 ;
        RECT 9.374 39.342 9.426 39.378 ;
        RECT 10.174 39.342 10.226 39.378 ;
        RECT 10.974 39.342 11.026 39.378 ;
        RECT 11.774 39.342 11.826 39.378 ;
        RECT 12.574 39.342 12.626 39.378 ;
        RECT 14.45 39.342 14.504 39.378 ;
        RECT 15.658 39.342 15.71 39.378 ;
        RECT 15.954 39.342 16.006 39.378 ;
        RECT 16.266 39.342 16.318 39.378 ;
        RECT 16.498 39.342 16.55 39.378 ;
        RECT 17.204 39.342 17.244 39.378 ;
        RECT 17.684 39.342 17.736 39.378 ;
        RECT 19.228 39.342 19.282 39.378 ;
        RECT 19.45 39.342 19.502 39.378 ;
        RECT 19.994 39.342 20.046 39.378 ;
        RECT 20.29 39.342 20.342 39.378 ;
        RECT 21.496 39.342 21.55 39.378 ;
        RECT 22.774 39.342 22.826 39.378 ;
        RECT 23.574 39.342 23.626 39.378 ;
        RECT 24.374 39.342 24.426 39.378 ;
        RECT 25.174 39.342 25.226 39.378 ;
        RECT 25.974 39.342 26.026 39.378 ;
        RECT 26.774 39.342 26.826 39.378 ;
        RECT 27.574 39.342 27.626 39.378 ;
        RECT 28.374 39.342 28.426 39.378 ;
        RECT 29.174 39.342 29.226 39.378 ;
        RECT 29.974 39.342 30.026 39.378 ;
        RECT 30.774 39.342 30.826 39.378 ;
        RECT 31.574 39.342 31.626 39.378 ;
        RECT 32.374 39.342 32.426 39.378 ;
        RECT 33.174 39.342 33.226 39.378 ;
        RECT 33.974 39.342 34.026 39.378 ;
        RECT 34.774 39.342 34.826 39.378 ;
        RECT 18.564 39.7075 18.636 39.7325 ;
        RECT 18.864 39.7075 18.936 39.7325 ;
        RECT 0.574 39.702 0.626 39.738 ;
        RECT 1.374 39.702 1.426 39.738 ;
        RECT 2.174 39.702 2.226 39.738 ;
        RECT 2.974 39.702 3.026 39.738 ;
        RECT 3.774 39.702 3.826 39.738 ;
        RECT 4.574 39.702 4.626 39.738 ;
        RECT 5.374 39.702 5.426 39.738 ;
        RECT 6.174 39.702 6.226 39.738 ;
        RECT 6.974 39.702 7.026 39.738 ;
        RECT 7.774 39.702 7.826 39.738 ;
        RECT 8.574 39.702 8.626 39.738 ;
        RECT 9.374 39.702 9.426 39.738 ;
        RECT 10.174 39.702 10.226 39.738 ;
        RECT 10.974 39.702 11.026 39.738 ;
        RECT 11.774 39.702 11.826 39.738 ;
        RECT 12.574 39.702 12.626 39.738 ;
        RECT 13.374 39.702 13.426 39.738 ;
        RECT 14.45 39.702 14.504 39.738 ;
        RECT 15.658 39.702 15.71 39.738 ;
        RECT 15.954 39.702 16.006 39.738 ;
        RECT 16.266 39.702 16.318 39.738 ;
        RECT 16.498 39.702 16.55 39.738 ;
        RECT 17.344 39.702 17.384 39.738 ;
        RECT 17.684 39.702 17.736 39.738 ;
        RECT 19.45 39.702 19.502 39.738 ;
        RECT 19.682 39.702 19.734 39.738 ;
        RECT 19.994 39.702 20.046 39.738 ;
        RECT 20.29 39.702 20.342 39.738 ;
        RECT 21.496 39.702 21.55 39.738 ;
        RECT 22.774 39.702 22.826 39.738 ;
        RECT 23.574 39.702 23.626 39.738 ;
        RECT 24.374 39.702 24.426 39.738 ;
        RECT 25.174 39.702 25.226 39.738 ;
        RECT 25.974 39.702 26.026 39.738 ;
        RECT 26.774 39.702 26.826 39.738 ;
        RECT 27.574 39.702 27.626 39.738 ;
        RECT 28.374 39.702 28.426 39.738 ;
        RECT 29.174 39.702 29.226 39.738 ;
        RECT 29.974 39.702 30.026 39.738 ;
        RECT 30.774 39.702 30.826 39.738 ;
        RECT 31.574 39.702 31.626 39.738 ;
        RECT 32.374 39.702 32.426 39.738 ;
        RECT 33.174 39.702 33.226 39.738 ;
        RECT 33.974 39.702 34.026 39.738 ;
        RECT 34.774 39.702 34.826 39.738 ;
        RECT 35.574 39.702 35.626 39.738 ;
        RECT 18.564 40.3075 18.636 40.3325 ;
        RECT 18.864 40.3075 18.936 40.3325 ;
        RECT 0.574 40.302 0.626 40.338 ;
        RECT 1.374 40.302 1.426 40.338 ;
        RECT 2.174 40.302 2.226 40.338 ;
        RECT 2.974 40.302 3.026 40.338 ;
        RECT 3.774 40.302 3.826 40.338 ;
        RECT 4.574 40.302 4.626 40.338 ;
        RECT 5.374 40.302 5.426 40.338 ;
        RECT 6.174 40.302 6.226 40.338 ;
        RECT 6.974 40.302 7.026 40.338 ;
        RECT 7.774 40.302 7.826 40.338 ;
        RECT 8.574 40.302 8.626 40.338 ;
        RECT 9.374 40.302 9.426 40.338 ;
        RECT 10.174 40.302 10.226 40.338 ;
        RECT 10.974 40.302 11.026 40.338 ;
        RECT 11.774 40.302 11.826 40.338 ;
        RECT 12.574 40.302 12.626 40.338 ;
        RECT 13.374 40.302 13.426 40.338 ;
        RECT 14.45 40.302 14.504 40.338 ;
        RECT 15.658 40.302 15.71 40.338 ;
        RECT 15.954 40.302 16.006 40.338 ;
        RECT 16.266 40.302 16.318 40.338 ;
        RECT 16.498 40.302 16.55 40.338 ;
        RECT 17.344 40.302 17.384 40.338 ;
        RECT 17.684 40.302 17.736 40.338 ;
        RECT 19.45 40.302 19.502 40.338 ;
        RECT 19.682 40.302 19.734 40.338 ;
        RECT 19.994 40.302 20.046 40.338 ;
        RECT 20.29 40.302 20.342 40.338 ;
        RECT 21.496 40.302 21.55 40.338 ;
        RECT 22.774 40.302 22.826 40.338 ;
        RECT 23.574 40.302 23.626 40.338 ;
        RECT 24.374 40.302 24.426 40.338 ;
        RECT 25.174 40.302 25.226 40.338 ;
        RECT 25.974 40.302 26.026 40.338 ;
        RECT 26.774 40.302 26.826 40.338 ;
        RECT 27.574 40.302 27.626 40.338 ;
        RECT 28.374 40.302 28.426 40.338 ;
        RECT 29.174 40.302 29.226 40.338 ;
        RECT 29.974 40.302 30.026 40.338 ;
        RECT 30.774 40.302 30.826 40.338 ;
        RECT 31.574 40.302 31.626 40.338 ;
        RECT 32.374 40.302 32.426 40.338 ;
        RECT 33.174 40.302 33.226 40.338 ;
        RECT 33.974 40.302 34.026 40.338 ;
        RECT 34.774 40.302 34.826 40.338 ;
        RECT 35.574 40.302 35.626 40.338 ;
        RECT 18.564 40.9075 18.636 40.9325 ;
        RECT 18.864 40.9075 18.936 40.9325 ;
        RECT 0.574 40.902 0.626 40.938 ;
        RECT 1.374 40.902 1.426 40.938 ;
        RECT 2.174 40.902 2.226 40.938 ;
        RECT 2.974 40.902 3.026 40.938 ;
        RECT 3.774 40.902 3.826 40.938 ;
        RECT 4.574 40.902 4.626 40.938 ;
        RECT 5.374 40.902 5.426 40.938 ;
        RECT 6.174 40.902 6.226 40.938 ;
        RECT 6.974 40.902 7.026 40.938 ;
        RECT 7.774 40.902 7.826 40.938 ;
        RECT 8.574 40.902 8.626 40.938 ;
        RECT 9.374 40.902 9.426 40.938 ;
        RECT 10.174 40.902 10.226 40.938 ;
        RECT 10.974 40.902 11.026 40.938 ;
        RECT 11.774 40.902 11.826 40.938 ;
        RECT 12.574 40.902 12.626 40.938 ;
        RECT 13.374 40.902 13.426 40.938 ;
        RECT 14.45 40.902 14.504 40.938 ;
        RECT 15.658 40.902 15.71 40.938 ;
        RECT 15.954 40.902 16.006 40.938 ;
        RECT 16.266 40.902 16.318 40.938 ;
        RECT 16.498 40.902 16.55 40.938 ;
        RECT 17.344 40.902 17.384 40.938 ;
        RECT 17.684 40.902 17.736 40.938 ;
        RECT 19.45 40.902 19.502 40.938 ;
        RECT 19.682 40.902 19.734 40.938 ;
        RECT 19.994 40.902 20.046 40.938 ;
        RECT 20.29 40.902 20.342 40.938 ;
        RECT 21.496 40.902 21.55 40.938 ;
        RECT 22.774 40.902 22.826 40.938 ;
        RECT 23.574 40.902 23.626 40.938 ;
        RECT 24.374 40.902 24.426 40.938 ;
        RECT 25.174 40.902 25.226 40.938 ;
        RECT 25.974 40.902 26.026 40.938 ;
        RECT 26.774 40.902 26.826 40.938 ;
        RECT 27.574 40.902 27.626 40.938 ;
        RECT 28.374 40.902 28.426 40.938 ;
        RECT 29.174 40.902 29.226 40.938 ;
        RECT 29.974 40.902 30.026 40.938 ;
        RECT 30.774 40.902 30.826 40.938 ;
        RECT 31.574 40.902 31.626 40.938 ;
        RECT 32.374 40.902 32.426 40.938 ;
        RECT 33.174 40.902 33.226 40.938 ;
        RECT 33.974 40.902 34.026 40.938 ;
        RECT 34.774 40.902 34.826 40.938 ;
        RECT 35.574 40.902 35.626 40.938 ;
        RECT 18.564 41.5075 18.636 41.5325 ;
        RECT 18.864 41.5075 18.936 41.5325 ;
        RECT 0.574 41.502 0.626 41.538 ;
        RECT 1.374 41.502 1.426 41.538 ;
        RECT 2.174 41.502 2.226 41.538 ;
        RECT 2.974 41.502 3.026 41.538 ;
        RECT 3.774 41.502 3.826 41.538 ;
        RECT 4.574 41.502 4.626 41.538 ;
        RECT 5.374 41.502 5.426 41.538 ;
        RECT 6.174 41.502 6.226 41.538 ;
        RECT 6.974 41.502 7.026 41.538 ;
        RECT 7.774 41.502 7.826 41.538 ;
        RECT 8.574 41.502 8.626 41.538 ;
        RECT 9.374 41.502 9.426 41.538 ;
        RECT 10.174 41.502 10.226 41.538 ;
        RECT 10.974 41.502 11.026 41.538 ;
        RECT 11.774 41.502 11.826 41.538 ;
        RECT 12.574 41.502 12.626 41.538 ;
        RECT 13.374 41.502 13.426 41.538 ;
        RECT 14.45 41.502 14.504 41.538 ;
        RECT 15.658 41.502 15.71 41.538 ;
        RECT 15.954 41.502 16.006 41.538 ;
        RECT 16.266 41.502 16.318 41.538 ;
        RECT 16.498 41.502 16.55 41.538 ;
        RECT 17.344 41.502 17.384 41.538 ;
        RECT 17.684 41.502 17.736 41.538 ;
        RECT 19.45 41.502 19.502 41.538 ;
        RECT 19.682 41.502 19.734 41.538 ;
        RECT 19.994 41.502 20.046 41.538 ;
        RECT 20.29 41.502 20.342 41.538 ;
        RECT 21.496 41.502 21.55 41.538 ;
        RECT 22.774 41.502 22.826 41.538 ;
        RECT 23.574 41.502 23.626 41.538 ;
        RECT 24.374 41.502 24.426 41.538 ;
        RECT 25.174 41.502 25.226 41.538 ;
        RECT 25.974 41.502 26.026 41.538 ;
        RECT 26.774 41.502 26.826 41.538 ;
        RECT 27.574 41.502 27.626 41.538 ;
        RECT 28.374 41.502 28.426 41.538 ;
        RECT 29.174 41.502 29.226 41.538 ;
        RECT 29.974 41.502 30.026 41.538 ;
        RECT 30.774 41.502 30.826 41.538 ;
        RECT 31.574 41.502 31.626 41.538 ;
        RECT 32.374 41.502 32.426 41.538 ;
        RECT 33.174 41.502 33.226 41.538 ;
        RECT 33.974 41.502 34.026 41.538 ;
        RECT 34.774 41.502 34.826 41.538 ;
        RECT 35.574 41.502 35.626 41.538 ;
        RECT 18.564 42.1075 18.636 42.1325 ;
        RECT 18.864 42.1075 18.936 42.1325 ;
        RECT 0.574 42.102 0.626 42.138 ;
        RECT 1.374 42.102 1.426 42.138 ;
        RECT 2.174 42.102 2.226 42.138 ;
        RECT 2.974 42.102 3.026 42.138 ;
        RECT 3.774 42.102 3.826 42.138 ;
        RECT 4.574 42.102 4.626 42.138 ;
        RECT 5.374 42.102 5.426 42.138 ;
        RECT 6.174 42.102 6.226 42.138 ;
        RECT 6.974 42.102 7.026 42.138 ;
        RECT 7.774 42.102 7.826 42.138 ;
        RECT 8.574 42.102 8.626 42.138 ;
        RECT 9.374 42.102 9.426 42.138 ;
        RECT 10.174 42.102 10.226 42.138 ;
        RECT 10.974 42.102 11.026 42.138 ;
        RECT 11.774 42.102 11.826 42.138 ;
        RECT 12.574 42.102 12.626 42.138 ;
        RECT 13.374 42.102 13.426 42.138 ;
        RECT 14.45 42.102 14.504 42.138 ;
        RECT 15.658 42.102 15.71 42.138 ;
        RECT 15.954 42.102 16.006 42.138 ;
        RECT 16.266 42.102 16.318 42.138 ;
        RECT 16.498 42.102 16.55 42.138 ;
        RECT 17.344 42.102 17.384 42.138 ;
        RECT 17.684 42.102 17.736 42.138 ;
        RECT 19.45 42.102 19.502 42.138 ;
        RECT 19.682 42.102 19.734 42.138 ;
        RECT 19.994 42.102 20.046 42.138 ;
        RECT 20.29 42.102 20.342 42.138 ;
        RECT 21.496 42.102 21.55 42.138 ;
        RECT 22.774 42.102 22.826 42.138 ;
        RECT 23.574 42.102 23.626 42.138 ;
        RECT 24.374 42.102 24.426 42.138 ;
        RECT 25.174 42.102 25.226 42.138 ;
        RECT 25.974 42.102 26.026 42.138 ;
        RECT 26.774 42.102 26.826 42.138 ;
        RECT 27.574 42.102 27.626 42.138 ;
        RECT 28.374 42.102 28.426 42.138 ;
        RECT 29.174 42.102 29.226 42.138 ;
        RECT 29.974 42.102 30.026 42.138 ;
        RECT 30.774 42.102 30.826 42.138 ;
        RECT 31.574 42.102 31.626 42.138 ;
        RECT 32.374 42.102 32.426 42.138 ;
        RECT 33.174 42.102 33.226 42.138 ;
        RECT 33.974 42.102 34.026 42.138 ;
        RECT 34.774 42.102 34.826 42.138 ;
        RECT 35.574 42.102 35.626 42.138 ;
        RECT 18.564 42.7075 18.636 42.7325 ;
        RECT 18.864 42.7075 18.936 42.7325 ;
        RECT 0.574 42.702 0.626 42.738 ;
        RECT 1.374 42.702 1.426 42.738 ;
        RECT 2.174 42.702 2.226 42.738 ;
        RECT 2.974 42.702 3.026 42.738 ;
        RECT 3.774 42.702 3.826 42.738 ;
        RECT 4.574 42.702 4.626 42.738 ;
        RECT 5.374 42.702 5.426 42.738 ;
        RECT 6.174 42.702 6.226 42.738 ;
        RECT 6.974 42.702 7.026 42.738 ;
        RECT 7.774 42.702 7.826 42.738 ;
        RECT 8.574 42.702 8.626 42.738 ;
        RECT 9.374 42.702 9.426 42.738 ;
        RECT 10.174 42.702 10.226 42.738 ;
        RECT 10.974 42.702 11.026 42.738 ;
        RECT 11.774 42.702 11.826 42.738 ;
        RECT 12.574 42.702 12.626 42.738 ;
        RECT 13.374 42.702 13.426 42.738 ;
        RECT 14.45 42.702 14.504 42.738 ;
        RECT 15.658 42.702 15.71 42.738 ;
        RECT 15.954 42.702 16.006 42.738 ;
        RECT 16.266 42.702 16.318 42.738 ;
        RECT 16.498 42.702 16.55 42.738 ;
        RECT 17.344 42.702 17.384 42.738 ;
        RECT 17.684 42.702 17.736 42.738 ;
        RECT 19.45 42.702 19.502 42.738 ;
        RECT 19.682 42.702 19.734 42.738 ;
        RECT 19.994 42.702 20.046 42.738 ;
        RECT 20.29 42.702 20.342 42.738 ;
        RECT 21.496 42.702 21.55 42.738 ;
        RECT 22.774 42.702 22.826 42.738 ;
        RECT 23.574 42.702 23.626 42.738 ;
        RECT 24.374 42.702 24.426 42.738 ;
        RECT 25.174 42.702 25.226 42.738 ;
        RECT 25.974 42.702 26.026 42.738 ;
        RECT 26.774 42.702 26.826 42.738 ;
        RECT 27.574 42.702 27.626 42.738 ;
        RECT 28.374 42.702 28.426 42.738 ;
        RECT 29.174 42.702 29.226 42.738 ;
        RECT 29.974 42.702 30.026 42.738 ;
        RECT 30.774 42.702 30.826 42.738 ;
        RECT 31.574 42.702 31.626 42.738 ;
        RECT 32.374 42.702 32.426 42.738 ;
        RECT 33.174 42.702 33.226 42.738 ;
        RECT 33.974 42.702 34.026 42.738 ;
        RECT 34.774 42.702 34.826 42.738 ;
        RECT 35.574 42.702 35.626 42.738 ;
        RECT 18.564 43.3075 18.636 43.3325 ;
        RECT 18.864 43.3075 18.936 43.3325 ;
        RECT 0.574 43.302 0.626 43.338 ;
        RECT 1.374 43.302 1.426 43.338 ;
        RECT 2.174 43.302 2.226 43.338 ;
        RECT 2.974 43.302 3.026 43.338 ;
        RECT 3.774 43.302 3.826 43.338 ;
        RECT 4.574 43.302 4.626 43.338 ;
        RECT 5.374 43.302 5.426 43.338 ;
        RECT 6.174 43.302 6.226 43.338 ;
        RECT 6.974 43.302 7.026 43.338 ;
        RECT 7.774 43.302 7.826 43.338 ;
        RECT 8.574 43.302 8.626 43.338 ;
        RECT 9.374 43.302 9.426 43.338 ;
        RECT 10.174 43.302 10.226 43.338 ;
        RECT 10.974 43.302 11.026 43.338 ;
        RECT 11.774 43.302 11.826 43.338 ;
        RECT 12.574 43.302 12.626 43.338 ;
        RECT 13.374 43.302 13.426 43.338 ;
        RECT 14.45 43.302 14.504 43.338 ;
        RECT 15.658 43.302 15.71 43.338 ;
        RECT 15.954 43.302 16.006 43.338 ;
        RECT 16.266 43.302 16.318 43.338 ;
        RECT 16.498 43.302 16.55 43.338 ;
        RECT 17.344 43.302 17.384 43.338 ;
        RECT 17.684 43.302 17.736 43.338 ;
        RECT 19.45 43.302 19.502 43.338 ;
        RECT 19.682 43.302 19.734 43.338 ;
        RECT 19.994 43.302 20.046 43.338 ;
        RECT 20.29 43.302 20.342 43.338 ;
        RECT 21.496 43.302 21.55 43.338 ;
        RECT 22.774 43.302 22.826 43.338 ;
        RECT 23.574 43.302 23.626 43.338 ;
        RECT 24.374 43.302 24.426 43.338 ;
        RECT 25.174 43.302 25.226 43.338 ;
        RECT 25.974 43.302 26.026 43.338 ;
        RECT 26.774 43.302 26.826 43.338 ;
        RECT 27.574 43.302 27.626 43.338 ;
        RECT 28.374 43.302 28.426 43.338 ;
        RECT 29.174 43.302 29.226 43.338 ;
        RECT 29.974 43.302 30.026 43.338 ;
        RECT 30.774 43.302 30.826 43.338 ;
        RECT 31.574 43.302 31.626 43.338 ;
        RECT 32.374 43.302 32.426 43.338 ;
        RECT 33.174 43.302 33.226 43.338 ;
        RECT 33.974 43.302 34.026 43.338 ;
        RECT 34.774 43.302 34.826 43.338 ;
        RECT 35.574 43.302 35.626 43.338 ;
        RECT 18.564 43.9075 18.636 43.9325 ;
        RECT 18.864 43.9075 18.936 43.9325 ;
        RECT 0.574 43.902 0.626 43.938 ;
        RECT 1.374 43.902 1.426 43.938 ;
        RECT 2.174 43.902 2.226 43.938 ;
        RECT 2.974 43.902 3.026 43.938 ;
        RECT 3.774 43.902 3.826 43.938 ;
        RECT 4.574 43.902 4.626 43.938 ;
        RECT 5.374 43.902 5.426 43.938 ;
        RECT 6.174 43.902 6.226 43.938 ;
        RECT 6.974 43.902 7.026 43.938 ;
        RECT 7.774 43.902 7.826 43.938 ;
        RECT 8.574 43.902 8.626 43.938 ;
        RECT 9.374 43.902 9.426 43.938 ;
        RECT 10.174 43.902 10.226 43.938 ;
        RECT 10.974 43.902 11.026 43.938 ;
        RECT 11.774 43.902 11.826 43.938 ;
        RECT 12.574 43.902 12.626 43.938 ;
        RECT 13.374 43.902 13.426 43.938 ;
        RECT 14.45 43.902 14.504 43.938 ;
        RECT 15.658 43.902 15.71 43.938 ;
        RECT 15.954 43.902 16.006 43.938 ;
        RECT 16.266 43.902 16.318 43.938 ;
        RECT 16.498 43.902 16.55 43.938 ;
        RECT 17.344 43.902 17.384 43.938 ;
        RECT 17.684 43.902 17.736 43.938 ;
        RECT 19.45 43.902 19.502 43.938 ;
        RECT 19.682 43.902 19.734 43.938 ;
        RECT 19.994 43.902 20.046 43.938 ;
        RECT 20.29 43.902 20.342 43.938 ;
        RECT 21.496 43.902 21.55 43.938 ;
        RECT 22.774 43.902 22.826 43.938 ;
        RECT 23.574 43.902 23.626 43.938 ;
        RECT 24.374 43.902 24.426 43.938 ;
        RECT 25.174 43.902 25.226 43.938 ;
        RECT 25.974 43.902 26.026 43.938 ;
        RECT 26.774 43.902 26.826 43.938 ;
        RECT 27.574 43.902 27.626 43.938 ;
        RECT 28.374 43.902 28.426 43.938 ;
        RECT 29.174 43.902 29.226 43.938 ;
        RECT 29.974 43.902 30.026 43.938 ;
        RECT 30.774 43.902 30.826 43.938 ;
        RECT 31.574 43.902 31.626 43.938 ;
        RECT 32.374 43.902 32.426 43.938 ;
        RECT 33.174 43.902 33.226 43.938 ;
        RECT 33.974 43.902 34.026 43.938 ;
        RECT 34.774 43.902 34.826 43.938 ;
        RECT 35.574 43.902 35.626 43.938 ;
        RECT 18.564 44.5075 18.636 44.5325 ;
        RECT 18.864 44.5075 18.936 44.5325 ;
        RECT 0.574 44.502 0.626 44.538 ;
        RECT 1.374 44.502 1.426 44.538 ;
        RECT 2.174 44.502 2.226 44.538 ;
        RECT 2.974 44.502 3.026 44.538 ;
        RECT 3.774 44.502 3.826 44.538 ;
        RECT 4.574 44.502 4.626 44.538 ;
        RECT 5.374 44.502 5.426 44.538 ;
        RECT 6.174 44.502 6.226 44.538 ;
        RECT 6.974 44.502 7.026 44.538 ;
        RECT 7.774 44.502 7.826 44.538 ;
        RECT 8.574 44.502 8.626 44.538 ;
        RECT 9.374 44.502 9.426 44.538 ;
        RECT 10.174 44.502 10.226 44.538 ;
        RECT 10.974 44.502 11.026 44.538 ;
        RECT 11.774 44.502 11.826 44.538 ;
        RECT 12.574 44.502 12.626 44.538 ;
        RECT 13.374 44.502 13.426 44.538 ;
        RECT 14.45 44.502 14.504 44.538 ;
        RECT 15.658 44.502 15.71 44.538 ;
        RECT 15.954 44.502 16.006 44.538 ;
        RECT 16.266 44.502 16.318 44.538 ;
        RECT 16.498 44.502 16.55 44.538 ;
        RECT 17.344 44.502 17.384 44.538 ;
        RECT 17.684 44.502 17.736 44.538 ;
        RECT 19.45 44.502 19.502 44.538 ;
        RECT 19.682 44.502 19.734 44.538 ;
        RECT 19.994 44.502 20.046 44.538 ;
        RECT 20.29 44.502 20.342 44.538 ;
        RECT 21.496 44.502 21.55 44.538 ;
        RECT 22.774 44.502 22.826 44.538 ;
        RECT 23.574 44.502 23.626 44.538 ;
        RECT 24.374 44.502 24.426 44.538 ;
        RECT 25.174 44.502 25.226 44.538 ;
        RECT 25.974 44.502 26.026 44.538 ;
        RECT 26.774 44.502 26.826 44.538 ;
        RECT 27.574 44.502 27.626 44.538 ;
        RECT 28.374 44.502 28.426 44.538 ;
        RECT 29.174 44.502 29.226 44.538 ;
        RECT 29.974 44.502 30.026 44.538 ;
        RECT 30.774 44.502 30.826 44.538 ;
        RECT 31.574 44.502 31.626 44.538 ;
        RECT 32.374 44.502 32.426 44.538 ;
        RECT 33.174 44.502 33.226 44.538 ;
        RECT 33.974 44.502 34.026 44.538 ;
        RECT 34.774 44.502 34.826 44.538 ;
        RECT 35.574 44.502 35.626 44.538 ;
        RECT 18.564 45.1075 18.636 45.1325 ;
        RECT 18.864 45.1075 18.936 45.1325 ;
        RECT 0.574 45.102 0.626 45.138 ;
        RECT 1.374 45.102 1.426 45.138 ;
        RECT 2.174 45.102 2.226 45.138 ;
        RECT 2.974 45.102 3.026 45.138 ;
        RECT 3.774 45.102 3.826 45.138 ;
        RECT 4.574 45.102 4.626 45.138 ;
        RECT 5.374 45.102 5.426 45.138 ;
        RECT 6.174 45.102 6.226 45.138 ;
        RECT 6.974 45.102 7.026 45.138 ;
        RECT 7.774 45.102 7.826 45.138 ;
        RECT 8.574 45.102 8.626 45.138 ;
        RECT 9.374 45.102 9.426 45.138 ;
        RECT 10.174 45.102 10.226 45.138 ;
        RECT 10.974 45.102 11.026 45.138 ;
        RECT 11.774 45.102 11.826 45.138 ;
        RECT 12.574 45.102 12.626 45.138 ;
        RECT 13.374 45.102 13.426 45.138 ;
        RECT 14.45 45.102 14.504 45.138 ;
        RECT 15.658 45.102 15.71 45.138 ;
        RECT 15.954 45.102 16.006 45.138 ;
        RECT 16.266 45.102 16.318 45.138 ;
        RECT 16.498 45.102 16.55 45.138 ;
        RECT 17.344 45.102 17.384 45.138 ;
        RECT 17.684 45.102 17.736 45.138 ;
        RECT 19.45 45.102 19.502 45.138 ;
        RECT 19.682 45.102 19.734 45.138 ;
        RECT 19.994 45.102 20.046 45.138 ;
        RECT 20.29 45.102 20.342 45.138 ;
        RECT 21.496 45.102 21.55 45.138 ;
        RECT 22.774 45.102 22.826 45.138 ;
        RECT 23.574 45.102 23.626 45.138 ;
        RECT 24.374 45.102 24.426 45.138 ;
        RECT 25.174 45.102 25.226 45.138 ;
        RECT 25.974 45.102 26.026 45.138 ;
        RECT 26.774 45.102 26.826 45.138 ;
        RECT 27.574 45.102 27.626 45.138 ;
        RECT 28.374 45.102 28.426 45.138 ;
        RECT 29.174 45.102 29.226 45.138 ;
        RECT 29.974 45.102 30.026 45.138 ;
        RECT 30.774 45.102 30.826 45.138 ;
        RECT 31.574 45.102 31.626 45.138 ;
        RECT 32.374 45.102 32.426 45.138 ;
        RECT 33.174 45.102 33.226 45.138 ;
        RECT 33.974 45.102 34.026 45.138 ;
        RECT 34.774 45.102 34.826 45.138 ;
        RECT 35.574 45.102 35.626 45.138 ;
        RECT 18.564 45.7075 18.636 45.7325 ;
        RECT 18.864 45.7075 18.936 45.7325 ;
        RECT 0.574 45.702 0.626 45.738 ;
        RECT 1.374 45.702 1.426 45.738 ;
        RECT 2.174 45.702 2.226 45.738 ;
        RECT 2.974 45.702 3.026 45.738 ;
        RECT 3.774 45.702 3.826 45.738 ;
        RECT 4.574 45.702 4.626 45.738 ;
        RECT 5.374 45.702 5.426 45.738 ;
        RECT 6.174 45.702 6.226 45.738 ;
        RECT 6.974 45.702 7.026 45.738 ;
        RECT 7.774 45.702 7.826 45.738 ;
        RECT 8.574 45.702 8.626 45.738 ;
        RECT 9.374 45.702 9.426 45.738 ;
        RECT 10.174 45.702 10.226 45.738 ;
        RECT 10.974 45.702 11.026 45.738 ;
        RECT 11.774 45.702 11.826 45.738 ;
        RECT 12.574 45.702 12.626 45.738 ;
        RECT 13.374 45.702 13.426 45.738 ;
        RECT 14.45 45.702 14.504 45.738 ;
        RECT 15.658 45.702 15.71 45.738 ;
        RECT 15.954 45.702 16.006 45.738 ;
        RECT 16.266 45.702 16.318 45.738 ;
        RECT 16.498 45.702 16.55 45.738 ;
        RECT 17.344 45.702 17.384 45.738 ;
        RECT 17.684 45.702 17.736 45.738 ;
        RECT 19.45 45.702 19.502 45.738 ;
        RECT 19.682 45.702 19.734 45.738 ;
        RECT 19.994 45.702 20.046 45.738 ;
        RECT 20.29 45.702 20.342 45.738 ;
        RECT 21.496 45.702 21.55 45.738 ;
        RECT 22.774 45.702 22.826 45.738 ;
        RECT 23.574 45.702 23.626 45.738 ;
        RECT 24.374 45.702 24.426 45.738 ;
        RECT 25.174 45.702 25.226 45.738 ;
        RECT 25.974 45.702 26.026 45.738 ;
        RECT 26.774 45.702 26.826 45.738 ;
        RECT 27.574 45.702 27.626 45.738 ;
        RECT 28.374 45.702 28.426 45.738 ;
        RECT 29.174 45.702 29.226 45.738 ;
        RECT 29.974 45.702 30.026 45.738 ;
        RECT 30.774 45.702 30.826 45.738 ;
        RECT 31.574 45.702 31.626 45.738 ;
        RECT 32.374 45.702 32.426 45.738 ;
        RECT 33.174 45.702 33.226 45.738 ;
        RECT 33.974 45.702 34.026 45.738 ;
        RECT 34.774 45.702 34.826 45.738 ;
        RECT 35.574 45.702 35.626 45.738 ;
        RECT 18.564 46.3075 18.636 46.3325 ;
        RECT 18.864 46.3075 18.936 46.3325 ;
        RECT 0.574 46.302 0.626 46.338 ;
        RECT 1.374 46.302 1.426 46.338 ;
        RECT 2.174 46.302 2.226 46.338 ;
        RECT 2.974 46.302 3.026 46.338 ;
        RECT 3.774 46.302 3.826 46.338 ;
        RECT 4.574 46.302 4.626 46.338 ;
        RECT 5.374 46.302 5.426 46.338 ;
        RECT 6.174 46.302 6.226 46.338 ;
        RECT 6.974 46.302 7.026 46.338 ;
        RECT 7.774 46.302 7.826 46.338 ;
        RECT 8.574 46.302 8.626 46.338 ;
        RECT 9.374 46.302 9.426 46.338 ;
        RECT 10.174 46.302 10.226 46.338 ;
        RECT 10.974 46.302 11.026 46.338 ;
        RECT 11.774 46.302 11.826 46.338 ;
        RECT 12.574 46.302 12.626 46.338 ;
        RECT 13.374 46.302 13.426 46.338 ;
        RECT 14.45 46.302 14.504 46.338 ;
        RECT 15.658 46.302 15.71 46.338 ;
        RECT 15.954 46.302 16.006 46.338 ;
        RECT 16.266 46.302 16.318 46.338 ;
        RECT 16.498 46.302 16.55 46.338 ;
        RECT 17.344 46.302 17.384 46.338 ;
        RECT 17.684 46.302 17.736 46.338 ;
        RECT 19.45 46.302 19.502 46.338 ;
        RECT 19.682 46.302 19.734 46.338 ;
        RECT 19.994 46.302 20.046 46.338 ;
        RECT 20.29 46.302 20.342 46.338 ;
        RECT 21.496 46.302 21.55 46.338 ;
        RECT 22.774 46.302 22.826 46.338 ;
        RECT 23.574 46.302 23.626 46.338 ;
        RECT 24.374 46.302 24.426 46.338 ;
        RECT 25.174 46.302 25.226 46.338 ;
        RECT 25.974 46.302 26.026 46.338 ;
        RECT 26.774 46.302 26.826 46.338 ;
        RECT 27.574 46.302 27.626 46.338 ;
        RECT 28.374 46.302 28.426 46.338 ;
        RECT 29.174 46.302 29.226 46.338 ;
        RECT 29.974 46.302 30.026 46.338 ;
        RECT 30.774 46.302 30.826 46.338 ;
        RECT 31.574 46.302 31.626 46.338 ;
        RECT 32.374 46.302 32.426 46.338 ;
        RECT 33.174 46.302 33.226 46.338 ;
        RECT 33.974 46.302 34.026 46.338 ;
        RECT 34.774 46.302 34.826 46.338 ;
        RECT 35.574 46.302 35.626 46.338 ;
        RECT 18.564 46.9075 18.636 46.9325 ;
        RECT 18.864 46.9075 18.936 46.9325 ;
        RECT 0.574 46.902 0.626 46.938 ;
        RECT 1.374 46.902 1.426 46.938 ;
        RECT 2.174 46.902 2.226 46.938 ;
        RECT 2.974 46.902 3.026 46.938 ;
        RECT 3.774 46.902 3.826 46.938 ;
        RECT 4.574 46.902 4.626 46.938 ;
        RECT 5.374 46.902 5.426 46.938 ;
        RECT 6.174 46.902 6.226 46.938 ;
        RECT 6.974 46.902 7.026 46.938 ;
        RECT 7.774 46.902 7.826 46.938 ;
        RECT 8.574 46.902 8.626 46.938 ;
        RECT 9.374 46.902 9.426 46.938 ;
        RECT 10.174 46.902 10.226 46.938 ;
        RECT 10.974 46.902 11.026 46.938 ;
        RECT 11.774 46.902 11.826 46.938 ;
        RECT 12.574 46.902 12.626 46.938 ;
        RECT 13.374 46.902 13.426 46.938 ;
        RECT 14.45 46.902 14.504 46.938 ;
        RECT 15.658 46.902 15.71 46.938 ;
        RECT 15.954 46.902 16.006 46.938 ;
        RECT 16.266 46.902 16.318 46.938 ;
        RECT 16.498 46.902 16.55 46.938 ;
        RECT 17.344 46.902 17.384 46.938 ;
        RECT 17.684 46.902 17.736 46.938 ;
        RECT 19.45 46.902 19.502 46.938 ;
        RECT 19.682 46.902 19.734 46.938 ;
        RECT 19.994 46.902 20.046 46.938 ;
        RECT 20.29 46.902 20.342 46.938 ;
        RECT 21.496 46.902 21.55 46.938 ;
        RECT 22.774 46.902 22.826 46.938 ;
        RECT 23.574 46.902 23.626 46.938 ;
        RECT 24.374 46.902 24.426 46.938 ;
        RECT 25.174 46.902 25.226 46.938 ;
        RECT 25.974 46.902 26.026 46.938 ;
        RECT 26.774 46.902 26.826 46.938 ;
        RECT 27.574 46.902 27.626 46.938 ;
        RECT 28.374 46.902 28.426 46.938 ;
        RECT 29.174 46.902 29.226 46.938 ;
        RECT 29.974 46.902 30.026 46.938 ;
        RECT 30.774 46.902 30.826 46.938 ;
        RECT 31.574 46.902 31.626 46.938 ;
        RECT 32.374 46.902 32.426 46.938 ;
        RECT 33.174 46.902 33.226 46.938 ;
        RECT 33.974 46.902 34.026 46.938 ;
        RECT 34.774 46.902 34.826 46.938 ;
        RECT 35.574 46.902 35.626 46.938 ;
        RECT 18.564 47.5075 18.636 47.5325 ;
        RECT 18.864 47.5075 18.936 47.5325 ;
        RECT 0.574 47.502 0.626 47.538 ;
        RECT 1.374 47.502 1.426 47.538 ;
        RECT 2.174 47.502 2.226 47.538 ;
        RECT 2.974 47.502 3.026 47.538 ;
        RECT 3.774 47.502 3.826 47.538 ;
        RECT 4.574 47.502 4.626 47.538 ;
        RECT 5.374 47.502 5.426 47.538 ;
        RECT 6.174 47.502 6.226 47.538 ;
        RECT 6.974 47.502 7.026 47.538 ;
        RECT 7.774 47.502 7.826 47.538 ;
        RECT 8.574 47.502 8.626 47.538 ;
        RECT 9.374 47.502 9.426 47.538 ;
        RECT 10.174 47.502 10.226 47.538 ;
        RECT 10.974 47.502 11.026 47.538 ;
        RECT 11.774 47.502 11.826 47.538 ;
        RECT 12.574 47.502 12.626 47.538 ;
        RECT 13.374 47.502 13.426 47.538 ;
        RECT 14.45 47.502 14.504 47.538 ;
        RECT 15.658 47.502 15.71 47.538 ;
        RECT 15.954 47.502 16.006 47.538 ;
        RECT 16.266 47.502 16.318 47.538 ;
        RECT 16.498 47.502 16.55 47.538 ;
        RECT 17.344 47.502 17.384 47.538 ;
        RECT 17.684 47.502 17.736 47.538 ;
        RECT 19.45 47.502 19.502 47.538 ;
        RECT 19.682 47.502 19.734 47.538 ;
        RECT 19.994 47.502 20.046 47.538 ;
        RECT 20.29 47.502 20.342 47.538 ;
        RECT 21.496 47.502 21.55 47.538 ;
        RECT 22.774 47.502 22.826 47.538 ;
        RECT 23.574 47.502 23.626 47.538 ;
        RECT 24.374 47.502 24.426 47.538 ;
        RECT 25.174 47.502 25.226 47.538 ;
        RECT 25.974 47.502 26.026 47.538 ;
        RECT 26.774 47.502 26.826 47.538 ;
        RECT 27.574 47.502 27.626 47.538 ;
        RECT 28.374 47.502 28.426 47.538 ;
        RECT 29.174 47.502 29.226 47.538 ;
        RECT 29.974 47.502 30.026 47.538 ;
        RECT 30.774 47.502 30.826 47.538 ;
        RECT 31.574 47.502 31.626 47.538 ;
        RECT 32.374 47.502 32.426 47.538 ;
        RECT 33.174 47.502 33.226 47.538 ;
        RECT 33.974 47.502 34.026 47.538 ;
        RECT 34.774 47.502 34.826 47.538 ;
        RECT 35.574 47.502 35.626 47.538 ;
        RECT 18.564 48.1075 18.636 48.1325 ;
        RECT 18.864 48.1075 18.936 48.1325 ;
        RECT 0.574 48.102 0.626 48.138 ;
        RECT 1.374 48.102 1.426 48.138 ;
        RECT 2.174 48.102 2.226 48.138 ;
        RECT 2.974 48.102 3.026 48.138 ;
        RECT 3.774 48.102 3.826 48.138 ;
        RECT 4.574 48.102 4.626 48.138 ;
        RECT 5.374 48.102 5.426 48.138 ;
        RECT 6.174 48.102 6.226 48.138 ;
        RECT 6.974 48.102 7.026 48.138 ;
        RECT 7.774 48.102 7.826 48.138 ;
        RECT 8.574 48.102 8.626 48.138 ;
        RECT 9.374 48.102 9.426 48.138 ;
        RECT 10.174 48.102 10.226 48.138 ;
        RECT 10.974 48.102 11.026 48.138 ;
        RECT 11.774 48.102 11.826 48.138 ;
        RECT 12.574 48.102 12.626 48.138 ;
        RECT 13.374 48.102 13.426 48.138 ;
        RECT 14.45 48.102 14.504 48.138 ;
        RECT 15.658 48.102 15.71 48.138 ;
        RECT 15.954 48.102 16.006 48.138 ;
        RECT 16.266 48.102 16.318 48.138 ;
        RECT 16.498 48.102 16.55 48.138 ;
        RECT 17.344 48.102 17.384 48.138 ;
        RECT 17.684 48.102 17.736 48.138 ;
        RECT 19.45 48.102 19.502 48.138 ;
        RECT 19.682 48.102 19.734 48.138 ;
        RECT 19.994 48.102 20.046 48.138 ;
        RECT 20.29 48.102 20.342 48.138 ;
        RECT 21.496 48.102 21.55 48.138 ;
        RECT 22.774 48.102 22.826 48.138 ;
        RECT 23.574 48.102 23.626 48.138 ;
        RECT 24.374 48.102 24.426 48.138 ;
        RECT 25.174 48.102 25.226 48.138 ;
        RECT 25.974 48.102 26.026 48.138 ;
        RECT 26.774 48.102 26.826 48.138 ;
        RECT 27.574 48.102 27.626 48.138 ;
        RECT 28.374 48.102 28.426 48.138 ;
        RECT 29.174 48.102 29.226 48.138 ;
        RECT 29.974 48.102 30.026 48.138 ;
        RECT 30.774 48.102 30.826 48.138 ;
        RECT 31.574 48.102 31.626 48.138 ;
        RECT 32.374 48.102 32.426 48.138 ;
        RECT 33.174 48.102 33.226 48.138 ;
        RECT 33.974 48.102 34.026 48.138 ;
        RECT 34.774 48.102 34.826 48.138 ;
        RECT 35.574 48.102 35.626 48.138 ;
        RECT 18.564 48.7075 18.636 48.7325 ;
        RECT 18.864 48.7075 18.936 48.7325 ;
        RECT 0.574 48.702 0.626 48.738 ;
        RECT 1.374 48.702 1.426 48.738 ;
        RECT 2.174 48.702 2.226 48.738 ;
        RECT 2.974 48.702 3.026 48.738 ;
        RECT 3.774 48.702 3.826 48.738 ;
        RECT 4.574 48.702 4.626 48.738 ;
        RECT 5.374 48.702 5.426 48.738 ;
        RECT 6.174 48.702 6.226 48.738 ;
        RECT 6.974 48.702 7.026 48.738 ;
        RECT 7.774 48.702 7.826 48.738 ;
        RECT 8.574 48.702 8.626 48.738 ;
        RECT 9.374 48.702 9.426 48.738 ;
        RECT 10.174 48.702 10.226 48.738 ;
        RECT 10.974 48.702 11.026 48.738 ;
        RECT 11.774 48.702 11.826 48.738 ;
        RECT 12.574 48.702 12.626 48.738 ;
        RECT 13.374 48.702 13.426 48.738 ;
        RECT 14.45 48.702 14.504 48.738 ;
        RECT 15.658 48.702 15.71 48.738 ;
        RECT 15.954 48.702 16.006 48.738 ;
        RECT 16.266 48.702 16.318 48.738 ;
        RECT 16.498 48.702 16.55 48.738 ;
        RECT 17.344 48.702 17.384 48.738 ;
        RECT 17.684 48.702 17.736 48.738 ;
        RECT 19.45 48.702 19.502 48.738 ;
        RECT 19.682 48.702 19.734 48.738 ;
        RECT 19.994 48.702 20.046 48.738 ;
        RECT 20.29 48.702 20.342 48.738 ;
        RECT 21.496 48.702 21.55 48.738 ;
        RECT 22.774 48.702 22.826 48.738 ;
        RECT 23.574 48.702 23.626 48.738 ;
        RECT 24.374 48.702 24.426 48.738 ;
        RECT 25.174 48.702 25.226 48.738 ;
        RECT 25.974 48.702 26.026 48.738 ;
        RECT 26.774 48.702 26.826 48.738 ;
        RECT 27.574 48.702 27.626 48.738 ;
        RECT 28.374 48.702 28.426 48.738 ;
        RECT 29.174 48.702 29.226 48.738 ;
        RECT 29.974 48.702 30.026 48.738 ;
        RECT 30.774 48.702 30.826 48.738 ;
        RECT 31.574 48.702 31.626 48.738 ;
        RECT 32.374 48.702 32.426 48.738 ;
        RECT 33.174 48.702 33.226 48.738 ;
        RECT 33.974 48.702 34.026 48.738 ;
        RECT 34.774 48.702 34.826 48.738 ;
        RECT 35.574 48.702 35.626 48.738 ;
        RECT 18.564 49.3075 18.636 49.3325 ;
        RECT 18.864 49.3075 18.936 49.3325 ;
        RECT 0.574 49.302 0.626 49.338 ;
        RECT 1.374 49.302 1.426 49.338 ;
        RECT 2.174 49.302 2.226 49.338 ;
        RECT 2.974 49.302 3.026 49.338 ;
        RECT 3.774 49.302 3.826 49.338 ;
        RECT 4.574 49.302 4.626 49.338 ;
        RECT 5.374 49.302 5.426 49.338 ;
        RECT 6.174 49.302 6.226 49.338 ;
        RECT 6.974 49.302 7.026 49.338 ;
        RECT 7.774 49.302 7.826 49.338 ;
        RECT 8.574 49.302 8.626 49.338 ;
        RECT 9.374 49.302 9.426 49.338 ;
        RECT 10.174 49.302 10.226 49.338 ;
        RECT 10.974 49.302 11.026 49.338 ;
        RECT 11.774 49.302 11.826 49.338 ;
        RECT 12.574 49.302 12.626 49.338 ;
        RECT 13.374 49.302 13.426 49.338 ;
        RECT 14.45 49.302 14.504 49.338 ;
        RECT 15.658 49.302 15.71 49.338 ;
        RECT 15.954 49.302 16.006 49.338 ;
        RECT 16.266 49.302 16.318 49.338 ;
        RECT 16.498 49.302 16.55 49.338 ;
        RECT 17.344 49.302 17.384 49.338 ;
        RECT 17.684 49.302 17.736 49.338 ;
        RECT 19.45 49.302 19.502 49.338 ;
        RECT 19.682 49.302 19.734 49.338 ;
        RECT 19.994 49.302 20.046 49.338 ;
        RECT 20.29 49.302 20.342 49.338 ;
        RECT 21.496 49.302 21.55 49.338 ;
        RECT 22.774 49.302 22.826 49.338 ;
        RECT 23.574 49.302 23.626 49.338 ;
        RECT 24.374 49.302 24.426 49.338 ;
        RECT 25.174 49.302 25.226 49.338 ;
        RECT 25.974 49.302 26.026 49.338 ;
        RECT 26.774 49.302 26.826 49.338 ;
        RECT 27.574 49.302 27.626 49.338 ;
        RECT 28.374 49.302 28.426 49.338 ;
        RECT 29.174 49.302 29.226 49.338 ;
        RECT 29.974 49.302 30.026 49.338 ;
        RECT 30.774 49.302 30.826 49.338 ;
        RECT 31.574 49.302 31.626 49.338 ;
        RECT 32.374 49.302 32.426 49.338 ;
        RECT 33.174 49.302 33.226 49.338 ;
        RECT 33.974 49.302 34.026 49.338 ;
        RECT 34.774 49.302 34.826 49.338 ;
        RECT 35.574 49.302 35.626 49.338 ;
        RECT 18.564 49.9075 18.636 49.9325 ;
        RECT 18.864 49.9075 18.936 49.9325 ;
        RECT 0.574 49.902 0.626 49.938 ;
        RECT 1.374 49.902 1.426 49.938 ;
        RECT 2.174 49.902 2.226 49.938 ;
        RECT 2.974 49.902 3.026 49.938 ;
        RECT 3.774 49.902 3.826 49.938 ;
        RECT 4.574 49.902 4.626 49.938 ;
        RECT 5.374 49.902 5.426 49.938 ;
        RECT 6.174 49.902 6.226 49.938 ;
        RECT 6.974 49.902 7.026 49.938 ;
        RECT 7.774 49.902 7.826 49.938 ;
        RECT 8.574 49.902 8.626 49.938 ;
        RECT 9.374 49.902 9.426 49.938 ;
        RECT 10.174 49.902 10.226 49.938 ;
        RECT 10.974 49.902 11.026 49.938 ;
        RECT 11.774 49.902 11.826 49.938 ;
        RECT 12.574 49.902 12.626 49.938 ;
        RECT 13.374 49.902 13.426 49.938 ;
        RECT 14.45 49.902 14.504 49.938 ;
        RECT 15.658 49.902 15.71 49.938 ;
        RECT 15.954 49.902 16.006 49.938 ;
        RECT 16.266 49.902 16.318 49.938 ;
        RECT 16.498 49.902 16.55 49.938 ;
        RECT 17.344 49.902 17.384 49.938 ;
        RECT 17.684 49.902 17.736 49.938 ;
        RECT 19.45 49.902 19.502 49.938 ;
        RECT 19.682 49.902 19.734 49.938 ;
        RECT 19.994 49.902 20.046 49.938 ;
        RECT 20.29 49.902 20.342 49.938 ;
        RECT 21.496 49.902 21.55 49.938 ;
        RECT 22.774 49.902 22.826 49.938 ;
        RECT 23.574 49.902 23.626 49.938 ;
        RECT 24.374 49.902 24.426 49.938 ;
        RECT 25.174 49.902 25.226 49.938 ;
        RECT 25.974 49.902 26.026 49.938 ;
        RECT 26.774 49.902 26.826 49.938 ;
        RECT 27.574 49.902 27.626 49.938 ;
        RECT 28.374 49.902 28.426 49.938 ;
        RECT 29.174 49.902 29.226 49.938 ;
        RECT 29.974 49.902 30.026 49.938 ;
        RECT 30.774 49.902 30.826 49.938 ;
        RECT 31.574 49.902 31.626 49.938 ;
        RECT 32.374 49.902 32.426 49.938 ;
        RECT 33.174 49.902 33.226 49.938 ;
        RECT 33.974 49.902 34.026 49.938 ;
        RECT 34.774 49.902 34.826 49.938 ;
        RECT 35.574 49.902 35.626 49.938 ;
        RECT 18.564 50.5075 18.636 50.5325 ;
        RECT 18.864 50.5075 18.936 50.5325 ;
        RECT 0.574 50.502 0.626 50.538 ;
        RECT 1.374 50.502 1.426 50.538 ;
        RECT 2.174 50.502 2.226 50.538 ;
        RECT 2.974 50.502 3.026 50.538 ;
        RECT 3.774 50.502 3.826 50.538 ;
        RECT 4.574 50.502 4.626 50.538 ;
        RECT 5.374 50.502 5.426 50.538 ;
        RECT 6.174 50.502 6.226 50.538 ;
        RECT 6.974 50.502 7.026 50.538 ;
        RECT 7.774 50.502 7.826 50.538 ;
        RECT 8.574 50.502 8.626 50.538 ;
        RECT 9.374 50.502 9.426 50.538 ;
        RECT 10.174 50.502 10.226 50.538 ;
        RECT 10.974 50.502 11.026 50.538 ;
        RECT 11.774 50.502 11.826 50.538 ;
        RECT 12.574 50.502 12.626 50.538 ;
        RECT 13.374 50.502 13.426 50.538 ;
        RECT 14.45 50.502 14.504 50.538 ;
        RECT 15.658 50.502 15.71 50.538 ;
        RECT 15.954 50.502 16.006 50.538 ;
        RECT 16.266 50.502 16.318 50.538 ;
        RECT 16.498 50.502 16.55 50.538 ;
        RECT 17.344 50.502 17.384 50.538 ;
        RECT 17.684 50.502 17.736 50.538 ;
        RECT 19.45 50.502 19.502 50.538 ;
        RECT 19.682 50.502 19.734 50.538 ;
        RECT 19.994 50.502 20.046 50.538 ;
        RECT 20.29 50.502 20.342 50.538 ;
        RECT 21.496 50.502 21.55 50.538 ;
        RECT 22.774 50.502 22.826 50.538 ;
        RECT 23.574 50.502 23.626 50.538 ;
        RECT 24.374 50.502 24.426 50.538 ;
        RECT 25.174 50.502 25.226 50.538 ;
        RECT 25.974 50.502 26.026 50.538 ;
        RECT 26.774 50.502 26.826 50.538 ;
        RECT 27.574 50.502 27.626 50.538 ;
        RECT 28.374 50.502 28.426 50.538 ;
        RECT 29.174 50.502 29.226 50.538 ;
        RECT 29.974 50.502 30.026 50.538 ;
        RECT 30.774 50.502 30.826 50.538 ;
        RECT 31.574 50.502 31.626 50.538 ;
        RECT 32.374 50.502 32.426 50.538 ;
        RECT 33.174 50.502 33.226 50.538 ;
        RECT 33.974 50.502 34.026 50.538 ;
        RECT 34.774 50.502 34.826 50.538 ;
        RECT 35.574 50.502 35.626 50.538 ;
        RECT 18.564 51.1075 18.636 51.1325 ;
        RECT 18.864 51.1075 18.936 51.1325 ;
        RECT 0.574 51.102 0.626 51.138 ;
        RECT 1.374 51.102 1.426 51.138 ;
        RECT 2.174 51.102 2.226 51.138 ;
        RECT 2.974 51.102 3.026 51.138 ;
        RECT 3.774 51.102 3.826 51.138 ;
        RECT 4.574 51.102 4.626 51.138 ;
        RECT 5.374 51.102 5.426 51.138 ;
        RECT 6.174 51.102 6.226 51.138 ;
        RECT 6.974 51.102 7.026 51.138 ;
        RECT 7.774 51.102 7.826 51.138 ;
        RECT 8.574 51.102 8.626 51.138 ;
        RECT 9.374 51.102 9.426 51.138 ;
        RECT 10.174 51.102 10.226 51.138 ;
        RECT 10.974 51.102 11.026 51.138 ;
        RECT 11.774 51.102 11.826 51.138 ;
        RECT 12.574 51.102 12.626 51.138 ;
        RECT 13.374 51.102 13.426 51.138 ;
        RECT 14.45 51.102 14.504 51.138 ;
        RECT 15.658 51.102 15.71 51.138 ;
        RECT 15.954 51.102 16.006 51.138 ;
        RECT 16.266 51.102 16.318 51.138 ;
        RECT 16.498 51.102 16.55 51.138 ;
        RECT 17.344 51.102 17.384 51.138 ;
        RECT 17.684 51.102 17.736 51.138 ;
        RECT 19.45 51.102 19.502 51.138 ;
        RECT 19.682 51.102 19.734 51.138 ;
        RECT 19.994 51.102 20.046 51.138 ;
        RECT 20.29 51.102 20.342 51.138 ;
        RECT 21.496 51.102 21.55 51.138 ;
        RECT 22.774 51.102 22.826 51.138 ;
        RECT 23.574 51.102 23.626 51.138 ;
        RECT 24.374 51.102 24.426 51.138 ;
        RECT 25.174 51.102 25.226 51.138 ;
        RECT 25.974 51.102 26.026 51.138 ;
        RECT 26.774 51.102 26.826 51.138 ;
        RECT 27.574 51.102 27.626 51.138 ;
        RECT 28.374 51.102 28.426 51.138 ;
        RECT 29.174 51.102 29.226 51.138 ;
        RECT 29.974 51.102 30.026 51.138 ;
        RECT 30.774 51.102 30.826 51.138 ;
        RECT 31.574 51.102 31.626 51.138 ;
        RECT 32.374 51.102 32.426 51.138 ;
        RECT 33.174 51.102 33.226 51.138 ;
        RECT 33.974 51.102 34.026 51.138 ;
        RECT 34.774 51.102 34.826 51.138 ;
        RECT 35.574 51.102 35.626 51.138 ;
        RECT 18.564 51.7075 18.636 51.7325 ;
        RECT 18.864 51.7075 18.936 51.7325 ;
        RECT 0.574 51.702 0.626 51.738 ;
        RECT 1.374 51.702 1.426 51.738 ;
        RECT 2.174 51.702 2.226 51.738 ;
        RECT 2.974 51.702 3.026 51.738 ;
        RECT 3.774 51.702 3.826 51.738 ;
        RECT 4.574 51.702 4.626 51.738 ;
        RECT 5.374 51.702 5.426 51.738 ;
        RECT 6.174 51.702 6.226 51.738 ;
        RECT 6.974 51.702 7.026 51.738 ;
        RECT 7.774 51.702 7.826 51.738 ;
        RECT 8.574 51.702 8.626 51.738 ;
        RECT 9.374 51.702 9.426 51.738 ;
        RECT 10.174 51.702 10.226 51.738 ;
        RECT 10.974 51.702 11.026 51.738 ;
        RECT 11.774 51.702 11.826 51.738 ;
        RECT 12.574 51.702 12.626 51.738 ;
        RECT 13.374 51.702 13.426 51.738 ;
        RECT 14.45 51.702 14.504 51.738 ;
        RECT 15.658 51.702 15.71 51.738 ;
        RECT 15.954 51.702 16.006 51.738 ;
        RECT 16.266 51.702 16.318 51.738 ;
        RECT 16.498 51.702 16.55 51.738 ;
        RECT 17.344 51.702 17.384 51.738 ;
        RECT 17.684 51.702 17.736 51.738 ;
        RECT 19.45 51.702 19.502 51.738 ;
        RECT 19.682 51.702 19.734 51.738 ;
        RECT 19.994 51.702 20.046 51.738 ;
        RECT 20.29 51.702 20.342 51.738 ;
        RECT 21.496 51.702 21.55 51.738 ;
        RECT 22.774 51.702 22.826 51.738 ;
        RECT 23.574 51.702 23.626 51.738 ;
        RECT 24.374 51.702 24.426 51.738 ;
        RECT 25.174 51.702 25.226 51.738 ;
        RECT 25.974 51.702 26.026 51.738 ;
        RECT 26.774 51.702 26.826 51.738 ;
        RECT 27.574 51.702 27.626 51.738 ;
        RECT 28.374 51.702 28.426 51.738 ;
        RECT 29.174 51.702 29.226 51.738 ;
        RECT 29.974 51.702 30.026 51.738 ;
        RECT 30.774 51.702 30.826 51.738 ;
        RECT 31.574 51.702 31.626 51.738 ;
        RECT 32.374 51.702 32.426 51.738 ;
        RECT 33.174 51.702 33.226 51.738 ;
        RECT 33.974 51.702 34.026 51.738 ;
        RECT 34.774 51.702 34.826 51.738 ;
        RECT 35.574 51.702 35.626 51.738 ;
        RECT 18.564 52.3075 18.636 52.3325 ;
        RECT 18.864 52.3075 18.936 52.3325 ;
        RECT 0.574 52.302 0.626 52.338 ;
        RECT 1.374 52.302 1.426 52.338 ;
        RECT 2.174 52.302 2.226 52.338 ;
        RECT 2.974 52.302 3.026 52.338 ;
        RECT 3.774 52.302 3.826 52.338 ;
        RECT 4.574 52.302 4.626 52.338 ;
        RECT 5.374 52.302 5.426 52.338 ;
        RECT 6.174 52.302 6.226 52.338 ;
        RECT 6.974 52.302 7.026 52.338 ;
        RECT 7.774 52.302 7.826 52.338 ;
        RECT 8.574 52.302 8.626 52.338 ;
        RECT 9.374 52.302 9.426 52.338 ;
        RECT 10.174 52.302 10.226 52.338 ;
        RECT 10.974 52.302 11.026 52.338 ;
        RECT 11.774 52.302 11.826 52.338 ;
        RECT 12.574 52.302 12.626 52.338 ;
        RECT 13.374 52.302 13.426 52.338 ;
        RECT 14.45 52.302 14.504 52.338 ;
        RECT 15.658 52.302 15.71 52.338 ;
        RECT 15.954 52.302 16.006 52.338 ;
        RECT 16.266 52.302 16.318 52.338 ;
        RECT 16.498 52.302 16.55 52.338 ;
        RECT 17.344 52.302 17.384 52.338 ;
        RECT 17.684 52.302 17.736 52.338 ;
        RECT 19.45 52.302 19.502 52.338 ;
        RECT 19.682 52.302 19.734 52.338 ;
        RECT 19.994 52.302 20.046 52.338 ;
        RECT 20.29 52.302 20.342 52.338 ;
        RECT 21.496 52.302 21.55 52.338 ;
        RECT 22.774 52.302 22.826 52.338 ;
        RECT 23.574 52.302 23.626 52.338 ;
        RECT 24.374 52.302 24.426 52.338 ;
        RECT 25.174 52.302 25.226 52.338 ;
        RECT 25.974 52.302 26.026 52.338 ;
        RECT 26.774 52.302 26.826 52.338 ;
        RECT 27.574 52.302 27.626 52.338 ;
        RECT 28.374 52.302 28.426 52.338 ;
        RECT 29.174 52.302 29.226 52.338 ;
        RECT 29.974 52.302 30.026 52.338 ;
        RECT 30.774 52.302 30.826 52.338 ;
        RECT 31.574 52.302 31.626 52.338 ;
        RECT 32.374 52.302 32.426 52.338 ;
        RECT 33.174 52.302 33.226 52.338 ;
        RECT 33.974 52.302 34.026 52.338 ;
        RECT 34.774 52.302 34.826 52.338 ;
        RECT 35.574 52.302 35.626 52.338 ;
        RECT 18.564 52.9075 18.636 52.9325 ;
        RECT 18.864 52.9075 18.936 52.9325 ;
        RECT 0.574 52.902 0.626 52.938 ;
        RECT 1.374 52.902 1.426 52.938 ;
        RECT 2.174 52.902 2.226 52.938 ;
        RECT 2.974 52.902 3.026 52.938 ;
        RECT 3.774 52.902 3.826 52.938 ;
        RECT 4.574 52.902 4.626 52.938 ;
        RECT 5.374 52.902 5.426 52.938 ;
        RECT 6.174 52.902 6.226 52.938 ;
        RECT 6.974 52.902 7.026 52.938 ;
        RECT 7.774 52.902 7.826 52.938 ;
        RECT 8.574 52.902 8.626 52.938 ;
        RECT 9.374 52.902 9.426 52.938 ;
        RECT 10.174 52.902 10.226 52.938 ;
        RECT 10.974 52.902 11.026 52.938 ;
        RECT 11.774 52.902 11.826 52.938 ;
        RECT 12.574 52.902 12.626 52.938 ;
        RECT 13.374 52.902 13.426 52.938 ;
        RECT 14.45 52.902 14.504 52.938 ;
        RECT 15.658 52.902 15.71 52.938 ;
        RECT 15.954 52.902 16.006 52.938 ;
        RECT 16.266 52.902 16.318 52.938 ;
        RECT 16.498 52.902 16.55 52.938 ;
        RECT 17.344 52.902 17.384 52.938 ;
        RECT 17.684 52.902 17.736 52.938 ;
        RECT 19.45 52.902 19.502 52.938 ;
        RECT 19.682 52.902 19.734 52.938 ;
        RECT 19.994 52.902 20.046 52.938 ;
        RECT 20.29 52.902 20.342 52.938 ;
        RECT 21.496 52.902 21.55 52.938 ;
        RECT 22.774 52.902 22.826 52.938 ;
        RECT 23.574 52.902 23.626 52.938 ;
        RECT 24.374 52.902 24.426 52.938 ;
        RECT 25.174 52.902 25.226 52.938 ;
        RECT 25.974 52.902 26.026 52.938 ;
        RECT 26.774 52.902 26.826 52.938 ;
        RECT 27.574 52.902 27.626 52.938 ;
        RECT 28.374 52.902 28.426 52.938 ;
        RECT 29.174 52.902 29.226 52.938 ;
        RECT 29.974 52.902 30.026 52.938 ;
        RECT 30.774 52.902 30.826 52.938 ;
        RECT 31.574 52.902 31.626 52.938 ;
        RECT 32.374 52.902 32.426 52.938 ;
        RECT 33.174 52.902 33.226 52.938 ;
        RECT 33.974 52.902 34.026 52.938 ;
        RECT 34.774 52.902 34.826 52.938 ;
        RECT 35.574 52.902 35.626 52.938 ;
        RECT 18.564 53.5075 18.636 53.5325 ;
        RECT 18.864 53.5075 18.936 53.5325 ;
        RECT 0.574 53.502 0.626 53.538 ;
        RECT 1.374 53.502 1.426 53.538 ;
        RECT 2.174 53.502 2.226 53.538 ;
        RECT 2.974 53.502 3.026 53.538 ;
        RECT 3.774 53.502 3.826 53.538 ;
        RECT 4.574 53.502 4.626 53.538 ;
        RECT 5.374 53.502 5.426 53.538 ;
        RECT 6.174 53.502 6.226 53.538 ;
        RECT 6.974 53.502 7.026 53.538 ;
        RECT 7.774 53.502 7.826 53.538 ;
        RECT 8.574 53.502 8.626 53.538 ;
        RECT 9.374 53.502 9.426 53.538 ;
        RECT 10.174 53.502 10.226 53.538 ;
        RECT 10.974 53.502 11.026 53.538 ;
        RECT 11.774 53.502 11.826 53.538 ;
        RECT 12.574 53.502 12.626 53.538 ;
        RECT 13.374 53.502 13.426 53.538 ;
        RECT 14.45 53.502 14.504 53.538 ;
        RECT 15.658 53.502 15.71 53.538 ;
        RECT 15.954 53.502 16.006 53.538 ;
        RECT 16.266 53.502 16.318 53.538 ;
        RECT 16.498 53.502 16.55 53.538 ;
        RECT 17.344 53.502 17.384 53.538 ;
        RECT 17.684 53.502 17.736 53.538 ;
        RECT 19.45 53.502 19.502 53.538 ;
        RECT 19.682 53.502 19.734 53.538 ;
        RECT 19.994 53.502 20.046 53.538 ;
        RECT 20.29 53.502 20.342 53.538 ;
        RECT 21.496 53.502 21.55 53.538 ;
        RECT 22.774 53.502 22.826 53.538 ;
        RECT 23.574 53.502 23.626 53.538 ;
        RECT 24.374 53.502 24.426 53.538 ;
        RECT 25.174 53.502 25.226 53.538 ;
        RECT 25.974 53.502 26.026 53.538 ;
        RECT 26.774 53.502 26.826 53.538 ;
        RECT 27.574 53.502 27.626 53.538 ;
        RECT 28.374 53.502 28.426 53.538 ;
        RECT 29.174 53.502 29.226 53.538 ;
        RECT 29.974 53.502 30.026 53.538 ;
        RECT 30.774 53.502 30.826 53.538 ;
        RECT 31.574 53.502 31.626 53.538 ;
        RECT 32.374 53.502 32.426 53.538 ;
        RECT 33.174 53.502 33.226 53.538 ;
        RECT 33.974 53.502 34.026 53.538 ;
        RECT 34.774 53.502 34.826 53.538 ;
        RECT 35.574 53.502 35.626 53.538 ;
        RECT 18.564 54.1075 18.636 54.1325 ;
        RECT 18.864 54.1075 18.936 54.1325 ;
        RECT 0.574 54.102 0.626 54.138 ;
        RECT 1.374 54.102 1.426 54.138 ;
        RECT 2.174 54.102 2.226 54.138 ;
        RECT 2.974 54.102 3.026 54.138 ;
        RECT 3.774 54.102 3.826 54.138 ;
        RECT 4.574 54.102 4.626 54.138 ;
        RECT 5.374 54.102 5.426 54.138 ;
        RECT 6.174 54.102 6.226 54.138 ;
        RECT 6.974 54.102 7.026 54.138 ;
        RECT 7.774 54.102 7.826 54.138 ;
        RECT 8.574 54.102 8.626 54.138 ;
        RECT 9.374 54.102 9.426 54.138 ;
        RECT 10.174 54.102 10.226 54.138 ;
        RECT 10.974 54.102 11.026 54.138 ;
        RECT 11.774 54.102 11.826 54.138 ;
        RECT 12.574 54.102 12.626 54.138 ;
        RECT 13.374 54.102 13.426 54.138 ;
        RECT 14.45 54.102 14.504 54.138 ;
        RECT 15.658 54.102 15.71 54.138 ;
        RECT 15.954 54.102 16.006 54.138 ;
        RECT 16.266 54.102 16.318 54.138 ;
        RECT 16.498 54.102 16.55 54.138 ;
        RECT 17.344 54.102 17.384 54.138 ;
        RECT 17.684 54.102 17.736 54.138 ;
        RECT 19.45 54.102 19.502 54.138 ;
        RECT 19.682 54.102 19.734 54.138 ;
        RECT 19.994 54.102 20.046 54.138 ;
        RECT 20.29 54.102 20.342 54.138 ;
        RECT 21.496 54.102 21.55 54.138 ;
        RECT 22.774 54.102 22.826 54.138 ;
        RECT 23.574 54.102 23.626 54.138 ;
        RECT 24.374 54.102 24.426 54.138 ;
        RECT 25.174 54.102 25.226 54.138 ;
        RECT 25.974 54.102 26.026 54.138 ;
        RECT 26.774 54.102 26.826 54.138 ;
        RECT 27.574 54.102 27.626 54.138 ;
        RECT 28.374 54.102 28.426 54.138 ;
        RECT 29.174 54.102 29.226 54.138 ;
        RECT 29.974 54.102 30.026 54.138 ;
        RECT 30.774 54.102 30.826 54.138 ;
        RECT 31.574 54.102 31.626 54.138 ;
        RECT 32.374 54.102 32.426 54.138 ;
        RECT 33.174 54.102 33.226 54.138 ;
        RECT 33.974 54.102 34.026 54.138 ;
        RECT 34.774 54.102 34.826 54.138 ;
        RECT 35.574 54.102 35.626 54.138 ;
        RECT 18.564 54.7075 18.636 54.7325 ;
        RECT 18.864 54.7075 18.936 54.7325 ;
        RECT 0.574 54.702 0.626 54.738 ;
        RECT 1.374 54.702 1.426 54.738 ;
        RECT 2.174 54.702 2.226 54.738 ;
        RECT 2.974 54.702 3.026 54.738 ;
        RECT 3.774 54.702 3.826 54.738 ;
        RECT 4.574 54.702 4.626 54.738 ;
        RECT 5.374 54.702 5.426 54.738 ;
        RECT 6.174 54.702 6.226 54.738 ;
        RECT 6.974 54.702 7.026 54.738 ;
        RECT 7.774 54.702 7.826 54.738 ;
        RECT 8.574 54.702 8.626 54.738 ;
        RECT 9.374 54.702 9.426 54.738 ;
        RECT 10.174 54.702 10.226 54.738 ;
        RECT 10.974 54.702 11.026 54.738 ;
        RECT 11.774 54.702 11.826 54.738 ;
        RECT 12.574 54.702 12.626 54.738 ;
        RECT 13.374 54.702 13.426 54.738 ;
        RECT 14.45 54.702 14.504 54.738 ;
        RECT 15.658 54.702 15.71 54.738 ;
        RECT 15.954 54.702 16.006 54.738 ;
        RECT 16.266 54.702 16.318 54.738 ;
        RECT 16.498 54.702 16.55 54.738 ;
        RECT 17.344 54.702 17.384 54.738 ;
        RECT 17.684 54.702 17.736 54.738 ;
        RECT 19.45 54.702 19.502 54.738 ;
        RECT 19.682 54.702 19.734 54.738 ;
        RECT 19.994 54.702 20.046 54.738 ;
        RECT 20.29 54.702 20.342 54.738 ;
        RECT 21.496 54.702 21.55 54.738 ;
        RECT 22.774 54.702 22.826 54.738 ;
        RECT 23.574 54.702 23.626 54.738 ;
        RECT 24.374 54.702 24.426 54.738 ;
        RECT 25.174 54.702 25.226 54.738 ;
        RECT 25.974 54.702 26.026 54.738 ;
        RECT 26.774 54.702 26.826 54.738 ;
        RECT 27.574 54.702 27.626 54.738 ;
        RECT 28.374 54.702 28.426 54.738 ;
        RECT 29.174 54.702 29.226 54.738 ;
        RECT 29.974 54.702 30.026 54.738 ;
        RECT 30.774 54.702 30.826 54.738 ;
        RECT 31.574 54.702 31.626 54.738 ;
        RECT 32.374 54.702 32.426 54.738 ;
        RECT 33.174 54.702 33.226 54.738 ;
        RECT 33.974 54.702 34.026 54.738 ;
        RECT 34.774 54.702 34.826 54.738 ;
        RECT 35.574 54.702 35.626 54.738 ;
        RECT 18.564 55.3075 18.636 55.3325 ;
        RECT 18.864 55.3075 18.936 55.3325 ;
        RECT 0.574 55.302 0.626 55.338 ;
        RECT 1.374 55.302 1.426 55.338 ;
        RECT 2.174 55.302 2.226 55.338 ;
        RECT 2.974 55.302 3.026 55.338 ;
        RECT 3.774 55.302 3.826 55.338 ;
        RECT 4.574 55.302 4.626 55.338 ;
        RECT 5.374 55.302 5.426 55.338 ;
        RECT 6.174 55.302 6.226 55.338 ;
        RECT 6.974 55.302 7.026 55.338 ;
        RECT 7.774 55.302 7.826 55.338 ;
        RECT 8.574 55.302 8.626 55.338 ;
        RECT 9.374 55.302 9.426 55.338 ;
        RECT 10.174 55.302 10.226 55.338 ;
        RECT 10.974 55.302 11.026 55.338 ;
        RECT 11.774 55.302 11.826 55.338 ;
        RECT 12.574 55.302 12.626 55.338 ;
        RECT 13.374 55.302 13.426 55.338 ;
        RECT 14.45 55.302 14.504 55.338 ;
        RECT 15.658 55.302 15.71 55.338 ;
        RECT 15.954 55.302 16.006 55.338 ;
        RECT 16.266 55.302 16.318 55.338 ;
        RECT 16.498 55.302 16.55 55.338 ;
        RECT 17.344 55.302 17.384 55.338 ;
        RECT 17.684 55.302 17.736 55.338 ;
        RECT 19.45 55.302 19.502 55.338 ;
        RECT 19.682 55.302 19.734 55.338 ;
        RECT 19.994 55.302 20.046 55.338 ;
        RECT 20.29 55.302 20.342 55.338 ;
        RECT 21.496 55.302 21.55 55.338 ;
        RECT 22.774 55.302 22.826 55.338 ;
        RECT 23.574 55.302 23.626 55.338 ;
        RECT 24.374 55.302 24.426 55.338 ;
        RECT 25.174 55.302 25.226 55.338 ;
        RECT 25.974 55.302 26.026 55.338 ;
        RECT 26.774 55.302 26.826 55.338 ;
        RECT 27.574 55.302 27.626 55.338 ;
        RECT 28.374 55.302 28.426 55.338 ;
        RECT 29.174 55.302 29.226 55.338 ;
        RECT 29.974 55.302 30.026 55.338 ;
        RECT 30.774 55.302 30.826 55.338 ;
        RECT 31.574 55.302 31.626 55.338 ;
        RECT 32.374 55.302 32.426 55.338 ;
        RECT 33.174 55.302 33.226 55.338 ;
        RECT 33.974 55.302 34.026 55.338 ;
        RECT 34.774 55.302 34.826 55.338 ;
        RECT 35.574 55.302 35.626 55.338 ;
        RECT 18.564 55.9075 18.636 55.9325 ;
        RECT 18.864 55.9075 18.936 55.9325 ;
        RECT 0.574 55.902 0.626 55.938 ;
        RECT 1.374 55.902 1.426 55.938 ;
        RECT 2.174 55.902 2.226 55.938 ;
        RECT 2.974 55.902 3.026 55.938 ;
        RECT 3.774 55.902 3.826 55.938 ;
        RECT 4.574 55.902 4.626 55.938 ;
        RECT 5.374 55.902 5.426 55.938 ;
        RECT 6.174 55.902 6.226 55.938 ;
        RECT 6.974 55.902 7.026 55.938 ;
        RECT 7.774 55.902 7.826 55.938 ;
        RECT 8.574 55.902 8.626 55.938 ;
        RECT 9.374 55.902 9.426 55.938 ;
        RECT 10.174 55.902 10.226 55.938 ;
        RECT 10.974 55.902 11.026 55.938 ;
        RECT 11.774 55.902 11.826 55.938 ;
        RECT 12.574 55.902 12.626 55.938 ;
        RECT 13.374 55.902 13.426 55.938 ;
        RECT 14.45 55.902 14.504 55.938 ;
        RECT 15.658 55.902 15.71 55.938 ;
        RECT 15.954 55.902 16.006 55.938 ;
        RECT 16.266 55.902 16.318 55.938 ;
        RECT 16.498 55.902 16.55 55.938 ;
        RECT 17.344 55.902 17.384 55.938 ;
        RECT 17.684 55.902 17.736 55.938 ;
        RECT 19.45 55.902 19.502 55.938 ;
        RECT 19.682 55.902 19.734 55.938 ;
        RECT 19.994 55.902 20.046 55.938 ;
        RECT 20.29 55.902 20.342 55.938 ;
        RECT 21.496 55.902 21.55 55.938 ;
        RECT 22.774 55.902 22.826 55.938 ;
        RECT 23.574 55.902 23.626 55.938 ;
        RECT 24.374 55.902 24.426 55.938 ;
        RECT 25.174 55.902 25.226 55.938 ;
        RECT 25.974 55.902 26.026 55.938 ;
        RECT 26.774 55.902 26.826 55.938 ;
        RECT 27.574 55.902 27.626 55.938 ;
        RECT 28.374 55.902 28.426 55.938 ;
        RECT 29.174 55.902 29.226 55.938 ;
        RECT 29.974 55.902 30.026 55.938 ;
        RECT 30.774 55.902 30.826 55.938 ;
        RECT 31.574 55.902 31.626 55.938 ;
        RECT 32.374 55.902 32.426 55.938 ;
        RECT 33.174 55.902 33.226 55.938 ;
        RECT 33.974 55.902 34.026 55.938 ;
        RECT 34.774 55.902 34.826 55.938 ;
        RECT 35.574 55.902 35.626 55.938 ;
        RECT 18.564 56.5075 18.636 56.5325 ;
        RECT 18.864 56.5075 18.936 56.5325 ;
        RECT 0.574 56.502 0.626 56.538 ;
        RECT 1.374 56.502 1.426 56.538 ;
        RECT 2.174 56.502 2.226 56.538 ;
        RECT 2.974 56.502 3.026 56.538 ;
        RECT 3.774 56.502 3.826 56.538 ;
        RECT 4.574 56.502 4.626 56.538 ;
        RECT 5.374 56.502 5.426 56.538 ;
        RECT 6.174 56.502 6.226 56.538 ;
        RECT 6.974 56.502 7.026 56.538 ;
        RECT 7.774 56.502 7.826 56.538 ;
        RECT 8.574 56.502 8.626 56.538 ;
        RECT 9.374 56.502 9.426 56.538 ;
        RECT 10.174 56.502 10.226 56.538 ;
        RECT 10.974 56.502 11.026 56.538 ;
        RECT 11.774 56.502 11.826 56.538 ;
        RECT 12.574 56.502 12.626 56.538 ;
        RECT 13.374 56.502 13.426 56.538 ;
        RECT 14.45 56.502 14.504 56.538 ;
        RECT 15.658 56.502 15.71 56.538 ;
        RECT 15.954 56.502 16.006 56.538 ;
        RECT 16.266 56.502 16.318 56.538 ;
        RECT 16.498 56.502 16.55 56.538 ;
        RECT 17.344 56.502 17.384 56.538 ;
        RECT 17.684 56.502 17.736 56.538 ;
        RECT 19.45 56.502 19.502 56.538 ;
        RECT 19.682 56.502 19.734 56.538 ;
        RECT 19.994 56.502 20.046 56.538 ;
        RECT 20.29 56.502 20.342 56.538 ;
        RECT 21.496 56.502 21.55 56.538 ;
        RECT 22.774 56.502 22.826 56.538 ;
        RECT 23.574 56.502 23.626 56.538 ;
        RECT 24.374 56.502 24.426 56.538 ;
        RECT 25.174 56.502 25.226 56.538 ;
        RECT 25.974 56.502 26.026 56.538 ;
        RECT 26.774 56.502 26.826 56.538 ;
        RECT 27.574 56.502 27.626 56.538 ;
        RECT 28.374 56.502 28.426 56.538 ;
        RECT 29.174 56.502 29.226 56.538 ;
        RECT 29.974 56.502 30.026 56.538 ;
        RECT 30.774 56.502 30.826 56.538 ;
        RECT 31.574 56.502 31.626 56.538 ;
        RECT 32.374 56.502 32.426 56.538 ;
        RECT 33.174 56.502 33.226 56.538 ;
        RECT 33.974 56.502 34.026 56.538 ;
        RECT 34.774 56.502 34.826 56.538 ;
        RECT 35.574 56.502 35.626 56.538 ;
        RECT 18.564 57.1075 18.636 57.1325 ;
        RECT 18.864 57.1075 18.936 57.1325 ;
        RECT 0.574 57.102 0.626 57.138 ;
        RECT 1.374 57.102 1.426 57.138 ;
        RECT 2.174 57.102 2.226 57.138 ;
        RECT 2.974 57.102 3.026 57.138 ;
        RECT 3.774 57.102 3.826 57.138 ;
        RECT 4.574 57.102 4.626 57.138 ;
        RECT 5.374 57.102 5.426 57.138 ;
        RECT 6.174 57.102 6.226 57.138 ;
        RECT 6.974 57.102 7.026 57.138 ;
        RECT 7.774 57.102 7.826 57.138 ;
        RECT 8.574 57.102 8.626 57.138 ;
        RECT 9.374 57.102 9.426 57.138 ;
        RECT 10.174 57.102 10.226 57.138 ;
        RECT 10.974 57.102 11.026 57.138 ;
        RECT 11.774 57.102 11.826 57.138 ;
        RECT 12.574 57.102 12.626 57.138 ;
        RECT 13.374 57.102 13.426 57.138 ;
        RECT 14.45 57.102 14.504 57.138 ;
        RECT 15.658 57.102 15.71 57.138 ;
        RECT 15.954 57.102 16.006 57.138 ;
        RECT 16.266 57.102 16.318 57.138 ;
        RECT 16.498 57.102 16.55 57.138 ;
        RECT 17.344 57.102 17.384 57.138 ;
        RECT 17.684 57.102 17.736 57.138 ;
        RECT 19.45 57.102 19.502 57.138 ;
        RECT 19.682 57.102 19.734 57.138 ;
        RECT 19.994 57.102 20.046 57.138 ;
        RECT 20.29 57.102 20.342 57.138 ;
        RECT 21.496 57.102 21.55 57.138 ;
        RECT 22.774 57.102 22.826 57.138 ;
        RECT 23.574 57.102 23.626 57.138 ;
        RECT 24.374 57.102 24.426 57.138 ;
        RECT 25.174 57.102 25.226 57.138 ;
        RECT 25.974 57.102 26.026 57.138 ;
        RECT 26.774 57.102 26.826 57.138 ;
        RECT 27.574 57.102 27.626 57.138 ;
        RECT 28.374 57.102 28.426 57.138 ;
        RECT 29.174 57.102 29.226 57.138 ;
        RECT 29.974 57.102 30.026 57.138 ;
        RECT 30.774 57.102 30.826 57.138 ;
        RECT 31.574 57.102 31.626 57.138 ;
        RECT 32.374 57.102 32.426 57.138 ;
        RECT 33.174 57.102 33.226 57.138 ;
        RECT 33.974 57.102 34.026 57.138 ;
        RECT 34.774 57.102 34.826 57.138 ;
        RECT 35.574 57.102 35.626 57.138 ;
        RECT 18.564 57.7075 18.636 57.7325 ;
        RECT 18.864 57.7075 18.936 57.7325 ;
        RECT 0.574 57.702 0.626 57.738 ;
        RECT 1.374 57.702 1.426 57.738 ;
        RECT 2.174 57.702 2.226 57.738 ;
        RECT 2.974 57.702 3.026 57.738 ;
        RECT 3.774 57.702 3.826 57.738 ;
        RECT 4.574 57.702 4.626 57.738 ;
        RECT 5.374 57.702 5.426 57.738 ;
        RECT 6.174 57.702 6.226 57.738 ;
        RECT 6.974 57.702 7.026 57.738 ;
        RECT 7.774 57.702 7.826 57.738 ;
        RECT 8.574 57.702 8.626 57.738 ;
        RECT 9.374 57.702 9.426 57.738 ;
        RECT 10.174 57.702 10.226 57.738 ;
        RECT 10.974 57.702 11.026 57.738 ;
        RECT 11.774 57.702 11.826 57.738 ;
        RECT 12.574 57.702 12.626 57.738 ;
        RECT 13.374 57.702 13.426 57.738 ;
        RECT 14.45 57.702 14.504 57.738 ;
        RECT 15.658 57.702 15.71 57.738 ;
        RECT 15.954 57.702 16.006 57.738 ;
        RECT 16.266 57.702 16.318 57.738 ;
        RECT 16.498 57.702 16.55 57.738 ;
        RECT 17.344 57.702 17.384 57.738 ;
        RECT 17.684 57.702 17.736 57.738 ;
        RECT 19.45 57.702 19.502 57.738 ;
        RECT 19.682 57.702 19.734 57.738 ;
        RECT 19.994 57.702 20.046 57.738 ;
        RECT 20.29 57.702 20.342 57.738 ;
        RECT 21.496 57.702 21.55 57.738 ;
        RECT 22.774 57.702 22.826 57.738 ;
        RECT 23.574 57.702 23.626 57.738 ;
        RECT 24.374 57.702 24.426 57.738 ;
        RECT 25.174 57.702 25.226 57.738 ;
        RECT 25.974 57.702 26.026 57.738 ;
        RECT 26.774 57.702 26.826 57.738 ;
        RECT 27.574 57.702 27.626 57.738 ;
        RECT 28.374 57.702 28.426 57.738 ;
        RECT 29.174 57.702 29.226 57.738 ;
        RECT 29.974 57.702 30.026 57.738 ;
        RECT 30.774 57.702 30.826 57.738 ;
        RECT 31.574 57.702 31.626 57.738 ;
        RECT 32.374 57.702 32.426 57.738 ;
        RECT 33.174 57.702 33.226 57.738 ;
        RECT 33.974 57.702 34.026 57.738 ;
        RECT 34.774 57.702 34.826 57.738 ;
        RECT 35.574 57.702 35.626 57.738 ;
        RECT 18.564 58.3075 18.636 58.3325 ;
        RECT 18.864 58.3075 18.936 58.3325 ;
        RECT 0.574 58.302 0.626 58.338 ;
        RECT 1.374 58.302 1.426 58.338 ;
        RECT 2.174 58.302 2.226 58.338 ;
        RECT 2.974 58.302 3.026 58.338 ;
        RECT 3.774 58.302 3.826 58.338 ;
        RECT 4.574 58.302 4.626 58.338 ;
        RECT 5.374 58.302 5.426 58.338 ;
        RECT 6.174 58.302 6.226 58.338 ;
        RECT 6.974 58.302 7.026 58.338 ;
        RECT 7.774 58.302 7.826 58.338 ;
        RECT 8.574 58.302 8.626 58.338 ;
        RECT 9.374 58.302 9.426 58.338 ;
        RECT 10.174 58.302 10.226 58.338 ;
        RECT 10.974 58.302 11.026 58.338 ;
        RECT 11.774 58.302 11.826 58.338 ;
        RECT 12.574 58.302 12.626 58.338 ;
        RECT 13.374 58.302 13.426 58.338 ;
        RECT 14.45 58.302 14.504 58.338 ;
        RECT 15.658 58.302 15.71 58.338 ;
        RECT 15.954 58.302 16.006 58.338 ;
        RECT 16.266 58.302 16.318 58.338 ;
        RECT 16.498 58.302 16.55 58.338 ;
        RECT 17.344 58.302 17.384 58.338 ;
        RECT 17.684 58.302 17.736 58.338 ;
        RECT 19.45 58.302 19.502 58.338 ;
        RECT 19.682 58.302 19.734 58.338 ;
        RECT 19.994 58.302 20.046 58.338 ;
        RECT 20.29 58.302 20.342 58.338 ;
        RECT 21.496 58.302 21.55 58.338 ;
        RECT 22.774 58.302 22.826 58.338 ;
        RECT 23.574 58.302 23.626 58.338 ;
        RECT 24.374 58.302 24.426 58.338 ;
        RECT 25.174 58.302 25.226 58.338 ;
        RECT 25.974 58.302 26.026 58.338 ;
        RECT 26.774 58.302 26.826 58.338 ;
        RECT 27.574 58.302 27.626 58.338 ;
        RECT 28.374 58.302 28.426 58.338 ;
        RECT 29.174 58.302 29.226 58.338 ;
        RECT 29.974 58.302 30.026 58.338 ;
        RECT 30.774 58.302 30.826 58.338 ;
        RECT 31.574 58.302 31.626 58.338 ;
        RECT 32.374 58.302 32.426 58.338 ;
        RECT 33.174 58.302 33.226 58.338 ;
        RECT 33.974 58.302 34.026 58.338 ;
        RECT 34.774 58.302 34.826 58.338 ;
        RECT 35.574 58.302 35.626 58.338 ;
        RECT 18.564 58.9075 18.636 58.9325 ;
        RECT 18.864 58.9075 18.936 58.9325 ;
        RECT 0.574 58.902 0.626 58.938 ;
        RECT 1.374 58.902 1.426 58.938 ;
        RECT 2.174 58.902 2.226 58.938 ;
        RECT 2.974 58.902 3.026 58.938 ;
        RECT 3.774 58.902 3.826 58.938 ;
        RECT 4.574 58.902 4.626 58.938 ;
        RECT 5.374 58.902 5.426 58.938 ;
        RECT 6.174 58.902 6.226 58.938 ;
        RECT 6.974 58.902 7.026 58.938 ;
        RECT 7.774 58.902 7.826 58.938 ;
        RECT 8.574 58.902 8.626 58.938 ;
        RECT 9.374 58.902 9.426 58.938 ;
        RECT 10.174 58.902 10.226 58.938 ;
        RECT 10.974 58.902 11.026 58.938 ;
        RECT 11.774 58.902 11.826 58.938 ;
        RECT 12.574 58.902 12.626 58.938 ;
        RECT 13.374 58.902 13.426 58.938 ;
        RECT 14.45 58.902 14.504 58.938 ;
        RECT 15.658 58.902 15.71 58.938 ;
        RECT 15.954 58.902 16.006 58.938 ;
        RECT 16.266 58.902 16.318 58.938 ;
        RECT 16.498 58.902 16.55 58.938 ;
        RECT 17.344 58.902 17.384 58.938 ;
        RECT 17.684 58.902 17.736 58.938 ;
        RECT 19.45 58.902 19.502 58.938 ;
        RECT 19.682 58.902 19.734 58.938 ;
        RECT 19.994 58.902 20.046 58.938 ;
        RECT 20.29 58.902 20.342 58.938 ;
        RECT 21.496 58.902 21.55 58.938 ;
        RECT 22.774 58.902 22.826 58.938 ;
        RECT 23.574 58.902 23.626 58.938 ;
        RECT 24.374 58.902 24.426 58.938 ;
        RECT 25.174 58.902 25.226 58.938 ;
        RECT 25.974 58.902 26.026 58.938 ;
        RECT 26.774 58.902 26.826 58.938 ;
        RECT 27.574 58.902 27.626 58.938 ;
        RECT 28.374 58.902 28.426 58.938 ;
        RECT 29.174 58.902 29.226 58.938 ;
        RECT 29.974 58.902 30.026 58.938 ;
        RECT 30.774 58.902 30.826 58.938 ;
        RECT 31.574 58.902 31.626 58.938 ;
        RECT 32.374 58.902 32.426 58.938 ;
        RECT 33.174 58.902 33.226 58.938 ;
        RECT 33.974 58.902 34.026 58.938 ;
        RECT 34.774 58.902 34.826 58.938 ;
        RECT 35.574 58.902 35.626 58.938 ;
        RECT 18.564 59.5075 18.636 59.5325 ;
        RECT 18.864 59.5075 18.936 59.5325 ;
        RECT 0.574 59.502 0.626 59.538 ;
        RECT 1.374 59.502 1.426 59.538 ;
        RECT 2.174 59.502 2.226 59.538 ;
        RECT 2.974 59.502 3.026 59.538 ;
        RECT 3.774 59.502 3.826 59.538 ;
        RECT 4.574 59.502 4.626 59.538 ;
        RECT 5.374 59.502 5.426 59.538 ;
        RECT 6.174 59.502 6.226 59.538 ;
        RECT 6.974 59.502 7.026 59.538 ;
        RECT 7.774 59.502 7.826 59.538 ;
        RECT 8.574 59.502 8.626 59.538 ;
        RECT 9.374 59.502 9.426 59.538 ;
        RECT 10.174 59.502 10.226 59.538 ;
        RECT 10.974 59.502 11.026 59.538 ;
        RECT 11.774 59.502 11.826 59.538 ;
        RECT 12.574 59.502 12.626 59.538 ;
        RECT 13.374 59.502 13.426 59.538 ;
        RECT 14.45 59.502 14.504 59.538 ;
        RECT 15.658 59.502 15.71 59.538 ;
        RECT 15.954 59.502 16.006 59.538 ;
        RECT 16.266 59.502 16.318 59.538 ;
        RECT 16.498 59.502 16.55 59.538 ;
        RECT 17.344 59.502 17.384 59.538 ;
        RECT 17.684 59.502 17.736 59.538 ;
        RECT 19.45 59.502 19.502 59.538 ;
        RECT 19.682 59.502 19.734 59.538 ;
        RECT 19.994 59.502 20.046 59.538 ;
        RECT 20.29 59.502 20.342 59.538 ;
        RECT 21.496 59.502 21.55 59.538 ;
        RECT 22.774 59.502 22.826 59.538 ;
        RECT 23.574 59.502 23.626 59.538 ;
        RECT 24.374 59.502 24.426 59.538 ;
        RECT 25.174 59.502 25.226 59.538 ;
        RECT 25.974 59.502 26.026 59.538 ;
        RECT 26.774 59.502 26.826 59.538 ;
        RECT 27.574 59.502 27.626 59.538 ;
        RECT 28.374 59.502 28.426 59.538 ;
        RECT 29.174 59.502 29.226 59.538 ;
        RECT 29.974 59.502 30.026 59.538 ;
        RECT 30.774 59.502 30.826 59.538 ;
        RECT 31.574 59.502 31.626 59.538 ;
        RECT 32.374 59.502 32.426 59.538 ;
        RECT 33.174 59.502 33.226 59.538 ;
        RECT 33.974 59.502 34.026 59.538 ;
        RECT 34.774 59.502 34.826 59.538 ;
        RECT 35.574 59.502 35.626 59.538 ;
        RECT 18.564 60.1075 18.636 60.1325 ;
        RECT 18.864 60.1075 18.936 60.1325 ;
        RECT 0.574 60.102 0.626 60.138 ;
        RECT 1.374 60.102 1.426 60.138 ;
        RECT 2.174 60.102 2.226 60.138 ;
        RECT 2.974 60.102 3.026 60.138 ;
        RECT 3.774 60.102 3.826 60.138 ;
        RECT 4.574 60.102 4.626 60.138 ;
        RECT 5.374 60.102 5.426 60.138 ;
        RECT 6.174 60.102 6.226 60.138 ;
        RECT 6.974 60.102 7.026 60.138 ;
        RECT 7.774 60.102 7.826 60.138 ;
        RECT 8.574 60.102 8.626 60.138 ;
        RECT 9.374 60.102 9.426 60.138 ;
        RECT 10.174 60.102 10.226 60.138 ;
        RECT 10.974 60.102 11.026 60.138 ;
        RECT 11.774 60.102 11.826 60.138 ;
        RECT 12.574 60.102 12.626 60.138 ;
        RECT 13.374 60.102 13.426 60.138 ;
        RECT 14.45 60.102 14.504 60.138 ;
        RECT 15.658 60.102 15.71 60.138 ;
        RECT 15.954 60.102 16.006 60.138 ;
        RECT 16.266 60.102 16.318 60.138 ;
        RECT 16.498 60.102 16.55 60.138 ;
        RECT 17.344 60.102 17.384 60.138 ;
        RECT 17.684 60.102 17.736 60.138 ;
        RECT 19.45 60.102 19.502 60.138 ;
        RECT 19.682 60.102 19.734 60.138 ;
        RECT 19.994 60.102 20.046 60.138 ;
        RECT 20.29 60.102 20.342 60.138 ;
        RECT 21.496 60.102 21.55 60.138 ;
        RECT 22.774 60.102 22.826 60.138 ;
        RECT 23.574 60.102 23.626 60.138 ;
        RECT 24.374 60.102 24.426 60.138 ;
        RECT 25.174 60.102 25.226 60.138 ;
        RECT 25.974 60.102 26.026 60.138 ;
        RECT 26.774 60.102 26.826 60.138 ;
        RECT 27.574 60.102 27.626 60.138 ;
        RECT 28.374 60.102 28.426 60.138 ;
        RECT 29.174 60.102 29.226 60.138 ;
        RECT 29.974 60.102 30.026 60.138 ;
        RECT 30.774 60.102 30.826 60.138 ;
        RECT 31.574 60.102 31.626 60.138 ;
        RECT 32.374 60.102 32.426 60.138 ;
        RECT 33.174 60.102 33.226 60.138 ;
        RECT 33.974 60.102 34.026 60.138 ;
        RECT 34.774 60.102 34.826 60.138 ;
        RECT 35.574 60.102 35.626 60.138 ;
        RECT 18.564 60.7075 18.636 60.7325 ;
        RECT 18.864 60.7075 18.936 60.7325 ;
        RECT 0.574 60.702 0.626 60.738 ;
        RECT 1.374 60.702 1.426 60.738 ;
        RECT 2.174 60.702 2.226 60.738 ;
        RECT 2.974 60.702 3.026 60.738 ;
        RECT 3.774 60.702 3.826 60.738 ;
        RECT 4.574 60.702 4.626 60.738 ;
        RECT 5.374 60.702 5.426 60.738 ;
        RECT 6.174 60.702 6.226 60.738 ;
        RECT 6.974 60.702 7.026 60.738 ;
        RECT 7.774 60.702 7.826 60.738 ;
        RECT 8.574 60.702 8.626 60.738 ;
        RECT 9.374 60.702 9.426 60.738 ;
        RECT 10.174 60.702 10.226 60.738 ;
        RECT 10.974 60.702 11.026 60.738 ;
        RECT 11.774 60.702 11.826 60.738 ;
        RECT 12.574 60.702 12.626 60.738 ;
        RECT 13.374 60.702 13.426 60.738 ;
        RECT 14.45 60.702 14.504 60.738 ;
        RECT 15.658 60.702 15.71 60.738 ;
        RECT 15.954 60.702 16.006 60.738 ;
        RECT 16.266 60.702 16.318 60.738 ;
        RECT 16.498 60.702 16.55 60.738 ;
        RECT 17.344 60.702 17.384 60.738 ;
        RECT 17.684 60.702 17.736 60.738 ;
        RECT 19.45 60.702 19.502 60.738 ;
        RECT 19.682 60.702 19.734 60.738 ;
        RECT 19.994 60.702 20.046 60.738 ;
        RECT 20.29 60.702 20.342 60.738 ;
        RECT 21.496 60.702 21.55 60.738 ;
        RECT 22.774 60.702 22.826 60.738 ;
        RECT 23.574 60.702 23.626 60.738 ;
        RECT 24.374 60.702 24.426 60.738 ;
        RECT 25.174 60.702 25.226 60.738 ;
        RECT 25.974 60.702 26.026 60.738 ;
        RECT 26.774 60.702 26.826 60.738 ;
        RECT 27.574 60.702 27.626 60.738 ;
        RECT 28.374 60.702 28.426 60.738 ;
        RECT 29.174 60.702 29.226 60.738 ;
        RECT 29.974 60.702 30.026 60.738 ;
        RECT 30.774 60.702 30.826 60.738 ;
        RECT 31.574 60.702 31.626 60.738 ;
        RECT 32.374 60.702 32.426 60.738 ;
        RECT 33.174 60.702 33.226 60.738 ;
        RECT 33.974 60.702 34.026 60.738 ;
        RECT 34.774 60.702 34.826 60.738 ;
        RECT 35.574 60.702 35.626 60.738 ;
        RECT 18.564 61.3075 18.636 61.3325 ;
        RECT 18.864 61.3075 18.936 61.3325 ;
        RECT 0.574 61.302 0.626 61.338 ;
        RECT 1.374 61.302 1.426 61.338 ;
        RECT 2.174 61.302 2.226 61.338 ;
        RECT 2.974 61.302 3.026 61.338 ;
        RECT 3.774 61.302 3.826 61.338 ;
        RECT 4.574 61.302 4.626 61.338 ;
        RECT 5.374 61.302 5.426 61.338 ;
        RECT 6.174 61.302 6.226 61.338 ;
        RECT 6.974 61.302 7.026 61.338 ;
        RECT 7.774 61.302 7.826 61.338 ;
        RECT 8.574 61.302 8.626 61.338 ;
        RECT 9.374 61.302 9.426 61.338 ;
        RECT 10.174 61.302 10.226 61.338 ;
        RECT 10.974 61.302 11.026 61.338 ;
        RECT 11.774 61.302 11.826 61.338 ;
        RECT 12.574 61.302 12.626 61.338 ;
        RECT 13.374 61.302 13.426 61.338 ;
        RECT 14.45 61.302 14.504 61.338 ;
        RECT 15.658 61.302 15.71 61.338 ;
        RECT 15.954 61.302 16.006 61.338 ;
        RECT 16.266 61.302 16.318 61.338 ;
        RECT 16.498 61.302 16.55 61.338 ;
        RECT 17.344 61.302 17.384 61.338 ;
        RECT 17.684 61.302 17.736 61.338 ;
        RECT 19.45 61.302 19.502 61.338 ;
        RECT 19.682 61.302 19.734 61.338 ;
        RECT 19.994 61.302 20.046 61.338 ;
        RECT 20.29 61.302 20.342 61.338 ;
        RECT 21.496 61.302 21.55 61.338 ;
        RECT 22.774 61.302 22.826 61.338 ;
        RECT 23.574 61.302 23.626 61.338 ;
        RECT 24.374 61.302 24.426 61.338 ;
        RECT 25.174 61.302 25.226 61.338 ;
        RECT 25.974 61.302 26.026 61.338 ;
        RECT 26.774 61.302 26.826 61.338 ;
        RECT 27.574 61.302 27.626 61.338 ;
        RECT 28.374 61.302 28.426 61.338 ;
        RECT 29.174 61.302 29.226 61.338 ;
        RECT 29.974 61.302 30.026 61.338 ;
        RECT 30.774 61.302 30.826 61.338 ;
        RECT 31.574 61.302 31.626 61.338 ;
        RECT 32.374 61.302 32.426 61.338 ;
        RECT 33.174 61.302 33.226 61.338 ;
        RECT 33.974 61.302 34.026 61.338 ;
        RECT 34.774 61.302 34.826 61.338 ;
        RECT 35.574 61.302 35.626 61.338 ;
        RECT 18.564 61.9075 18.636 61.9325 ;
        RECT 18.864 61.9075 18.936 61.9325 ;
        RECT 0.574 61.902 0.626 61.938 ;
        RECT 1.374 61.902 1.426 61.938 ;
        RECT 2.174 61.902 2.226 61.938 ;
        RECT 2.974 61.902 3.026 61.938 ;
        RECT 3.774 61.902 3.826 61.938 ;
        RECT 4.574 61.902 4.626 61.938 ;
        RECT 5.374 61.902 5.426 61.938 ;
        RECT 6.174 61.902 6.226 61.938 ;
        RECT 6.974 61.902 7.026 61.938 ;
        RECT 7.774 61.902 7.826 61.938 ;
        RECT 8.574 61.902 8.626 61.938 ;
        RECT 9.374 61.902 9.426 61.938 ;
        RECT 10.174 61.902 10.226 61.938 ;
        RECT 10.974 61.902 11.026 61.938 ;
        RECT 11.774 61.902 11.826 61.938 ;
        RECT 12.574 61.902 12.626 61.938 ;
        RECT 13.374 61.902 13.426 61.938 ;
        RECT 14.45 61.902 14.504 61.938 ;
        RECT 15.658 61.902 15.71 61.938 ;
        RECT 15.954 61.902 16.006 61.938 ;
        RECT 16.266 61.902 16.318 61.938 ;
        RECT 16.498 61.902 16.55 61.938 ;
        RECT 17.344 61.902 17.384 61.938 ;
        RECT 17.684 61.902 17.736 61.938 ;
        RECT 19.45 61.902 19.502 61.938 ;
        RECT 19.682 61.902 19.734 61.938 ;
        RECT 19.994 61.902 20.046 61.938 ;
        RECT 20.29 61.902 20.342 61.938 ;
        RECT 21.496 61.902 21.55 61.938 ;
        RECT 22.774 61.902 22.826 61.938 ;
        RECT 23.574 61.902 23.626 61.938 ;
        RECT 24.374 61.902 24.426 61.938 ;
        RECT 25.174 61.902 25.226 61.938 ;
        RECT 25.974 61.902 26.026 61.938 ;
        RECT 26.774 61.902 26.826 61.938 ;
        RECT 27.574 61.902 27.626 61.938 ;
        RECT 28.374 61.902 28.426 61.938 ;
        RECT 29.174 61.902 29.226 61.938 ;
        RECT 29.974 61.902 30.026 61.938 ;
        RECT 30.774 61.902 30.826 61.938 ;
        RECT 31.574 61.902 31.626 61.938 ;
        RECT 32.374 61.902 32.426 61.938 ;
        RECT 33.174 61.902 33.226 61.938 ;
        RECT 33.974 61.902 34.026 61.938 ;
        RECT 34.774 61.902 34.826 61.938 ;
        RECT 35.574 61.902 35.626 61.938 ;
        RECT 18.564 62.5075 18.636 62.5325 ;
        RECT 18.864 62.5075 18.936 62.5325 ;
        RECT 0.574 62.502 0.626 62.538 ;
        RECT 1.374 62.502 1.426 62.538 ;
        RECT 2.174 62.502 2.226 62.538 ;
        RECT 2.974 62.502 3.026 62.538 ;
        RECT 3.774 62.502 3.826 62.538 ;
        RECT 4.574 62.502 4.626 62.538 ;
        RECT 5.374 62.502 5.426 62.538 ;
        RECT 6.174 62.502 6.226 62.538 ;
        RECT 6.974 62.502 7.026 62.538 ;
        RECT 7.774 62.502 7.826 62.538 ;
        RECT 8.574 62.502 8.626 62.538 ;
        RECT 9.374 62.502 9.426 62.538 ;
        RECT 10.174 62.502 10.226 62.538 ;
        RECT 10.974 62.502 11.026 62.538 ;
        RECT 11.774 62.502 11.826 62.538 ;
        RECT 12.574 62.502 12.626 62.538 ;
        RECT 13.374 62.502 13.426 62.538 ;
        RECT 14.45 62.502 14.504 62.538 ;
        RECT 15.658 62.502 15.71 62.538 ;
        RECT 15.954 62.502 16.006 62.538 ;
        RECT 16.266 62.502 16.318 62.538 ;
        RECT 16.498 62.502 16.55 62.538 ;
        RECT 17.344 62.502 17.384 62.538 ;
        RECT 17.684 62.502 17.736 62.538 ;
        RECT 19.45 62.502 19.502 62.538 ;
        RECT 19.682 62.502 19.734 62.538 ;
        RECT 19.994 62.502 20.046 62.538 ;
        RECT 20.29 62.502 20.342 62.538 ;
        RECT 21.496 62.502 21.55 62.538 ;
        RECT 22.774 62.502 22.826 62.538 ;
        RECT 23.574 62.502 23.626 62.538 ;
        RECT 24.374 62.502 24.426 62.538 ;
        RECT 25.174 62.502 25.226 62.538 ;
        RECT 25.974 62.502 26.026 62.538 ;
        RECT 26.774 62.502 26.826 62.538 ;
        RECT 27.574 62.502 27.626 62.538 ;
        RECT 28.374 62.502 28.426 62.538 ;
        RECT 29.174 62.502 29.226 62.538 ;
        RECT 29.974 62.502 30.026 62.538 ;
        RECT 30.774 62.502 30.826 62.538 ;
        RECT 31.574 62.502 31.626 62.538 ;
        RECT 32.374 62.502 32.426 62.538 ;
        RECT 33.174 62.502 33.226 62.538 ;
        RECT 33.974 62.502 34.026 62.538 ;
        RECT 34.774 62.502 34.826 62.538 ;
        RECT 35.574 62.502 35.626 62.538 ;
        RECT 18.564 63.1075 18.636 63.1325 ;
        RECT 18.864 63.1075 18.936 63.1325 ;
        RECT 0.574 63.102 0.626 63.138 ;
        RECT 1.374 63.102 1.426 63.138 ;
        RECT 2.174 63.102 2.226 63.138 ;
        RECT 2.974 63.102 3.026 63.138 ;
        RECT 3.774 63.102 3.826 63.138 ;
        RECT 4.574 63.102 4.626 63.138 ;
        RECT 5.374 63.102 5.426 63.138 ;
        RECT 6.174 63.102 6.226 63.138 ;
        RECT 6.974 63.102 7.026 63.138 ;
        RECT 7.774 63.102 7.826 63.138 ;
        RECT 8.574 63.102 8.626 63.138 ;
        RECT 9.374 63.102 9.426 63.138 ;
        RECT 10.174 63.102 10.226 63.138 ;
        RECT 10.974 63.102 11.026 63.138 ;
        RECT 11.774 63.102 11.826 63.138 ;
        RECT 12.574 63.102 12.626 63.138 ;
        RECT 13.374 63.102 13.426 63.138 ;
        RECT 14.45 63.102 14.504 63.138 ;
        RECT 15.658 63.102 15.71 63.138 ;
        RECT 15.954 63.102 16.006 63.138 ;
        RECT 16.266 63.102 16.318 63.138 ;
        RECT 16.498 63.102 16.55 63.138 ;
        RECT 17.344 63.102 17.384 63.138 ;
        RECT 17.684 63.102 17.736 63.138 ;
        RECT 19.45 63.102 19.502 63.138 ;
        RECT 19.682 63.102 19.734 63.138 ;
        RECT 19.994 63.102 20.046 63.138 ;
        RECT 20.29 63.102 20.342 63.138 ;
        RECT 21.496 63.102 21.55 63.138 ;
        RECT 22.774 63.102 22.826 63.138 ;
        RECT 23.574 63.102 23.626 63.138 ;
        RECT 24.374 63.102 24.426 63.138 ;
        RECT 25.174 63.102 25.226 63.138 ;
        RECT 25.974 63.102 26.026 63.138 ;
        RECT 26.774 63.102 26.826 63.138 ;
        RECT 27.574 63.102 27.626 63.138 ;
        RECT 28.374 63.102 28.426 63.138 ;
        RECT 29.174 63.102 29.226 63.138 ;
        RECT 29.974 63.102 30.026 63.138 ;
        RECT 30.774 63.102 30.826 63.138 ;
        RECT 31.574 63.102 31.626 63.138 ;
        RECT 32.374 63.102 32.426 63.138 ;
        RECT 33.174 63.102 33.226 63.138 ;
        RECT 33.974 63.102 34.026 63.138 ;
        RECT 34.774 63.102 34.826 63.138 ;
        RECT 35.574 63.102 35.626 63.138 ;
        RECT 18.564 63.7075 18.636 63.7325 ;
        RECT 18.864 63.7075 18.936 63.7325 ;
        RECT 0.574 63.702 0.626 63.738 ;
        RECT 1.374 63.702 1.426 63.738 ;
        RECT 2.174 63.702 2.226 63.738 ;
        RECT 2.974 63.702 3.026 63.738 ;
        RECT 3.774 63.702 3.826 63.738 ;
        RECT 4.574 63.702 4.626 63.738 ;
        RECT 5.374 63.702 5.426 63.738 ;
        RECT 6.174 63.702 6.226 63.738 ;
        RECT 6.974 63.702 7.026 63.738 ;
        RECT 7.774 63.702 7.826 63.738 ;
        RECT 8.574 63.702 8.626 63.738 ;
        RECT 9.374 63.702 9.426 63.738 ;
        RECT 10.174 63.702 10.226 63.738 ;
        RECT 10.974 63.702 11.026 63.738 ;
        RECT 11.774 63.702 11.826 63.738 ;
        RECT 12.574 63.702 12.626 63.738 ;
        RECT 13.374 63.702 13.426 63.738 ;
        RECT 14.45 63.702 14.504 63.738 ;
        RECT 15.658 63.702 15.71 63.738 ;
        RECT 15.954 63.702 16.006 63.738 ;
        RECT 16.266 63.702 16.318 63.738 ;
        RECT 16.498 63.702 16.55 63.738 ;
        RECT 17.344 63.702 17.384 63.738 ;
        RECT 17.684 63.702 17.736 63.738 ;
        RECT 19.45 63.702 19.502 63.738 ;
        RECT 19.682 63.702 19.734 63.738 ;
        RECT 19.994 63.702 20.046 63.738 ;
        RECT 20.29 63.702 20.342 63.738 ;
        RECT 21.496 63.702 21.55 63.738 ;
        RECT 22.774 63.702 22.826 63.738 ;
        RECT 23.574 63.702 23.626 63.738 ;
        RECT 24.374 63.702 24.426 63.738 ;
        RECT 25.174 63.702 25.226 63.738 ;
        RECT 25.974 63.702 26.026 63.738 ;
        RECT 26.774 63.702 26.826 63.738 ;
        RECT 27.574 63.702 27.626 63.738 ;
        RECT 28.374 63.702 28.426 63.738 ;
        RECT 29.174 63.702 29.226 63.738 ;
        RECT 29.974 63.702 30.026 63.738 ;
        RECT 30.774 63.702 30.826 63.738 ;
        RECT 31.574 63.702 31.626 63.738 ;
        RECT 32.374 63.702 32.426 63.738 ;
        RECT 33.174 63.702 33.226 63.738 ;
        RECT 33.974 63.702 34.026 63.738 ;
        RECT 34.774 63.702 34.826 63.738 ;
        RECT 35.574 63.702 35.626 63.738 ;
        RECT 18.564 64.3075 18.636 64.3325 ;
        RECT 18.864 64.3075 18.936 64.3325 ;
        RECT 0.574 64.302 0.626 64.338 ;
        RECT 1.374 64.302 1.426 64.338 ;
        RECT 2.174 64.302 2.226 64.338 ;
        RECT 2.974 64.302 3.026 64.338 ;
        RECT 3.774 64.302 3.826 64.338 ;
        RECT 4.574 64.302 4.626 64.338 ;
        RECT 5.374 64.302 5.426 64.338 ;
        RECT 6.174 64.302 6.226 64.338 ;
        RECT 6.974 64.302 7.026 64.338 ;
        RECT 7.774 64.302 7.826 64.338 ;
        RECT 8.574 64.302 8.626 64.338 ;
        RECT 9.374 64.302 9.426 64.338 ;
        RECT 10.174 64.302 10.226 64.338 ;
        RECT 10.974 64.302 11.026 64.338 ;
        RECT 11.774 64.302 11.826 64.338 ;
        RECT 12.574 64.302 12.626 64.338 ;
        RECT 13.374 64.302 13.426 64.338 ;
        RECT 14.45 64.302 14.504 64.338 ;
        RECT 15.658 64.302 15.71 64.338 ;
        RECT 15.954 64.302 16.006 64.338 ;
        RECT 16.266 64.302 16.318 64.338 ;
        RECT 16.498 64.302 16.55 64.338 ;
        RECT 17.344 64.302 17.384 64.338 ;
        RECT 17.684 64.302 17.736 64.338 ;
        RECT 19.45 64.302 19.502 64.338 ;
        RECT 19.682 64.302 19.734 64.338 ;
        RECT 19.994 64.302 20.046 64.338 ;
        RECT 20.29 64.302 20.342 64.338 ;
        RECT 21.496 64.302 21.55 64.338 ;
        RECT 22.774 64.302 22.826 64.338 ;
        RECT 23.574 64.302 23.626 64.338 ;
        RECT 24.374 64.302 24.426 64.338 ;
        RECT 25.174 64.302 25.226 64.338 ;
        RECT 25.974 64.302 26.026 64.338 ;
        RECT 26.774 64.302 26.826 64.338 ;
        RECT 27.574 64.302 27.626 64.338 ;
        RECT 28.374 64.302 28.426 64.338 ;
        RECT 29.174 64.302 29.226 64.338 ;
        RECT 29.974 64.302 30.026 64.338 ;
        RECT 30.774 64.302 30.826 64.338 ;
        RECT 31.574 64.302 31.626 64.338 ;
        RECT 32.374 64.302 32.426 64.338 ;
        RECT 33.174 64.302 33.226 64.338 ;
        RECT 33.974 64.302 34.026 64.338 ;
        RECT 34.774 64.302 34.826 64.338 ;
        RECT 35.574 64.302 35.626 64.338 ;
        RECT 18.564 64.9075 18.636 64.9325 ;
        RECT 18.864 64.9075 18.936 64.9325 ;
        RECT 0.574 64.902 0.626 64.938 ;
        RECT 1.374 64.902 1.426 64.938 ;
        RECT 2.174 64.902 2.226 64.938 ;
        RECT 2.974 64.902 3.026 64.938 ;
        RECT 3.774 64.902 3.826 64.938 ;
        RECT 4.574 64.902 4.626 64.938 ;
        RECT 5.374 64.902 5.426 64.938 ;
        RECT 6.174 64.902 6.226 64.938 ;
        RECT 6.974 64.902 7.026 64.938 ;
        RECT 7.774 64.902 7.826 64.938 ;
        RECT 8.574 64.902 8.626 64.938 ;
        RECT 9.374 64.902 9.426 64.938 ;
        RECT 10.174 64.902 10.226 64.938 ;
        RECT 10.974 64.902 11.026 64.938 ;
        RECT 11.774 64.902 11.826 64.938 ;
        RECT 12.574 64.902 12.626 64.938 ;
        RECT 13.374 64.902 13.426 64.938 ;
        RECT 14.45 64.902 14.504 64.938 ;
        RECT 15.658 64.902 15.71 64.938 ;
        RECT 15.954 64.902 16.006 64.938 ;
        RECT 16.266 64.902 16.318 64.938 ;
        RECT 16.498 64.902 16.55 64.938 ;
        RECT 17.344 64.902 17.384 64.938 ;
        RECT 17.684 64.902 17.736 64.938 ;
        RECT 19.45 64.902 19.502 64.938 ;
        RECT 19.682 64.902 19.734 64.938 ;
        RECT 19.994 64.902 20.046 64.938 ;
        RECT 20.29 64.902 20.342 64.938 ;
        RECT 21.496 64.902 21.55 64.938 ;
        RECT 22.774 64.902 22.826 64.938 ;
        RECT 23.574 64.902 23.626 64.938 ;
        RECT 24.374 64.902 24.426 64.938 ;
        RECT 25.174 64.902 25.226 64.938 ;
        RECT 25.974 64.902 26.026 64.938 ;
        RECT 26.774 64.902 26.826 64.938 ;
        RECT 27.574 64.902 27.626 64.938 ;
        RECT 28.374 64.902 28.426 64.938 ;
        RECT 29.174 64.902 29.226 64.938 ;
        RECT 29.974 64.902 30.026 64.938 ;
        RECT 30.774 64.902 30.826 64.938 ;
        RECT 31.574 64.902 31.626 64.938 ;
        RECT 32.374 64.902 32.426 64.938 ;
        RECT 33.174 64.902 33.226 64.938 ;
        RECT 33.974 64.902 34.026 64.938 ;
        RECT 34.774 64.902 34.826 64.938 ;
        RECT 35.574 64.902 35.626 64.938 ;
        RECT 18.564 65.5075 18.636 65.5325 ;
        RECT 18.864 65.5075 18.936 65.5325 ;
        RECT 0.574 65.502 0.626 65.538 ;
        RECT 1.374 65.502 1.426 65.538 ;
        RECT 2.174 65.502 2.226 65.538 ;
        RECT 2.974 65.502 3.026 65.538 ;
        RECT 3.774 65.502 3.826 65.538 ;
        RECT 4.574 65.502 4.626 65.538 ;
        RECT 5.374 65.502 5.426 65.538 ;
        RECT 6.174 65.502 6.226 65.538 ;
        RECT 6.974 65.502 7.026 65.538 ;
        RECT 7.774 65.502 7.826 65.538 ;
        RECT 8.574 65.502 8.626 65.538 ;
        RECT 9.374 65.502 9.426 65.538 ;
        RECT 10.174 65.502 10.226 65.538 ;
        RECT 10.974 65.502 11.026 65.538 ;
        RECT 11.774 65.502 11.826 65.538 ;
        RECT 12.574 65.502 12.626 65.538 ;
        RECT 13.374 65.502 13.426 65.538 ;
        RECT 14.45 65.502 14.504 65.538 ;
        RECT 15.658 65.502 15.71 65.538 ;
        RECT 15.954 65.502 16.006 65.538 ;
        RECT 16.266 65.502 16.318 65.538 ;
        RECT 16.498 65.502 16.55 65.538 ;
        RECT 17.344 65.502 17.384 65.538 ;
        RECT 17.684 65.502 17.736 65.538 ;
        RECT 19.45 65.502 19.502 65.538 ;
        RECT 19.682 65.502 19.734 65.538 ;
        RECT 19.994 65.502 20.046 65.538 ;
        RECT 20.29 65.502 20.342 65.538 ;
        RECT 21.496 65.502 21.55 65.538 ;
        RECT 22.774 65.502 22.826 65.538 ;
        RECT 23.574 65.502 23.626 65.538 ;
        RECT 24.374 65.502 24.426 65.538 ;
        RECT 25.174 65.502 25.226 65.538 ;
        RECT 25.974 65.502 26.026 65.538 ;
        RECT 26.774 65.502 26.826 65.538 ;
        RECT 27.574 65.502 27.626 65.538 ;
        RECT 28.374 65.502 28.426 65.538 ;
        RECT 29.174 65.502 29.226 65.538 ;
        RECT 29.974 65.502 30.026 65.538 ;
        RECT 30.774 65.502 30.826 65.538 ;
        RECT 31.574 65.502 31.626 65.538 ;
        RECT 32.374 65.502 32.426 65.538 ;
        RECT 33.174 65.502 33.226 65.538 ;
        RECT 33.974 65.502 34.026 65.538 ;
        RECT 34.774 65.502 34.826 65.538 ;
        RECT 35.574 65.502 35.626 65.538 ;
        RECT 18.564 66.1075 18.636 66.1325 ;
        RECT 18.864 66.1075 18.936 66.1325 ;
        RECT 0.574 66.102 0.626 66.138 ;
        RECT 1.374 66.102 1.426 66.138 ;
        RECT 2.174 66.102 2.226 66.138 ;
        RECT 2.974 66.102 3.026 66.138 ;
        RECT 3.774 66.102 3.826 66.138 ;
        RECT 4.574 66.102 4.626 66.138 ;
        RECT 5.374 66.102 5.426 66.138 ;
        RECT 6.174 66.102 6.226 66.138 ;
        RECT 6.974 66.102 7.026 66.138 ;
        RECT 7.774 66.102 7.826 66.138 ;
        RECT 8.574 66.102 8.626 66.138 ;
        RECT 9.374 66.102 9.426 66.138 ;
        RECT 10.174 66.102 10.226 66.138 ;
        RECT 10.974 66.102 11.026 66.138 ;
        RECT 11.774 66.102 11.826 66.138 ;
        RECT 12.574 66.102 12.626 66.138 ;
        RECT 13.374 66.102 13.426 66.138 ;
        RECT 14.45 66.102 14.504 66.138 ;
        RECT 15.658 66.102 15.71 66.138 ;
        RECT 15.954 66.102 16.006 66.138 ;
        RECT 16.266 66.102 16.318 66.138 ;
        RECT 16.498 66.102 16.55 66.138 ;
        RECT 17.344 66.102 17.384 66.138 ;
        RECT 17.684 66.102 17.736 66.138 ;
        RECT 19.45 66.102 19.502 66.138 ;
        RECT 19.682 66.102 19.734 66.138 ;
        RECT 19.994 66.102 20.046 66.138 ;
        RECT 20.29 66.102 20.342 66.138 ;
        RECT 21.496 66.102 21.55 66.138 ;
        RECT 22.774 66.102 22.826 66.138 ;
        RECT 23.574 66.102 23.626 66.138 ;
        RECT 24.374 66.102 24.426 66.138 ;
        RECT 25.174 66.102 25.226 66.138 ;
        RECT 25.974 66.102 26.026 66.138 ;
        RECT 26.774 66.102 26.826 66.138 ;
        RECT 27.574 66.102 27.626 66.138 ;
        RECT 28.374 66.102 28.426 66.138 ;
        RECT 29.174 66.102 29.226 66.138 ;
        RECT 29.974 66.102 30.026 66.138 ;
        RECT 30.774 66.102 30.826 66.138 ;
        RECT 31.574 66.102 31.626 66.138 ;
        RECT 32.374 66.102 32.426 66.138 ;
        RECT 33.174 66.102 33.226 66.138 ;
        RECT 33.974 66.102 34.026 66.138 ;
        RECT 34.774 66.102 34.826 66.138 ;
        RECT 35.574 66.102 35.626 66.138 ;
        RECT 18.564 66.7075 18.636 66.7325 ;
        RECT 18.864 66.7075 18.936 66.7325 ;
        RECT 0.574 66.702 0.626 66.738 ;
        RECT 1.374 66.702 1.426 66.738 ;
        RECT 2.174 66.702 2.226 66.738 ;
        RECT 2.974 66.702 3.026 66.738 ;
        RECT 3.774 66.702 3.826 66.738 ;
        RECT 4.574 66.702 4.626 66.738 ;
        RECT 5.374 66.702 5.426 66.738 ;
        RECT 6.174 66.702 6.226 66.738 ;
        RECT 6.974 66.702 7.026 66.738 ;
        RECT 7.774 66.702 7.826 66.738 ;
        RECT 8.574 66.702 8.626 66.738 ;
        RECT 9.374 66.702 9.426 66.738 ;
        RECT 10.174 66.702 10.226 66.738 ;
        RECT 10.974 66.702 11.026 66.738 ;
        RECT 11.774 66.702 11.826 66.738 ;
        RECT 12.574 66.702 12.626 66.738 ;
        RECT 13.374 66.702 13.426 66.738 ;
        RECT 14.45 66.702 14.504 66.738 ;
        RECT 15.658 66.702 15.71 66.738 ;
        RECT 15.954 66.702 16.006 66.738 ;
        RECT 16.266 66.702 16.318 66.738 ;
        RECT 16.498 66.702 16.55 66.738 ;
        RECT 17.344 66.702 17.384 66.738 ;
        RECT 17.684 66.702 17.736 66.738 ;
        RECT 19.45 66.702 19.502 66.738 ;
        RECT 19.682 66.702 19.734 66.738 ;
        RECT 19.994 66.702 20.046 66.738 ;
        RECT 20.29 66.702 20.342 66.738 ;
        RECT 21.496 66.702 21.55 66.738 ;
        RECT 22.774 66.702 22.826 66.738 ;
        RECT 23.574 66.702 23.626 66.738 ;
        RECT 24.374 66.702 24.426 66.738 ;
        RECT 25.174 66.702 25.226 66.738 ;
        RECT 25.974 66.702 26.026 66.738 ;
        RECT 26.774 66.702 26.826 66.738 ;
        RECT 27.574 66.702 27.626 66.738 ;
        RECT 28.374 66.702 28.426 66.738 ;
        RECT 29.174 66.702 29.226 66.738 ;
        RECT 29.974 66.702 30.026 66.738 ;
        RECT 30.774 66.702 30.826 66.738 ;
        RECT 31.574 66.702 31.626 66.738 ;
        RECT 32.374 66.702 32.426 66.738 ;
        RECT 33.174 66.702 33.226 66.738 ;
        RECT 33.974 66.702 34.026 66.738 ;
        RECT 34.774 66.702 34.826 66.738 ;
        RECT 35.574 66.702 35.626 66.738 ;
        RECT 18.564 67.3075 18.636 67.3325 ;
        RECT 18.864 67.3075 18.936 67.3325 ;
        RECT 0.574 67.302 0.626 67.338 ;
        RECT 1.374 67.302 1.426 67.338 ;
        RECT 2.174 67.302 2.226 67.338 ;
        RECT 2.974 67.302 3.026 67.338 ;
        RECT 3.774 67.302 3.826 67.338 ;
        RECT 4.574 67.302 4.626 67.338 ;
        RECT 5.374 67.302 5.426 67.338 ;
        RECT 6.174 67.302 6.226 67.338 ;
        RECT 6.974 67.302 7.026 67.338 ;
        RECT 7.774 67.302 7.826 67.338 ;
        RECT 8.574 67.302 8.626 67.338 ;
        RECT 9.374 67.302 9.426 67.338 ;
        RECT 10.174 67.302 10.226 67.338 ;
        RECT 10.974 67.302 11.026 67.338 ;
        RECT 11.774 67.302 11.826 67.338 ;
        RECT 12.574 67.302 12.626 67.338 ;
        RECT 13.374 67.302 13.426 67.338 ;
        RECT 14.45 67.302 14.504 67.338 ;
        RECT 15.658 67.302 15.71 67.338 ;
        RECT 15.954 67.302 16.006 67.338 ;
        RECT 16.266 67.302 16.318 67.338 ;
        RECT 16.498 67.302 16.55 67.338 ;
        RECT 17.344 67.302 17.384 67.338 ;
        RECT 17.684 67.302 17.736 67.338 ;
        RECT 19.45 67.302 19.502 67.338 ;
        RECT 19.682 67.302 19.734 67.338 ;
        RECT 19.994 67.302 20.046 67.338 ;
        RECT 20.29 67.302 20.342 67.338 ;
        RECT 21.496 67.302 21.55 67.338 ;
        RECT 22.774 67.302 22.826 67.338 ;
        RECT 23.574 67.302 23.626 67.338 ;
        RECT 24.374 67.302 24.426 67.338 ;
        RECT 25.174 67.302 25.226 67.338 ;
        RECT 25.974 67.302 26.026 67.338 ;
        RECT 26.774 67.302 26.826 67.338 ;
        RECT 27.574 67.302 27.626 67.338 ;
        RECT 28.374 67.302 28.426 67.338 ;
        RECT 29.174 67.302 29.226 67.338 ;
        RECT 29.974 67.302 30.026 67.338 ;
        RECT 30.774 67.302 30.826 67.338 ;
        RECT 31.574 67.302 31.626 67.338 ;
        RECT 32.374 67.302 32.426 67.338 ;
        RECT 33.174 67.302 33.226 67.338 ;
        RECT 33.974 67.302 34.026 67.338 ;
        RECT 34.774 67.302 34.826 67.338 ;
        RECT 35.574 67.302 35.626 67.338 ;
        RECT 18.564 67.9075 18.636 67.9325 ;
        RECT 18.864 67.9075 18.936 67.9325 ;
        RECT 0.574 67.902 0.626 67.938 ;
        RECT 1.374 67.902 1.426 67.938 ;
        RECT 2.174 67.902 2.226 67.938 ;
        RECT 2.974 67.902 3.026 67.938 ;
        RECT 3.774 67.902 3.826 67.938 ;
        RECT 4.574 67.902 4.626 67.938 ;
        RECT 5.374 67.902 5.426 67.938 ;
        RECT 6.174 67.902 6.226 67.938 ;
        RECT 6.974 67.902 7.026 67.938 ;
        RECT 7.774 67.902 7.826 67.938 ;
        RECT 8.574 67.902 8.626 67.938 ;
        RECT 9.374 67.902 9.426 67.938 ;
        RECT 10.174 67.902 10.226 67.938 ;
        RECT 10.974 67.902 11.026 67.938 ;
        RECT 11.774 67.902 11.826 67.938 ;
        RECT 12.574 67.902 12.626 67.938 ;
        RECT 13.374 67.902 13.426 67.938 ;
        RECT 14.45 67.902 14.504 67.938 ;
        RECT 15.658 67.902 15.71 67.938 ;
        RECT 15.954 67.902 16.006 67.938 ;
        RECT 16.266 67.902 16.318 67.938 ;
        RECT 16.498 67.902 16.55 67.938 ;
        RECT 17.344 67.902 17.384 67.938 ;
        RECT 17.684 67.902 17.736 67.938 ;
        RECT 19.45 67.902 19.502 67.938 ;
        RECT 19.682 67.902 19.734 67.938 ;
        RECT 19.994 67.902 20.046 67.938 ;
        RECT 20.29 67.902 20.342 67.938 ;
        RECT 21.496 67.902 21.55 67.938 ;
        RECT 22.774 67.902 22.826 67.938 ;
        RECT 23.574 67.902 23.626 67.938 ;
        RECT 24.374 67.902 24.426 67.938 ;
        RECT 25.174 67.902 25.226 67.938 ;
        RECT 25.974 67.902 26.026 67.938 ;
        RECT 26.774 67.902 26.826 67.938 ;
        RECT 27.574 67.902 27.626 67.938 ;
        RECT 28.374 67.902 28.426 67.938 ;
        RECT 29.174 67.902 29.226 67.938 ;
        RECT 29.974 67.902 30.026 67.938 ;
        RECT 30.774 67.902 30.826 67.938 ;
        RECT 31.574 67.902 31.626 67.938 ;
        RECT 32.374 67.902 32.426 67.938 ;
        RECT 33.174 67.902 33.226 67.938 ;
        RECT 33.974 67.902 34.026 67.938 ;
        RECT 34.774 67.902 34.826 67.938 ;
        RECT 35.574 67.902 35.626 67.938 ;
        RECT 18.564 68.5075 18.636 68.5325 ;
        RECT 18.864 68.5075 18.936 68.5325 ;
        RECT 0.574 68.502 0.626 68.538 ;
        RECT 1.374 68.502 1.426 68.538 ;
        RECT 2.174 68.502 2.226 68.538 ;
        RECT 2.974 68.502 3.026 68.538 ;
        RECT 3.774 68.502 3.826 68.538 ;
        RECT 4.574 68.502 4.626 68.538 ;
        RECT 5.374 68.502 5.426 68.538 ;
        RECT 6.174 68.502 6.226 68.538 ;
        RECT 6.974 68.502 7.026 68.538 ;
        RECT 7.774 68.502 7.826 68.538 ;
        RECT 8.574 68.502 8.626 68.538 ;
        RECT 9.374 68.502 9.426 68.538 ;
        RECT 10.174 68.502 10.226 68.538 ;
        RECT 10.974 68.502 11.026 68.538 ;
        RECT 11.774 68.502 11.826 68.538 ;
        RECT 12.574 68.502 12.626 68.538 ;
        RECT 13.374 68.502 13.426 68.538 ;
        RECT 14.45 68.502 14.504 68.538 ;
        RECT 15.658 68.502 15.71 68.538 ;
        RECT 15.954 68.502 16.006 68.538 ;
        RECT 16.266 68.502 16.318 68.538 ;
        RECT 16.498 68.502 16.55 68.538 ;
        RECT 17.344 68.502 17.384 68.538 ;
        RECT 17.684 68.502 17.736 68.538 ;
        RECT 19.45 68.502 19.502 68.538 ;
        RECT 19.682 68.502 19.734 68.538 ;
        RECT 19.994 68.502 20.046 68.538 ;
        RECT 20.29 68.502 20.342 68.538 ;
        RECT 21.496 68.502 21.55 68.538 ;
        RECT 22.774 68.502 22.826 68.538 ;
        RECT 23.574 68.502 23.626 68.538 ;
        RECT 24.374 68.502 24.426 68.538 ;
        RECT 25.174 68.502 25.226 68.538 ;
        RECT 25.974 68.502 26.026 68.538 ;
        RECT 26.774 68.502 26.826 68.538 ;
        RECT 27.574 68.502 27.626 68.538 ;
        RECT 28.374 68.502 28.426 68.538 ;
        RECT 29.174 68.502 29.226 68.538 ;
        RECT 29.974 68.502 30.026 68.538 ;
        RECT 30.774 68.502 30.826 68.538 ;
        RECT 31.574 68.502 31.626 68.538 ;
        RECT 32.374 68.502 32.426 68.538 ;
        RECT 33.174 68.502 33.226 68.538 ;
        RECT 33.974 68.502 34.026 68.538 ;
        RECT 34.774 68.502 34.826 68.538 ;
        RECT 35.574 68.502 35.626 68.538 ;
        RECT 18.564 69.1075 18.636 69.1325 ;
        RECT 18.864 69.1075 18.936 69.1325 ;
        RECT 0.574 69.102 0.626 69.138 ;
        RECT 1.374 69.102 1.426 69.138 ;
        RECT 2.174 69.102 2.226 69.138 ;
        RECT 2.974 69.102 3.026 69.138 ;
        RECT 3.774 69.102 3.826 69.138 ;
        RECT 4.574 69.102 4.626 69.138 ;
        RECT 5.374 69.102 5.426 69.138 ;
        RECT 6.174 69.102 6.226 69.138 ;
        RECT 6.974 69.102 7.026 69.138 ;
        RECT 7.774 69.102 7.826 69.138 ;
        RECT 8.574 69.102 8.626 69.138 ;
        RECT 9.374 69.102 9.426 69.138 ;
        RECT 10.174 69.102 10.226 69.138 ;
        RECT 10.974 69.102 11.026 69.138 ;
        RECT 11.774 69.102 11.826 69.138 ;
        RECT 12.574 69.102 12.626 69.138 ;
        RECT 13.374 69.102 13.426 69.138 ;
        RECT 14.45 69.102 14.504 69.138 ;
        RECT 15.658 69.102 15.71 69.138 ;
        RECT 15.954 69.102 16.006 69.138 ;
        RECT 16.266 69.102 16.318 69.138 ;
        RECT 16.498 69.102 16.55 69.138 ;
        RECT 17.344 69.102 17.384 69.138 ;
        RECT 17.684 69.102 17.736 69.138 ;
        RECT 19.45 69.102 19.502 69.138 ;
        RECT 19.682 69.102 19.734 69.138 ;
        RECT 19.994 69.102 20.046 69.138 ;
        RECT 20.29 69.102 20.342 69.138 ;
        RECT 21.496 69.102 21.55 69.138 ;
        RECT 22.774 69.102 22.826 69.138 ;
        RECT 23.574 69.102 23.626 69.138 ;
        RECT 24.374 69.102 24.426 69.138 ;
        RECT 25.174 69.102 25.226 69.138 ;
        RECT 25.974 69.102 26.026 69.138 ;
        RECT 26.774 69.102 26.826 69.138 ;
        RECT 27.574 69.102 27.626 69.138 ;
        RECT 28.374 69.102 28.426 69.138 ;
        RECT 29.174 69.102 29.226 69.138 ;
        RECT 29.974 69.102 30.026 69.138 ;
        RECT 30.774 69.102 30.826 69.138 ;
        RECT 31.574 69.102 31.626 69.138 ;
        RECT 32.374 69.102 32.426 69.138 ;
        RECT 33.174 69.102 33.226 69.138 ;
        RECT 33.974 69.102 34.026 69.138 ;
        RECT 34.774 69.102 34.826 69.138 ;
        RECT 35.574 69.102 35.626 69.138 ;
        RECT 18.564 69.7075 18.636 69.7325 ;
        RECT 18.864 69.7075 18.936 69.7325 ;
        RECT 0.574 69.702 0.626 69.738 ;
        RECT 1.374 69.702 1.426 69.738 ;
        RECT 2.174 69.702 2.226 69.738 ;
        RECT 2.974 69.702 3.026 69.738 ;
        RECT 3.774 69.702 3.826 69.738 ;
        RECT 4.574 69.702 4.626 69.738 ;
        RECT 5.374 69.702 5.426 69.738 ;
        RECT 6.174 69.702 6.226 69.738 ;
        RECT 6.974 69.702 7.026 69.738 ;
        RECT 7.774 69.702 7.826 69.738 ;
        RECT 8.574 69.702 8.626 69.738 ;
        RECT 9.374 69.702 9.426 69.738 ;
        RECT 10.174 69.702 10.226 69.738 ;
        RECT 10.974 69.702 11.026 69.738 ;
        RECT 11.774 69.702 11.826 69.738 ;
        RECT 12.574 69.702 12.626 69.738 ;
        RECT 13.374 69.702 13.426 69.738 ;
        RECT 14.45 69.702 14.504 69.738 ;
        RECT 15.658 69.702 15.71 69.738 ;
        RECT 15.954 69.702 16.006 69.738 ;
        RECT 16.266 69.702 16.318 69.738 ;
        RECT 16.498 69.702 16.55 69.738 ;
        RECT 17.344 69.702 17.384 69.738 ;
        RECT 17.684 69.702 17.736 69.738 ;
        RECT 19.45 69.702 19.502 69.738 ;
        RECT 19.682 69.702 19.734 69.738 ;
        RECT 19.994 69.702 20.046 69.738 ;
        RECT 20.29 69.702 20.342 69.738 ;
        RECT 21.496 69.702 21.55 69.738 ;
        RECT 22.774 69.702 22.826 69.738 ;
        RECT 23.574 69.702 23.626 69.738 ;
        RECT 24.374 69.702 24.426 69.738 ;
        RECT 25.174 69.702 25.226 69.738 ;
        RECT 25.974 69.702 26.026 69.738 ;
        RECT 26.774 69.702 26.826 69.738 ;
        RECT 27.574 69.702 27.626 69.738 ;
        RECT 28.374 69.702 28.426 69.738 ;
        RECT 29.174 69.702 29.226 69.738 ;
        RECT 29.974 69.702 30.026 69.738 ;
        RECT 30.774 69.702 30.826 69.738 ;
        RECT 31.574 69.702 31.626 69.738 ;
        RECT 32.374 69.702 32.426 69.738 ;
        RECT 33.174 69.702 33.226 69.738 ;
        RECT 33.974 69.702 34.026 69.738 ;
        RECT 34.774 69.702 34.826 69.738 ;
        RECT 35.574 69.702 35.626 69.738 ;
        RECT 18.564 70.3075 18.636 70.3325 ;
        RECT 18.864 70.3075 18.936 70.3325 ;
        RECT 0.574 70.302 0.626 70.338 ;
        RECT 1.374 70.302 1.426 70.338 ;
        RECT 2.174 70.302 2.226 70.338 ;
        RECT 2.974 70.302 3.026 70.338 ;
        RECT 3.774 70.302 3.826 70.338 ;
        RECT 4.574 70.302 4.626 70.338 ;
        RECT 5.374 70.302 5.426 70.338 ;
        RECT 6.174 70.302 6.226 70.338 ;
        RECT 6.974 70.302 7.026 70.338 ;
        RECT 7.774 70.302 7.826 70.338 ;
        RECT 8.574 70.302 8.626 70.338 ;
        RECT 9.374 70.302 9.426 70.338 ;
        RECT 10.174 70.302 10.226 70.338 ;
        RECT 10.974 70.302 11.026 70.338 ;
        RECT 11.774 70.302 11.826 70.338 ;
        RECT 12.574 70.302 12.626 70.338 ;
        RECT 13.374 70.302 13.426 70.338 ;
        RECT 14.45 70.302 14.504 70.338 ;
        RECT 15.658 70.302 15.71 70.338 ;
        RECT 15.954 70.302 16.006 70.338 ;
        RECT 16.266 70.302 16.318 70.338 ;
        RECT 16.498 70.302 16.55 70.338 ;
        RECT 17.344 70.302 17.384 70.338 ;
        RECT 17.684 70.302 17.736 70.338 ;
        RECT 19.45 70.302 19.502 70.338 ;
        RECT 19.682 70.302 19.734 70.338 ;
        RECT 19.994 70.302 20.046 70.338 ;
        RECT 20.29 70.302 20.342 70.338 ;
        RECT 21.496 70.302 21.55 70.338 ;
        RECT 22.774 70.302 22.826 70.338 ;
        RECT 23.574 70.302 23.626 70.338 ;
        RECT 24.374 70.302 24.426 70.338 ;
        RECT 25.174 70.302 25.226 70.338 ;
        RECT 25.974 70.302 26.026 70.338 ;
        RECT 26.774 70.302 26.826 70.338 ;
        RECT 27.574 70.302 27.626 70.338 ;
        RECT 28.374 70.302 28.426 70.338 ;
        RECT 29.174 70.302 29.226 70.338 ;
        RECT 29.974 70.302 30.026 70.338 ;
        RECT 30.774 70.302 30.826 70.338 ;
        RECT 31.574 70.302 31.626 70.338 ;
        RECT 32.374 70.302 32.426 70.338 ;
        RECT 33.174 70.302 33.226 70.338 ;
        RECT 33.974 70.302 34.026 70.338 ;
        RECT 34.774 70.302 34.826 70.338 ;
        RECT 35.574 70.302 35.626 70.338 ;
        RECT 18.564 70.9075 18.636 70.9325 ;
        RECT 18.864 70.9075 18.936 70.9325 ;
        RECT 0.574 70.902 0.626 70.938 ;
        RECT 1.374 70.902 1.426 70.938 ;
        RECT 2.174 70.902 2.226 70.938 ;
        RECT 2.974 70.902 3.026 70.938 ;
        RECT 3.774 70.902 3.826 70.938 ;
        RECT 4.574 70.902 4.626 70.938 ;
        RECT 5.374 70.902 5.426 70.938 ;
        RECT 6.174 70.902 6.226 70.938 ;
        RECT 6.974 70.902 7.026 70.938 ;
        RECT 7.774 70.902 7.826 70.938 ;
        RECT 8.574 70.902 8.626 70.938 ;
        RECT 9.374 70.902 9.426 70.938 ;
        RECT 10.174 70.902 10.226 70.938 ;
        RECT 10.974 70.902 11.026 70.938 ;
        RECT 11.774 70.902 11.826 70.938 ;
        RECT 12.574 70.902 12.626 70.938 ;
        RECT 13.374 70.902 13.426 70.938 ;
        RECT 14.45 70.902 14.504 70.938 ;
        RECT 15.658 70.902 15.71 70.938 ;
        RECT 15.954 70.902 16.006 70.938 ;
        RECT 16.266 70.902 16.318 70.938 ;
        RECT 16.498 70.902 16.55 70.938 ;
        RECT 17.344 70.902 17.384 70.938 ;
        RECT 17.684 70.902 17.736 70.938 ;
        RECT 19.45 70.902 19.502 70.938 ;
        RECT 19.682 70.902 19.734 70.938 ;
        RECT 19.994 70.902 20.046 70.938 ;
        RECT 20.29 70.902 20.342 70.938 ;
        RECT 21.496 70.902 21.55 70.938 ;
        RECT 22.774 70.902 22.826 70.938 ;
        RECT 23.574 70.902 23.626 70.938 ;
        RECT 24.374 70.902 24.426 70.938 ;
        RECT 25.174 70.902 25.226 70.938 ;
        RECT 25.974 70.902 26.026 70.938 ;
        RECT 26.774 70.902 26.826 70.938 ;
        RECT 27.574 70.902 27.626 70.938 ;
        RECT 28.374 70.902 28.426 70.938 ;
        RECT 29.174 70.902 29.226 70.938 ;
        RECT 29.974 70.902 30.026 70.938 ;
        RECT 30.774 70.902 30.826 70.938 ;
        RECT 31.574 70.902 31.626 70.938 ;
        RECT 32.374 70.902 32.426 70.938 ;
        RECT 33.174 70.902 33.226 70.938 ;
        RECT 33.974 70.902 34.026 70.938 ;
        RECT 34.774 70.902 34.826 70.938 ;
        RECT 35.574 70.902 35.626 70.938 ;
        RECT 18.564 71.5075 18.636 71.5325 ;
        RECT 18.864 71.5075 18.936 71.5325 ;
        RECT 0.574 71.502 0.626 71.538 ;
        RECT 1.374 71.502 1.426 71.538 ;
        RECT 2.174 71.502 2.226 71.538 ;
        RECT 2.974 71.502 3.026 71.538 ;
        RECT 3.774 71.502 3.826 71.538 ;
        RECT 4.574 71.502 4.626 71.538 ;
        RECT 5.374 71.502 5.426 71.538 ;
        RECT 6.174 71.502 6.226 71.538 ;
        RECT 6.974 71.502 7.026 71.538 ;
        RECT 7.774 71.502 7.826 71.538 ;
        RECT 8.574 71.502 8.626 71.538 ;
        RECT 9.374 71.502 9.426 71.538 ;
        RECT 10.174 71.502 10.226 71.538 ;
        RECT 10.974 71.502 11.026 71.538 ;
        RECT 11.774 71.502 11.826 71.538 ;
        RECT 12.574 71.502 12.626 71.538 ;
        RECT 13.374 71.502 13.426 71.538 ;
        RECT 14.45 71.502 14.504 71.538 ;
        RECT 15.658 71.502 15.71 71.538 ;
        RECT 15.954 71.502 16.006 71.538 ;
        RECT 16.266 71.502 16.318 71.538 ;
        RECT 16.498 71.502 16.55 71.538 ;
        RECT 17.344 71.502 17.384 71.538 ;
        RECT 17.684 71.502 17.736 71.538 ;
        RECT 19.45 71.502 19.502 71.538 ;
        RECT 19.682 71.502 19.734 71.538 ;
        RECT 19.994 71.502 20.046 71.538 ;
        RECT 20.29 71.502 20.342 71.538 ;
        RECT 21.496 71.502 21.55 71.538 ;
        RECT 22.774 71.502 22.826 71.538 ;
        RECT 23.574 71.502 23.626 71.538 ;
        RECT 24.374 71.502 24.426 71.538 ;
        RECT 25.174 71.502 25.226 71.538 ;
        RECT 25.974 71.502 26.026 71.538 ;
        RECT 26.774 71.502 26.826 71.538 ;
        RECT 27.574 71.502 27.626 71.538 ;
        RECT 28.374 71.502 28.426 71.538 ;
        RECT 29.174 71.502 29.226 71.538 ;
        RECT 29.974 71.502 30.026 71.538 ;
        RECT 30.774 71.502 30.826 71.538 ;
        RECT 31.574 71.502 31.626 71.538 ;
        RECT 32.374 71.502 32.426 71.538 ;
        RECT 33.174 71.502 33.226 71.538 ;
        RECT 33.974 71.502 34.026 71.538 ;
        RECT 34.774 71.502 34.826 71.538 ;
        RECT 35.574 71.502 35.626 71.538 ;
        RECT 18.564 72.1075 18.636 72.1325 ;
        RECT 18.864 72.1075 18.936 72.1325 ;
        RECT 0.574 72.102 0.626 72.138 ;
        RECT 1.374 72.102 1.426 72.138 ;
        RECT 2.174 72.102 2.226 72.138 ;
        RECT 2.974 72.102 3.026 72.138 ;
        RECT 3.774 72.102 3.826 72.138 ;
        RECT 4.574 72.102 4.626 72.138 ;
        RECT 5.374 72.102 5.426 72.138 ;
        RECT 6.174 72.102 6.226 72.138 ;
        RECT 6.974 72.102 7.026 72.138 ;
        RECT 7.774 72.102 7.826 72.138 ;
        RECT 8.574 72.102 8.626 72.138 ;
        RECT 9.374 72.102 9.426 72.138 ;
        RECT 10.174 72.102 10.226 72.138 ;
        RECT 10.974 72.102 11.026 72.138 ;
        RECT 11.774 72.102 11.826 72.138 ;
        RECT 12.574 72.102 12.626 72.138 ;
        RECT 13.374 72.102 13.426 72.138 ;
        RECT 14.45 72.102 14.504 72.138 ;
        RECT 15.658 72.102 15.71 72.138 ;
        RECT 15.954 72.102 16.006 72.138 ;
        RECT 16.266 72.102 16.318 72.138 ;
        RECT 16.498 72.102 16.55 72.138 ;
        RECT 17.344 72.102 17.384 72.138 ;
        RECT 17.684 72.102 17.736 72.138 ;
        RECT 19.45 72.102 19.502 72.138 ;
        RECT 19.682 72.102 19.734 72.138 ;
        RECT 19.994 72.102 20.046 72.138 ;
        RECT 20.29 72.102 20.342 72.138 ;
        RECT 21.496 72.102 21.55 72.138 ;
        RECT 22.774 72.102 22.826 72.138 ;
        RECT 23.574 72.102 23.626 72.138 ;
        RECT 24.374 72.102 24.426 72.138 ;
        RECT 25.174 72.102 25.226 72.138 ;
        RECT 25.974 72.102 26.026 72.138 ;
        RECT 26.774 72.102 26.826 72.138 ;
        RECT 27.574 72.102 27.626 72.138 ;
        RECT 28.374 72.102 28.426 72.138 ;
        RECT 29.174 72.102 29.226 72.138 ;
        RECT 29.974 72.102 30.026 72.138 ;
        RECT 30.774 72.102 30.826 72.138 ;
        RECT 31.574 72.102 31.626 72.138 ;
        RECT 32.374 72.102 32.426 72.138 ;
        RECT 33.174 72.102 33.226 72.138 ;
        RECT 33.974 72.102 34.026 72.138 ;
        RECT 34.774 72.102 34.826 72.138 ;
        RECT 35.574 72.102 35.626 72.138 ;
      LAYER m5 ;
        RECT 17.344 0.5695 17.384 32.14 ;
        RECT 16.882 32.353 16.936 39.1925 ;
        RECT 19.228 31.84 19.282 39.68 ;
        RECT 17.204 31.82 17.244 39.7 ;
        RECT 18.216 31.82 18.256 39.7 ;
        RECT 0.574 0.5695 0.626 72.1505 ;
        RECT 1.374 0.5695 1.426 72.1505 ;
        RECT 2.174 0.5695 2.226 72.1505 ;
        RECT 2.974 0.5695 3.026 72.1505 ;
        RECT 3.774 0.5695 3.826 72.1505 ;
        RECT 4.574 0.5695 4.626 72.1505 ;
        RECT 5.374 0.5695 5.426 72.1505 ;
        RECT 6.174 0.5695 6.226 72.1505 ;
        RECT 6.974 0.5695 7.026 72.1505 ;
        RECT 7.774 0.5695 7.826 72.1505 ;
        RECT 8.574 0.5695 8.626 72.1505 ;
        RECT 9.374 0.5695 9.426 72.1505 ;
        RECT 10.174 0.5695 10.226 72.1505 ;
        RECT 10.974 0.5695 11.026 72.1505 ;
        RECT 11.774 0.5695 11.826 72.1505 ;
        RECT 12.574 0.5695 12.626 72.1505 ;
        RECT 13.374 0.5695 13.426 72.1505 ;
        RECT 14.45 0.5695 14.504 72.1505 ;
        RECT 15.658 0.5695 15.71 72.1505 ;
        RECT 15.954 0.5695 16.006 72.1505 ;
        RECT 16.266 0.5695 16.318 72.1505 ;
        RECT 16.498 0.5695 16.55 72.1505 ;
        RECT 17.344 39.38 17.384 72.1505 ;
        RECT 17.684 0.5695 17.736 72.1505 ;
        RECT 18.564 0.5695 18.636 72.1505 ;
        RECT 18.864 0.5695 18.936 72.1505 ;
        RECT 19.45 0.5695 19.502 72.1505 ;
        RECT 19.682 0.5695 19.734 72.1505 ;
        RECT 19.994 0.5695 20.046 72.1505 ;
        RECT 20.29 0.5695 20.342 72.1505 ;
        RECT 21.496 0.5695 21.55 72.1505 ;
        RECT 22.774 0.5695 22.826 72.1505 ;
        RECT 23.574 0.5695 23.626 72.1505 ;
        RECT 24.374 0.5695 24.426 72.1505 ;
        RECT 25.174 0.5695 25.226 72.1505 ;
        RECT 25.974 0.5695 26.026 72.1505 ;
        RECT 26.774 0.5695 26.826 72.1505 ;
        RECT 27.574 0.5695 27.626 72.1505 ;
        RECT 28.374 0.5695 28.426 72.1505 ;
        RECT 29.174 0.5695 29.226 72.1505 ;
        RECT 29.974 0.5695 30.026 72.1505 ;
        RECT 30.774 0.5695 30.826 72.1505 ;
        RECT 31.574 0.5695 31.626 72.1505 ;
        RECT 32.374 0.5695 32.426 72.1505 ;
        RECT 33.174 0.5695 33.226 72.1505 ;
        RECT 33.974 0.5695 34.026 72.1505 ;
        RECT 34.774 0.5695 34.826 72.1505 ;
        RECT 35.574 0.5695 35.626 72.1505 ;
    END
  END vss
  OBS
    LAYER m0 ;
      RECT 0 0 36.3 72.72 ;
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 36.316 72.734 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 36.32 72.74 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 36.3705 72.758 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 36.335 72.79 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 36.37 72.758 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 72.1505 36.359 72.81 ;
      RECT 17.036 72.1 17.344 72.1505 ;
      RECT 17.384 72.1 17.684 72.1505 ;
      RECT 17.036 70.94 17.136 72.1 ;
      RECT 17.176 70.94 17.344 72.1 ;
      RECT 17.384 70.94 17.412 72.1 ;
      RECT 17.452 70.94 17.684 72.1 ;
      RECT 17.036 70.9 17.344 70.94 ;
      RECT 17.384 70.9 17.684 70.94 ;
      RECT 17.036 69.74 17.136 70.9 ;
      RECT 17.176 69.74 17.344 70.9 ;
      RECT 17.384 69.74 17.412 70.9 ;
      RECT 17.452 69.74 17.684 70.9 ;
      RECT 17.036 69.7 17.344 69.74 ;
      RECT 17.384 69.7 17.684 69.74 ;
      RECT 17.036 68.54 17.136 69.7 ;
      RECT 17.176 68.54 17.344 69.7 ;
      RECT 17.384 68.54 17.412 69.7 ;
      RECT 17.452 68.54 17.684 69.7 ;
      RECT 17.036 68.5 17.344 68.54 ;
      RECT 17.384 68.5 17.684 68.54 ;
      RECT 17.036 67.34 17.136 68.5 ;
      RECT 17.176 67.34 17.344 68.5 ;
      RECT 17.384 67.34 17.412 68.5 ;
      RECT 17.452 67.34 17.684 68.5 ;
      RECT 17.036 67.3 17.344 67.34 ;
      RECT 17.384 67.3 17.684 67.34 ;
      RECT 17.036 66.14 17.136 67.3 ;
      RECT 17.176 66.14 17.344 67.3 ;
      RECT 17.384 66.14 17.412 67.3 ;
      RECT 17.452 66.14 17.684 67.3 ;
      RECT 17.036 66.1 17.344 66.14 ;
      RECT 17.384 66.1 17.684 66.14 ;
      RECT 17.036 64.94 17.136 66.1 ;
      RECT 17.176 64.94 17.344 66.1 ;
      RECT 17.384 64.94 17.412 66.1 ;
      RECT 17.452 64.94 17.684 66.1 ;
      RECT 17.036 64.9 17.344 64.94 ;
      RECT 17.384 64.9 17.684 64.94 ;
      RECT 17.036 63.74 17.136 64.9 ;
      RECT 17.176 63.74 17.344 64.9 ;
      RECT 17.384 63.74 17.412 64.9 ;
      RECT 17.452 63.74 17.684 64.9 ;
      RECT 17.036 63.7 17.344 63.74 ;
      RECT 17.384 63.7 17.684 63.74 ;
      RECT 17.036 62.54 17.136 63.7 ;
      RECT 17.176 62.54 17.344 63.7 ;
      RECT 17.384 62.54 17.412 63.7 ;
      RECT 17.452 62.54 17.684 63.7 ;
      RECT 17.036 62.5 17.344 62.54 ;
      RECT 17.384 62.5 17.684 62.54 ;
      RECT 17.036 61.34 17.136 62.5 ;
      RECT 17.176 61.34 17.344 62.5 ;
      RECT 17.384 61.34 17.412 62.5 ;
      RECT 17.452 61.34 17.684 62.5 ;
      RECT 17.036 61.3 17.344 61.34 ;
      RECT 17.384 61.3 17.684 61.34 ;
      RECT 17.036 60.14 17.136 61.3 ;
      RECT 17.176 60.14 17.344 61.3 ;
      RECT 17.384 60.14 17.412 61.3 ;
      RECT 17.452 60.14 17.684 61.3 ;
      RECT 17.036 60.1 17.344 60.14 ;
      RECT 17.384 60.1 17.684 60.14 ;
      RECT 17.036 58.94 17.136 60.1 ;
      RECT 17.176 58.94 17.344 60.1 ;
      RECT 17.384 58.94 17.412 60.1 ;
      RECT 17.452 58.94 17.684 60.1 ;
      RECT 17.036 58.9 17.344 58.94 ;
      RECT 17.384 58.9 17.684 58.94 ;
      RECT 17.036 57.74 17.136 58.9 ;
      RECT 17.176 57.74 17.344 58.9 ;
      RECT 17.384 57.74 17.412 58.9 ;
      RECT 17.452 57.74 17.684 58.9 ;
      RECT 17.036 57.7 17.344 57.74 ;
      RECT 17.384 57.7 17.684 57.74 ;
      RECT 17.036 56.54 17.136 57.7 ;
      RECT 17.176 56.54 17.344 57.7 ;
      RECT 17.384 56.54 17.412 57.7 ;
      RECT 17.452 56.54 17.684 57.7 ;
      RECT 17.036 56.5 17.344 56.54 ;
      RECT 17.384 56.5 17.684 56.54 ;
      RECT 17.036 55.34 17.136 56.5 ;
      RECT 17.176 55.34 17.344 56.5 ;
      RECT 17.384 55.34 17.412 56.5 ;
      RECT 17.452 55.34 17.684 56.5 ;
      RECT 17.036 55.3 17.344 55.34 ;
      RECT 17.384 55.3 17.684 55.34 ;
      RECT 17.036 54.14 17.136 55.3 ;
      RECT 17.176 54.14 17.344 55.3 ;
      RECT 17.384 54.14 17.412 55.3 ;
      RECT 17.452 54.14 17.684 55.3 ;
      RECT 17.036 54.1 17.344 54.14 ;
      RECT 17.384 54.1 17.684 54.14 ;
      RECT 17.036 52.94 17.136 54.1 ;
      RECT 17.176 52.94 17.344 54.1 ;
      RECT 17.384 52.94 17.412 54.1 ;
      RECT 17.452 52.94 17.684 54.1 ;
      RECT 17.036 52.9 17.344 52.94 ;
      RECT 17.384 52.9 17.684 52.94 ;
      RECT 17.036 51.74 17.136 52.9 ;
      RECT 17.176 51.74 17.344 52.9 ;
      RECT 17.384 51.74 17.412 52.9 ;
      RECT 17.452 51.74 17.684 52.9 ;
      RECT 17.036 51.7 17.344 51.74 ;
      RECT 17.384 51.7 17.684 51.74 ;
      RECT 17.036 50.54 17.136 51.7 ;
      RECT 17.176 50.54 17.344 51.7 ;
      RECT 17.384 50.54 17.412 51.7 ;
      RECT 17.452 50.54 17.684 51.7 ;
      RECT 17.036 50.5 17.344 50.54 ;
      RECT 17.384 50.5 17.684 50.54 ;
      RECT 17.036 49.34 17.136 50.5 ;
      RECT 17.176 49.34 17.344 50.5 ;
      RECT 17.384 49.34 17.412 50.5 ;
      RECT 17.452 49.34 17.684 50.5 ;
      RECT 17.036 49.3 17.344 49.34 ;
      RECT 17.384 49.3 17.684 49.34 ;
      RECT 17.036 48.14 17.136 49.3 ;
      RECT 17.176 48.14 17.344 49.3 ;
      RECT 17.384 48.14 17.412 49.3 ;
      RECT 17.452 48.14 17.684 49.3 ;
      RECT 17.036 48.1 17.344 48.14 ;
      RECT 17.384 48.1 17.684 48.14 ;
      RECT 17.036 46.94 17.136 48.1 ;
      RECT 17.176 46.94 17.344 48.1 ;
      RECT 17.384 46.94 17.412 48.1 ;
      RECT 17.452 46.94 17.684 48.1 ;
      RECT 17.036 46.9 17.344 46.94 ;
      RECT 17.384 46.9 17.684 46.94 ;
      RECT 17.036 45.74 17.136 46.9 ;
      RECT 17.176 45.74 17.344 46.9 ;
      RECT 17.384 45.74 17.412 46.9 ;
      RECT 17.452 45.74 17.684 46.9 ;
      RECT 17.036 45.7 17.344 45.74 ;
      RECT 17.384 45.7 17.684 45.74 ;
      RECT 17.036 44.54 17.136 45.7 ;
      RECT 17.176 44.54 17.344 45.7 ;
      RECT 17.384 44.54 17.412 45.7 ;
      RECT 17.452 44.54 17.684 45.7 ;
      RECT 17.036 44.5 17.344 44.54 ;
      RECT 17.384 44.5 17.684 44.54 ;
      RECT 17.036 43.34 17.136 44.5 ;
      RECT 17.176 43.34 17.344 44.5 ;
      RECT 17.384 43.34 17.412 44.5 ;
      RECT 17.452 43.34 17.684 44.5 ;
      RECT 17.036 43.3 17.344 43.34 ;
      RECT 17.384 43.3 17.684 43.34 ;
      RECT 17.036 42.14 17.136 43.3 ;
      RECT 17.176 42.14 17.344 43.3 ;
      RECT 17.384 42.14 17.412 43.3 ;
      RECT 17.452 42.14 17.684 43.3 ;
      RECT 17.036 42.1 17.344 42.14 ;
      RECT 17.384 42.1 17.684 42.14 ;
      RECT 17.036 40.94 17.136 42.1 ;
      RECT 17.176 40.94 17.344 42.1 ;
      RECT 17.384 40.94 17.412 42.1 ;
      RECT 17.452 40.94 17.684 42.1 ;
      RECT 17.036 40.9 17.344 40.94 ;
      RECT 17.384 40.9 17.684 40.94 ;
      RECT 20.046 72.12 20.29 72.1505 ;
      RECT 17.036 39.74 17.136 40.9 ;
      RECT 17.176 39.74 17.344 40.9 ;
      RECT 17.384 39.74 17.412 40.9 ;
      RECT 17.452 39.74 17.684 40.9 ;
      RECT 19.036 39.72 19.45 72.1505 ;
      RECT 18.188 39.7 18.356 72.1505 ;
      RECT 17.036 39.7 17.344 39.74 ;
      RECT 17.384 39.38 17.684 39.74 ;
      RECT 17.244 39.38 17.344 39.7 ;
      RECT 17.244 39.34 17.684 39.38 ;
      RECT 26.826 72.12 27.574 72.1505 ;
      RECT 31.626 72.12 32.374 72.1505 ;
      RECT 32.426 72.12 33.174 72.1505 ;
      RECT 33.226 72.12 33.974 72.1505 ;
      RECT 34.026 72.12 34.774 72.1505 ;
      RECT 34.826 72.12 35.574 72.1505 ;
      RECT 27.626 72.12 28.374 72.1505 ;
      RECT 28.426 72.12 29.174 72.1505 ;
      RECT 29.226 72.12 29.974 72.1505 ;
      RECT 30.026 72.12 30.774 72.1505 ;
      RECT 30.826 72.12 31.574 72.1505 ;
      RECT 22.826 72.12 23.574 72.1505 ;
      RECT 23.626 72.12 24.374 72.1505 ;
      RECT 24.426 72.12 25.174 72.1505 ;
      RECT 25.226 72.12 25.974 72.1505 ;
      RECT 26.026 72.12 26.774 72.1505 ;
      RECT 19.036 39.68 19.31 39.72 ;
      RECT 8.626 72.12 9.374 72.1505 ;
      RECT 15.71 72.12 15.954 72.1505 ;
      RECT 9.426 72.12 10.174 72.1505 ;
      RECT 10.226 72.12 10.974 72.1505 ;
      RECT 11.026 72.12 11.774 72.1505 ;
      RECT 11.826 72.12 12.574 72.1505 ;
      RECT 12.626 72.12 13.374 72.1505 ;
      RECT 3.826 72.12 4.574 72.1505 ;
      RECT 4.626 72.12 5.374 72.1505 ;
      RECT 5.426 72.12 6.174 72.1505 ;
      RECT 6.226 72.12 6.974 72.1505 ;
      RECT 7.026 72.12 7.774 72.1505 ;
      RECT 7.826 72.12 8.574 72.1505 ;
      RECT 0.626 72.12 1.374 72.1505 ;
      RECT 1.426 72.12 2.174 72.1505 ;
      RECT 2.226 72.12 2.974 72.1505 ;
      RECT 3.026 72.12 3.774 72.1505 ;
      RECT 16.854 39.1925 16.964 72.1505 ;
      RECT 17.452 38.93 17.684 39.34 ;
      RECT 17.036 38.81 17.204 39.7 ;
      RECT 17.244 38.81 17.412 39.34 ;
      RECT 17.52 38.81 17.684 38.93 ;
      RECT 17.452 37.97 17.48 38.93 ;
      RECT 17.52 37.97 17.548 38.81 ;
      RECT 17.452 37.93 17.548 37.97 ;
      RECT 17.036 37.85 17.136 38.81 ;
      RECT 17.176 37.85 17.204 38.81 ;
      RECT 17.244 37.85 17.344 38.81 ;
      RECT 17.384 37.85 17.412 38.81 ;
      RECT 17.588 37.85 17.616 38.81 ;
      RECT 17.656 37.85 17.684 38.81 ;
      RECT 17.52 37.85 17.548 37.93 ;
      RECT 31.626 38.5695 31.974 72.12 ;
      RECT 34.026 38.5695 34.374 72.12 ;
      RECT 34.826 38.5695 35.174 72.12 ;
      RECT 32.426 38.5695 32.774 72.12 ;
      RECT 33.226 38.5695 33.574 72.12 ;
      RECT 29.226 38.5695 29.574 72.12 ;
      RECT 30.026 38.5695 30.374 72.12 ;
      RECT 30.826 38.5695 31.174 72.12 ;
      RECT 27.626 38.5695 27.974 72.12 ;
      RECT 28.426 38.5695 28.774 72.12 ;
      RECT 25.226 38.5695 25.574 72.12 ;
      RECT 26.026 38.5695 26.374 72.12 ;
      RECT 26.826 38.5695 27.174 72.12 ;
      RECT 22.826 38.5695 23.174 72.12 ;
      RECT 23.626 38.5695 23.974 72.12 ;
      RECT 24.426 38.5695 24.774 72.12 ;
      RECT 20.342 38.199 20.47 72.1505 ;
      RECT 20.522 38.199 20.63 72.1505 ;
      RECT 15.37 38.199 15.478 72.1505 ;
      RECT 15.53 38.199 15.658 72.1505 ;
      RECT 11.026 38.5695 11.374 72.12 ;
      RECT 11.826 38.5695 12.174 72.12 ;
      RECT 12.626 38.5695 12.974 72.12 ;
      RECT 9.426 38.5695 9.774 72.12 ;
      RECT 10.226 38.5695 10.574 72.12 ;
      RECT 7.026 38.5695 7.374 72.12 ;
      RECT 7.826 38.5695 8.174 72.12 ;
      RECT 8.626 38.5695 8.974 72.12 ;
      RECT 4.626 38.5695 4.974 72.12 ;
      RECT 5.426 38.5695 5.774 72.12 ;
      RECT 6.226 38.5695 6.574 72.12 ;
      RECT 2.226 38.5695 2.574 72.12 ;
      RECT 3.026 38.5695 3.374 72.12 ;
      RECT 3.826 38.5695 4.174 72.12 ;
      RECT 0.626 38.5695 0.974 72.12 ;
      RECT 1.426 38.5695 1.774 72.12 ;
      RECT 17.036 37.81 17.204 37.85 ;
      RECT 17.244 37.81 17.412 37.85 ;
      RECT 17.452 36.97 17.48 37.93 ;
      RECT 17.52 36.97 17.548 37.81 ;
      RECT 17.916 37.81 18.148 72.1505 ;
      RECT 18.396 37.81 18.564 72.1505 ;
      RECT 17.036 36.85 17.136 37.81 ;
      RECT 17.176 36.85 17.204 37.81 ;
      RECT 17.244 36.85 17.344 37.81 ;
      RECT 17.384 36.85 17.412 37.81 ;
      RECT 17.452 36.85 17.548 36.97 ;
      RECT 17.52 37.81 17.684 37.85 ;
      RECT 17.588 36.85 17.616 37.81 ;
      RECT 17.656 36.85 17.684 37.81 ;
      RECT 17.916 36.85 17.944 37.81 ;
      RECT 17.984 36.85 18.012 37.81 ;
      RECT 18.052 36.85 18.08 37.81 ;
      RECT 18.12 36.85 18.148 37.81 ;
      RECT 17.036 36.81 17.204 36.85 ;
      RECT 17.244 36.81 17.412 36.85 ;
      RECT 17.452 36.81 17.684 36.85 ;
      RECT 17.036 35.85 17.136 36.81 ;
      RECT 17.176 35.85 17.204 36.81 ;
      RECT 17.244 35.85 17.344 36.81 ;
      RECT 17.384 35.85 17.412 36.81 ;
      RECT 17.452 35.85 17.616 36.81 ;
      RECT 17.656 35.85 17.684 36.81 ;
      RECT 17.036 35.26 17.204 35.85 ;
      RECT 17.452 35.26 17.684 35.85 ;
      RECT 18.396 36.85 18.424 37.81 ;
      RECT 18.464 36.85 18.564 37.81 ;
      RECT 17.244 35.14 17.412 35.85 ;
      RECT 17.036 35.14 17.136 35.26 ;
      RECT 17.52 35.14 17.684 35.26 ;
      RECT 17.916 35.14 18.148 36.85 ;
      RECT 17.176 34.3 17.204 35.26 ;
      RECT 17.452 34.3 17.48 35.26 ;
      RECT 17.108 34.3 17.136 35.14 ;
      RECT 17.52 34.3 17.616 35.14 ;
      RECT 17.108 34.26 17.204 34.3 ;
      RECT 17.452 34.26 17.616 34.3 ;
      RECT 18.256 35.14 18.356 39.7 ;
      RECT 17.036 34.18 17.064 35.14 ;
      RECT 17.244 34.18 17.272 35.14 ;
      RECT 17.316 34.18 17.344 35.14 ;
      RECT 17.384 34.18 17.412 35.14 ;
      RECT 17.108 34.18 17.136 34.26 ;
      RECT 17.656 34.18 17.684 35.14 ;
      RECT 17.916 34.18 18.012 35.14 ;
      RECT 18.052 34.18 18.148 35.14 ;
      RECT 18.256 34.18 18.284 35.14 ;
      RECT 18.328 34.18 18.356 35.14 ;
      RECT 17.244 34.14 17.412 34.18 ;
      RECT 17.52 34.18 17.616 34.26 ;
      RECT 17.916 34.14 18.148 34.18 ;
      RECT 17.176 33.3 17.204 34.26 ;
      RECT 17.452 33.3 17.48 34.26 ;
      RECT 17.036 33.3 17.136 34.18 ;
      RECT 18.256 34.14 18.356 34.18 ;
      RECT 17.244 33.18 17.272 34.14 ;
      RECT 17.316 33.18 17.412 34.14 ;
      RECT 17.52 33.3 17.684 34.18 ;
      RECT 17.916 33.18 17.944 34.14 ;
      RECT 17.984 33.18 18.012 34.14 ;
      RECT 18.052 33.18 18.148 34.14 ;
      RECT 18.256 33.18 18.284 34.14 ;
      RECT 18.328 33.18 18.356 34.14 ;
      RECT 18.256 33.14 18.356 33.18 ;
      RECT 17.452 33.14 17.684 33.3 ;
      RECT 17.244 33.14 17.412 33.18 ;
      RECT 31.706 32.9505 31.974 38.5695 ;
      RECT 34.106 32.9505 34.374 38.5695 ;
      RECT 34.826 32.9505 34.854 38.5695 ;
      RECT 34.906 32.9505 35.174 38.5695 ;
      RECT 32.426 32.9505 32.454 38.5695 ;
      RECT 32.506 32.9505 32.774 38.5695 ;
      RECT 33.226 32.9505 33.254 38.5695 ;
      RECT 33.306 32.9505 33.574 38.5695 ;
      RECT 34.026 32.9505 34.054 38.5695 ;
      RECT 29.306 32.9505 29.574 38.5695 ;
      RECT 30.026 32.9505 30.054 38.5695 ;
      RECT 30.106 32.9505 30.374 38.5695 ;
      RECT 30.826 32.9505 30.854 38.5695 ;
      RECT 30.906 32.9505 31.174 38.5695 ;
      RECT 31.626 32.9505 31.654 38.5695 ;
      RECT 27.626 32.9505 27.654 38.5695 ;
      RECT 27.706 32.9505 27.974 38.5695 ;
      RECT 28.426 32.9505 28.454 38.5695 ;
      RECT 28.506 32.9505 28.774 38.5695 ;
      RECT 29.226 32.9505 29.254 38.5695 ;
      RECT 25.226 32.9505 25.254 38.5695 ;
      RECT 25.306 32.9505 25.574 38.5695 ;
      RECT 26.026 32.9505 26.054 38.5695 ;
      RECT 26.106 32.9505 26.374 38.5695 ;
      RECT 26.826 32.9505 26.854 38.5695 ;
      RECT 26.906 32.9505 27.174 38.5695 ;
      RECT 22.826 32.9505 22.854 38.5695 ;
      RECT 22.906 32.9505 23.174 38.5695 ;
      RECT 23.626 32.9505 23.654 38.5695 ;
      RECT 23.706 32.9505 23.974 38.5695 ;
      RECT 24.426 32.9505 24.454 38.5695 ;
      RECT 24.506 32.9505 24.774 38.5695 ;
      RECT 20.342 32.8595 20.63 38.199 ;
      RECT 16.854 32.353 16.882 39.1925 ;
      RECT 16.936 32.353 16.964 39.1925 ;
      RECT 15.37 32.8595 15.658 38.199 ;
      RECT 11.106 32.9505 11.374 38.5695 ;
      RECT 11.826 32.9505 11.854 38.5695 ;
      RECT 11.906 32.9505 12.174 38.5695 ;
      RECT 12.626 32.9505 12.654 38.5695 ;
      RECT 12.706 32.9505 12.974 38.5695 ;
      RECT 9.426 32.9505 9.454 38.5695 ;
      RECT 9.506 32.9505 9.774 38.5695 ;
      RECT 10.226 32.9505 10.254 38.5695 ;
      RECT 10.306 32.9505 10.574 38.5695 ;
      RECT 11.026 32.9505 11.054 38.5695 ;
      RECT 7.026 32.9505 7.054 38.5695 ;
      RECT 7.106 32.9505 7.374 38.5695 ;
      RECT 7.826 32.9505 7.854 38.5695 ;
      RECT 7.906 32.9505 8.174 38.5695 ;
      RECT 8.626 32.9505 8.654 38.5695 ;
      RECT 8.706 32.9505 8.974 38.5695 ;
      RECT 4.626 32.9505 4.654 38.5695 ;
      RECT 4.706 32.9505 4.974 38.5695 ;
      RECT 5.426 32.9505 5.454 38.5695 ;
      RECT 5.506 32.9505 5.774 38.5695 ;
      RECT 6.226 32.9505 6.254 38.5695 ;
      RECT 6.306 32.9505 6.574 38.5695 ;
      RECT 2.226 32.9505 2.254 38.5695 ;
      RECT 2.306 32.9505 2.574 38.5695 ;
      RECT 3.026 32.9505 3.054 38.5695 ;
      RECT 3.106 32.9505 3.374 38.5695 ;
      RECT 3.826 32.9505 3.854 38.5695 ;
      RECT 3.906 32.9505 4.174 38.5695 ;
      RECT 0.626 32.9505 0.654 38.5695 ;
      RECT 0.706 32.9505 0.974 38.5695 ;
      RECT 1.426 32.9505 1.454 38.5695 ;
      RECT 1.506 32.9505 1.774 38.5695 ;
      RECT 17.244 32.18 17.344 33.14 ;
      RECT 17.384 32.18 17.412 33.14 ;
      RECT 17.452 32.18 17.548 33.14 ;
      RECT 17.588 32.18 17.616 33.14 ;
      RECT 17.656 32.18 17.684 33.14 ;
      RECT 18.256 32.18 18.284 33.14 ;
      RECT 18.328 32.18 18.356 33.14 ;
      RECT 17.244 32.14 17.684 32.18 ;
      RECT 19.036 31.84 19.228 39.68 ;
      RECT 19.282 31.84 19.31 39.68 ;
      RECT 18.188 31.82 18.216 39.7 ;
      RECT 18.256 31.82 18.356 32.18 ;
      RECT 17.036 31.82 17.204 33.3 ;
      RECT 17.244 31.82 17.344 32.14 ;
      RECT 17.384 31.78 17.684 32.14 ;
      RECT 17.036 31.78 17.344 31.82 ;
      RECT 17.036 30.62 17.136 31.78 ;
      RECT 17.176 30.62 17.344 31.78 ;
      RECT 17.384 30.62 17.412 31.78 ;
      RECT 17.452 30.62 17.684 31.78 ;
      RECT 17.384 30.58 17.684 30.62 ;
      RECT 17.036 30.58 17.344 30.62 ;
      RECT 17.036 29.42 17.136 30.58 ;
      RECT 17.176 29.42 17.344 30.58 ;
      RECT 17.384 29.42 17.412 30.58 ;
      RECT 17.452 29.42 17.684 30.58 ;
      RECT 17.384 29.38 17.684 29.42 ;
      RECT 17.036 29.38 17.344 29.42 ;
      RECT 17.036 28.22 17.136 29.38 ;
      RECT 17.176 28.22 17.344 29.38 ;
      RECT 17.384 28.22 17.412 29.38 ;
      RECT 17.452 28.22 17.684 29.38 ;
      RECT 17.384 28.18 17.684 28.22 ;
      RECT 17.036 28.18 17.344 28.22 ;
      RECT 17.036 27.02 17.136 28.18 ;
      RECT 17.176 27.02 17.344 28.18 ;
      RECT 17.384 27.02 17.412 28.18 ;
      RECT 17.452 27.02 17.684 28.18 ;
      RECT 17.384 26.98 17.684 27.02 ;
      RECT 17.036 26.98 17.344 27.02 ;
      RECT 17.036 25.82 17.136 26.98 ;
      RECT 17.176 25.82 17.344 26.98 ;
      RECT 17.384 25.82 17.412 26.98 ;
      RECT 17.452 25.82 17.684 26.98 ;
      RECT 17.384 25.78 17.684 25.82 ;
      RECT 17.036 25.78 17.344 25.82 ;
      RECT 17.036 24.62 17.136 25.78 ;
      RECT 17.176 24.62 17.344 25.78 ;
      RECT 17.384 24.62 17.412 25.78 ;
      RECT 17.452 24.62 17.684 25.78 ;
      RECT 17.384 24.58 17.684 24.62 ;
      RECT 17.036 24.58 17.344 24.62 ;
      RECT 17.036 23.42 17.136 24.58 ;
      RECT 17.176 23.42 17.344 24.58 ;
      RECT 17.384 23.42 17.412 24.58 ;
      RECT 17.452 23.42 17.684 24.58 ;
      RECT 17.384 23.38 17.684 23.42 ;
      RECT 17.036 23.38 17.344 23.42 ;
      RECT 17.036 22.22 17.136 23.38 ;
      RECT 17.176 22.22 17.344 23.38 ;
      RECT 17.384 22.22 17.412 23.38 ;
      RECT 17.452 22.22 17.684 23.38 ;
      RECT 17.384 22.18 17.684 22.22 ;
      RECT 17.036 22.18 17.344 22.22 ;
      RECT 17.036 21.02 17.136 22.18 ;
      RECT 17.176 21.02 17.344 22.18 ;
      RECT 17.384 21.02 17.412 22.18 ;
      RECT 17.452 21.02 17.684 22.18 ;
      RECT 17.384 20.98 17.684 21.02 ;
      RECT 17.036 20.98 17.344 21.02 ;
      RECT 17.036 19.82 17.136 20.98 ;
      RECT 17.176 19.82 17.344 20.98 ;
      RECT 17.384 19.82 17.412 20.98 ;
      RECT 17.452 19.82 17.684 20.98 ;
      RECT 17.384 19.78 17.684 19.82 ;
      RECT 17.036 19.78 17.344 19.82 ;
      RECT 17.036 18.62 17.136 19.78 ;
      RECT 17.176 18.62 17.344 19.78 ;
      RECT 17.384 18.62 17.412 19.78 ;
      RECT 17.452 18.62 17.684 19.78 ;
      RECT 17.384 18.58 17.684 18.62 ;
      RECT 17.036 18.58 17.344 18.62 ;
      RECT 17.036 17.42 17.136 18.58 ;
      RECT 17.176 17.42 17.344 18.58 ;
      RECT 17.384 17.42 17.412 18.58 ;
      RECT 17.452 17.42 17.684 18.58 ;
      RECT 17.384 17.38 17.684 17.42 ;
      RECT 17.036 17.38 17.344 17.42 ;
      RECT 17.036 16.22 17.136 17.38 ;
      RECT 17.176 16.22 17.344 17.38 ;
      RECT 17.384 16.22 17.412 17.38 ;
      RECT 17.452 16.22 17.684 17.38 ;
      RECT 17.384 16.18 17.684 16.22 ;
      RECT 17.036 16.18 17.344 16.22 ;
      RECT 17.036 15.02 17.136 16.18 ;
      RECT 17.176 15.02 17.344 16.18 ;
      RECT 17.384 15.02 17.412 16.18 ;
      RECT 17.452 15.02 17.684 16.18 ;
      RECT 17.384 14.98 17.684 15.02 ;
      RECT 17.036 14.98 17.344 15.02 ;
      RECT 17.036 13.82 17.136 14.98 ;
      RECT 17.176 13.82 17.344 14.98 ;
      RECT 17.384 13.82 17.412 14.98 ;
      RECT 17.452 13.82 17.684 14.98 ;
      RECT 17.384 13.78 17.684 13.82 ;
      RECT 17.036 13.78 17.344 13.82 ;
      RECT 17.036 12.62 17.136 13.78 ;
      RECT 17.176 12.62 17.344 13.78 ;
      RECT 17.384 12.62 17.412 13.78 ;
      RECT 17.452 12.62 17.684 13.78 ;
      RECT 17.384 12.58 17.684 12.62 ;
      RECT 17.036 12.58 17.344 12.62 ;
      RECT 17.036 11.42 17.136 12.58 ;
      RECT 17.176 11.42 17.344 12.58 ;
      RECT 17.384 11.42 17.412 12.58 ;
      RECT 17.452 11.42 17.684 12.58 ;
      RECT 17.384 11.38 17.684 11.42 ;
      RECT 17.036 11.38 17.344 11.42 ;
      RECT 17.036 10.22 17.136 11.38 ;
      RECT 17.176 10.22 17.344 11.38 ;
      RECT 17.384 10.22 17.412 11.38 ;
      RECT 17.452 10.22 17.684 11.38 ;
      RECT 17.384 10.18 17.684 10.22 ;
      RECT 17.036 10.18 17.344 10.22 ;
      RECT 17.036 9.02 17.136 10.18 ;
      RECT 17.176 9.02 17.344 10.18 ;
      RECT 17.384 9.02 17.412 10.18 ;
      RECT 17.452 9.02 17.684 10.18 ;
      RECT 17.384 8.98 17.684 9.02 ;
      RECT 17.036 8.98 17.344 9.02 ;
      RECT 17.036 7.82 17.136 8.98 ;
      RECT 17.176 7.82 17.344 8.98 ;
      RECT 17.384 7.82 17.412 8.98 ;
      RECT 17.452 7.82 17.684 8.98 ;
      RECT 17.384 7.78 17.684 7.82 ;
      RECT 17.036 7.78 17.344 7.82 ;
      RECT 17.036 6.62 17.136 7.78 ;
      RECT 17.176 6.62 17.344 7.78 ;
      RECT 17.384 6.62 17.412 7.78 ;
      RECT 17.452 6.62 17.684 7.78 ;
      RECT 17.384 6.58 17.684 6.62 ;
      RECT 17.036 6.58 17.344 6.62 ;
      RECT 17.036 5.42 17.136 6.58 ;
      RECT 17.176 5.42 17.344 6.58 ;
      RECT 17.384 5.42 17.412 6.58 ;
      RECT 17.452 5.42 17.684 6.58 ;
      RECT 17.384 5.38 17.684 5.42 ;
      RECT 17.036 5.38 17.344 5.42 ;
      RECT 17.036 4.22 17.136 5.38 ;
      RECT 17.176 4.22 17.344 5.38 ;
      RECT 17.384 4.22 17.412 5.38 ;
      RECT 17.452 4.22 17.684 5.38 ;
      RECT 17.384 4.18 17.684 4.22 ;
      RECT 17.036 4.18 17.344 4.22 ;
      RECT 17.036 3.02 17.136 4.18 ;
      RECT 17.176 3.02 17.344 4.18 ;
      RECT 17.384 3.02 17.412 4.18 ;
      RECT 17.452 3.02 17.684 4.18 ;
      RECT 17.384 2.98 17.684 3.02 ;
      RECT 17.036 2.98 17.344 3.02 ;
      RECT 17.036 1.82 17.136 2.98 ;
      RECT 17.176 1.82 17.344 2.98 ;
      RECT 17.384 1.82 17.412 2.98 ;
      RECT 17.452 1.82 17.684 2.98 ;
      RECT 17.384 1.78 17.684 1.82 ;
      RECT 17.036 1.78 17.344 1.82 ;
      RECT 19.35 31.8 19.45 39.72 ;
      RECT 19.036 31.8 19.31 31.84 ;
      RECT 17.452 0.62 17.684 1.78 ;
      RECT 17.036 0.62 17.136 1.78 ;
      RECT 17.176 0.62 17.344 1.78 ;
      RECT 17.384 0.62 17.412 1.78 ;
      RECT 27.226 0.6 27.574 72.12 ;
      RECT 31.626 0.6 31.974 32.9505 ;
      RECT 34.026 0.6 34.374 32.9505 ;
      RECT 34.426 0.6 34.774 72.12 ;
      RECT 35.226 0.6 35.574 72.12 ;
      RECT 34.826 0.6 35.174 32.9505 ;
      RECT 32.026 0.6 32.374 72.12 ;
      RECT 32.826 0.6 33.174 72.12 ;
      RECT 33.626 0.6 33.974 72.12 ;
      RECT 32.426 0.6 32.774 32.9505 ;
      RECT 33.226 0.6 33.574 32.9505 ;
      RECT 29.226 0.6 29.574 32.9505 ;
      RECT 29.626 0.6 29.974 72.12 ;
      RECT 30.426 0.6 30.774 72.12 ;
      RECT 31.226 0.6 31.574 72.12 ;
      RECT 30.026 0.6 30.374 32.9505 ;
      RECT 30.826 0.6 31.174 32.9505 ;
      RECT 28.026 0.6 28.374 72.12 ;
      RECT 28.826 0.6 29.174 72.12 ;
      RECT 27.626 0.6 27.974 32.9505 ;
      RECT 28.426 0.6 28.774 32.9505 ;
      RECT 24.826 0.6 25.174 72.12 ;
      RECT 25.626 0.6 25.974 72.12 ;
      RECT 26.426 0.6 26.774 72.12 ;
      RECT 25.226 0.6 25.574 32.9505 ;
      RECT 26.026 0.6 26.374 32.9505 ;
      RECT 26.826 0.6 27.174 32.9505 ;
      RECT 23.226 0.6 23.574 72.12 ;
      RECT 24.026 0.6 24.374 72.12 ;
      RECT 22.826 0.6 23.174 32.9505 ;
      RECT 23.626 0.6 23.974 32.9505 ;
      RECT 24.426 0.6 24.774 32.9505 ;
      RECT 20.046 0.6 20.074 72.12 ;
      RECT 20.126 0.6 20.29 72.12 ;
      RECT 9.026 0.6 9.374 72.12 ;
      RECT 15.71 0.6 15.874 72.12 ;
      RECT 15.926 0.6 15.954 72.12 ;
      RECT 11.026 0.6 11.374 32.9505 ;
      RECT 11.426 0.6 11.774 72.12 ;
      RECT 12.226 0.6 12.574 72.12 ;
      RECT 13.026 0.6 13.374 72.12 ;
      RECT 11.826 0.6 12.174 32.9505 ;
      RECT 12.626 0.6 12.974 32.9505 ;
      RECT 9.826 0.6 10.174 72.12 ;
      RECT 10.626 0.6 10.974 72.12 ;
      RECT 9.426 0.6 9.774 32.9505 ;
      RECT 10.226 0.6 10.574 32.9505 ;
      RECT 4.226 0.6 4.574 72.12 ;
      RECT 6.626 0.6 6.974 72.12 ;
      RECT 7.426 0.6 7.774 72.12 ;
      RECT 8.226 0.6 8.574 72.12 ;
      RECT 7.026 0.6 7.374 32.9505 ;
      RECT 7.826 0.6 8.174 32.9505 ;
      RECT 8.626 0.6 8.974 32.9505 ;
      RECT 5.026 0.6 5.374 72.12 ;
      RECT 5.826 0.6 6.174 72.12 ;
      RECT 4.626 0.6 4.974 32.9505 ;
      RECT 5.426 0.6 5.774 32.9505 ;
      RECT 6.226 0.6 6.574 32.9505 ;
      RECT 2.626 0.6 2.974 72.12 ;
      RECT 3.426 0.6 3.774 72.12 ;
      RECT 2.226 0.6 2.574 32.9505 ;
      RECT 3.026 0.6 3.374 32.9505 ;
      RECT 3.826 0.6 4.174 32.9505 ;
      RECT 1.026 0.6 1.374 72.12 ;
      RECT 1.826 0.6 2.174 72.12 ;
      RECT 0.626 0.6 0.974 32.9505 ;
      RECT 1.426 0.6 1.774 32.9505 ;
      RECT -0.059 -0.09 36.359 0.5695 ;
      RECT 26.826 0.5695 27.574 0.6 ;
      RECT 31.626 0.5695 32.374 0.6 ;
      RECT 34.026 0.5695 34.774 0.6 ;
      RECT 35.626 0.5695 36.359 72.1505 ;
      RECT 34.826 0.5695 35.574 0.6 ;
      RECT 32.426 0.5695 33.174 0.6 ;
      RECT 33.226 0.5695 33.974 0.6 ;
      RECT 29.226 0.5695 29.974 0.6 ;
      RECT 30.026 0.5695 30.774 0.6 ;
      RECT 30.826 0.5695 31.574 0.6 ;
      RECT 27.626 0.5695 28.374 0.6 ;
      RECT 28.426 0.5695 29.174 0.6 ;
      RECT 21.95 0.5695 22.774 72.1505 ;
      RECT 24.426 0.5695 25.174 0.6 ;
      RECT 25.226 0.5695 25.974 0.6 ;
      RECT 26.026 0.5695 26.774 0.6 ;
      RECT 22.826 0.5695 23.574 0.6 ;
      RECT 23.626 0.5695 24.374 0.6 ;
      RECT 20.342 0.5695 20.47 32.8595 ;
      RECT 20.682 0.5695 21.014 72.1505 ;
      RECT 21.068 0.5695 21.496 72.1505 ;
      RECT 21.55 0.5695 21.65 72.1505 ;
      RECT 21.704 0.5695 21.896 72.1505 ;
      RECT 20.522 0.5695 20.63 32.8595 ;
      RECT 18.636 0.5695 18.664 72.1505 ;
      RECT 18.736 0.5695 18.864 72.1505 ;
      RECT 18.936 0.5695 18.964 72.1505 ;
      RECT 19.502 0.5695 19.682 72.1505 ;
      RECT 19.734 0.5695 19.914 72.1505 ;
      RECT 19.966 0.5695 19.994 72.1505 ;
      RECT 18.396 0.5695 18.564 36.85 ;
      RECT 18.188 0.5695 18.356 31.82 ;
      RECT 19.036 0.5695 19.45 31.8 ;
      RECT 20.046 0.5695 20.29 0.6 ;
      RECT 8.626 0.5695 9.374 0.6 ;
      RECT 13.426 0.5695 14.05 72.1505 ;
      RECT 15.71 0.5695 15.954 0.6 ;
      RECT 17.384 0.5695 17.684 0.62 ;
      RECT 17.736 0.5695 17.844 72.1505 ;
      RECT 17.916 0.5695 18.148 33.18 ;
      RECT 17.036 0.5695 17.344 0.62 ;
      RECT 16.006 0.5695 16.034 72.1505 ;
      RECT 16.086 0.5695 16.266 72.1505 ;
      RECT 16.318 0.5695 16.498 72.1505 ;
      RECT 16.55 0.5695 16.8 72.1505 ;
      RECT 16.854 0.5695 16.964 32.353 ;
      RECT 14.104 0.5695 14.296 72.1505 ;
      RECT 14.35 0.5695 14.45 72.1505 ;
      RECT 14.504 0.5695 14.932 72.1505 ;
      RECT 14.986 0.5695 15.318 72.1505 ;
      RECT 15.37 0.5695 15.478 32.8595 ;
      RECT 15.53 0.5695 15.658 32.8595 ;
      RECT 11.026 0.5695 11.774 0.6 ;
      RECT 11.826 0.5695 12.574 0.6 ;
      RECT 12.626 0.5695 13.374 0.6 ;
      RECT 9.426 0.5695 10.174 0.6 ;
      RECT 10.226 0.5695 10.974 0.6 ;
      RECT 3.826 0.5695 4.574 0.6 ;
      RECT 6.226 0.5695 6.974 0.6 ;
      RECT 7.026 0.5695 7.774 0.6 ;
      RECT 7.826 0.5695 8.574 0.6 ;
      RECT 4.626 0.5695 5.374 0.6 ;
      RECT 5.426 0.5695 6.174 0.6 ;
      RECT 2.226 0.5695 2.974 0.6 ;
      RECT 3.026 0.5695 3.774 0.6 ;
      RECT -0.059 0.5695 0.574 72.1505 ;
      RECT 0.626 0.5695 1.374 0.6 ;
      RECT 1.426 0.5695 2.174 0.6 ;
    LAYER v4 ;
      RECT 21.978 72.102 22.022 72.138 ;
      RECT 21.096 72.102 21.14 72.138 ;
      RECT 14.86 72.102 14.904 72.138 ;
      RECT 13.978 72.102 14.022 72.138 ;
      RECT 35.494 71.878 35.546 71.914 ;
      RECT 35.094 71.878 35.146 71.914 ;
      RECT 34.694 71.878 34.746 71.914 ;
      RECT 34.294 71.878 34.346 71.914 ;
      RECT 33.894 71.878 33.946 71.914 ;
      RECT 33.494 71.878 33.546 71.914 ;
      RECT 33.094 71.878 33.146 71.914 ;
      RECT 32.694 71.878 32.746 71.914 ;
      RECT 32.294 71.878 32.346 71.914 ;
      RECT 31.894 71.878 31.946 71.914 ;
      RECT 31.494 71.878 31.546 71.914 ;
      RECT 31.094 71.878 31.146 71.914 ;
      RECT 30.694 71.878 30.746 71.914 ;
      RECT 30.294 71.878 30.346 71.914 ;
      RECT 29.894 71.878 29.946 71.914 ;
      RECT 29.494 71.878 29.546 71.914 ;
      RECT 29.094 71.878 29.146 71.914 ;
      RECT 28.694 71.878 28.746 71.914 ;
      RECT 28.294 71.878 28.346 71.914 ;
      RECT 27.894 71.878 27.946 71.914 ;
      RECT 27.494 71.878 27.546 71.914 ;
      RECT 27.094 71.878 27.146 71.914 ;
      RECT 26.694 71.878 26.746 71.914 ;
      RECT 26.294 71.878 26.346 71.914 ;
      RECT 25.894 71.878 25.946 71.914 ;
      RECT 25.494 71.878 25.546 71.914 ;
      RECT 25.094 71.878 25.146 71.914 ;
      RECT 24.694 71.878 24.746 71.914 ;
      RECT 24.294 71.878 24.346 71.914 ;
      RECT 23.894 71.878 23.946 71.914 ;
      RECT 23.494 71.878 23.546 71.914 ;
      RECT 23.094 71.878 23.146 71.914 ;
      RECT 21.814 71.878 21.868 71.914 ;
      RECT 19.838 71.878 19.886 71.914 ;
      RECT 19.53 71.878 19.578 71.914 ;
      RECT 16.882 71.878 16.936 71.914 ;
      RECT 16.422 71.878 16.47 71.914 ;
      RECT 16.114 71.878 16.162 71.914 ;
      RECT 14.132 71.878 14.186 71.914 ;
      RECT 13.294 71.878 13.346 71.914 ;
      RECT 12.894 71.878 12.946 71.914 ;
      RECT 12.494 71.878 12.546 71.914 ;
      RECT 12.094 71.878 12.146 71.914 ;
      RECT 11.694 71.878 11.746 71.914 ;
      RECT 11.294 71.878 11.346 71.914 ;
      RECT 10.894 71.878 10.946 71.914 ;
      RECT 10.494 71.878 10.546 71.914 ;
      RECT 10.094 71.878 10.146 71.914 ;
      RECT 9.694 71.878 9.746 71.914 ;
      RECT 9.294 71.878 9.346 71.914 ;
      RECT 8.894 71.878 8.946 71.914 ;
      RECT 8.494 71.878 8.546 71.914 ;
      RECT 8.094 71.878 8.146 71.914 ;
      RECT 7.694 71.878 7.746 71.914 ;
      RECT 7.294 71.878 7.346 71.914 ;
      RECT 6.894 71.878 6.946 71.914 ;
      RECT 6.494 71.878 6.546 71.914 ;
      RECT 6.094 71.878 6.146 71.914 ;
      RECT 5.694 71.878 5.746 71.914 ;
      RECT 5.294 71.878 5.346 71.914 ;
      RECT 4.894 71.878 4.946 71.914 ;
      RECT 4.494 71.878 4.546 71.914 ;
      RECT 4.094 71.878 4.146 71.914 ;
      RECT 3.694 71.878 3.746 71.914 ;
      RECT 3.294 71.878 3.346 71.914 ;
      RECT 2.894 71.878 2.946 71.914 ;
      RECT 2.494 71.878 2.546 71.914 ;
      RECT 2.094 71.878 2.146 71.914 ;
      RECT 1.694 71.878 1.746 71.914 ;
      RECT 1.294 71.878 1.346 71.914 ;
      RECT 0.894 71.878 0.946 71.914 ;
      RECT 21.414 71.802 21.468 71.838 ;
      RECT 14.532 71.802 14.586 71.838 ;
      RECT 19.606 71.649 19.654 71.685 ;
      RECT 18.08 71.649 18.12 71.685 ;
      RECT 16.718 71.649 16.772 71.685 ;
      RECT 16.346 71.649 16.394 71.685 ;
      RECT 20.37 71.6545 20.442 71.6795 ;
      RECT 18.764 71.6545 18.836 71.6795 ;
      RECT 15.558 71.6545 15.63 71.6795 ;
      RECT 21.978 71.502 22.022 71.538 ;
      RECT 13.978 71.502 14.022 71.538 ;
      RECT 18.764 71.5075 18.836 71.5325 ;
      RECT 19.762 71.355 19.81 71.391 ;
      RECT 17.616 71.355 17.656 71.391 ;
      RECT 16.19 71.355 16.238 71.391 ;
      RECT 35.254 71.126 35.306 71.162 ;
      RECT 34.854 71.126 34.906 71.162 ;
      RECT 34.454 71.126 34.506 71.162 ;
      RECT 34.054 71.126 34.106 71.162 ;
      RECT 33.654 71.126 33.706 71.162 ;
      RECT 33.254 71.126 33.306 71.162 ;
      RECT 32.854 71.126 32.906 71.162 ;
      RECT 32.454 71.126 32.506 71.162 ;
      RECT 32.054 71.126 32.106 71.162 ;
      RECT 31.654 71.126 31.706 71.162 ;
      RECT 31.254 71.126 31.306 71.162 ;
      RECT 30.854 71.126 30.906 71.162 ;
      RECT 30.454 71.126 30.506 71.162 ;
      RECT 30.054 71.126 30.106 71.162 ;
      RECT 29.654 71.126 29.706 71.162 ;
      RECT 29.254 71.126 29.306 71.162 ;
      RECT 28.854 71.126 28.906 71.162 ;
      RECT 28.454 71.126 28.506 71.162 ;
      RECT 28.054 71.126 28.106 71.162 ;
      RECT 27.654 71.126 27.706 71.162 ;
      RECT 27.254 71.126 27.306 71.162 ;
      RECT 26.854 71.126 26.906 71.162 ;
      RECT 26.454 71.126 26.506 71.162 ;
      RECT 26.054 71.126 26.106 71.162 ;
      RECT 25.654 71.126 25.706 71.162 ;
      RECT 25.254 71.126 25.306 71.162 ;
      RECT 24.854 71.126 24.906 71.162 ;
      RECT 24.454 71.126 24.506 71.162 ;
      RECT 24.054 71.126 24.106 71.162 ;
      RECT 23.654 71.126 23.706 71.162 ;
      RECT 23.254 71.126 23.306 71.162 ;
      RECT 22.854 71.126 22.906 71.162 ;
      RECT 22.694 71.126 22.746 71.162 ;
      RECT 21.732 71.126 21.786 71.162 ;
      RECT 14.214 71.126 14.268 71.162 ;
      RECT 13.054 71.126 13.106 71.162 ;
      RECT 12.654 71.126 12.706 71.162 ;
      RECT 12.254 71.126 12.306 71.162 ;
      RECT 11.854 71.126 11.906 71.162 ;
      RECT 11.454 71.126 11.506 71.162 ;
      RECT 11.054 71.126 11.106 71.162 ;
      RECT 10.654 71.126 10.706 71.162 ;
      RECT 10.254 71.126 10.306 71.162 ;
      RECT 9.854 71.126 9.906 71.162 ;
      RECT 9.454 71.126 9.506 71.162 ;
      RECT 9.054 71.126 9.106 71.162 ;
      RECT 8.654 71.126 8.706 71.162 ;
      RECT 8.254 71.126 8.306 71.162 ;
      RECT 7.854 71.126 7.906 71.162 ;
      RECT 7.454 71.126 7.506 71.162 ;
      RECT 7.054 71.126 7.106 71.162 ;
      RECT 6.654 71.126 6.706 71.162 ;
      RECT 6.254 71.126 6.306 71.162 ;
      RECT 5.854 71.126 5.906 71.162 ;
      RECT 5.454 71.126 5.506 71.162 ;
      RECT 5.054 71.126 5.106 71.162 ;
      RECT 4.654 71.126 4.706 71.162 ;
      RECT 4.254 71.126 4.306 71.162 ;
      RECT 3.854 71.126 3.906 71.162 ;
      RECT 3.454 71.126 3.506 71.162 ;
      RECT 3.054 71.126 3.106 71.162 ;
      RECT 2.654 71.126 2.706 71.162 ;
      RECT 2.254 71.126 2.306 71.162 ;
      RECT 1.854 71.126 1.906 71.162 ;
      RECT 1.454 71.126 1.506 71.162 ;
      RECT 1.054 71.126 1.106 71.162 ;
      RECT 0.654 71.126 0.706 71.162 ;
      RECT 21.978 70.902 22.022 70.938 ;
      RECT 21.096 70.902 21.14 70.938 ;
      RECT 14.86 70.902 14.904 70.938 ;
      RECT 13.978 70.902 14.022 70.938 ;
      RECT 35.494 70.678 35.546 70.714 ;
      RECT 35.094 70.678 35.146 70.714 ;
      RECT 34.694 70.678 34.746 70.714 ;
      RECT 34.294 70.678 34.346 70.714 ;
      RECT 33.894 70.678 33.946 70.714 ;
      RECT 33.494 70.678 33.546 70.714 ;
      RECT 33.094 70.678 33.146 70.714 ;
      RECT 32.694 70.678 32.746 70.714 ;
      RECT 32.294 70.678 32.346 70.714 ;
      RECT 31.894 70.678 31.946 70.714 ;
      RECT 31.494 70.678 31.546 70.714 ;
      RECT 31.094 70.678 31.146 70.714 ;
      RECT 30.694 70.678 30.746 70.714 ;
      RECT 30.294 70.678 30.346 70.714 ;
      RECT 29.894 70.678 29.946 70.714 ;
      RECT 29.494 70.678 29.546 70.714 ;
      RECT 29.094 70.678 29.146 70.714 ;
      RECT 28.694 70.678 28.746 70.714 ;
      RECT 28.294 70.678 28.346 70.714 ;
      RECT 27.894 70.678 27.946 70.714 ;
      RECT 27.494 70.678 27.546 70.714 ;
      RECT 27.094 70.678 27.146 70.714 ;
      RECT 26.694 70.678 26.746 70.714 ;
      RECT 26.294 70.678 26.346 70.714 ;
      RECT 25.894 70.678 25.946 70.714 ;
      RECT 25.494 70.678 25.546 70.714 ;
      RECT 25.094 70.678 25.146 70.714 ;
      RECT 24.694 70.678 24.746 70.714 ;
      RECT 24.294 70.678 24.346 70.714 ;
      RECT 23.894 70.678 23.946 70.714 ;
      RECT 23.494 70.678 23.546 70.714 ;
      RECT 23.094 70.678 23.146 70.714 ;
      RECT 21.814 70.678 21.868 70.714 ;
      RECT 19.838 70.678 19.886 70.714 ;
      RECT 19.53 70.678 19.578 70.714 ;
      RECT 16.882 70.678 16.936 70.714 ;
      RECT 16.422 70.678 16.47 70.714 ;
      RECT 16.114 70.678 16.162 70.714 ;
      RECT 14.132 70.678 14.186 70.714 ;
      RECT 13.294 70.678 13.346 70.714 ;
      RECT 12.894 70.678 12.946 70.714 ;
      RECT 12.494 70.678 12.546 70.714 ;
      RECT 12.094 70.678 12.146 70.714 ;
      RECT 11.694 70.678 11.746 70.714 ;
      RECT 11.294 70.678 11.346 70.714 ;
      RECT 10.894 70.678 10.946 70.714 ;
      RECT 10.494 70.678 10.546 70.714 ;
      RECT 10.094 70.678 10.146 70.714 ;
      RECT 9.694 70.678 9.746 70.714 ;
      RECT 9.294 70.678 9.346 70.714 ;
      RECT 8.894 70.678 8.946 70.714 ;
      RECT 8.494 70.678 8.546 70.714 ;
      RECT 8.094 70.678 8.146 70.714 ;
      RECT 7.694 70.678 7.746 70.714 ;
      RECT 7.294 70.678 7.346 70.714 ;
      RECT 6.894 70.678 6.946 70.714 ;
      RECT 6.494 70.678 6.546 70.714 ;
      RECT 6.094 70.678 6.146 70.714 ;
      RECT 5.694 70.678 5.746 70.714 ;
      RECT 5.294 70.678 5.346 70.714 ;
      RECT 4.894 70.678 4.946 70.714 ;
      RECT 4.494 70.678 4.546 70.714 ;
      RECT 4.094 70.678 4.146 70.714 ;
      RECT 3.694 70.678 3.746 70.714 ;
      RECT 3.294 70.678 3.346 70.714 ;
      RECT 2.894 70.678 2.946 70.714 ;
      RECT 2.494 70.678 2.546 70.714 ;
      RECT 2.094 70.678 2.146 70.714 ;
      RECT 1.694 70.678 1.746 70.714 ;
      RECT 1.294 70.678 1.346 70.714 ;
      RECT 0.894 70.678 0.946 70.714 ;
      RECT 21.414 70.602 21.468 70.638 ;
      RECT 14.532 70.602 14.586 70.638 ;
      RECT 19.606 70.449 19.654 70.485 ;
      RECT 18.08 70.449 18.12 70.485 ;
      RECT 16.718 70.449 16.772 70.485 ;
      RECT 16.346 70.449 16.394 70.485 ;
      RECT 20.37 70.4545 20.442 70.4795 ;
      RECT 18.764 70.4545 18.836 70.4795 ;
      RECT 15.558 70.4545 15.63 70.4795 ;
      RECT 21.978 70.302 22.022 70.338 ;
      RECT 13.978 70.302 14.022 70.338 ;
      RECT 18.764 70.3075 18.836 70.3325 ;
      RECT 19.762 70.155 19.81 70.191 ;
      RECT 17.616 70.155 17.656 70.191 ;
      RECT 16.19 70.155 16.238 70.191 ;
      RECT 35.254 69.926 35.306 69.962 ;
      RECT 34.854 69.926 34.906 69.962 ;
      RECT 34.454 69.926 34.506 69.962 ;
      RECT 34.054 69.926 34.106 69.962 ;
      RECT 33.654 69.926 33.706 69.962 ;
      RECT 33.254 69.926 33.306 69.962 ;
      RECT 32.854 69.926 32.906 69.962 ;
      RECT 32.454 69.926 32.506 69.962 ;
      RECT 32.054 69.926 32.106 69.962 ;
      RECT 31.654 69.926 31.706 69.962 ;
      RECT 31.254 69.926 31.306 69.962 ;
      RECT 30.854 69.926 30.906 69.962 ;
      RECT 30.454 69.926 30.506 69.962 ;
      RECT 30.054 69.926 30.106 69.962 ;
      RECT 29.654 69.926 29.706 69.962 ;
      RECT 29.254 69.926 29.306 69.962 ;
      RECT 28.854 69.926 28.906 69.962 ;
      RECT 28.454 69.926 28.506 69.962 ;
      RECT 28.054 69.926 28.106 69.962 ;
      RECT 27.654 69.926 27.706 69.962 ;
      RECT 27.254 69.926 27.306 69.962 ;
      RECT 26.854 69.926 26.906 69.962 ;
      RECT 26.454 69.926 26.506 69.962 ;
      RECT 26.054 69.926 26.106 69.962 ;
      RECT 25.654 69.926 25.706 69.962 ;
      RECT 25.254 69.926 25.306 69.962 ;
      RECT 24.854 69.926 24.906 69.962 ;
      RECT 24.454 69.926 24.506 69.962 ;
      RECT 24.054 69.926 24.106 69.962 ;
      RECT 23.654 69.926 23.706 69.962 ;
      RECT 23.254 69.926 23.306 69.962 ;
      RECT 22.854 69.926 22.906 69.962 ;
      RECT 22.694 69.926 22.746 69.962 ;
      RECT 21.732 69.926 21.786 69.962 ;
      RECT 14.214 69.926 14.268 69.962 ;
      RECT 13.054 69.926 13.106 69.962 ;
      RECT 12.654 69.926 12.706 69.962 ;
      RECT 12.254 69.926 12.306 69.962 ;
      RECT 11.854 69.926 11.906 69.962 ;
      RECT 11.454 69.926 11.506 69.962 ;
      RECT 11.054 69.926 11.106 69.962 ;
      RECT 10.654 69.926 10.706 69.962 ;
      RECT 10.254 69.926 10.306 69.962 ;
      RECT 9.854 69.926 9.906 69.962 ;
      RECT 9.454 69.926 9.506 69.962 ;
      RECT 9.054 69.926 9.106 69.962 ;
      RECT 8.654 69.926 8.706 69.962 ;
      RECT 8.254 69.926 8.306 69.962 ;
      RECT 7.854 69.926 7.906 69.962 ;
      RECT 7.454 69.926 7.506 69.962 ;
      RECT 7.054 69.926 7.106 69.962 ;
      RECT 6.654 69.926 6.706 69.962 ;
      RECT 6.254 69.926 6.306 69.962 ;
      RECT 5.854 69.926 5.906 69.962 ;
      RECT 5.454 69.926 5.506 69.962 ;
      RECT 5.054 69.926 5.106 69.962 ;
      RECT 4.654 69.926 4.706 69.962 ;
      RECT 4.254 69.926 4.306 69.962 ;
      RECT 3.854 69.926 3.906 69.962 ;
      RECT 3.454 69.926 3.506 69.962 ;
      RECT 3.054 69.926 3.106 69.962 ;
      RECT 2.654 69.926 2.706 69.962 ;
      RECT 2.254 69.926 2.306 69.962 ;
      RECT 1.854 69.926 1.906 69.962 ;
      RECT 1.454 69.926 1.506 69.962 ;
      RECT 1.054 69.926 1.106 69.962 ;
      RECT 0.654 69.926 0.706 69.962 ;
      RECT 21.978 69.702 22.022 69.738 ;
      RECT 21.096 69.702 21.14 69.738 ;
      RECT 14.86 69.702 14.904 69.738 ;
      RECT 13.978 69.702 14.022 69.738 ;
      RECT 35.494 69.478 35.546 69.514 ;
      RECT 35.094 69.478 35.146 69.514 ;
      RECT 34.694 69.478 34.746 69.514 ;
      RECT 34.294 69.478 34.346 69.514 ;
      RECT 33.894 69.478 33.946 69.514 ;
      RECT 33.494 69.478 33.546 69.514 ;
      RECT 33.094 69.478 33.146 69.514 ;
      RECT 32.694 69.478 32.746 69.514 ;
      RECT 32.294 69.478 32.346 69.514 ;
      RECT 31.894 69.478 31.946 69.514 ;
      RECT 31.494 69.478 31.546 69.514 ;
      RECT 31.094 69.478 31.146 69.514 ;
      RECT 30.694 69.478 30.746 69.514 ;
      RECT 30.294 69.478 30.346 69.514 ;
      RECT 29.894 69.478 29.946 69.514 ;
      RECT 29.494 69.478 29.546 69.514 ;
      RECT 29.094 69.478 29.146 69.514 ;
      RECT 28.694 69.478 28.746 69.514 ;
      RECT 28.294 69.478 28.346 69.514 ;
      RECT 27.894 69.478 27.946 69.514 ;
      RECT 27.494 69.478 27.546 69.514 ;
      RECT 27.094 69.478 27.146 69.514 ;
      RECT 26.694 69.478 26.746 69.514 ;
      RECT 26.294 69.478 26.346 69.514 ;
      RECT 25.894 69.478 25.946 69.514 ;
      RECT 25.494 69.478 25.546 69.514 ;
      RECT 25.094 69.478 25.146 69.514 ;
      RECT 24.694 69.478 24.746 69.514 ;
      RECT 24.294 69.478 24.346 69.514 ;
      RECT 23.894 69.478 23.946 69.514 ;
      RECT 23.494 69.478 23.546 69.514 ;
      RECT 23.094 69.478 23.146 69.514 ;
      RECT 21.814 69.478 21.868 69.514 ;
      RECT 19.838 69.478 19.886 69.514 ;
      RECT 19.53 69.478 19.578 69.514 ;
      RECT 16.882 69.478 16.936 69.514 ;
      RECT 16.422 69.478 16.47 69.514 ;
      RECT 16.114 69.478 16.162 69.514 ;
      RECT 14.132 69.478 14.186 69.514 ;
      RECT 13.294 69.478 13.346 69.514 ;
      RECT 12.894 69.478 12.946 69.514 ;
      RECT 12.494 69.478 12.546 69.514 ;
      RECT 12.094 69.478 12.146 69.514 ;
      RECT 11.694 69.478 11.746 69.514 ;
      RECT 11.294 69.478 11.346 69.514 ;
      RECT 10.894 69.478 10.946 69.514 ;
      RECT 10.494 69.478 10.546 69.514 ;
      RECT 10.094 69.478 10.146 69.514 ;
      RECT 9.694 69.478 9.746 69.514 ;
      RECT 9.294 69.478 9.346 69.514 ;
      RECT 8.894 69.478 8.946 69.514 ;
      RECT 8.494 69.478 8.546 69.514 ;
      RECT 8.094 69.478 8.146 69.514 ;
      RECT 7.694 69.478 7.746 69.514 ;
      RECT 7.294 69.478 7.346 69.514 ;
      RECT 6.894 69.478 6.946 69.514 ;
      RECT 6.494 69.478 6.546 69.514 ;
      RECT 6.094 69.478 6.146 69.514 ;
      RECT 5.694 69.478 5.746 69.514 ;
      RECT 5.294 69.478 5.346 69.514 ;
      RECT 4.894 69.478 4.946 69.514 ;
      RECT 4.494 69.478 4.546 69.514 ;
      RECT 4.094 69.478 4.146 69.514 ;
      RECT 3.694 69.478 3.746 69.514 ;
      RECT 3.294 69.478 3.346 69.514 ;
      RECT 2.894 69.478 2.946 69.514 ;
      RECT 2.494 69.478 2.546 69.514 ;
      RECT 2.094 69.478 2.146 69.514 ;
      RECT 1.694 69.478 1.746 69.514 ;
      RECT 1.294 69.478 1.346 69.514 ;
      RECT 0.894 69.478 0.946 69.514 ;
      RECT 21.414 69.402 21.468 69.438 ;
      RECT 14.532 69.402 14.586 69.438 ;
      RECT 19.606 69.249 19.654 69.285 ;
      RECT 18.08 69.249 18.12 69.285 ;
      RECT 16.718 69.249 16.772 69.285 ;
      RECT 16.346 69.249 16.394 69.285 ;
      RECT 20.37 69.2545 20.442 69.2795 ;
      RECT 18.764 69.2545 18.836 69.2795 ;
      RECT 15.558 69.2545 15.63 69.2795 ;
      RECT 21.978 69.102 22.022 69.138 ;
      RECT 13.978 69.102 14.022 69.138 ;
      RECT 18.764 69.1075 18.836 69.1325 ;
      RECT 19.762 68.955 19.81 68.991 ;
      RECT 17.616 68.955 17.656 68.991 ;
      RECT 16.19 68.955 16.238 68.991 ;
      RECT 35.254 68.726 35.306 68.762 ;
      RECT 34.854 68.726 34.906 68.762 ;
      RECT 34.454 68.726 34.506 68.762 ;
      RECT 34.054 68.726 34.106 68.762 ;
      RECT 33.654 68.726 33.706 68.762 ;
      RECT 33.254 68.726 33.306 68.762 ;
      RECT 32.854 68.726 32.906 68.762 ;
      RECT 32.454 68.726 32.506 68.762 ;
      RECT 32.054 68.726 32.106 68.762 ;
      RECT 31.654 68.726 31.706 68.762 ;
      RECT 31.254 68.726 31.306 68.762 ;
      RECT 30.854 68.726 30.906 68.762 ;
      RECT 30.454 68.726 30.506 68.762 ;
      RECT 30.054 68.726 30.106 68.762 ;
      RECT 29.654 68.726 29.706 68.762 ;
      RECT 29.254 68.726 29.306 68.762 ;
      RECT 28.854 68.726 28.906 68.762 ;
      RECT 28.454 68.726 28.506 68.762 ;
      RECT 28.054 68.726 28.106 68.762 ;
      RECT 27.654 68.726 27.706 68.762 ;
      RECT 27.254 68.726 27.306 68.762 ;
      RECT 26.854 68.726 26.906 68.762 ;
      RECT 26.454 68.726 26.506 68.762 ;
      RECT 26.054 68.726 26.106 68.762 ;
      RECT 25.654 68.726 25.706 68.762 ;
      RECT 25.254 68.726 25.306 68.762 ;
      RECT 24.854 68.726 24.906 68.762 ;
      RECT 24.454 68.726 24.506 68.762 ;
      RECT 24.054 68.726 24.106 68.762 ;
      RECT 23.654 68.726 23.706 68.762 ;
      RECT 23.254 68.726 23.306 68.762 ;
      RECT 22.854 68.726 22.906 68.762 ;
      RECT 22.694 68.726 22.746 68.762 ;
      RECT 21.732 68.726 21.786 68.762 ;
      RECT 14.214 68.726 14.268 68.762 ;
      RECT 13.054 68.726 13.106 68.762 ;
      RECT 12.654 68.726 12.706 68.762 ;
      RECT 12.254 68.726 12.306 68.762 ;
      RECT 11.854 68.726 11.906 68.762 ;
      RECT 11.454 68.726 11.506 68.762 ;
      RECT 11.054 68.726 11.106 68.762 ;
      RECT 10.654 68.726 10.706 68.762 ;
      RECT 10.254 68.726 10.306 68.762 ;
      RECT 9.854 68.726 9.906 68.762 ;
      RECT 9.454 68.726 9.506 68.762 ;
      RECT 9.054 68.726 9.106 68.762 ;
      RECT 8.654 68.726 8.706 68.762 ;
      RECT 8.254 68.726 8.306 68.762 ;
      RECT 7.854 68.726 7.906 68.762 ;
      RECT 7.454 68.726 7.506 68.762 ;
      RECT 7.054 68.726 7.106 68.762 ;
      RECT 6.654 68.726 6.706 68.762 ;
      RECT 6.254 68.726 6.306 68.762 ;
      RECT 5.854 68.726 5.906 68.762 ;
      RECT 5.454 68.726 5.506 68.762 ;
      RECT 5.054 68.726 5.106 68.762 ;
      RECT 4.654 68.726 4.706 68.762 ;
      RECT 4.254 68.726 4.306 68.762 ;
      RECT 3.854 68.726 3.906 68.762 ;
      RECT 3.454 68.726 3.506 68.762 ;
      RECT 3.054 68.726 3.106 68.762 ;
      RECT 2.654 68.726 2.706 68.762 ;
      RECT 2.254 68.726 2.306 68.762 ;
      RECT 1.854 68.726 1.906 68.762 ;
      RECT 1.454 68.726 1.506 68.762 ;
      RECT 1.054 68.726 1.106 68.762 ;
      RECT 0.654 68.726 0.706 68.762 ;
      RECT 21.978 68.502 22.022 68.538 ;
      RECT 21.096 68.502 21.14 68.538 ;
      RECT 14.86 68.502 14.904 68.538 ;
      RECT 13.978 68.502 14.022 68.538 ;
      RECT 35.494 68.278 35.546 68.314 ;
      RECT 35.094 68.278 35.146 68.314 ;
      RECT 34.694 68.278 34.746 68.314 ;
      RECT 34.294 68.278 34.346 68.314 ;
      RECT 33.894 68.278 33.946 68.314 ;
      RECT 33.494 68.278 33.546 68.314 ;
      RECT 33.094 68.278 33.146 68.314 ;
      RECT 32.694 68.278 32.746 68.314 ;
      RECT 32.294 68.278 32.346 68.314 ;
      RECT 31.894 68.278 31.946 68.314 ;
      RECT 31.494 68.278 31.546 68.314 ;
      RECT 31.094 68.278 31.146 68.314 ;
      RECT 30.694 68.278 30.746 68.314 ;
      RECT 30.294 68.278 30.346 68.314 ;
      RECT 29.894 68.278 29.946 68.314 ;
      RECT 29.494 68.278 29.546 68.314 ;
      RECT 29.094 68.278 29.146 68.314 ;
      RECT 28.694 68.278 28.746 68.314 ;
      RECT 28.294 68.278 28.346 68.314 ;
      RECT 27.894 68.278 27.946 68.314 ;
      RECT 27.494 68.278 27.546 68.314 ;
      RECT 27.094 68.278 27.146 68.314 ;
      RECT 26.694 68.278 26.746 68.314 ;
      RECT 26.294 68.278 26.346 68.314 ;
      RECT 25.894 68.278 25.946 68.314 ;
      RECT 25.494 68.278 25.546 68.314 ;
      RECT 25.094 68.278 25.146 68.314 ;
      RECT 24.694 68.278 24.746 68.314 ;
      RECT 24.294 68.278 24.346 68.314 ;
      RECT 23.894 68.278 23.946 68.314 ;
      RECT 23.494 68.278 23.546 68.314 ;
      RECT 23.094 68.278 23.146 68.314 ;
      RECT 21.814 68.278 21.868 68.314 ;
      RECT 19.838 68.278 19.886 68.314 ;
      RECT 19.53 68.278 19.578 68.314 ;
      RECT 16.882 68.278 16.936 68.314 ;
      RECT 16.422 68.278 16.47 68.314 ;
      RECT 16.114 68.278 16.162 68.314 ;
      RECT 14.132 68.278 14.186 68.314 ;
      RECT 13.294 68.278 13.346 68.314 ;
      RECT 12.894 68.278 12.946 68.314 ;
      RECT 12.494 68.278 12.546 68.314 ;
      RECT 12.094 68.278 12.146 68.314 ;
      RECT 11.694 68.278 11.746 68.314 ;
      RECT 11.294 68.278 11.346 68.314 ;
      RECT 10.894 68.278 10.946 68.314 ;
      RECT 10.494 68.278 10.546 68.314 ;
      RECT 10.094 68.278 10.146 68.314 ;
      RECT 9.694 68.278 9.746 68.314 ;
      RECT 9.294 68.278 9.346 68.314 ;
      RECT 8.894 68.278 8.946 68.314 ;
      RECT 8.494 68.278 8.546 68.314 ;
      RECT 8.094 68.278 8.146 68.314 ;
      RECT 7.694 68.278 7.746 68.314 ;
      RECT 7.294 68.278 7.346 68.314 ;
      RECT 6.894 68.278 6.946 68.314 ;
      RECT 6.494 68.278 6.546 68.314 ;
      RECT 6.094 68.278 6.146 68.314 ;
      RECT 5.694 68.278 5.746 68.314 ;
      RECT 5.294 68.278 5.346 68.314 ;
      RECT 4.894 68.278 4.946 68.314 ;
      RECT 4.494 68.278 4.546 68.314 ;
      RECT 4.094 68.278 4.146 68.314 ;
      RECT 3.694 68.278 3.746 68.314 ;
      RECT 3.294 68.278 3.346 68.314 ;
      RECT 2.894 68.278 2.946 68.314 ;
      RECT 2.494 68.278 2.546 68.314 ;
      RECT 2.094 68.278 2.146 68.314 ;
      RECT 1.694 68.278 1.746 68.314 ;
      RECT 1.294 68.278 1.346 68.314 ;
      RECT 0.894 68.278 0.946 68.314 ;
      RECT 21.414 68.202 21.468 68.238 ;
      RECT 14.532 68.202 14.586 68.238 ;
      RECT 19.606 68.049 19.654 68.085 ;
      RECT 18.08 68.049 18.12 68.085 ;
      RECT 16.718 68.049 16.772 68.085 ;
      RECT 16.346 68.049 16.394 68.085 ;
      RECT 20.37 68.0545 20.442 68.0795 ;
      RECT 18.764 68.0545 18.836 68.0795 ;
      RECT 15.558 68.0545 15.63 68.0795 ;
      RECT 21.978 67.902 22.022 67.938 ;
      RECT 13.978 67.902 14.022 67.938 ;
      RECT 18.764 67.9075 18.836 67.9325 ;
      RECT 19.762 67.755 19.81 67.791 ;
      RECT 17.616 67.755 17.656 67.791 ;
      RECT 16.19 67.755 16.238 67.791 ;
      RECT 35.254 67.526 35.306 67.562 ;
      RECT 34.854 67.526 34.906 67.562 ;
      RECT 34.454 67.526 34.506 67.562 ;
      RECT 34.054 67.526 34.106 67.562 ;
      RECT 33.654 67.526 33.706 67.562 ;
      RECT 33.254 67.526 33.306 67.562 ;
      RECT 32.854 67.526 32.906 67.562 ;
      RECT 32.454 67.526 32.506 67.562 ;
      RECT 32.054 67.526 32.106 67.562 ;
      RECT 31.654 67.526 31.706 67.562 ;
      RECT 31.254 67.526 31.306 67.562 ;
      RECT 30.854 67.526 30.906 67.562 ;
      RECT 30.454 67.526 30.506 67.562 ;
      RECT 30.054 67.526 30.106 67.562 ;
      RECT 29.654 67.526 29.706 67.562 ;
      RECT 29.254 67.526 29.306 67.562 ;
      RECT 28.854 67.526 28.906 67.562 ;
      RECT 28.454 67.526 28.506 67.562 ;
      RECT 28.054 67.526 28.106 67.562 ;
      RECT 27.654 67.526 27.706 67.562 ;
      RECT 27.254 67.526 27.306 67.562 ;
      RECT 26.854 67.526 26.906 67.562 ;
      RECT 26.454 67.526 26.506 67.562 ;
      RECT 26.054 67.526 26.106 67.562 ;
      RECT 25.654 67.526 25.706 67.562 ;
      RECT 25.254 67.526 25.306 67.562 ;
      RECT 24.854 67.526 24.906 67.562 ;
      RECT 24.454 67.526 24.506 67.562 ;
      RECT 24.054 67.526 24.106 67.562 ;
      RECT 23.654 67.526 23.706 67.562 ;
      RECT 23.254 67.526 23.306 67.562 ;
      RECT 22.854 67.526 22.906 67.562 ;
      RECT 22.694 67.526 22.746 67.562 ;
      RECT 21.732 67.526 21.786 67.562 ;
      RECT 14.214 67.526 14.268 67.562 ;
      RECT 13.054 67.526 13.106 67.562 ;
      RECT 12.654 67.526 12.706 67.562 ;
      RECT 12.254 67.526 12.306 67.562 ;
      RECT 11.854 67.526 11.906 67.562 ;
      RECT 11.454 67.526 11.506 67.562 ;
      RECT 11.054 67.526 11.106 67.562 ;
      RECT 10.654 67.526 10.706 67.562 ;
      RECT 10.254 67.526 10.306 67.562 ;
      RECT 9.854 67.526 9.906 67.562 ;
      RECT 9.454 67.526 9.506 67.562 ;
      RECT 9.054 67.526 9.106 67.562 ;
      RECT 8.654 67.526 8.706 67.562 ;
      RECT 8.254 67.526 8.306 67.562 ;
      RECT 7.854 67.526 7.906 67.562 ;
      RECT 7.454 67.526 7.506 67.562 ;
      RECT 7.054 67.526 7.106 67.562 ;
      RECT 6.654 67.526 6.706 67.562 ;
      RECT 6.254 67.526 6.306 67.562 ;
      RECT 5.854 67.526 5.906 67.562 ;
      RECT 5.454 67.526 5.506 67.562 ;
      RECT 5.054 67.526 5.106 67.562 ;
      RECT 4.654 67.526 4.706 67.562 ;
      RECT 4.254 67.526 4.306 67.562 ;
      RECT 3.854 67.526 3.906 67.562 ;
      RECT 3.454 67.526 3.506 67.562 ;
      RECT 3.054 67.526 3.106 67.562 ;
      RECT 2.654 67.526 2.706 67.562 ;
      RECT 2.254 67.526 2.306 67.562 ;
      RECT 1.854 67.526 1.906 67.562 ;
      RECT 1.454 67.526 1.506 67.562 ;
      RECT 1.054 67.526 1.106 67.562 ;
      RECT 0.654 67.526 0.706 67.562 ;
      RECT 21.978 67.302 22.022 67.338 ;
      RECT 21.096 67.302 21.14 67.338 ;
      RECT 14.86 67.302 14.904 67.338 ;
      RECT 13.978 67.302 14.022 67.338 ;
      RECT 35.494 67.078 35.546 67.114 ;
      RECT 35.094 67.078 35.146 67.114 ;
      RECT 34.694 67.078 34.746 67.114 ;
      RECT 34.294 67.078 34.346 67.114 ;
      RECT 33.894 67.078 33.946 67.114 ;
      RECT 33.494 67.078 33.546 67.114 ;
      RECT 33.094 67.078 33.146 67.114 ;
      RECT 32.694 67.078 32.746 67.114 ;
      RECT 32.294 67.078 32.346 67.114 ;
      RECT 31.894 67.078 31.946 67.114 ;
      RECT 31.494 67.078 31.546 67.114 ;
      RECT 31.094 67.078 31.146 67.114 ;
      RECT 30.694 67.078 30.746 67.114 ;
      RECT 30.294 67.078 30.346 67.114 ;
      RECT 29.894 67.078 29.946 67.114 ;
      RECT 29.494 67.078 29.546 67.114 ;
      RECT 29.094 67.078 29.146 67.114 ;
      RECT 28.694 67.078 28.746 67.114 ;
      RECT 28.294 67.078 28.346 67.114 ;
      RECT 27.894 67.078 27.946 67.114 ;
      RECT 27.494 67.078 27.546 67.114 ;
      RECT 27.094 67.078 27.146 67.114 ;
      RECT 26.694 67.078 26.746 67.114 ;
      RECT 26.294 67.078 26.346 67.114 ;
      RECT 25.894 67.078 25.946 67.114 ;
      RECT 25.494 67.078 25.546 67.114 ;
      RECT 25.094 67.078 25.146 67.114 ;
      RECT 24.694 67.078 24.746 67.114 ;
      RECT 24.294 67.078 24.346 67.114 ;
      RECT 23.894 67.078 23.946 67.114 ;
      RECT 23.494 67.078 23.546 67.114 ;
      RECT 23.094 67.078 23.146 67.114 ;
      RECT 21.814 67.078 21.868 67.114 ;
      RECT 19.838 67.078 19.886 67.114 ;
      RECT 19.53 67.078 19.578 67.114 ;
      RECT 16.882 67.078 16.936 67.114 ;
      RECT 16.422 67.078 16.47 67.114 ;
      RECT 16.114 67.078 16.162 67.114 ;
      RECT 14.132 67.078 14.186 67.114 ;
      RECT 13.294 67.078 13.346 67.114 ;
      RECT 12.894 67.078 12.946 67.114 ;
      RECT 12.494 67.078 12.546 67.114 ;
      RECT 12.094 67.078 12.146 67.114 ;
      RECT 11.694 67.078 11.746 67.114 ;
      RECT 11.294 67.078 11.346 67.114 ;
      RECT 10.894 67.078 10.946 67.114 ;
      RECT 10.494 67.078 10.546 67.114 ;
      RECT 10.094 67.078 10.146 67.114 ;
      RECT 9.694 67.078 9.746 67.114 ;
      RECT 9.294 67.078 9.346 67.114 ;
      RECT 8.894 67.078 8.946 67.114 ;
      RECT 8.494 67.078 8.546 67.114 ;
      RECT 8.094 67.078 8.146 67.114 ;
      RECT 7.694 67.078 7.746 67.114 ;
      RECT 7.294 67.078 7.346 67.114 ;
      RECT 6.894 67.078 6.946 67.114 ;
      RECT 6.494 67.078 6.546 67.114 ;
      RECT 6.094 67.078 6.146 67.114 ;
      RECT 5.694 67.078 5.746 67.114 ;
      RECT 5.294 67.078 5.346 67.114 ;
      RECT 4.894 67.078 4.946 67.114 ;
      RECT 4.494 67.078 4.546 67.114 ;
      RECT 4.094 67.078 4.146 67.114 ;
      RECT 3.694 67.078 3.746 67.114 ;
      RECT 3.294 67.078 3.346 67.114 ;
      RECT 2.894 67.078 2.946 67.114 ;
      RECT 2.494 67.078 2.546 67.114 ;
      RECT 2.094 67.078 2.146 67.114 ;
      RECT 1.694 67.078 1.746 67.114 ;
      RECT 1.294 67.078 1.346 67.114 ;
      RECT 0.894 67.078 0.946 67.114 ;
      RECT 21.414 67.002 21.468 67.038 ;
      RECT 14.532 67.002 14.586 67.038 ;
      RECT 19.606 66.849 19.654 66.885 ;
      RECT 18.08 66.849 18.12 66.885 ;
      RECT 16.718 66.849 16.772 66.885 ;
      RECT 16.346 66.849 16.394 66.885 ;
      RECT 20.37 66.8545 20.442 66.8795 ;
      RECT 18.764 66.8545 18.836 66.8795 ;
      RECT 15.558 66.8545 15.63 66.8795 ;
      RECT 21.978 66.702 22.022 66.738 ;
      RECT 13.978 66.702 14.022 66.738 ;
      RECT 18.764 66.7075 18.836 66.7325 ;
      RECT 19.762 66.555 19.81 66.591 ;
      RECT 17.616 66.555 17.656 66.591 ;
      RECT 16.19 66.555 16.238 66.591 ;
      RECT 35.254 66.326 35.306 66.362 ;
      RECT 34.854 66.326 34.906 66.362 ;
      RECT 34.454 66.326 34.506 66.362 ;
      RECT 34.054 66.326 34.106 66.362 ;
      RECT 33.654 66.326 33.706 66.362 ;
      RECT 33.254 66.326 33.306 66.362 ;
      RECT 32.854 66.326 32.906 66.362 ;
      RECT 32.454 66.326 32.506 66.362 ;
      RECT 32.054 66.326 32.106 66.362 ;
      RECT 31.654 66.326 31.706 66.362 ;
      RECT 31.254 66.326 31.306 66.362 ;
      RECT 30.854 66.326 30.906 66.362 ;
      RECT 30.454 66.326 30.506 66.362 ;
      RECT 30.054 66.326 30.106 66.362 ;
      RECT 29.654 66.326 29.706 66.362 ;
      RECT 29.254 66.326 29.306 66.362 ;
      RECT 28.854 66.326 28.906 66.362 ;
      RECT 28.454 66.326 28.506 66.362 ;
      RECT 28.054 66.326 28.106 66.362 ;
      RECT 27.654 66.326 27.706 66.362 ;
      RECT 27.254 66.326 27.306 66.362 ;
      RECT 26.854 66.326 26.906 66.362 ;
      RECT 26.454 66.326 26.506 66.362 ;
      RECT 26.054 66.326 26.106 66.362 ;
      RECT 25.654 66.326 25.706 66.362 ;
      RECT 25.254 66.326 25.306 66.362 ;
      RECT 24.854 66.326 24.906 66.362 ;
      RECT 24.454 66.326 24.506 66.362 ;
      RECT 24.054 66.326 24.106 66.362 ;
      RECT 23.654 66.326 23.706 66.362 ;
      RECT 23.254 66.326 23.306 66.362 ;
      RECT 22.854 66.326 22.906 66.362 ;
      RECT 22.694 66.326 22.746 66.362 ;
      RECT 21.732 66.326 21.786 66.362 ;
      RECT 14.214 66.326 14.268 66.362 ;
      RECT 13.054 66.326 13.106 66.362 ;
      RECT 12.654 66.326 12.706 66.362 ;
      RECT 12.254 66.326 12.306 66.362 ;
      RECT 11.854 66.326 11.906 66.362 ;
      RECT 11.454 66.326 11.506 66.362 ;
      RECT 11.054 66.326 11.106 66.362 ;
      RECT 10.654 66.326 10.706 66.362 ;
      RECT 10.254 66.326 10.306 66.362 ;
      RECT 9.854 66.326 9.906 66.362 ;
      RECT 9.454 66.326 9.506 66.362 ;
      RECT 9.054 66.326 9.106 66.362 ;
      RECT 8.654 66.326 8.706 66.362 ;
      RECT 8.254 66.326 8.306 66.362 ;
      RECT 7.854 66.326 7.906 66.362 ;
      RECT 7.454 66.326 7.506 66.362 ;
      RECT 7.054 66.326 7.106 66.362 ;
      RECT 6.654 66.326 6.706 66.362 ;
      RECT 6.254 66.326 6.306 66.362 ;
      RECT 5.854 66.326 5.906 66.362 ;
      RECT 5.454 66.326 5.506 66.362 ;
      RECT 5.054 66.326 5.106 66.362 ;
      RECT 4.654 66.326 4.706 66.362 ;
      RECT 4.254 66.326 4.306 66.362 ;
      RECT 3.854 66.326 3.906 66.362 ;
      RECT 3.454 66.326 3.506 66.362 ;
      RECT 3.054 66.326 3.106 66.362 ;
      RECT 2.654 66.326 2.706 66.362 ;
      RECT 2.254 66.326 2.306 66.362 ;
      RECT 1.854 66.326 1.906 66.362 ;
      RECT 1.454 66.326 1.506 66.362 ;
      RECT 1.054 66.326 1.106 66.362 ;
      RECT 0.654 66.326 0.706 66.362 ;
      RECT 21.978 66.102 22.022 66.138 ;
      RECT 21.096 66.102 21.14 66.138 ;
      RECT 14.86 66.102 14.904 66.138 ;
      RECT 13.978 66.102 14.022 66.138 ;
      RECT 35.494 65.878 35.546 65.914 ;
      RECT 35.094 65.878 35.146 65.914 ;
      RECT 34.694 65.878 34.746 65.914 ;
      RECT 34.294 65.878 34.346 65.914 ;
      RECT 33.894 65.878 33.946 65.914 ;
      RECT 33.494 65.878 33.546 65.914 ;
      RECT 33.094 65.878 33.146 65.914 ;
      RECT 32.694 65.878 32.746 65.914 ;
      RECT 32.294 65.878 32.346 65.914 ;
      RECT 31.894 65.878 31.946 65.914 ;
      RECT 31.494 65.878 31.546 65.914 ;
      RECT 31.094 65.878 31.146 65.914 ;
      RECT 30.694 65.878 30.746 65.914 ;
      RECT 30.294 65.878 30.346 65.914 ;
      RECT 29.894 65.878 29.946 65.914 ;
      RECT 29.494 65.878 29.546 65.914 ;
      RECT 29.094 65.878 29.146 65.914 ;
      RECT 28.694 65.878 28.746 65.914 ;
      RECT 28.294 65.878 28.346 65.914 ;
      RECT 27.894 65.878 27.946 65.914 ;
      RECT 27.494 65.878 27.546 65.914 ;
      RECT 27.094 65.878 27.146 65.914 ;
      RECT 26.694 65.878 26.746 65.914 ;
      RECT 26.294 65.878 26.346 65.914 ;
      RECT 25.894 65.878 25.946 65.914 ;
      RECT 25.494 65.878 25.546 65.914 ;
      RECT 25.094 65.878 25.146 65.914 ;
      RECT 24.694 65.878 24.746 65.914 ;
      RECT 24.294 65.878 24.346 65.914 ;
      RECT 23.894 65.878 23.946 65.914 ;
      RECT 23.494 65.878 23.546 65.914 ;
      RECT 23.094 65.878 23.146 65.914 ;
      RECT 21.814 65.878 21.868 65.914 ;
      RECT 19.838 65.878 19.886 65.914 ;
      RECT 19.53 65.878 19.578 65.914 ;
      RECT 16.882 65.878 16.936 65.914 ;
      RECT 16.422 65.878 16.47 65.914 ;
      RECT 16.114 65.878 16.162 65.914 ;
      RECT 14.132 65.878 14.186 65.914 ;
      RECT 13.294 65.878 13.346 65.914 ;
      RECT 12.894 65.878 12.946 65.914 ;
      RECT 12.494 65.878 12.546 65.914 ;
      RECT 12.094 65.878 12.146 65.914 ;
      RECT 11.694 65.878 11.746 65.914 ;
      RECT 11.294 65.878 11.346 65.914 ;
      RECT 10.894 65.878 10.946 65.914 ;
      RECT 10.494 65.878 10.546 65.914 ;
      RECT 10.094 65.878 10.146 65.914 ;
      RECT 9.694 65.878 9.746 65.914 ;
      RECT 9.294 65.878 9.346 65.914 ;
      RECT 8.894 65.878 8.946 65.914 ;
      RECT 8.494 65.878 8.546 65.914 ;
      RECT 8.094 65.878 8.146 65.914 ;
      RECT 7.694 65.878 7.746 65.914 ;
      RECT 7.294 65.878 7.346 65.914 ;
      RECT 6.894 65.878 6.946 65.914 ;
      RECT 6.494 65.878 6.546 65.914 ;
      RECT 6.094 65.878 6.146 65.914 ;
      RECT 5.694 65.878 5.746 65.914 ;
      RECT 5.294 65.878 5.346 65.914 ;
      RECT 4.894 65.878 4.946 65.914 ;
      RECT 4.494 65.878 4.546 65.914 ;
      RECT 4.094 65.878 4.146 65.914 ;
      RECT 3.694 65.878 3.746 65.914 ;
      RECT 3.294 65.878 3.346 65.914 ;
      RECT 2.894 65.878 2.946 65.914 ;
      RECT 2.494 65.878 2.546 65.914 ;
      RECT 2.094 65.878 2.146 65.914 ;
      RECT 1.694 65.878 1.746 65.914 ;
      RECT 1.294 65.878 1.346 65.914 ;
      RECT 0.894 65.878 0.946 65.914 ;
      RECT 21.414 65.802 21.468 65.838 ;
      RECT 14.532 65.802 14.586 65.838 ;
      RECT 19.606 65.649 19.654 65.685 ;
      RECT 18.08 65.649 18.12 65.685 ;
      RECT 16.718 65.649 16.772 65.685 ;
      RECT 16.346 65.649 16.394 65.685 ;
      RECT 20.37 65.6545 20.442 65.6795 ;
      RECT 18.764 65.6545 18.836 65.6795 ;
      RECT 15.558 65.6545 15.63 65.6795 ;
      RECT 21.978 65.502 22.022 65.538 ;
      RECT 13.978 65.502 14.022 65.538 ;
      RECT 18.764 65.5075 18.836 65.5325 ;
      RECT 19.762 65.355 19.81 65.391 ;
      RECT 17.616 65.355 17.656 65.391 ;
      RECT 16.19 65.355 16.238 65.391 ;
      RECT 35.254 65.126 35.306 65.162 ;
      RECT 34.854 65.126 34.906 65.162 ;
      RECT 34.454 65.126 34.506 65.162 ;
      RECT 34.054 65.126 34.106 65.162 ;
      RECT 33.654 65.126 33.706 65.162 ;
      RECT 33.254 65.126 33.306 65.162 ;
      RECT 32.854 65.126 32.906 65.162 ;
      RECT 32.454 65.126 32.506 65.162 ;
      RECT 32.054 65.126 32.106 65.162 ;
      RECT 31.654 65.126 31.706 65.162 ;
      RECT 31.254 65.126 31.306 65.162 ;
      RECT 30.854 65.126 30.906 65.162 ;
      RECT 30.454 65.126 30.506 65.162 ;
      RECT 30.054 65.126 30.106 65.162 ;
      RECT 29.654 65.126 29.706 65.162 ;
      RECT 29.254 65.126 29.306 65.162 ;
      RECT 28.854 65.126 28.906 65.162 ;
      RECT 28.454 65.126 28.506 65.162 ;
      RECT 28.054 65.126 28.106 65.162 ;
      RECT 27.654 65.126 27.706 65.162 ;
      RECT 27.254 65.126 27.306 65.162 ;
      RECT 26.854 65.126 26.906 65.162 ;
      RECT 26.454 65.126 26.506 65.162 ;
      RECT 26.054 65.126 26.106 65.162 ;
      RECT 25.654 65.126 25.706 65.162 ;
      RECT 25.254 65.126 25.306 65.162 ;
      RECT 24.854 65.126 24.906 65.162 ;
      RECT 24.454 65.126 24.506 65.162 ;
      RECT 24.054 65.126 24.106 65.162 ;
      RECT 23.654 65.126 23.706 65.162 ;
      RECT 23.254 65.126 23.306 65.162 ;
      RECT 22.854 65.126 22.906 65.162 ;
      RECT 22.694 65.126 22.746 65.162 ;
      RECT 21.732 65.126 21.786 65.162 ;
      RECT 14.214 65.126 14.268 65.162 ;
      RECT 13.054 65.126 13.106 65.162 ;
      RECT 12.654 65.126 12.706 65.162 ;
      RECT 12.254 65.126 12.306 65.162 ;
      RECT 11.854 65.126 11.906 65.162 ;
      RECT 11.454 65.126 11.506 65.162 ;
      RECT 11.054 65.126 11.106 65.162 ;
      RECT 10.654 65.126 10.706 65.162 ;
      RECT 10.254 65.126 10.306 65.162 ;
      RECT 9.854 65.126 9.906 65.162 ;
      RECT 9.454 65.126 9.506 65.162 ;
      RECT 9.054 65.126 9.106 65.162 ;
      RECT 8.654 65.126 8.706 65.162 ;
      RECT 8.254 65.126 8.306 65.162 ;
      RECT 7.854 65.126 7.906 65.162 ;
      RECT 7.454 65.126 7.506 65.162 ;
      RECT 7.054 65.126 7.106 65.162 ;
      RECT 6.654 65.126 6.706 65.162 ;
      RECT 6.254 65.126 6.306 65.162 ;
      RECT 5.854 65.126 5.906 65.162 ;
      RECT 5.454 65.126 5.506 65.162 ;
      RECT 5.054 65.126 5.106 65.162 ;
      RECT 4.654 65.126 4.706 65.162 ;
      RECT 4.254 65.126 4.306 65.162 ;
      RECT 3.854 65.126 3.906 65.162 ;
      RECT 3.454 65.126 3.506 65.162 ;
      RECT 3.054 65.126 3.106 65.162 ;
      RECT 2.654 65.126 2.706 65.162 ;
      RECT 2.254 65.126 2.306 65.162 ;
      RECT 1.854 65.126 1.906 65.162 ;
      RECT 1.454 65.126 1.506 65.162 ;
      RECT 1.054 65.126 1.106 65.162 ;
      RECT 0.654 65.126 0.706 65.162 ;
      RECT 21.978 64.902 22.022 64.938 ;
      RECT 21.096 64.902 21.14 64.938 ;
      RECT 14.86 64.902 14.904 64.938 ;
      RECT 13.978 64.902 14.022 64.938 ;
      RECT 35.494 64.678 35.546 64.714 ;
      RECT 35.094 64.678 35.146 64.714 ;
      RECT 34.694 64.678 34.746 64.714 ;
      RECT 34.294 64.678 34.346 64.714 ;
      RECT 33.894 64.678 33.946 64.714 ;
      RECT 33.494 64.678 33.546 64.714 ;
      RECT 33.094 64.678 33.146 64.714 ;
      RECT 32.694 64.678 32.746 64.714 ;
      RECT 32.294 64.678 32.346 64.714 ;
      RECT 31.894 64.678 31.946 64.714 ;
      RECT 31.494 64.678 31.546 64.714 ;
      RECT 31.094 64.678 31.146 64.714 ;
      RECT 30.694 64.678 30.746 64.714 ;
      RECT 30.294 64.678 30.346 64.714 ;
      RECT 29.894 64.678 29.946 64.714 ;
      RECT 29.494 64.678 29.546 64.714 ;
      RECT 29.094 64.678 29.146 64.714 ;
      RECT 28.694 64.678 28.746 64.714 ;
      RECT 28.294 64.678 28.346 64.714 ;
      RECT 27.894 64.678 27.946 64.714 ;
      RECT 27.494 64.678 27.546 64.714 ;
      RECT 27.094 64.678 27.146 64.714 ;
      RECT 26.694 64.678 26.746 64.714 ;
      RECT 26.294 64.678 26.346 64.714 ;
      RECT 25.894 64.678 25.946 64.714 ;
      RECT 25.494 64.678 25.546 64.714 ;
      RECT 25.094 64.678 25.146 64.714 ;
      RECT 24.694 64.678 24.746 64.714 ;
      RECT 24.294 64.678 24.346 64.714 ;
      RECT 23.894 64.678 23.946 64.714 ;
      RECT 23.494 64.678 23.546 64.714 ;
      RECT 23.094 64.678 23.146 64.714 ;
      RECT 21.814 64.678 21.868 64.714 ;
      RECT 19.838 64.678 19.886 64.714 ;
      RECT 19.53 64.678 19.578 64.714 ;
      RECT 16.882 64.678 16.936 64.714 ;
      RECT 16.422 64.678 16.47 64.714 ;
      RECT 16.114 64.678 16.162 64.714 ;
      RECT 14.132 64.678 14.186 64.714 ;
      RECT 13.294 64.678 13.346 64.714 ;
      RECT 12.894 64.678 12.946 64.714 ;
      RECT 12.494 64.678 12.546 64.714 ;
      RECT 12.094 64.678 12.146 64.714 ;
      RECT 11.694 64.678 11.746 64.714 ;
      RECT 11.294 64.678 11.346 64.714 ;
      RECT 10.894 64.678 10.946 64.714 ;
      RECT 10.494 64.678 10.546 64.714 ;
      RECT 10.094 64.678 10.146 64.714 ;
      RECT 9.694 64.678 9.746 64.714 ;
      RECT 9.294 64.678 9.346 64.714 ;
      RECT 8.894 64.678 8.946 64.714 ;
      RECT 8.494 64.678 8.546 64.714 ;
      RECT 8.094 64.678 8.146 64.714 ;
      RECT 7.694 64.678 7.746 64.714 ;
      RECT 7.294 64.678 7.346 64.714 ;
      RECT 6.894 64.678 6.946 64.714 ;
      RECT 6.494 64.678 6.546 64.714 ;
      RECT 6.094 64.678 6.146 64.714 ;
      RECT 5.694 64.678 5.746 64.714 ;
      RECT 5.294 64.678 5.346 64.714 ;
      RECT 4.894 64.678 4.946 64.714 ;
      RECT 4.494 64.678 4.546 64.714 ;
      RECT 4.094 64.678 4.146 64.714 ;
      RECT 3.694 64.678 3.746 64.714 ;
      RECT 3.294 64.678 3.346 64.714 ;
      RECT 2.894 64.678 2.946 64.714 ;
      RECT 2.494 64.678 2.546 64.714 ;
      RECT 2.094 64.678 2.146 64.714 ;
      RECT 1.694 64.678 1.746 64.714 ;
      RECT 1.294 64.678 1.346 64.714 ;
      RECT 0.894 64.678 0.946 64.714 ;
      RECT 21.414 64.602 21.468 64.638 ;
      RECT 14.532 64.602 14.586 64.638 ;
      RECT 19.606 64.449 19.654 64.485 ;
      RECT 18.08 64.449 18.12 64.485 ;
      RECT 16.718 64.449 16.772 64.485 ;
      RECT 16.346 64.449 16.394 64.485 ;
      RECT 20.37 64.4545 20.442 64.4795 ;
      RECT 18.764 64.4545 18.836 64.4795 ;
      RECT 15.558 64.4545 15.63 64.4795 ;
      RECT 21.978 64.302 22.022 64.338 ;
      RECT 13.978 64.302 14.022 64.338 ;
      RECT 18.764 64.3075 18.836 64.3325 ;
      RECT 19.762 64.155 19.81 64.191 ;
      RECT 17.616 64.155 17.656 64.191 ;
      RECT 16.19 64.155 16.238 64.191 ;
      RECT 35.254 63.926 35.306 63.962 ;
      RECT 34.854 63.926 34.906 63.962 ;
      RECT 34.454 63.926 34.506 63.962 ;
      RECT 34.054 63.926 34.106 63.962 ;
      RECT 33.654 63.926 33.706 63.962 ;
      RECT 33.254 63.926 33.306 63.962 ;
      RECT 32.854 63.926 32.906 63.962 ;
      RECT 32.454 63.926 32.506 63.962 ;
      RECT 32.054 63.926 32.106 63.962 ;
      RECT 31.654 63.926 31.706 63.962 ;
      RECT 31.254 63.926 31.306 63.962 ;
      RECT 30.854 63.926 30.906 63.962 ;
      RECT 30.454 63.926 30.506 63.962 ;
      RECT 30.054 63.926 30.106 63.962 ;
      RECT 29.654 63.926 29.706 63.962 ;
      RECT 29.254 63.926 29.306 63.962 ;
      RECT 28.854 63.926 28.906 63.962 ;
      RECT 28.454 63.926 28.506 63.962 ;
      RECT 28.054 63.926 28.106 63.962 ;
      RECT 27.654 63.926 27.706 63.962 ;
      RECT 27.254 63.926 27.306 63.962 ;
      RECT 26.854 63.926 26.906 63.962 ;
      RECT 26.454 63.926 26.506 63.962 ;
      RECT 26.054 63.926 26.106 63.962 ;
      RECT 25.654 63.926 25.706 63.962 ;
      RECT 25.254 63.926 25.306 63.962 ;
      RECT 24.854 63.926 24.906 63.962 ;
      RECT 24.454 63.926 24.506 63.962 ;
      RECT 24.054 63.926 24.106 63.962 ;
      RECT 23.654 63.926 23.706 63.962 ;
      RECT 23.254 63.926 23.306 63.962 ;
      RECT 22.854 63.926 22.906 63.962 ;
      RECT 22.694 63.926 22.746 63.962 ;
      RECT 21.732 63.926 21.786 63.962 ;
      RECT 14.214 63.926 14.268 63.962 ;
      RECT 13.054 63.926 13.106 63.962 ;
      RECT 12.654 63.926 12.706 63.962 ;
      RECT 12.254 63.926 12.306 63.962 ;
      RECT 11.854 63.926 11.906 63.962 ;
      RECT 11.454 63.926 11.506 63.962 ;
      RECT 11.054 63.926 11.106 63.962 ;
      RECT 10.654 63.926 10.706 63.962 ;
      RECT 10.254 63.926 10.306 63.962 ;
      RECT 9.854 63.926 9.906 63.962 ;
      RECT 9.454 63.926 9.506 63.962 ;
      RECT 9.054 63.926 9.106 63.962 ;
      RECT 8.654 63.926 8.706 63.962 ;
      RECT 8.254 63.926 8.306 63.962 ;
      RECT 7.854 63.926 7.906 63.962 ;
      RECT 7.454 63.926 7.506 63.962 ;
      RECT 7.054 63.926 7.106 63.962 ;
      RECT 6.654 63.926 6.706 63.962 ;
      RECT 6.254 63.926 6.306 63.962 ;
      RECT 5.854 63.926 5.906 63.962 ;
      RECT 5.454 63.926 5.506 63.962 ;
      RECT 5.054 63.926 5.106 63.962 ;
      RECT 4.654 63.926 4.706 63.962 ;
      RECT 4.254 63.926 4.306 63.962 ;
      RECT 3.854 63.926 3.906 63.962 ;
      RECT 3.454 63.926 3.506 63.962 ;
      RECT 3.054 63.926 3.106 63.962 ;
      RECT 2.654 63.926 2.706 63.962 ;
      RECT 2.254 63.926 2.306 63.962 ;
      RECT 1.854 63.926 1.906 63.962 ;
      RECT 1.454 63.926 1.506 63.962 ;
      RECT 1.054 63.926 1.106 63.962 ;
      RECT 0.654 63.926 0.706 63.962 ;
      RECT 21.978 63.702 22.022 63.738 ;
      RECT 21.096 63.702 21.14 63.738 ;
      RECT 14.86 63.702 14.904 63.738 ;
      RECT 13.978 63.702 14.022 63.738 ;
      RECT 35.494 63.478 35.546 63.514 ;
      RECT 35.094 63.478 35.146 63.514 ;
      RECT 34.694 63.478 34.746 63.514 ;
      RECT 34.294 63.478 34.346 63.514 ;
      RECT 33.894 63.478 33.946 63.514 ;
      RECT 33.494 63.478 33.546 63.514 ;
      RECT 33.094 63.478 33.146 63.514 ;
      RECT 32.694 63.478 32.746 63.514 ;
      RECT 32.294 63.478 32.346 63.514 ;
      RECT 31.894 63.478 31.946 63.514 ;
      RECT 31.494 63.478 31.546 63.514 ;
      RECT 31.094 63.478 31.146 63.514 ;
      RECT 30.694 63.478 30.746 63.514 ;
      RECT 30.294 63.478 30.346 63.514 ;
      RECT 29.894 63.478 29.946 63.514 ;
      RECT 29.494 63.478 29.546 63.514 ;
      RECT 29.094 63.478 29.146 63.514 ;
      RECT 28.694 63.478 28.746 63.514 ;
      RECT 28.294 63.478 28.346 63.514 ;
      RECT 27.894 63.478 27.946 63.514 ;
      RECT 27.494 63.478 27.546 63.514 ;
      RECT 27.094 63.478 27.146 63.514 ;
      RECT 26.694 63.478 26.746 63.514 ;
      RECT 26.294 63.478 26.346 63.514 ;
      RECT 25.894 63.478 25.946 63.514 ;
      RECT 25.494 63.478 25.546 63.514 ;
      RECT 25.094 63.478 25.146 63.514 ;
      RECT 24.694 63.478 24.746 63.514 ;
      RECT 24.294 63.478 24.346 63.514 ;
      RECT 23.894 63.478 23.946 63.514 ;
      RECT 23.494 63.478 23.546 63.514 ;
      RECT 23.094 63.478 23.146 63.514 ;
      RECT 21.814 63.478 21.868 63.514 ;
      RECT 19.838 63.478 19.886 63.514 ;
      RECT 19.53 63.478 19.578 63.514 ;
      RECT 16.882 63.478 16.936 63.514 ;
      RECT 16.422 63.478 16.47 63.514 ;
      RECT 16.114 63.478 16.162 63.514 ;
      RECT 14.132 63.478 14.186 63.514 ;
      RECT 13.294 63.478 13.346 63.514 ;
      RECT 12.894 63.478 12.946 63.514 ;
      RECT 12.494 63.478 12.546 63.514 ;
      RECT 12.094 63.478 12.146 63.514 ;
      RECT 11.694 63.478 11.746 63.514 ;
      RECT 11.294 63.478 11.346 63.514 ;
      RECT 10.894 63.478 10.946 63.514 ;
      RECT 10.494 63.478 10.546 63.514 ;
      RECT 10.094 63.478 10.146 63.514 ;
      RECT 9.694 63.478 9.746 63.514 ;
      RECT 9.294 63.478 9.346 63.514 ;
      RECT 8.894 63.478 8.946 63.514 ;
      RECT 8.494 63.478 8.546 63.514 ;
      RECT 8.094 63.478 8.146 63.514 ;
      RECT 7.694 63.478 7.746 63.514 ;
      RECT 7.294 63.478 7.346 63.514 ;
      RECT 6.894 63.478 6.946 63.514 ;
      RECT 6.494 63.478 6.546 63.514 ;
      RECT 6.094 63.478 6.146 63.514 ;
      RECT 5.694 63.478 5.746 63.514 ;
      RECT 5.294 63.478 5.346 63.514 ;
      RECT 4.894 63.478 4.946 63.514 ;
      RECT 4.494 63.478 4.546 63.514 ;
      RECT 4.094 63.478 4.146 63.514 ;
      RECT 3.694 63.478 3.746 63.514 ;
      RECT 3.294 63.478 3.346 63.514 ;
      RECT 2.894 63.478 2.946 63.514 ;
      RECT 2.494 63.478 2.546 63.514 ;
      RECT 2.094 63.478 2.146 63.514 ;
      RECT 1.694 63.478 1.746 63.514 ;
      RECT 1.294 63.478 1.346 63.514 ;
      RECT 0.894 63.478 0.946 63.514 ;
      RECT 21.414 63.402 21.468 63.438 ;
      RECT 14.532 63.402 14.586 63.438 ;
      RECT 19.606 63.249 19.654 63.285 ;
      RECT 18.08 63.249 18.12 63.285 ;
      RECT 16.718 63.249 16.772 63.285 ;
      RECT 16.346 63.249 16.394 63.285 ;
      RECT 20.37 63.2545 20.442 63.2795 ;
      RECT 18.764 63.2545 18.836 63.2795 ;
      RECT 15.558 63.2545 15.63 63.2795 ;
      RECT 21.978 63.102 22.022 63.138 ;
      RECT 13.978 63.102 14.022 63.138 ;
      RECT 18.764 63.1075 18.836 63.1325 ;
      RECT 19.762 62.955 19.81 62.991 ;
      RECT 17.616 62.955 17.656 62.991 ;
      RECT 16.19 62.955 16.238 62.991 ;
      RECT 35.254 62.726 35.306 62.762 ;
      RECT 34.854 62.726 34.906 62.762 ;
      RECT 34.454 62.726 34.506 62.762 ;
      RECT 34.054 62.726 34.106 62.762 ;
      RECT 33.654 62.726 33.706 62.762 ;
      RECT 33.254 62.726 33.306 62.762 ;
      RECT 32.854 62.726 32.906 62.762 ;
      RECT 32.454 62.726 32.506 62.762 ;
      RECT 32.054 62.726 32.106 62.762 ;
      RECT 31.654 62.726 31.706 62.762 ;
      RECT 31.254 62.726 31.306 62.762 ;
      RECT 30.854 62.726 30.906 62.762 ;
      RECT 30.454 62.726 30.506 62.762 ;
      RECT 30.054 62.726 30.106 62.762 ;
      RECT 29.654 62.726 29.706 62.762 ;
      RECT 29.254 62.726 29.306 62.762 ;
      RECT 28.854 62.726 28.906 62.762 ;
      RECT 28.454 62.726 28.506 62.762 ;
      RECT 28.054 62.726 28.106 62.762 ;
      RECT 27.654 62.726 27.706 62.762 ;
      RECT 27.254 62.726 27.306 62.762 ;
      RECT 26.854 62.726 26.906 62.762 ;
      RECT 26.454 62.726 26.506 62.762 ;
      RECT 26.054 62.726 26.106 62.762 ;
      RECT 25.654 62.726 25.706 62.762 ;
      RECT 25.254 62.726 25.306 62.762 ;
      RECT 24.854 62.726 24.906 62.762 ;
      RECT 24.454 62.726 24.506 62.762 ;
      RECT 24.054 62.726 24.106 62.762 ;
      RECT 23.654 62.726 23.706 62.762 ;
      RECT 23.254 62.726 23.306 62.762 ;
      RECT 22.854 62.726 22.906 62.762 ;
      RECT 22.694 62.726 22.746 62.762 ;
      RECT 21.732 62.726 21.786 62.762 ;
      RECT 14.214 62.726 14.268 62.762 ;
      RECT 13.054 62.726 13.106 62.762 ;
      RECT 12.654 62.726 12.706 62.762 ;
      RECT 12.254 62.726 12.306 62.762 ;
      RECT 11.854 62.726 11.906 62.762 ;
      RECT 11.454 62.726 11.506 62.762 ;
      RECT 11.054 62.726 11.106 62.762 ;
      RECT 10.654 62.726 10.706 62.762 ;
      RECT 10.254 62.726 10.306 62.762 ;
      RECT 9.854 62.726 9.906 62.762 ;
      RECT 9.454 62.726 9.506 62.762 ;
      RECT 9.054 62.726 9.106 62.762 ;
      RECT 8.654 62.726 8.706 62.762 ;
      RECT 8.254 62.726 8.306 62.762 ;
      RECT 7.854 62.726 7.906 62.762 ;
      RECT 7.454 62.726 7.506 62.762 ;
      RECT 7.054 62.726 7.106 62.762 ;
      RECT 6.654 62.726 6.706 62.762 ;
      RECT 6.254 62.726 6.306 62.762 ;
      RECT 5.854 62.726 5.906 62.762 ;
      RECT 5.454 62.726 5.506 62.762 ;
      RECT 5.054 62.726 5.106 62.762 ;
      RECT 4.654 62.726 4.706 62.762 ;
      RECT 4.254 62.726 4.306 62.762 ;
      RECT 3.854 62.726 3.906 62.762 ;
      RECT 3.454 62.726 3.506 62.762 ;
      RECT 3.054 62.726 3.106 62.762 ;
      RECT 2.654 62.726 2.706 62.762 ;
      RECT 2.254 62.726 2.306 62.762 ;
      RECT 1.854 62.726 1.906 62.762 ;
      RECT 1.454 62.726 1.506 62.762 ;
      RECT 1.054 62.726 1.106 62.762 ;
      RECT 0.654 62.726 0.706 62.762 ;
      RECT 21.978 62.502 22.022 62.538 ;
      RECT 21.096 62.502 21.14 62.538 ;
      RECT 14.86 62.502 14.904 62.538 ;
      RECT 13.978 62.502 14.022 62.538 ;
      RECT 35.494 62.278 35.546 62.314 ;
      RECT 35.094 62.278 35.146 62.314 ;
      RECT 34.694 62.278 34.746 62.314 ;
      RECT 34.294 62.278 34.346 62.314 ;
      RECT 33.894 62.278 33.946 62.314 ;
      RECT 33.494 62.278 33.546 62.314 ;
      RECT 33.094 62.278 33.146 62.314 ;
      RECT 32.694 62.278 32.746 62.314 ;
      RECT 32.294 62.278 32.346 62.314 ;
      RECT 31.894 62.278 31.946 62.314 ;
      RECT 31.494 62.278 31.546 62.314 ;
      RECT 31.094 62.278 31.146 62.314 ;
      RECT 30.694 62.278 30.746 62.314 ;
      RECT 30.294 62.278 30.346 62.314 ;
      RECT 29.894 62.278 29.946 62.314 ;
      RECT 29.494 62.278 29.546 62.314 ;
      RECT 29.094 62.278 29.146 62.314 ;
      RECT 28.694 62.278 28.746 62.314 ;
      RECT 28.294 62.278 28.346 62.314 ;
      RECT 27.894 62.278 27.946 62.314 ;
      RECT 27.494 62.278 27.546 62.314 ;
      RECT 27.094 62.278 27.146 62.314 ;
      RECT 26.694 62.278 26.746 62.314 ;
      RECT 26.294 62.278 26.346 62.314 ;
      RECT 25.894 62.278 25.946 62.314 ;
      RECT 25.494 62.278 25.546 62.314 ;
      RECT 25.094 62.278 25.146 62.314 ;
      RECT 24.694 62.278 24.746 62.314 ;
      RECT 24.294 62.278 24.346 62.314 ;
      RECT 23.894 62.278 23.946 62.314 ;
      RECT 23.494 62.278 23.546 62.314 ;
      RECT 23.094 62.278 23.146 62.314 ;
      RECT 21.814 62.278 21.868 62.314 ;
      RECT 19.838 62.278 19.886 62.314 ;
      RECT 19.53 62.278 19.578 62.314 ;
      RECT 16.882 62.278 16.936 62.314 ;
      RECT 16.422 62.278 16.47 62.314 ;
      RECT 16.114 62.278 16.162 62.314 ;
      RECT 14.132 62.278 14.186 62.314 ;
      RECT 13.294 62.278 13.346 62.314 ;
      RECT 12.894 62.278 12.946 62.314 ;
      RECT 12.494 62.278 12.546 62.314 ;
      RECT 12.094 62.278 12.146 62.314 ;
      RECT 11.694 62.278 11.746 62.314 ;
      RECT 11.294 62.278 11.346 62.314 ;
      RECT 10.894 62.278 10.946 62.314 ;
      RECT 10.494 62.278 10.546 62.314 ;
      RECT 10.094 62.278 10.146 62.314 ;
      RECT 9.694 62.278 9.746 62.314 ;
      RECT 9.294 62.278 9.346 62.314 ;
      RECT 8.894 62.278 8.946 62.314 ;
      RECT 8.494 62.278 8.546 62.314 ;
      RECT 8.094 62.278 8.146 62.314 ;
      RECT 7.694 62.278 7.746 62.314 ;
      RECT 7.294 62.278 7.346 62.314 ;
      RECT 6.894 62.278 6.946 62.314 ;
      RECT 6.494 62.278 6.546 62.314 ;
      RECT 6.094 62.278 6.146 62.314 ;
      RECT 5.694 62.278 5.746 62.314 ;
      RECT 5.294 62.278 5.346 62.314 ;
      RECT 4.894 62.278 4.946 62.314 ;
      RECT 4.494 62.278 4.546 62.314 ;
      RECT 4.094 62.278 4.146 62.314 ;
      RECT 3.694 62.278 3.746 62.314 ;
      RECT 3.294 62.278 3.346 62.314 ;
      RECT 2.894 62.278 2.946 62.314 ;
      RECT 2.494 62.278 2.546 62.314 ;
      RECT 2.094 62.278 2.146 62.314 ;
      RECT 1.694 62.278 1.746 62.314 ;
      RECT 1.294 62.278 1.346 62.314 ;
      RECT 0.894 62.278 0.946 62.314 ;
      RECT 21.414 62.202 21.468 62.238 ;
      RECT 14.532 62.202 14.586 62.238 ;
      RECT 19.606 62.049 19.654 62.085 ;
      RECT 18.08 62.049 18.12 62.085 ;
      RECT 16.718 62.049 16.772 62.085 ;
      RECT 16.346 62.049 16.394 62.085 ;
      RECT 20.37 62.0545 20.442 62.0795 ;
      RECT 18.764 62.0545 18.836 62.0795 ;
      RECT 15.558 62.0545 15.63 62.0795 ;
      RECT 21.978 61.902 22.022 61.938 ;
      RECT 13.978 61.902 14.022 61.938 ;
      RECT 18.764 61.9075 18.836 61.9325 ;
      RECT 19.762 61.755 19.81 61.791 ;
      RECT 17.616 61.755 17.656 61.791 ;
      RECT 16.19 61.755 16.238 61.791 ;
      RECT 35.254 61.526 35.306 61.562 ;
      RECT 34.854 61.526 34.906 61.562 ;
      RECT 34.454 61.526 34.506 61.562 ;
      RECT 34.054 61.526 34.106 61.562 ;
      RECT 33.654 61.526 33.706 61.562 ;
      RECT 33.254 61.526 33.306 61.562 ;
      RECT 32.854 61.526 32.906 61.562 ;
      RECT 32.454 61.526 32.506 61.562 ;
      RECT 32.054 61.526 32.106 61.562 ;
      RECT 31.654 61.526 31.706 61.562 ;
      RECT 31.254 61.526 31.306 61.562 ;
      RECT 30.854 61.526 30.906 61.562 ;
      RECT 30.454 61.526 30.506 61.562 ;
      RECT 30.054 61.526 30.106 61.562 ;
      RECT 29.654 61.526 29.706 61.562 ;
      RECT 29.254 61.526 29.306 61.562 ;
      RECT 28.854 61.526 28.906 61.562 ;
      RECT 28.454 61.526 28.506 61.562 ;
      RECT 28.054 61.526 28.106 61.562 ;
      RECT 27.654 61.526 27.706 61.562 ;
      RECT 27.254 61.526 27.306 61.562 ;
      RECT 26.854 61.526 26.906 61.562 ;
      RECT 26.454 61.526 26.506 61.562 ;
      RECT 26.054 61.526 26.106 61.562 ;
      RECT 25.654 61.526 25.706 61.562 ;
      RECT 25.254 61.526 25.306 61.562 ;
      RECT 24.854 61.526 24.906 61.562 ;
      RECT 24.454 61.526 24.506 61.562 ;
      RECT 24.054 61.526 24.106 61.562 ;
      RECT 23.654 61.526 23.706 61.562 ;
      RECT 23.254 61.526 23.306 61.562 ;
      RECT 22.854 61.526 22.906 61.562 ;
      RECT 22.694 61.526 22.746 61.562 ;
      RECT 21.732 61.526 21.786 61.562 ;
      RECT 14.214 61.526 14.268 61.562 ;
      RECT 13.054 61.526 13.106 61.562 ;
      RECT 12.654 61.526 12.706 61.562 ;
      RECT 12.254 61.526 12.306 61.562 ;
      RECT 11.854 61.526 11.906 61.562 ;
      RECT 11.454 61.526 11.506 61.562 ;
      RECT 11.054 61.526 11.106 61.562 ;
      RECT 10.654 61.526 10.706 61.562 ;
      RECT 10.254 61.526 10.306 61.562 ;
      RECT 9.854 61.526 9.906 61.562 ;
      RECT 9.454 61.526 9.506 61.562 ;
      RECT 9.054 61.526 9.106 61.562 ;
      RECT 8.654 61.526 8.706 61.562 ;
      RECT 8.254 61.526 8.306 61.562 ;
      RECT 7.854 61.526 7.906 61.562 ;
      RECT 7.454 61.526 7.506 61.562 ;
      RECT 7.054 61.526 7.106 61.562 ;
      RECT 6.654 61.526 6.706 61.562 ;
      RECT 6.254 61.526 6.306 61.562 ;
      RECT 5.854 61.526 5.906 61.562 ;
      RECT 5.454 61.526 5.506 61.562 ;
      RECT 5.054 61.526 5.106 61.562 ;
      RECT 4.654 61.526 4.706 61.562 ;
      RECT 4.254 61.526 4.306 61.562 ;
      RECT 3.854 61.526 3.906 61.562 ;
      RECT 3.454 61.526 3.506 61.562 ;
      RECT 3.054 61.526 3.106 61.562 ;
      RECT 2.654 61.526 2.706 61.562 ;
      RECT 2.254 61.526 2.306 61.562 ;
      RECT 1.854 61.526 1.906 61.562 ;
      RECT 1.454 61.526 1.506 61.562 ;
      RECT 1.054 61.526 1.106 61.562 ;
      RECT 0.654 61.526 0.706 61.562 ;
      RECT 21.978 61.302 22.022 61.338 ;
      RECT 21.096 61.302 21.14 61.338 ;
      RECT 14.86 61.302 14.904 61.338 ;
      RECT 13.978 61.302 14.022 61.338 ;
      RECT 35.494 61.078 35.546 61.114 ;
      RECT 35.094 61.078 35.146 61.114 ;
      RECT 34.694 61.078 34.746 61.114 ;
      RECT 34.294 61.078 34.346 61.114 ;
      RECT 33.894 61.078 33.946 61.114 ;
      RECT 33.494 61.078 33.546 61.114 ;
      RECT 33.094 61.078 33.146 61.114 ;
      RECT 32.694 61.078 32.746 61.114 ;
      RECT 32.294 61.078 32.346 61.114 ;
      RECT 31.894 61.078 31.946 61.114 ;
      RECT 31.494 61.078 31.546 61.114 ;
      RECT 31.094 61.078 31.146 61.114 ;
      RECT 30.694 61.078 30.746 61.114 ;
      RECT 30.294 61.078 30.346 61.114 ;
      RECT 29.894 61.078 29.946 61.114 ;
      RECT 29.494 61.078 29.546 61.114 ;
      RECT 29.094 61.078 29.146 61.114 ;
      RECT 28.694 61.078 28.746 61.114 ;
      RECT 28.294 61.078 28.346 61.114 ;
      RECT 27.894 61.078 27.946 61.114 ;
      RECT 27.494 61.078 27.546 61.114 ;
      RECT 27.094 61.078 27.146 61.114 ;
      RECT 26.694 61.078 26.746 61.114 ;
      RECT 26.294 61.078 26.346 61.114 ;
      RECT 25.894 61.078 25.946 61.114 ;
      RECT 25.494 61.078 25.546 61.114 ;
      RECT 25.094 61.078 25.146 61.114 ;
      RECT 24.694 61.078 24.746 61.114 ;
      RECT 24.294 61.078 24.346 61.114 ;
      RECT 23.894 61.078 23.946 61.114 ;
      RECT 23.494 61.078 23.546 61.114 ;
      RECT 23.094 61.078 23.146 61.114 ;
      RECT 21.814 61.078 21.868 61.114 ;
      RECT 19.838 61.078 19.886 61.114 ;
      RECT 19.53 61.078 19.578 61.114 ;
      RECT 16.882 61.078 16.936 61.114 ;
      RECT 16.422 61.078 16.47 61.114 ;
      RECT 16.114 61.078 16.162 61.114 ;
      RECT 14.132 61.078 14.186 61.114 ;
      RECT 13.294 61.078 13.346 61.114 ;
      RECT 12.894 61.078 12.946 61.114 ;
      RECT 12.494 61.078 12.546 61.114 ;
      RECT 12.094 61.078 12.146 61.114 ;
      RECT 11.694 61.078 11.746 61.114 ;
      RECT 11.294 61.078 11.346 61.114 ;
      RECT 10.894 61.078 10.946 61.114 ;
      RECT 10.494 61.078 10.546 61.114 ;
      RECT 10.094 61.078 10.146 61.114 ;
      RECT 9.694 61.078 9.746 61.114 ;
      RECT 9.294 61.078 9.346 61.114 ;
      RECT 8.894 61.078 8.946 61.114 ;
      RECT 8.494 61.078 8.546 61.114 ;
      RECT 8.094 61.078 8.146 61.114 ;
      RECT 7.694 61.078 7.746 61.114 ;
      RECT 7.294 61.078 7.346 61.114 ;
      RECT 6.894 61.078 6.946 61.114 ;
      RECT 6.494 61.078 6.546 61.114 ;
      RECT 6.094 61.078 6.146 61.114 ;
      RECT 5.694 61.078 5.746 61.114 ;
      RECT 5.294 61.078 5.346 61.114 ;
      RECT 4.894 61.078 4.946 61.114 ;
      RECT 4.494 61.078 4.546 61.114 ;
      RECT 4.094 61.078 4.146 61.114 ;
      RECT 3.694 61.078 3.746 61.114 ;
      RECT 3.294 61.078 3.346 61.114 ;
      RECT 2.894 61.078 2.946 61.114 ;
      RECT 2.494 61.078 2.546 61.114 ;
      RECT 2.094 61.078 2.146 61.114 ;
      RECT 1.694 61.078 1.746 61.114 ;
      RECT 1.294 61.078 1.346 61.114 ;
      RECT 0.894 61.078 0.946 61.114 ;
      RECT 21.414 61.002 21.468 61.038 ;
      RECT 14.532 61.002 14.586 61.038 ;
      RECT 19.606 60.849 19.654 60.885 ;
      RECT 18.08 60.849 18.12 60.885 ;
      RECT 16.718 60.849 16.772 60.885 ;
      RECT 16.346 60.849 16.394 60.885 ;
      RECT 20.37 60.8545 20.442 60.8795 ;
      RECT 18.764 60.8545 18.836 60.8795 ;
      RECT 15.558 60.8545 15.63 60.8795 ;
      RECT 21.978 60.702 22.022 60.738 ;
      RECT 13.978 60.702 14.022 60.738 ;
      RECT 18.764 60.7075 18.836 60.7325 ;
      RECT 19.762 60.555 19.81 60.591 ;
      RECT 17.616 60.555 17.656 60.591 ;
      RECT 16.19 60.555 16.238 60.591 ;
      RECT 35.254 60.326 35.306 60.362 ;
      RECT 34.854 60.326 34.906 60.362 ;
      RECT 34.454 60.326 34.506 60.362 ;
      RECT 34.054 60.326 34.106 60.362 ;
      RECT 33.654 60.326 33.706 60.362 ;
      RECT 33.254 60.326 33.306 60.362 ;
      RECT 32.854 60.326 32.906 60.362 ;
      RECT 32.454 60.326 32.506 60.362 ;
      RECT 32.054 60.326 32.106 60.362 ;
      RECT 31.654 60.326 31.706 60.362 ;
      RECT 31.254 60.326 31.306 60.362 ;
      RECT 30.854 60.326 30.906 60.362 ;
      RECT 30.454 60.326 30.506 60.362 ;
      RECT 30.054 60.326 30.106 60.362 ;
      RECT 29.654 60.326 29.706 60.362 ;
      RECT 29.254 60.326 29.306 60.362 ;
      RECT 28.854 60.326 28.906 60.362 ;
      RECT 28.454 60.326 28.506 60.362 ;
      RECT 28.054 60.326 28.106 60.362 ;
      RECT 27.654 60.326 27.706 60.362 ;
      RECT 27.254 60.326 27.306 60.362 ;
      RECT 26.854 60.326 26.906 60.362 ;
      RECT 26.454 60.326 26.506 60.362 ;
      RECT 26.054 60.326 26.106 60.362 ;
      RECT 25.654 60.326 25.706 60.362 ;
      RECT 25.254 60.326 25.306 60.362 ;
      RECT 24.854 60.326 24.906 60.362 ;
      RECT 24.454 60.326 24.506 60.362 ;
      RECT 24.054 60.326 24.106 60.362 ;
      RECT 23.654 60.326 23.706 60.362 ;
      RECT 23.254 60.326 23.306 60.362 ;
      RECT 22.854 60.326 22.906 60.362 ;
      RECT 22.694 60.326 22.746 60.362 ;
      RECT 21.732 60.326 21.786 60.362 ;
      RECT 14.214 60.326 14.268 60.362 ;
      RECT 13.054 60.326 13.106 60.362 ;
      RECT 12.654 60.326 12.706 60.362 ;
      RECT 12.254 60.326 12.306 60.362 ;
      RECT 11.854 60.326 11.906 60.362 ;
      RECT 11.454 60.326 11.506 60.362 ;
      RECT 11.054 60.326 11.106 60.362 ;
      RECT 10.654 60.326 10.706 60.362 ;
      RECT 10.254 60.326 10.306 60.362 ;
      RECT 9.854 60.326 9.906 60.362 ;
      RECT 9.454 60.326 9.506 60.362 ;
      RECT 9.054 60.326 9.106 60.362 ;
      RECT 8.654 60.326 8.706 60.362 ;
      RECT 8.254 60.326 8.306 60.362 ;
      RECT 7.854 60.326 7.906 60.362 ;
      RECT 7.454 60.326 7.506 60.362 ;
      RECT 7.054 60.326 7.106 60.362 ;
      RECT 6.654 60.326 6.706 60.362 ;
      RECT 6.254 60.326 6.306 60.362 ;
      RECT 5.854 60.326 5.906 60.362 ;
      RECT 5.454 60.326 5.506 60.362 ;
      RECT 5.054 60.326 5.106 60.362 ;
      RECT 4.654 60.326 4.706 60.362 ;
      RECT 4.254 60.326 4.306 60.362 ;
      RECT 3.854 60.326 3.906 60.362 ;
      RECT 3.454 60.326 3.506 60.362 ;
      RECT 3.054 60.326 3.106 60.362 ;
      RECT 2.654 60.326 2.706 60.362 ;
      RECT 2.254 60.326 2.306 60.362 ;
      RECT 1.854 60.326 1.906 60.362 ;
      RECT 1.454 60.326 1.506 60.362 ;
      RECT 1.054 60.326 1.106 60.362 ;
      RECT 0.654 60.326 0.706 60.362 ;
      RECT 21.978 60.102 22.022 60.138 ;
      RECT 21.096 60.102 21.14 60.138 ;
      RECT 14.86 60.102 14.904 60.138 ;
      RECT 13.978 60.102 14.022 60.138 ;
      RECT 35.494 59.878 35.546 59.914 ;
      RECT 35.094 59.878 35.146 59.914 ;
      RECT 34.694 59.878 34.746 59.914 ;
      RECT 34.294 59.878 34.346 59.914 ;
      RECT 33.894 59.878 33.946 59.914 ;
      RECT 33.494 59.878 33.546 59.914 ;
      RECT 33.094 59.878 33.146 59.914 ;
      RECT 32.694 59.878 32.746 59.914 ;
      RECT 32.294 59.878 32.346 59.914 ;
      RECT 31.894 59.878 31.946 59.914 ;
      RECT 31.494 59.878 31.546 59.914 ;
      RECT 31.094 59.878 31.146 59.914 ;
      RECT 30.694 59.878 30.746 59.914 ;
      RECT 30.294 59.878 30.346 59.914 ;
      RECT 29.894 59.878 29.946 59.914 ;
      RECT 29.494 59.878 29.546 59.914 ;
      RECT 29.094 59.878 29.146 59.914 ;
      RECT 28.694 59.878 28.746 59.914 ;
      RECT 28.294 59.878 28.346 59.914 ;
      RECT 27.894 59.878 27.946 59.914 ;
      RECT 27.494 59.878 27.546 59.914 ;
      RECT 27.094 59.878 27.146 59.914 ;
      RECT 26.694 59.878 26.746 59.914 ;
      RECT 26.294 59.878 26.346 59.914 ;
      RECT 25.894 59.878 25.946 59.914 ;
      RECT 25.494 59.878 25.546 59.914 ;
      RECT 25.094 59.878 25.146 59.914 ;
      RECT 24.694 59.878 24.746 59.914 ;
      RECT 24.294 59.878 24.346 59.914 ;
      RECT 23.894 59.878 23.946 59.914 ;
      RECT 23.494 59.878 23.546 59.914 ;
      RECT 23.094 59.878 23.146 59.914 ;
      RECT 21.814 59.878 21.868 59.914 ;
      RECT 19.838 59.878 19.886 59.914 ;
      RECT 19.53 59.878 19.578 59.914 ;
      RECT 16.882 59.878 16.936 59.914 ;
      RECT 16.422 59.878 16.47 59.914 ;
      RECT 16.114 59.878 16.162 59.914 ;
      RECT 14.132 59.878 14.186 59.914 ;
      RECT 13.294 59.878 13.346 59.914 ;
      RECT 12.894 59.878 12.946 59.914 ;
      RECT 12.494 59.878 12.546 59.914 ;
      RECT 12.094 59.878 12.146 59.914 ;
      RECT 11.694 59.878 11.746 59.914 ;
      RECT 11.294 59.878 11.346 59.914 ;
      RECT 10.894 59.878 10.946 59.914 ;
      RECT 10.494 59.878 10.546 59.914 ;
      RECT 10.094 59.878 10.146 59.914 ;
      RECT 9.694 59.878 9.746 59.914 ;
      RECT 9.294 59.878 9.346 59.914 ;
      RECT 8.894 59.878 8.946 59.914 ;
      RECT 8.494 59.878 8.546 59.914 ;
      RECT 8.094 59.878 8.146 59.914 ;
      RECT 7.694 59.878 7.746 59.914 ;
      RECT 7.294 59.878 7.346 59.914 ;
      RECT 6.894 59.878 6.946 59.914 ;
      RECT 6.494 59.878 6.546 59.914 ;
      RECT 6.094 59.878 6.146 59.914 ;
      RECT 5.694 59.878 5.746 59.914 ;
      RECT 5.294 59.878 5.346 59.914 ;
      RECT 4.894 59.878 4.946 59.914 ;
      RECT 4.494 59.878 4.546 59.914 ;
      RECT 4.094 59.878 4.146 59.914 ;
      RECT 3.694 59.878 3.746 59.914 ;
      RECT 3.294 59.878 3.346 59.914 ;
      RECT 2.894 59.878 2.946 59.914 ;
      RECT 2.494 59.878 2.546 59.914 ;
      RECT 2.094 59.878 2.146 59.914 ;
      RECT 1.694 59.878 1.746 59.914 ;
      RECT 1.294 59.878 1.346 59.914 ;
      RECT 0.894 59.878 0.946 59.914 ;
      RECT 21.414 59.802 21.468 59.838 ;
      RECT 14.532 59.802 14.586 59.838 ;
      RECT 19.606 59.649 19.654 59.685 ;
      RECT 18.08 59.649 18.12 59.685 ;
      RECT 16.718 59.649 16.772 59.685 ;
      RECT 16.346 59.649 16.394 59.685 ;
      RECT 20.37 59.6545 20.442 59.6795 ;
      RECT 18.764 59.6545 18.836 59.6795 ;
      RECT 15.558 59.6545 15.63 59.6795 ;
      RECT 21.978 59.502 22.022 59.538 ;
      RECT 13.978 59.502 14.022 59.538 ;
      RECT 18.764 59.5075 18.836 59.5325 ;
      RECT 19.762 59.355 19.81 59.391 ;
      RECT 17.616 59.355 17.656 59.391 ;
      RECT 16.19 59.355 16.238 59.391 ;
      RECT 35.254 59.126 35.306 59.162 ;
      RECT 34.854 59.126 34.906 59.162 ;
      RECT 34.454 59.126 34.506 59.162 ;
      RECT 34.054 59.126 34.106 59.162 ;
      RECT 33.654 59.126 33.706 59.162 ;
      RECT 33.254 59.126 33.306 59.162 ;
      RECT 32.854 59.126 32.906 59.162 ;
      RECT 32.454 59.126 32.506 59.162 ;
      RECT 32.054 59.126 32.106 59.162 ;
      RECT 31.654 59.126 31.706 59.162 ;
      RECT 31.254 59.126 31.306 59.162 ;
      RECT 30.854 59.126 30.906 59.162 ;
      RECT 30.454 59.126 30.506 59.162 ;
      RECT 30.054 59.126 30.106 59.162 ;
      RECT 29.654 59.126 29.706 59.162 ;
      RECT 29.254 59.126 29.306 59.162 ;
      RECT 28.854 59.126 28.906 59.162 ;
      RECT 28.454 59.126 28.506 59.162 ;
      RECT 28.054 59.126 28.106 59.162 ;
      RECT 27.654 59.126 27.706 59.162 ;
      RECT 27.254 59.126 27.306 59.162 ;
      RECT 26.854 59.126 26.906 59.162 ;
      RECT 26.454 59.126 26.506 59.162 ;
      RECT 26.054 59.126 26.106 59.162 ;
      RECT 25.654 59.126 25.706 59.162 ;
      RECT 25.254 59.126 25.306 59.162 ;
      RECT 24.854 59.126 24.906 59.162 ;
      RECT 24.454 59.126 24.506 59.162 ;
      RECT 24.054 59.126 24.106 59.162 ;
      RECT 23.654 59.126 23.706 59.162 ;
      RECT 23.254 59.126 23.306 59.162 ;
      RECT 22.854 59.126 22.906 59.162 ;
      RECT 22.694 59.126 22.746 59.162 ;
      RECT 21.732 59.126 21.786 59.162 ;
      RECT 14.214 59.126 14.268 59.162 ;
      RECT 13.054 59.126 13.106 59.162 ;
      RECT 12.654 59.126 12.706 59.162 ;
      RECT 12.254 59.126 12.306 59.162 ;
      RECT 11.854 59.126 11.906 59.162 ;
      RECT 11.454 59.126 11.506 59.162 ;
      RECT 11.054 59.126 11.106 59.162 ;
      RECT 10.654 59.126 10.706 59.162 ;
      RECT 10.254 59.126 10.306 59.162 ;
      RECT 9.854 59.126 9.906 59.162 ;
      RECT 9.454 59.126 9.506 59.162 ;
      RECT 9.054 59.126 9.106 59.162 ;
      RECT 8.654 59.126 8.706 59.162 ;
      RECT 8.254 59.126 8.306 59.162 ;
      RECT 7.854 59.126 7.906 59.162 ;
      RECT 7.454 59.126 7.506 59.162 ;
      RECT 7.054 59.126 7.106 59.162 ;
      RECT 6.654 59.126 6.706 59.162 ;
      RECT 6.254 59.126 6.306 59.162 ;
      RECT 5.854 59.126 5.906 59.162 ;
      RECT 5.454 59.126 5.506 59.162 ;
      RECT 5.054 59.126 5.106 59.162 ;
      RECT 4.654 59.126 4.706 59.162 ;
      RECT 4.254 59.126 4.306 59.162 ;
      RECT 3.854 59.126 3.906 59.162 ;
      RECT 3.454 59.126 3.506 59.162 ;
      RECT 3.054 59.126 3.106 59.162 ;
      RECT 2.654 59.126 2.706 59.162 ;
      RECT 2.254 59.126 2.306 59.162 ;
      RECT 1.854 59.126 1.906 59.162 ;
      RECT 1.454 59.126 1.506 59.162 ;
      RECT 1.054 59.126 1.106 59.162 ;
      RECT 0.654 59.126 0.706 59.162 ;
      RECT 21.978 58.902 22.022 58.938 ;
      RECT 21.096 58.902 21.14 58.938 ;
      RECT 14.86 58.902 14.904 58.938 ;
      RECT 13.978 58.902 14.022 58.938 ;
      RECT 35.494 58.678 35.546 58.714 ;
      RECT 35.094 58.678 35.146 58.714 ;
      RECT 34.694 58.678 34.746 58.714 ;
      RECT 34.294 58.678 34.346 58.714 ;
      RECT 33.894 58.678 33.946 58.714 ;
      RECT 33.494 58.678 33.546 58.714 ;
      RECT 33.094 58.678 33.146 58.714 ;
      RECT 32.694 58.678 32.746 58.714 ;
      RECT 32.294 58.678 32.346 58.714 ;
      RECT 31.894 58.678 31.946 58.714 ;
      RECT 31.494 58.678 31.546 58.714 ;
      RECT 31.094 58.678 31.146 58.714 ;
      RECT 30.694 58.678 30.746 58.714 ;
      RECT 30.294 58.678 30.346 58.714 ;
      RECT 29.894 58.678 29.946 58.714 ;
      RECT 29.494 58.678 29.546 58.714 ;
      RECT 29.094 58.678 29.146 58.714 ;
      RECT 28.694 58.678 28.746 58.714 ;
      RECT 28.294 58.678 28.346 58.714 ;
      RECT 27.894 58.678 27.946 58.714 ;
      RECT 27.494 58.678 27.546 58.714 ;
      RECT 27.094 58.678 27.146 58.714 ;
      RECT 26.694 58.678 26.746 58.714 ;
      RECT 26.294 58.678 26.346 58.714 ;
      RECT 25.894 58.678 25.946 58.714 ;
      RECT 25.494 58.678 25.546 58.714 ;
      RECT 25.094 58.678 25.146 58.714 ;
      RECT 24.694 58.678 24.746 58.714 ;
      RECT 24.294 58.678 24.346 58.714 ;
      RECT 23.894 58.678 23.946 58.714 ;
      RECT 23.494 58.678 23.546 58.714 ;
      RECT 23.094 58.678 23.146 58.714 ;
      RECT 21.814 58.678 21.868 58.714 ;
      RECT 19.838 58.678 19.886 58.714 ;
      RECT 19.53 58.678 19.578 58.714 ;
      RECT 16.882 58.678 16.936 58.714 ;
      RECT 16.422 58.678 16.47 58.714 ;
      RECT 16.114 58.678 16.162 58.714 ;
      RECT 14.132 58.678 14.186 58.714 ;
      RECT 13.294 58.678 13.346 58.714 ;
      RECT 12.894 58.678 12.946 58.714 ;
      RECT 12.494 58.678 12.546 58.714 ;
      RECT 12.094 58.678 12.146 58.714 ;
      RECT 11.694 58.678 11.746 58.714 ;
      RECT 11.294 58.678 11.346 58.714 ;
      RECT 10.894 58.678 10.946 58.714 ;
      RECT 10.494 58.678 10.546 58.714 ;
      RECT 10.094 58.678 10.146 58.714 ;
      RECT 9.694 58.678 9.746 58.714 ;
      RECT 9.294 58.678 9.346 58.714 ;
      RECT 8.894 58.678 8.946 58.714 ;
      RECT 8.494 58.678 8.546 58.714 ;
      RECT 8.094 58.678 8.146 58.714 ;
      RECT 7.694 58.678 7.746 58.714 ;
      RECT 7.294 58.678 7.346 58.714 ;
      RECT 6.894 58.678 6.946 58.714 ;
      RECT 6.494 58.678 6.546 58.714 ;
      RECT 6.094 58.678 6.146 58.714 ;
      RECT 5.694 58.678 5.746 58.714 ;
      RECT 5.294 58.678 5.346 58.714 ;
      RECT 4.894 58.678 4.946 58.714 ;
      RECT 4.494 58.678 4.546 58.714 ;
      RECT 4.094 58.678 4.146 58.714 ;
      RECT 3.694 58.678 3.746 58.714 ;
      RECT 3.294 58.678 3.346 58.714 ;
      RECT 2.894 58.678 2.946 58.714 ;
      RECT 2.494 58.678 2.546 58.714 ;
      RECT 2.094 58.678 2.146 58.714 ;
      RECT 1.694 58.678 1.746 58.714 ;
      RECT 1.294 58.678 1.346 58.714 ;
      RECT 0.894 58.678 0.946 58.714 ;
      RECT 21.414 58.602 21.468 58.638 ;
      RECT 14.532 58.602 14.586 58.638 ;
      RECT 19.606 58.449 19.654 58.485 ;
      RECT 18.08 58.449 18.12 58.485 ;
      RECT 16.718 58.449 16.772 58.485 ;
      RECT 16.346 58.449 16.394 58.485 ;
      RECT 20.37 58.4545 20.442 58.4795 ;
      RECT 18.764 58.4545 18.836 58.4795 ;
      RECT 15.558 58.4545 15.63 58.4795 ;
      RECT 21.978 58.302 22.022 58.338 ;
      RECT 13.978 58.302 14.022 58.338 ;
      RECT 18.764 58.3075 18.836 58.3325 ;
      RECT 19.762 58.155 19.81 58.191 ;
      RECT 17.616 58.155 17.656 58.191 ;
      RECT 16.19 58.155 16.238 58.191 ;
      RECT 35.254 57.926 35.306 57.962 ;
      RECT 34.854 57.926 34.906 57.962 ;
      RECT 34.454 57.926 34.506 57.962 ;
      RECT 34.054 57.926 34.106 57.962 ;
      RECT 33.654 57.926 33.706 57.962 ;
      RECT 33.254 57.926 33.306 57.962 ;
      RECT 32.854 57.926 32.906 57.962 ;
      RECT 32.454 57.926 32.506 57.962 ;
      RECT 32.054 57.926 32.106 57.962 ;
      RECT 31.654 57.926 31.706 57.962 ;
      RECT 31.254 57.926 31.306 57.962 ;
      RECT 30.854 57.926 30.906 57.962 ;
      RECT 30.454 57.926 30.506 57.962 ;
      RECT 30.054 57.926 30.106 57.962 ;
      RECT 29.654 57.926 29.706 57.962 ;
      RECT 29.254 57.926 29.306 57.962 ;
      RECT 28.854 57.926 28.906 57.962 ;
      RECT 28.454 57.926 28.506 57.962 ;
      RECT 28.054 57.926 28.106 57.962 ;
      RECT 27.654 57.926 27.706 57.962 ;
      RECT 27.254 57.926 27.306 57.962 ;
      RECT 26.854 57.926 26.906 57.962 ;
      RECT 26.454 57.926 26.506 57.962 ;
      RECT 26.054 57.926 26.106 57.962 ;
      RECT 25.654 57.926 25.706 57.962 ;
      RECT 25.254 57.926 25.306 57.962 ;
      RECT 24.854 57.926 24.906 57.962 ;
      RECT 24.454 57.926 24.506 57.962 ;
      RECT 24.054 57.926 24.106 57.962 ;
      RECT 23.654 57.926 23.706 57.962 ;
      RECT 23.254 57.926 23.306 57.962 ;
      RECT 22.854 57.926 22.906 57.962 ;
      RECT 22.694 57.926 22.746 57.962 ;
      RECT 21.732 57.926 21.786 57.962 ;
      RECT 14.214 57.926 14.268 57.962 ;
      RECT 13.054 57.926 13.106 57.962 ;
      RECT 12.654 57.926 12.706 57.962 ;
      RECT 12.254 57.926 12.306 57.962 ;
      RECT 11.854 57.926 11.906 57.962 ;
      RECT 11.454 57.926 11.506 57.962 ;
      RECT 11.054 57.926 11.106 57.962 ;
      RECT 10.654 57.926 10.706 57.962 ;
      RECT 10.254 57.926 10.306 57.962 ;
      RECT 9.854 57.926 9.906 57.962 ;
      RECT 9.454 57.926 9.506 57.962 ;
      RECT 9.054 57.926 9.106 57.962 ;
      RECT 8.654 57.926 8.706 57.962 ;
      RECT 8.254 57.926 8.306 57.962 ;
      RECT 7.854 57.926 7.906 57.962 ;
      RECT 7.454 57.926 7.506 57.962 ;
      RECT 7.054 57.926 7.106 57.962 ;
      RECT 6.654 57.926 6.706 57.962 ;
      RECT 6.254 57.926 6.306 57.962 ;
      RECT 5.854 57.926 5.906 57.962 ;
      RECT 5.454 57.926 5.506 57.962 ;
      RECT 5.054 57.926 5.106 57.962 ;
      RECT 4.654 57.926 4.706 57.962 ;
      RECT 4.254 57.926 4.306 57.962 ;
      RECT 3.854 57.926 3.906 57.962 ;
      RECT 3.454 57.926 3.506 57.962 ;
      RECT 3.054 57.926 3.106 57.962 ;
      RECT 2.654 57.926 2.706 57.962 ;
      RECT 2.254 57.926 2.306 57.962 ;
      RECT 1.854 57.926 1.906 57.962 ;
      RECT 1.454 57.926 1.506 57.962 ;
      RECT 1.054 57.926 1.106 57.962 ;
      RECT 0.654 57.926 0.706 57.962 ;
      RECT 21.978 57.702 22.022 57.738 ;
      RECT 21.096 57.702 21.14 57.738 ;
      RECT 14.86 57.702 14.904 57.738 ;
      RECT 13.978 57.702 14.022 57.738 ;
      RECT 35.494 57.478 35.546 57.514 ;
      RECT 35.094 57.478 35.146 57.514 ;
      RECT 34.694 57.478 34.746 57.514 ;
      RECT 34.294 57.478 34.346 57.514 ;
      RECT 33.894 57.478 33.946 57.514 ;
      RECT 33.494 57.478 33.546 57.514 ;
      RECT 33.094 57.478 33.146 57.514 ;
      RECT 32.694 57.478 32.746 57.514 ;
      RECT 32.294 57.478 32.346 57.514 ;
      RECT 31.894 57.478 31.946 57.514 ;
      RECT 31.494 57.478 31.546 57.514 ;
      RECT 31.094 57.478 31.146 57.514 ;
      RECT 30.694 57.478 30.746 57.514 ;
      RECT 30.294 57.478 30.346 57.514 ;
      RECT 29.894 57.478 29.946 57.514 ;
      RECT 29.494 57.478 29.546 57.514 ;
      RECT 29.094 57.478 29.146 57.514 ;
      RECT 28.694 57.478 28.746 57.514 ;
      RECT 28.294 57.478 28.346 57.514 ;
      RECT 27.894 57.478 27.946 57.514 ;
      RECT 27.494 57.478 27.546 57.514 ;
      RECT 27.094 57.478 27.146 57.514 ;
      RECT 26.694 57.478 26.746 57.514 ;
      RECT 26.294 57.478 26.346 57.514 ;
      RECT 25.894 57.478 25.946 57.514 ;
      RECT 25.494 57.478 25.546 57.514 ;
      RECT 25.094 57.478 25.146 57.514 ;
      RECT 24.694 57.478 24.746 57.514 ;
      RECT 24.294 57.478 24.346 57.514 ;
      RECT 23.894 57.478 23.946 57.514 ;
      RECT 23.494 57.478 23.546 57.514 ;
      RECT 23.094 57.478 23.146 57.514 ;
      RECT 21.814 57.478 21.868 57.514 ;
      RECT 19.838 57.478 19.886 57.514 ;
      RECT 19.53 57.478 19.578 57.514 ;
      RECT 16.882 57.478 16.936 57.514 ;
      RECT 16.422 57.478 16.47 57.514 ;
      RECT 16.114 57.478 16.162 57.514 ;
      RECT 14.132 57.478 14.186 57.514 ;
      RECT 13.294 57.478 13.346 57.514 ;
      RECT 12.894 57.478 12.946 57.514 ;
      RECT 12.494 57.478 12.546 57.514 ;
      RECT 12.094 57.478 12.146 57.514 ;
      RECT 11.694 57.478 11.746 57.514 ;
      RECT 11.294 57.478 11.346 57.514 ;
      RECT 10.894 57.478 10.946 57.514 ;
      RECT 10.494 57.478 10.546 57.514 ;
      RECT 10.094 57.478 10.146 57.514 ;
      RECT 9.694 57.478 9.746 57.514 ;
      RECT 9.294 57.478 9.346 57.514 ;
      RECT 8.894 57.478 8.946 57.514 ;
      RECT 8.494 57.478 8.546 57.514 ;
      RECT 8.094 57.478 8.146 57.514 ;
      RECT 7.694 57.478 7.746 57.514 ;
      RECT 7.294 57.478 7.346 57.514 ;
      RECT 6.894 57.478 6.946 57.514 ;
      RECT 6.494 57.478 6.546 57.514 ;
      RECT 6.094 57.478 6.146 57.514 ;
      RECT 5.694 57.478 5.746 57.514 ;
      RECT 5.294 57.478 5.346 57.514 ;
      RECT 4.894 57.478 4.946 57.514 ;
      RECT 4.494 57.478 4.546 57.514 ;
      RECT 4.094 57.478 4.146 57.514 ;
      RECT 3.694 57.478 3.746 57.514 ;
      RECT 3.294 57.478 3.346 57.514 ;
      RECT 2.894 57.478 2.946 57.514 ;
      RECT 2.494 57.478 2.546 57.514 ;
      RECT 2.094 57.478 2.146 57.514 ;
      RECT 1.694 57.478 1.746 57.514 ;
      RECT 1.294 57.478 1.346 57.514 ;
      RECT 0.894 57.478 0.946 57.514 ;
      RECT 21.414 57.402 21.468 57.438 ;
      RECT 14.532 57.402 14.586 57.438 ;
      RECT 19.606 57.249 19.654 57.285 ;
      RECT 18.08 57.249 18.12 57.285 ;
      RECT 16.718 57.249 16.772 57.285 ;
      RECT 16.346 57.249 16.394 57.285 ;
      RECT 20.37 57.2545 20.442 57.2795 ;
      RECT 18.764 57.2545 18.836 57.2795 ;
      RECT 15.558 57.2545 15.63 57.2795 ;
      RECT 21.978 57.102 22.022 57.138 ;
      RECT 13.978 57.102 14.022 57.138 ;
      RECT 18.764 57.1075 18.836 57.1325 ;
      RECT 19.762 56.955 19.81 56.991 ;
      RECT 17.616 56.955 17.656 56.991 ;
      RECT 16.19 56.955 16.238 56.991 ;
      RECT 35.254 56.726 35.306 56.762 ;
      RECT 34.854 56.726 34.906 56.762 ;
      RECT 34.454 56.726 34.506 56.762 ;
      RECT 34.054 56.726 34.106 56.762 ;
      RECT 33.654 56.726 33.706 56.762 ;
      RECT 33.254 56.726 33.306 56.762 ;
      RECT 32.854 56.726 32.906 56.762 ;
      RECT 32.454 56.726 32.506 56.762 ;
      RECT 32.054 56.726 32.106 56.762 ;
      RECT 31.654 56.726 31.706 56.762 ;
      RECT 31.254 56.726 31.306 56.762 ;
      RECT 30.854 56.726 30.906 56.762 ;
      RECT 30.454 56.726 30.506 56.762 ;
      RECT 30.054 56.726 30.106 56.762 ;
      RECT 29.654 56.726 29.706 56.762 ;
      RECT 29.254 56.726 29.306 56.762 ;
      RECT 28.854 56.726 28.906 56.762 ;
      RECT 28.454 56.726 28.506 56.762 ;
      RECT 28.054 56.726 28.106 56.762 ;
      RECT 27.654 56.726 27.706 56.762 ;
      RECT 27.254 56.726 27.306 56.762 ;
      RECT 26.854 56.726 26.906 56.762 ;
      RECT 26.454 56.726 26.506 56.762 ;
      RECT 26.054 56.726 26.106 56.762 ;
      RECT 25.654 56.726 25.706 56.762 ;
      RECT 25.254 56.726 25.306 56.762 ;
      RECT 24.854 56.726 24.906 56.762 ;
      RECT 24.454 56.726 24.506 56.762 ;
      RECT 24.054 56.726 24.106 56.762 ;
      RECT 23.654 56.726 23.706 56.762 ;
      RECT 23.254 56.726 23.306 56.762 ;
      RECT 22.854 56.726 22.906 56.762 ;
      RECT 22.694 56.726 22.746 56.762 ;
      RECT 21.732 56.726 21.786 56.762 ;
      RECT 14.214 56.726 14.268 56.762 ;
      RECT 13.054 56.726 13.106 56.762 ;
      RECT 12.654 56.726 12.706 56.762 ;
      RECT 12.254 56.726 12.306 56.762 ;
      RECT 11.854 56.726 11.906 56.762 ;
      RECT 11.454 56.726 11.506 56.762 ;
      RECT 11.054 56.726 11.106 56.762 ;
      RECT 10.654 56.726 10.706 56.762 ;
      RECT 10.254 56.726 10.306 56.762 ;
      RECT 9.854 56.726 9.906 56.762 ;
      RECT 9.454 56.726 9.506 56.762 ;
      RECT 9.054 56.726 9.106 56.762 ;
      RECT 8.654 56.726 8.706 56.762 ;
      RECT 8.254 56.726 8.306 56.762 ;
      RECT 7.854 56.726 7.906 56.762 ;
      RECT 7.454 56.726 7.506 56.762 ;
      RECT 7.054 56.726 7.106 56.762 ;
      RECT 6.654 56.726 6.706 56.762 ;
      RECT 6.254 56.726 6.306 56.762 ;
      RECT 5.854 56.726 5.906 56.762 ;
      RECT 5.454 56.726 5.506 56.762 ;
      RECT 5.054 56.726 5.106 56.762 ;
      RECT 4.654 56.726 4.706 56.762 ;
      RECT 4.254 56.726 4.306 56.762 ;
      RECT 3.854 56.726 3.906 56.762 ;
      RECT 3.454 56.726 3.506 56.762 ;
      RECT 3.054 56.726 3.106 56.762 ;
      RECT 2.654 56.726 2.706 56.762 ;
      RECT 2.254 56.726 2.306 56.762 ;
      RECT 1.854 56.726 1.906 56.762 ;
      RECT 1.454 56.726 1.506 56.762 ;
      RECT 1.054 56.726 1.106 56.762 ;
      RECT 0.654 56.726 0.706 56.762 ;
      RECT 21.978 56.502 22.022 56.538 ;
      RECT 21.096 56.502 21.14 56.538 ;
      RECT 14.86 56.502 14.904 56.538 ;
      RECT 13.978 56.502 14.022 56.538 ;
      RECT 35.494 56.278 35.546 56.314 ;
      RECT 35.094 56.278 35.146 56.314 ;
      RECT 34.694 56.278 34.746 56.314 ;
      RECT 34.294 56.278 34.346 56.314 ;
      RECT 33.894 56.278 33.946 56.314 ;
      RECT 33.494 56.278 33.546 56.314 ;
      RECT 33.094 56.278 33.146 56.314 ;
      RECT 32.694 56.278 32.746 56.314 ;
      RECT 32.294 56.278 32.346 56.314 ;
      RECT 31.894 56.278 31.946 56.314 ;
      RECT 31.494 56.278 31.546 56.314 ;
      RECT 31.094 56.278 31.146 56.314 ;
      RECT 30.694 56.278 30.746 56.314 ;
      RECT 30.294 56.278 30.346 56.314 ;
      RECT 29.894 56.278 29.946 56.314 ;
      RECT 29.494 56.278 29.546 56.314 ;
      RECT 29.094 56.278 29.146 56.314 ;
      RECT 28.694 56.278 28.746 56.314 ;
      RECT 28.294 56.278 28.346 56.314 ;
      RECT 27.894 56.278 27.946 56.314 ;
      RECT 27.494 56.278 27.546 56.314 ;
      RECT 27.094 56.278 27.146 56.314 ;
      RECT 26.694 56.278 26.746 56.314 ;
      RECT 26.294 56.278 26.346 56.314 ;
      RECT 25.894 56.278 25.946 56.314 ;
      RECT 25.494 56.278 25.546 56.314 ;
      RECT 25.094 56.278 25.146 56.314 ;
      RECT 24.694 56.278 24.746 56.314 ;
      RECT 24.294 56.278 24.346 56.314 ;
      RECT 23.894 56.278 23.946 56.314 ;
      RECT 23.494 56.278 23.546 56.314 ;
      RECT 23.094 56.278 23.146 56.314 ;
      RECT 21.814 56.278 21.868 56.314 ;
      RECT 19.838 56.278 19.886 56.314 ;
      RECT 19.53 56.278 19.578 56.314 ;
      RECT 16.882 56.278 16.936 56.314 ;
      RECT 16.422 56.278 16.47 56.314 ;
      RECT 16.114 56.278 16.162 56.314 ;
      RECT 14.132 56.278 14.186 56.314 ;
      RECT 13.294 56.278 13.346 56.314 ;
      RECT 12.894 56.278 12.946 56.314 ;
      RECT 12.494 56.278 12.546 56.314 ;
      RECT 12.094 56.278 12.146 56.314 ;
      RECT 11.694 56.278 11.746 56.314 ;
      RECT 11.294 56.278 11.346 56.314 ;
      RECT 10.894 56.278 10.946 56.314 ;
      RECT 10.494 56.278 10.546 56.314 ;
      RECT 10.094 56.278 10.146 56.314 ;
      RECT 9.694 56.278 9.746 56.314 ;
      RECT 9.294 56.278 9.346 56.314 ;
      RECT 8.894 56.278 8.946 56.314 ;
      RECT 8.494 56.278 8.546 56.314 ;
      RECT 8.094 56.278 8.146 56.314 ;
      RECT 7.694 56.278 7.746 56.314 ;
      RECT 7.294 56.278 7.346 56.314 ;
      RECT 6.894 56.278 6.946 56.314 ;
      RECT 6.494 56.278 6.546 56.314 ;
      RECT 6.094 56.278 6.146 56.314 ;
      RECT 5.694 56.278 5.746 56.314 ;
      RECT 5.294 56.278 5.346 56.314 ;
      RECT 4.894 56.278 4.946 56.314 ;
      RECT 4.494 56.278 4.546 56.314 ;
      RECT 4.094 56.278 4.146 56.314 ;
      RECT 3.694 56.278 3.746 56.314 ;
      RECT 3.294 56.278 3.346 56.314 ;
      RECT 2.894 56.278 2.946 56.314 ;
      RECT 2.494 56.278 2.546 56.314 ;
      RECT 2.094 56.278 2.146 56.314 ;
      RECT 1.694 56.278 1.746 56.314 ;
      RECT 1.294 56.278 1.346 56.314 ;
      RECT 0.894 56.278 0.946 56.314 ;
      RECT 21.414 56.202 21.468 56.238 ;
      RECT 14.532 56.202 14.586 56.238 ;
      RECT 19.606 56.049 19.654 56.085 ;
      RECT 18.08 56.049 18.12 56.085 ;
      RECT 16.718 56.049 16.772 56.085 ;
      RECT 16.346 56.049 16.394 56.085 ;
      RECT 20.37 56.0545 20.442 56.0795 ;
      RECT 18.764 56.0545 18.836 56.0795 ;
      RECT 15.558 56.0545 15.63 56.0795 ;
      RECT 21.978 55.902 22.022 55.938 ;
      RECT 13.978 55.902 14.022 55.938 ;
      RECT 18.764 55.9075 18.836 55.9325 ;
      RECT 19.762 55.755 19.81 55.791 ;
      RECT 17.616 55.755 17.656 55.791 ;
      RECT 16.19 55.755 16.238 55.791 ;
      RECT 35.254 55.526 35.306 55.562 ;
      RECT 34.854 55.526 34.906 55.562 ;
      RECT 34.454 55.526 34.506 55.562 ;
      RECT 34.054 55.526 34.106 55.562 ;
      RECT 33.654 55.526 33.706 55.562 ;
      RECT 33.254 55.526 33.306 55.562 ;
      RECT 32.854 55.526 32.906 55.562 ;
      RECT 32.454 55.526 32.506 55.562 ;
      RECT 32.054 55.526 32.106 55.562 ;
      RECT 31.654 55.526 31.706 55.562 ;
      RECT 31.254 55.526 31.306 55.562 ;
      RECT 30.854 55.526 30.906 55.562 ;
      RECT 30.454 55.526 30.506 55.562 ;
      RECT 30.054 55.526 30.106 55.562 ;
      RECT 29.654 55.526 29.706 55.562 ;
      RECT 29.254 55.526 29.306 55.562 ;
      RECT 28.854 55.526 28.906 55.562 ;
      RECT 28.454 55.526 28.506 55.562 ;
      RECT 28.054 55.526 28.106 55.562 ;
      RECT 27.654 55.526 27.706 55.562 ;
      RECT 27.254 55.526 27.306 55.562 ;
      RECT 26.854 55.526 26.906 55.562 ;
      RECT 26.454 55.526 26.506 55.562 ;
      RECT 26.054 55.526 26.106 55.562 ;
      RECT 25.654 55.526 25.706 55.562 ;
      RECT 25.254 55.526 25.306 55.562 ;
      RECT 24.854 55.526 24.906 55.562 ;
      RECT 24.454 55.526 24.506 55.562 ;
      RECT 24.054 55.526 24.106 55.562 ;
      RECT 23.654 55.526 23.706 55.562 ;
      RECT 23.254 55.526 23.306 55.562 ;
      RECT 22.854 55.526 22.906 55.562 ;
      RECT 22.694 55.526 22.746 55.562 ;
      RECT 21.732 55.526 21.786 55.562 ;
      RECT 14.214 55.526 14.268 55.562 ;
      RECT 13.054 55.526 13.106 55.562 ;
      RECT 12.654 55.526 12.706 55.562 ;
      RECT 12.254 55.526 12.306 55.562 ;
      RECT 11.854 55.526 11.906 55.562 ;
      RECT 11.454 55.526 11.506 55.562 ;
      RECT 11.054 55.526 11.106 55.562 ;
      RECT 10.654 55.526 10.706 55.562 ;
      RECT 10.254 55.526 10.306 55.562 ;
      RECT 9.854 55.526 9.906 55.562 ;
      RECT 9.454 55.526 9.506 55.562 ;
      RECT 9.054 55.526 9.106 55.562 ;
      RECT 8.654 55.526 8.706 55.562 ;
      RECT 8.254 55.526 8.306 55.562 ;
      RECT 7.854 55.526 7.906 55.562 ;
      RECT 7.454 55.526 7.506 55.562 ;
      RECT 7.054 55.526 7.106 55.562 ;
      RECT 6.654 55.526 6.706 55.562 ;
      RECT 6.254 55.526 6.306 55.562 ;
      RECT 5.854 55.526 5.906 55.562 ;
      RECT 5.454 55.526 5.506 55.562 ;
      RECT 5.054 55.526 5.106 55.562 ;
      RECT 4.654 55.526 4.706 55.562 ;
      RECT 4.254 55.526 4.306 55.562 ;
      RECT 3.854 55.526 3.906 55.562 ;
      RECT 3.454 55.526 3.506 55.562 ;
      RECT 3.054 55.526 3.106 55.562 ;
      RECT 2.654 55.526 2.706 55.562 ;
      RECT 2.254 55.526 2.306 55.562 ;
      RECT 1.854 55.526 1.906 55.562 ;
      RECT 1.454 55.526 1.506 55.562 ;
      RECT 1.054 55.526 1.106 55.562 ;
      RECT 0.654 55.526 0.706 55.562 ;
      RECT 21.978 55.302 22.022 55.338 ;
      RECT 21.096 55.302 21.14 55.338 ;
      RECT 14.86 55.302 14.904 55.338 ;
      RECT 13.978 55.302 14.022 55.338 ;
      RECT 35.494 55.078 35.546 55.114 ;
      RECT 35.094 55.078 35.146 55.114 ;
      RECT 34.694 55.078 34.746 55.114 ;
      RECT 34.294 55.078 34.346 55.114 ;
      RECT 33.894 55.078 33.946 55.114 ;
      RECT 33.494 55.078 33.546 55.114 ;
      RECT 33.094 55.078 33.146 55.114 ;
      RECT 32.694 55.078 32.746 55.114 ;
      RECT 32.294 55.078 32.346 55.114 ;
      RECT 31.894 55.078 31.946 55.114 ;
      RECT 31.494 55.078 31.546 55.114 ;
      RECT 31.094 55.078 31.146 55.114 ;
      RECT 30.694 55.078 30.746 55.114 ;
      RECT 30.294 55.078 30.346 55.114 ;
      RECT 29.894 55.078 29.946 55.114 ;
      RECT 29.494 55.078 29.546 55.114 ;
      RECT 29.094 55.078 29.146 55.114 ;
      RECT 28.694 55.078 28.746 55.114 ;
      RECT 28.294 55.078 28.346 55.114 ;
      RECT 27.894 55.078 27.946 55.114 ;
      RECT 27.494 55.078 27.546 55.114 ;
      RECT 27.094 55.078 27.146 55.114 ;
      RECT 26.694 55.078 26.746 55.114 ;
      RECT 26.294 55.078 26.346 55.114 ;
      RECT 25.894 55.078 25.946 55.114 ;
      RECT 25.494 55.078 25.546 55.114 ;
      RECT 25.094 55.078 25.146 55.114 ;
      RECT 24.694 55.078 24.746 55.114 ;
      RECT 24.294 55.078 24.346 55.114 ;
      RECT 23.894 55.078 23.946 55.114 ;
      RECT 23.494 55.078 23.546 55.114 ;
      RECT 23.094 55.078 23.146 55.114 ;
      RECT 21.814 55.078 21.868 55.114 ;
      RECT 19.838 55.078 19.886 55.114 ;
      RECT 19.53 55.078 19.578 55.114 ;
      RECT 16.882 55.078 16.936 55.114 ;
      RECT 16.422 55.078 16.47 55.114 ;
      RECT 16.114 55.078 16.162 55.114 ;
      RECT 14.132 55.078 14.186 55.114 ;
      RECT 13.294 55.078 13.346 55.114 ;
      RECT 12.894 55.078 12.946 55.114 ;
      RECT 12.494 55.078 12.546 55.114 ;
      RECT 12.094 55.078 12.146 55.114 ;
      RECT 11.694 55.078 11.746 55.114 ;
      RECT 11.294 55.078 11.346 55.114 ;
      RECT 10.894 55.078 10.946 55.114 ;
      RECT 10.494 55.078 10.546 55.114 ;
      RECT 10.094 55.078 10.146 55.114 ;
      RECT 9.694 55.078 9.746 55.114 ;
      RECT 9.294 55.078 9.346 55.114 ;
      RECT 8.894 55.078 8.946 55.114 ;
      RECT 8.494 55.078 8.546 55.114 ;
      RECT 8.094 55.078 8.146 55.114 ;
      RECT 7.694 55.078 7.746 55.114 ;
      RECT 7.294 55.078 7.346 55.114 ;
      RECT 6.894 55.078 6.946 55.114 ;
      RECT 6.494 55.078 6.546 55.114 ;
      RECT 6.094 55.078 6.146 55.114 ;
      RECT 5.694 55.078 5.746 55.114 ;
      RECT 5.294 55.078 5.346 55.114 ;
      RECT 4.894 55.078 4.946 55.114 ;
      RECT 4.494 55.078 4.546 55.114 ;
      RECT 4.094 55.078 4.146 55.114 ;
      RECT 3.694 55.078 3.746 55.114 ;
      RECT 3.294 55.078 3.346 55.114 ;
      RECT 2.894 55.078 2.946 55.114 ;
      RECT 2.494 55.078 2.546 55.114 ;
      RECT 2.094 55.078 2.146 55.114 ;
      RECT 1.694 55.078 1.746 55.114 ;
      RECT 1.294 55.078 1.346 55.114 ;
      RECT 0.894 55.078 0.946 55.114 ;
      RECT 21.414 55.002 21.468 55.038 ;
      RECT 14.532 55.002 14.586 55.038 ;
      RECT 19.606 54.849 19.654 54.885 ;
      RECT 18.08 54.849 18.12 54.885 ;
      RECT 16.718 54.849 16.772 54.885 ;
      RECT 16.346 54.849 16.394 54.885 ;
      RECT 20.37 54.8545 20.442 54.8795 ;
      RECT 18.764 54.8545 18.836 54.8795 ;
      RECT 15.558 54.8545 15.63 54.8795 ;
      RECT 21.978 54.702 22.022 54.738 ;
      RECT 13.978 54.702 14.022 54.738 ;
      RECT 18.764 54.7075 18.836 54.7325 ;
      RECT 19.762 54.555 19.81 54.591 ;
      RECT 17.616 54.555 17.656 54.591 ;
      RECT 16.19 54.555 16.238 54.591 ;
      RECT 35.254 54.326 35.306 54.362 ;
      RECT 34.854 54.326 34.906 54.362 ;
      RECT 34.454 54.326 34.506 54.362 ;
      RECT 34.054 54.326 34.106 54.362 ;
      RECT 33.654 54.326 33.706 54.362 ;
      RECT 33.254 54.326 33.306 54.362 ;
      RECT 32.854 54.326 32.906 54.362 ;
      RECT 32.454 54.326 32.506 54.362 ;
      RECT 32.054 54.326 32.106 54.362 ;
      RECT 31.654 54.326 31.706 54.362 ;
      RECT 31.254 54.326 31.306 54.362 ;
      RECT 30.854 54.326 30.906 54.362 ;
      RECT 30.454 54.326 30.506 54.362 ;
      RECT 30.054 54.326 30.106 54.362 ;
      RECT 29.654 54.326 29.706 54.362 ;
      RECT 29.254 54.326 29.306 54.362 ;
      RECT 28.854 54.326 28.906 54.362 ;
      RECT 28.454 54.326 28.506 54.362 ;
      RECT 28.054 54.326 28.106 54.362 ;
      RECT 27.654 54.326 27.706 54.362 ;
      RECT 27.254 54.326 27.306 54.362 ;
      RECT 26.854 54.326 26.906 54.362 ;
      RECT 26.454 54.326 26.506 54.362 ;
      RECT 26.054 54.326 26.106 54.362 ;
      RECT 25.654 54.326 25.706 54.362 ;
      RECT 25.254 54.326 25.306 54.362 ;
      RECT 24.854 54.326 24.906 54.362 ;
      RECT 24.454 54.326 24.506 54.362 ;
      RECT 24.054 54.326 24.106 54.362 ;
      RECT 23.654 54.326 23.706 54.362 ;
      RECT 23.254 54.326 23.306 54.362 ;
      RECT 22.854 54.326 22.906 54.362 ;
      RECT 22.694 54.326 22.746 54.362 ;
      RECT 21.732 54.326 21.786 54.362 ;
      RECT 14.214 54.326 14.268 54.362 ;
      RECT 13.054 54.326 13.106 54.362 ;
      RECT 12.654 54.326 12.706 54.362 ;
      RECT 12.254 54.326 12.306 54.362 ;
      RECT 11.854 54.326 11.906 54.362 ;
      RECT 11.454 54.326 11.506 54.362 ;
      RECT 11.054 54.326 11.106 54.362 ;
      RECT 10.654 54.326 10.706 54.362 ;
      RECT 10.254 54.326 10.306 54.362 ;
      RECT 9.854 54.326 9.906 54.362 ;
      RECT 9.454 54.326 9.506 54.362 ;
      RECT 9.054 54.326 9.106 54.362 ;
      RECT 8.654 54.326 8.706 54.362 ;
      RECT 8.254 54.326 8.306 54.362 ;
      RECT 7.854 54.326 7.906 54.362 ;
      RECT 7.454 54.326 7.506 54.362 ;
      RECT 7.054 54.326 7.106 54.362 ;
      RECT 6.654 54.326 6.706 54.362 ;
      RECT 6.254 54.326 6.306 54.362 ;
      RECT 5.854 54.326 5.906 54.362 ;
      RECT 5.454 54.326 5.506 54.362 ;
      RECT 5.054 54.326 5.106 54.362 ;
      RECT 4.654 54.326 4.706 54.362 ;
      RECT 4.254 54.326 4.306 54.362 ;
      RECT 3.854 54.326 3.906 54.362 ;
      RECT 3.454 54.326 3.506 54.362 ;
      RECT 3.054 54.326 3.106 54.362 ;
      RECT 2.654 54.326 2.706 54.362 ;
      RECT 2.254 54.326 2.306 54.362 ;
      RECT 1.854 54.326 1.906 54.362 ;
      RECT 1.454 54.326 1.506 54.362 ;
      RECT 1.054 54.326 1.106 54.362 ;
      RECT 0.654 54.326 0.706 54.362 ;
      RECT 21.978 54.102 22.022 54.138 ;
      RECT 21.096 54.102 21.14 54.138 ;
      RECT 14.86 54.102 14.904 54.138 ;
      RECT 13.978 54.102 14.022 54.138 ;
      RECT 35.494 53.878 35.546 53.914 ;
      RECT 35.094 53.878 35.146 53.914 ;
      RECT 34.694 53.878 34.746 53.914 ;
      RECT 34.294 53.878 34.346 53.914 ;
      RECT 33.894 53.878 33.946 53.914 ;
      RECT 33.494 53.878 33.546 53.914 ;
      RECT 33.094 53.878 33.146 53.914 ;
      RECT 32.694 53.878 32.746 53.914 ;
      RECT 32.294 53.878 32.346 53.914 ;
      RECT 31.894 53.878 31.946 53.914 ;
      RECT 31.494 53.878 31.546 53.914 ;
      RECT 31.094 53.878 31.146 53.914 ;
      RECT 30.694 53.878 30.746 53.914 ;
      RECT 30.294 53.878 30.346 53.914 ;
      RECT 29.894 53.878 29.946 53.914 ;
      RECT 29.494 53.878 29.546 53.914 ;
      RECT 29.094 53.878 29.146 53.914 ;
      RECT 28.694 53.878 28.746 53.914 ;
      RECT 28.294 53.878 28.346 53.914 ;
      RECT 27.894 53.878 27.946 53.914 ;
      RECT 27.494 53.878 27.546 53.914 ;
      RECT 27.094 53.878 27.146 53.914 ;
      RECT 26.694 53.878 26.746 53.914 ;
      RECT 26.294 53.878 26.346 53.914 ;
      RECT 25.894 53.878 25.946 53.914 ;
      RECT 25.494 53.878 25.546 53.914 ;
      RECT 25.094 53.878 25.146 53.914 ;
      RECT 24.694 53.878 24.746 53.914 ;
      RECT 24.294 53.878 24.346 53.914 ;
      RECT 23.894 53.878 23.946 53.914 ;
      RECT 23.494 53.878 23.546 53.914 ;
      RECT 23.094 53.878 23.146 53.914 ;
      RECT 21.814 53.878 21.868 53.914 ;
      RECT 19.838 53.878 19.886 53.914 ;
      RECT 19.53 53.878 19.578 53.914 ;
      RECT 16.882 53.878 16.936 53.914 ;
      RECT 16.422 53.878 16.47 53.914 ;
      RECT 16.114 53.878 16.162 53.914 ;
      RECT 14.132 53.878 14.186 53.914 ;
      RECT 13.294 53.878 13.346 53.914 ;
      RECT 12.894 53.878 12.946 53.914 ;
      RECT 12.494 53.878 12.546 53.914 ;
      RECT 12.094 53.878 12.146 53.914 ;
      RECT 11.694 53.878 11.746 53.914 ;
      RECT 11.294 53.878 11.346 53.914 ;
      RECT 10.894 53.878 10.946 53.914 ;
      RECT 10.494 53.878 10.546 53.914 ;
      RECT 10.094 53.878 10.146 53.914 ;
      RECT 9.694 53.878 9.746 53.914 ;
      RECT 9.294 53.878 9.346 53.914 ;
      RECT 8.894 53.878 8.946 53.914 ;
      RECT 8.494 53.878 8.546 53.914 ;
      RECT 8.094 53.878 8.146 53.914 ;
      RECT 7.694 53.878 7.746 53.914 ;
      RECT 7.294 53.878 7.346 53.914 ;
      RECT 6.894 53.878 6.946 53.914 ;
      RECT 6.494 53.878 6.546 53.914 ;
      RECT 6.094 53.878 6.146 53.914 ;
      RECT 5.694 53.878 5.746 53.914 ;
      RECT 5.294 53.878 5.346 53.914 ;
      RECT 4.894 53.878 4.946 53.914 ;
      RECT 4.494 53.878 4.546 53.914 ;
      RECT 4.094 53.878 4.146 53.914 ;
      RECT 3.694 53.878 3.746 53.914 ;
      RECT 3.294 53.878 3.346 53.914 ;
      RECT 2.894 53.878 2.946 53.914 ;
      RECT 2.494 53.878 2.546 53.914 ;
      RECT 2.094 53.878 2.146 53.914 ;
      RECT 1.694 53.878 1.746 53.914 ;
      RECT 1.294 53.878 1.346 53.914 ;
      RECT 0.894 53.878 0.946 53.914 ;
      RECT 21.414 53.802 21.468 53.838 ;
      RECT 14.532 53.802 14.586 53.838 ;
      RECT 19.606 53.649 19.654 53.685 ;
      RECT 18.08 53.649 18.12 53.685 ;
      RECT 16.718 53.649 16.772 53.685 ;
      RECT 16.346 53.649 16.394 53.685 ;
      RECT 20.37 53.6545 20.442 53.6795 ;
      RECT 18.764 53.6545 18.836 53.6795 ;
      RECT 15.558 53.6545 15.63 53.6795 ;
      RECT 21.978 53.502 22.022 53.538 ;
      RECT 13.978 53.502 14.022 53.538 ;
      RECT 18.764 53.5075 18.836 53.5325 ;
      RECT 19.762 53.355 19.81 53.391 ;
      RECT 17.616 53.355 17.656 53.391 ;
      RECT 16.19 53.355 16.238 53.391 ;
      RECT 35.254 53.126 35.306 53.162 ;
      RECT 34.854 53.126 34.906 53.162 ;
      RECT 34.454 53.126 34.506 53.162 ;
      RECT 34.054 53.126 34.106 53.162 ;
      RECT 33.654 53.126 33.706 53.162 ;
      RECT 33.254 53.126 33.306 53.162 ;
      RECT 32.854 53.126 32.906 53.162 ;
      RECT 32.454 53.126 32.506 53.162 ;
      RECT 32.054 53.126 32.106 53.162 ;
      RECT 31.654 53.126 31.706 53.162 ;
      RECT 31.254 53.126 31.306 53.162 ;
      RECT 30.854 53.126 30.906 53.162 ;
      RECT 30.454 53.126 30.506 53.162 ;
      RECT 30.054 53.126 30.106 53.162 ;
      RECT 29.654 53.126 29.706 53.162 ;
      RECT 29.254 53.126 29.306 53.162 ;
      RECT 28.854 53.126 28.906 53.162 ;
      RECT 28.454 53.126 28.506 53.162 ;
      RECT 28.054 53.126 28.106 53.162 ;
      RECT 27.654 53.126 27.706 53.162 ;
      RECT 27.254 53.126 27.306 53.162 ;
      RECT 26.854 53.126 26.906 53.162 ;
      RECT 26.454 53.126 26.506 53.162 ;
      RECT 26.054 53.126 26.106 53.162 ;
      RECT 25.654 53.126 25.706 53.162 ;
      RECT 25.254 53.126 25.306 53.162 ;
      RECT 24.854 53.126 24.906 53.162 ;
      RECT 24.454 53.126 24.506 53.162 ;
      RECT 24.054 53.126 24.106 53.162 ;
      RECT 23.654 53.126 23.706 53.162 ;
      RECT 23.254 53.126 23.306 53.162 ;
      RECT 22.854 53.126 22.906 53.162 ;
      RECT 22.694 53.126 22.746 53.162 ;
      RECT 21.732 53.126 21.786 53.162 ;
      RECT 14.214 53.126 14.268 53.162 ;
      RECT 13.054 53.126 13.106 53.162 ;
      RECT 12.654 53.126 12.706 53.162 ;
      RECT 12.254 53.126 12.306 53.162 ;
      RECT 11.854 53.126 11.906 53.162 ;
      RECT 11.454 53.126 11.506 53.162 ;
      RECT 11.054 53.126 11.106 53.162 ;
      RECT 10.654 53.126 10.706 53.162 ;
      RECT 10.254 53.126 10.306 53.162 ;
      RECT 9.854 53.126 9.906 53.162 ;
      RECT 9.454 53.126 9.506 53.162 ;
      RECT 9.054 53.126 9.106 53.162 ;
      RECT 8.654 53.126 8.706 53.162 ;
      RECT 8.254 53.126 8.306 53.162 ;
      RECT 7.854 53.126 7.906 53.162 ;
      RECT 7.454 53.126 7.506 53.162 ;
      RECT 7.054 53.126 7.106 53.162 ;
      RECT 6.654 53.126 6.706 53.162 ;
      RECT 6.254 53.126 6.306 53.162 ;
      RECT 5.854 53.126 5.906 53.162 ;
      RECT 5.454 53.126 5.506 53.162 ;
      RECT 5.054 53.126 5.106 53.162 ;
      RECT 4.654 53.126 4.706 53.162 ;
      RECT 4.254 53.126 4.306 53.162 ;
      RECT 3.854 53.126 3.906 53.162 ;
      RECT 3.454 53.126 3.506 53.162 ;
      RECT 3.054 53.126 3.106 53.162 ;
      RECT 2.654 53.126 2.706 53.162 ;
      RECT 2.254 53.126 2.306 53.162 ;
      RECT 1.854 53.126 1.906 53.162 ;
      RECT 1.454 53.126 1.506 53.162 ;
      RECT 1.054 53.126 1.106 53.162 ;
      RECT 0.654 53.126 0.706 53.162 ;
      RECT 21.978 52.902 22.022 52.938 ;
      RECT 21.096 52.902 21.14 52.938 ;
      RECT 14.86 52.902 14.904 52.938 ;
      RECT 13.978 52.902 14.022 52.938 ;
      RECT 35.494 52.678 35.546 52.714 ;
      RECT 35.094 52.678 35.146 52.714 ;
      RECT 34.694 52.678 34.746 52.714 ;
      RECT 34.294 52.678 34.346 52.714 ;
      RECT 33.894 52.678 33.946 52.714 ;
      RECT 33.494 52.678 33.546 52.714 ;
      RECT 33.094 52.678 33.146 52.714 ;
      RECT 32.694 52.678 32.746 52.714 ;
      RECT 32.294 52.678 32.346 52.714 ;
      RECT 31.894 52.678 31.946 52.714 ;
      RECT 31.494 52.678 31.546 52.714 ;
      RECT 31.094 52.678 31.146 52.714 ;
      RECT 30.694 52.678 30.746 52.714 ;
      RECT 30.294 52.678 30.346 52.714 ;
      RECT 29.894 52.678 29.946 52.714 ;
      RECT 29.494 52.678 29.546 52.714 ;
      RECT 29.094 52.678 29.146 52.714 ;
      RECT 28.694 52.678 28.746 52.714 ;
      RECT 28.294 52.678 28.346 52.714 ;
      RECT 27.894 52.678 27.946 52.714 ;
      RECT 27.494 52.678 27.546 52.714 ;
      RECT 27.094 52.678 27.146 52.714 ;
      RECT 26.694 52.678 26.746 52.714 ;
      RECT 26.294 52.678 26.346 52.714 ;
      RECT 25.894 52.678 25.946 52.714 ;
      RECT 25.494 52.678 25.546 52.714 ;
      RECT 25.094 52.678 25.146 52.714 ;
      RECT 24.694 52.678 24.746 52.714 ;
      RECT 24.294 52.678 24.346 52.714 ;
      RECT 23.894 52.678 23.946 52.714 ;
      RECT 23.494 52.678 23.546 52.714 ;
      RECT 23.094 52.678 23.146 52.714 ;
      RECT 21.814 52.678 21.868 52.714 ;
      RECT 19.838 52.678 19.886 52.714 ;
      RECT 19.53 52.678 19.578 52.714 ;
      RECT 16.882 52.678 16.936 52.714 ;
      RECT 16.422 52.678 16.47 52.714 ;
      RECT 16.114 52.678 16.162 52.714 ;
      RECT 14.132 52.678 14.186 52.714 ;
      RECT 13.294 52.678 13.346 52.714 ;
      RECT 12.894 52.678 12.946 52.714 ;
      RECT 12.494 52.678 12.546 52.714 ;
      RECT 12.094 52.678 12.146 52.714 ;
      RECT 11.694 52.678 11.746 52.714 ;
      RECT 11.294 52.678 11.346 52.714 ;
      RECT 10.894 52.678 10.946 52.714 ;
      RECT 10.494 52.678 10.546 52.714 ;
      RECT 10.094 52.678 10.146 52.714 ;
      RECT 9.694 52.678 9.746 52.714 ;
      RECT 9.294 52.678 9.346 52.714 ;
      RECT 8.894 52.678 8.946 52.714 ;
      RECT 8.494 52.678 8.546 52.714 ;
      RECT 8.094 52.678 8.146 52.714 ;
      RECT 7.694 52.678 7.746 52.714 ;
      RECT 7.294 52.678 7.346 52.714 ;
      RECT 6.894 52.678 6.946 52.714 ;
      RECT 6.494 52.678 6.546 52.714 ;
      RECT 6.094 52.678 6.146 52.714 ;
      RECT 5.694 52.678 5.746 52.714 ;
      RECT 5.294 52.678 5.346 52.714 ;
      RECT 4.894 52.678 4.946 52.714 ;
      RECT 4.494 52.678 4.546 52.714 ;
      RECT 4.094 52.678 4.146 52.714 ;
      RECT 3.694 52.678 3.746 52.714 ;
      RECT 3.294 52.678 3.346 52.714 ;
      RECT 2.894 52.678 2.946 52.714 ;
      RECT 2.494 52.678 2.546 52.714 ;
      RECT 2.094 52.678 2.146 52.714 ;
      RECT 1.694 52.678 1.746 52.714 ;
      RECT 1.294 52.678 1.346 52.714 ;
      RECT 0.894 52.678 0.946 52.714 ;
      RECT 21.414 52.602 21.468 52.638 ;
      RECT 14.532 52.602 14.586 52.638 ;
      RECT 19.606 52.449 19.654 52.485 ;
      RECT 18.08 52.449 18.12 52.485 ;
      RECT 16.718 52.449 16.772 52.485 ;
      RECT 16.346 52.449 16.394 52.485 ;
      RECT 20.37 52.4545 20.442 52.4795 ;
      RECT 18.764 52.4545 18.836 52.4795 ;
      RECT 15.558 52.4545 15.63 52.4795 ;
      RECT 21.978 52.302 22.022 52.338 ;
      RECT 13.978 52.302 14.022 52.338 ;
      RECT 18.764 52.3075 18.836 52.3325 ;
      RECT 19.762 52.155 19.81 52.191 ;
      RECT 17.616 52.155 17.656 52.191 ;
      RECT 16.19 52.155 16.238 52.191 ;
      RECT 35.254 51.926 35.306 51.962 ;
      RECT 34.854 51.926 34.906 51.962 ;
      RECT 34.454 51.926 34.506 51.962 ;
      RECT 34.054 51.926 34.106 51.962 ;
      RECT 33.654 51.926 33.706 51.962 ;
      RECT 33.254 51.926 33.306 51.962 ;
      RECT 32.854 51.926 32.906 51.962 ;
      RECT 32.454 51.926 32.506 51.962 ;
      RECT 32.054 51.926 32.106 51.962 ;
      RECT 31.654 51.926 31.706 51.962 ;
      RECT 31.254 51.926 31.306 51.962 ;
      RECT 30.854 51.926 30.906 51.962 ;
      RECT 30.454 51.926 30.506 51.962 ;
      RECT 30.054 51.926 30.106 51.962 ;
      RECT 29.654 51.926 29.706 51.962 ;
      RECT 29.254 51.926 29.306 51.962 ;
      RECT 28.854 51.926 28.906 51.962 ;
      RECT 28.454 51.926 28.506 51.962 ;
      RECT 28.054 51.926 28.106 51.962 ;
      RECT 27.654 51.926 27.706 51.962 ;
      RECT 27.254 51.926 27.306 51.962 ;
      RECT 26.854 51.926 26.906 51.962 ;
      RECT 26.454 51.926 26.506 51.962 ;
      RECT 26.054 51.926 26.106 51.962 ;
      RECT 25.654 51.926 25.706 51.962 ;
      RECT 25.254 51.926 25.306 51.962 ;
      RECT 24.854 51.926 24.906 51.962 ;
      RECT 24.454 51.926 24.506 51.962 ;
      RECT 24.054 51.926 24.106 51.962 ;
      RECT 23.654 51.926 23.706 51.962 ;
      RECT 23.254 51.926 23.306 51.962 ;
      RECT 22.854 51.926 22.906 51.962 ;
      RECT 22.694 51.926 22.746 51.962 ;
      RECT 21.732 51.926 21.786 51.962 ;
      RECT 14.214 51.926 14.268 51.962 ;
      RECT 13.054 51.926 13.106 51.962 ;
      RECT 12.654 51.926 12.706 51.962 ;
      RECT 12.254 51.926 12.306 51.962 ;
      RECT 11.854 51.926 11.906 51.962 ;
      RECT 11.454 51.926 11.506 51.962 ;
      RECT 11.054 51.926 11.106 51.962 ;
      RECT 10.654 51.926 10.706 51.962 ;
      RECT 10.254 51.926 10.306 51.962 ;
      RECT 9.854 51.926 9.906 51.962 ;
      RECT 9.454 51.926 9.506 51.962 ;
      RECT 9.054 51.926 9.106 51.962 ;
      RECT 8.654 51.926 8.706 51.962 ;
      RECT 8.254 51.926 8.306 51.962 ;
      RECT 7.854 51.926 7.906 51.962 ;
      RECT 7.454 51.926 7.506 51.962 ;
      RECT 7.054 51.926 7.106 51.962 ;
      RECT 6.654 51.926 6.706 51.962 ;
      RECT 6.254 51.926 6.306 51.962 ;
      RECT 5.854 51.926 5.906 51.962 ;
      RECT 5.454 51.926 5.506 51.962 ;
      RECT 5.054 51.926 5.106 51.962 ;
      RECT 4.654 51.926 4.706 51.962 ;
      RECT 4.254 51.926 4.306 51.962 ;
      RECT 3.854 51.926 3.906 51.962 ;
      RECT 3.454 51.926 3.506 51.962 ;
      RECT 3.054 51.926 3.106 51.962 ;
      RECT 2.654 51.926 2.706 51.962 ;
      RECT 2.254 51.926 2.306 51.962 ;
      RECT 1.854 51.926 1.906 51.962 ;
      RECT 1.454 51.926 1.506 51.962 ;
      RECT 1.054 51.926 1.106 51.962 ;
      RECT 0.654 51.926 0.706 51.962 ;
      RECT 21.978 51.702 22.022 51.738 ;
      RECT 21.096 51.702 21.14 51.738 ;
      RECT 14.86 51.702 14.904 51.738 ;
      RECT 13.978 51.702 14.022 51.738 ;
      RECT 35.494 51.478 35.546 51.514 ;
      RECT 35.094 51.478 35.146 51.514 ;
      RECT 34.694 51.478 34.746 51.514 ;
      RECT 34.294 51.478 34.346 51.514 ;
      RECT 33.894 51.478 33.946 51.514 ;
      RECT 33.494 51.478 33.546 51.514 ;
      RECT 33.094 51.478 33.146 51.514 ;
      RECT 32.694 51.478 32.746 51.514 ;
      RECT 32.294 51.478 32.346 51.514 ;
      RECT 31.894 51.478 31.946 51.514 ;
      RECT 31.494 51.478 31.546 51.514 ;
      RECT 31.094 51.478 31.146 51.514 ;
      RECT 30.694 51.478 30.746 51.514 ;
      RECT 30.294 51.478 30.346 51.514 ;
      RECT 29.894 51.478 29.946 51.514 ;
      RECT 29.494 51.478 29.546 51.514 ;
      RECT 29.094 51.478 29.146 51.514 ;
      RECT 28.694 51.478 28.746 51.514 ;
      RECT 28.294 51.478 28.346 51.514 ;
      RECT 27.894 51.478 27.946 51.514 ;
      RECT 27.494 51.478 27.546 51.514 ;
      RECT 27.094 51.478 27.146 51.514 ;
      RECT 26.694 51.478 26.746 51.514 ;
      RECT 26.294 51.478 26.346 51.514 ;
      RECT 25.894 51.478 25.946 51.514 ;
      RECT 25.494 51.478 25.546 51.514 ;
      RECT 25.094 51.478 25.146 51.514 ;
      RECT 24.694 51.478 24.746 51.514 ;
      RECT 24.294 51.478 24.346 51.514 ;
      RECT 23.894 51.478 23.946 51.514 ;
      RECT 23.494 51.478 23.546 51.514 ;
      RECT 23.094 51.478 23.146 51.514 ;
      RECT 21.814 51.478 21.868 51.514 ;
      RECT 19.838 51.478 19.886 51.514 ;
      RECT 19.53 51.478 19.578 51.514 ;
      RECT 16.882 51.478 16.936 51.514 ;
      RECT 16.422 51.478 16.47 51.514 ;
      RECT 16.114 51.478 16.162 51.514 ;
      RECT 14.132 51.478 14.186 51.514 ;
      RECT 13.294 51.478 13.346 51.514 ;
      RECT 12.894 51.478 12.946 51.514 ;
      RECT 12.494 51.478 12.546 51.514 ;
      RECT 12.094 51.478 12.146 51.514 ;
      RECT 11.694 51.478 11.746 51.514 ;
      RECT 11.294 51.478 11.346 51.514 ;
      RECT 10.894 51.478 10.946 51.514 ;
      RECT 10.494 51.478 10.546 51.514 ;
      RECT 10.094 51.478 10.146 51.514 ;
      RECT 9.694 51.478 9.746 51.514 ;
      RECT 9.294 51.478 9.346 51.514 ;
      RECT 8.894 51.478 8.946 51.514 ;
      RECT 8.494 51.478 8.546 51.514 ;
      RECT 8.094 51.478 8.146 51.514 ;
      RECT 7.694 51.478 7.746 51.514 ;
      RECT 7.294 51.478 7.346 51.514 ;
      RECT 6.894 51.478 6.946 51.514 ;
      RECT 6.494 51.478 6.546 51.514 ;
      RECT 6.094 51.478 6.146 51.514 ;
      RECT 5.694 51.478 5.746 51.514 ;
      RECT 5.294 51.478 5.346 51.514 ;
      RECT 4.894 51.478 4.946 51.514 ;
      RECT 4.494 51.478 4.546 51.514 ;
      RECT 4.094 51.478 4.146 51.514 ;
      RECT 3.694 51.478 3.746 51.514 ;
      RECT 3.294 51.478 3.346 51.514 ;
      RECT 2.894 51.478 2.946 51.514 ;
      RECT 2.494 51.478 2.546 51.514 ;
      RECT 2.094 51.478 2.146 51.514 ;
      RECT 1.694 51.478 1.746 51.514 ;
      RECT 1.294 51.478 1.346 51.514 ;
      RECT 0.894 51.478 0.946 51.514 ;
      RECT 21.414 51.402 21.468 51.438 ;
      RECT 14.532 51.402 14.586 51.438 ;
      RECT 19.606 51.249 19.654 51.285 ;
      RECT 18.08 51.249 18.12 51.285 ;
      RECT 16.718 51.249 16.772 51.285 ;
      RECT 16.346 51.249 16.394 51.285 ;
      RECT 20.37 51.2545 20.442 51.2795 ;
      RECT 18.764 51.2545 18.836 51.2795 ;
      RECT 15.558 51.2545 15.63 51.2795 ;
      RECT 21.978 51.102 22.022 51.138 ;
      RECT 13.978 51.102 14.022 51.138 ;
      RECT 18.764 51.1075 18.836 51.1325 ;
      RECT 19.762 50.955 19.81 50.991 ;
      RECT 17.616 50.955 17.656 50.991 ;
      RECT 16.19 50.955 16.238 50.991 ;
      RECT 35.254 50.726 35.306 50.762 ;
      RECT 34.854 50.726 34.906 50.762 ;
      RECT 34.454 50.726 34.506 50.762 ;
      RECT 34.054 50.726 34.106 50.762 ;
      RECT 33.654 50.726 33.706 50.762 ;
      RECT 33.254 50.726 33.306 50.762 ;
      RECT 32.854 50.726 32.906 50.762 ;
      RECT 32.454 50.726 32.506 50.762 ;
      RECT 32.054 50.726 32.106 50.762 ;
      RECT 31.654 50.726 31.706 50.762 ;
      RECT 31.254 50.726 31.306 50.762 ;
      RECT 30.854 50.726 30.906 50.762 ;
      RECT 30.454 50.726 30.506 50.762 ;
      RECT 30.054 50.726 30.106 50.762 ;
      RECT 29.654 50.726 29.706 50.762 ;
      RECT 29.254 50.726 29.306 50.762 ;
      RECT 28.854 50.726 28.906 50.762 ;
      RECT 28.454 50.726 28.506 50.762 ;
      RECT 28.054 50.726 28.106 50.762 ;
      RECT 27.654 50.726 27.706 50.762 ;
      RECT 27.254 50.726 27.306 50.762 ;
      RECT 26.854 50.726 26.906 50.762 ;
      RECT 26.454 50.726 26.506 50.762 ;
      RECT 26.054 50.726 26.106 50.762 ;
      RECT 25.654 50.726 25.706 50.762 ;
      RECT 25.254 50.726 25.306 50.762 ;
      RECT 24.854 50.726 24.906 50.762 ;
      RECT 24.454 50.726 24.506 50.762 ;
      RECT 24.054 50.726 24.106 50.762 ;
      RECT 23.654 50.726 23.706 50.762 ;
      RECT 23.254 50.726 23.306 50.762 ;
      RECT 22.854 50.726 22.906 50.762 ;
      RECT 22.694 50.726 22.746 50.762 ;
      RECT 21.732 50.726 21.786 50.762 ;
      RECT 14.214 50.726 14.268 50.762 ;
      RECT 13.054 50.726 13.106 50.762 ;
      RECT 12.654 50.726 12.706 50.762 ;
      RECT 12.254 50.726 12.306 50.762 ;
      RECT 11.854 50.726 11.906 50.762 ;
      RECT 11.454 50.726 11.506 50.762 ;
      RECT 11.054 50.726 11.106 50.762 ;
      RECT 10.654 50.726 10.706 50.762 ;
      RECT 10.254 50.726 10.306 50.762 ;
      RECT 9.854 50.726 9.906 50.762 ;
      RECT 9.454 50.726 9.506 50.762 ;
      RECT 9.054 50.726 9.106 50.762 ;
      RECT 8.654 50.726 8.706 50.762 ;
      RECT 8.254 50.726 8.306 50.762 ;
      RECT 7.854 50.726 7.906 50.762 ;
      RECT 7.454 50.726 7.506 50.762 ;
      RECT 7.054 50.726 7.106 50.762 ;
      RECT 6.654 50.726 6.706 50.762 ;
      RECT 6.254 50.726 6.306 50.762 ;
      RECT 5.854 50.726 5.906 50.762 ;
      RECT 5.454 50.726 5.506 50.762 ;
      RECT 5.054 50.726 5.106 50.762 ;
      RECT 4.654 50.726 4.706 50.762 ;
      RECT 4.254 50.726 4.306 50.762 ;
      RECT 3.854 50.726 3.906 50.762 ;
      RECT 3.454 50.726 3.506 50.762 ;
      RECT 3.054 50.726 3.106 50.762 ;
      RECT 2.654 50.726 2.706 50.762 ;
      RECT 2.254 50.726 2.306 50.762 ;
      RECT 1.854 50.726 1.906 50.762 ;
      RECT 1.454 50.726 1.506 50.762 ;
      RECT 1.054 50.726 1.106 50.762 ;
      RECT 0.654 50.726 0.706 50.762 ;
      RECT 21.978 50.502 22.022 50.538 ;
      RECT 21.096 50.502 21.14 50.538 ;
      RECT 14.86 50.502 14.904 50.538 ;
      RECT 13.978 50.502 14.022 50.538 ;
      RECT 35.494 50.278 35.546 50.314 ;
      RECT 35.094 50.278 35.146 50.314 ;
      RECT 34.694 50.278 34.746 50.314 ;
      RECT 34.294 50.278 34.346 50.314 ;
      RECT 33.894 50.278 33.946 50.314 ;
      RECT 33.494 50.278 33.546 50.314 ;
      RECT 33.094 50.278 33.146 50.314 ;
      RECT 32.694 50.278 32.746 50.314 ;
      RECT 32.294 50.278 32.346 50.314 ;
      RECT 31.894 50.278 31.946 50.314 ;
      RECT 31.494 50.278 31.546 50.314 ;
      RECT 31.094 50.278 31.146 50.314 ;
      RECT 30.694 50.278 30.746 50.314 ;
      RECT 30.294 50.278 30.346 50.314 ;
      RECT 29.894 50.278 29.946 50.314 ;
      RECT 29.494 50.278 29.546 50.314 ;
      RECT 29.094 50.278 29.146 50.314 ;
      RECT 28.694 50.278 28.746 50.314 ;
      RECT 28.294 50.278 28.346 50.314 ;
      RECT 27.894 50.278 27.946 50.314 ;
      RECT 27.494 50.278 27.546 50.314 ;
      RECT 27.094 50.278 27.146 50.314 ;
      RECT 26.694 50.278 26.746 50.314 ;
      RECT 26.294 50.278 26.346 50.314 ;
      RECT 25.894 50.278 25.946 50.314 ;
      RECT 25.494 50.278 25.546 50.314 ;
      RECT 25.094 50.278 25.146 50.314 ;
      RECT 24.694 50.278 24.746 50.314 ;
      RECT 24.294 50.278 24.346 50.314 ;
      RECT 23.894 50.278 23.946 50.314 ;
      RECT 23.494 50.278 23.546 50.314 ;
      RECT 23.094 50.278 23.146 50.314 ;
      RECT 21.814 50.278 21.868 50.314 ;
      RECT 19.838 50.278 19.886 50.314 ;
      RECT 19.53 50.278 19.578 50.314 ;
      RECT 16.882 50.278 16.936 50.314 ;
      RECT 16.422 50.278 16.47 50.314 ;
      RECT 16.114 50.278 16.162 50.314 ;
      RECT 14.132 50.278 14.186 50.314 ;
      RECT 13.294 50.278 13.346 50.314 ;
      RECT 12.894 50.278 12.946 50.314 ;
      RECT 12.494 50.278 12.546 50.314 ;
      RECT 12.094 50.278 12.146 50.314 ;
      RECT 11.694 50.278 11.746 50.314 ;
      RECT 11.294 50.278 11.346 50.314 ;
      RECT 10.894 50.278 10.946 50.314 ;
      RECT 10.494 50.278 10.546 50.314 ;
      RECT 10.094 50.278 10.146 50.314 ;
      RECT 9.694 50.278 9.746 50.314 ;
      RECT 9.294 50.278 9.346 50.314 ;
      RECT 8.894 50.278 8.946 50.314 ;
      RECT 8.494 50.278 8.546 50.314 ;
      RECT 8.094 50.278 8.146 50.314 ;
      RECT 7.694 50.278 7.746 50.314 ;
      RECT 7.294 50.278 7.346 50.314 ;
      RECT 6.894 50.278 6.946 50.314 ;
      RECT 6.494 50.278 6.546 50.314 ;
      RECT 6.094 50.278 6.146 50.314 ;
      RECT 5.694 50.278 5.746 50.314 ;
      RECT 5.294 50.278 5.346 50.314 ;
      RECT 4.894 50.278 4.946 50.314 ;
      RECT 4.494 50.278 4.546 50.314 ;
      RECT 4.094 50.278 4.146 50.314 ;
      RECT 3.694 50.278 3.746 50.314 ;
      RECT 3.294 50.278 3.346 50.314 ;
      RECT 2.894 50.278 2.946 50.314 ;
      RECT 2.494 50.278 2.546 50.314 ;
      RECT 2.094 50.278 2.146 50.314 ;
      RECT 1.694 50.278 1.746 50.314 ;
      RECT 1.294 50.278 1.346 50.314 ;
      RECT 0.894 50.278 0.946 50.314 ;
      RECT 21.414 50.202 21.468 50.238 ;
      RECT 14.532 50.202 14.586 50.238 ;
      RECT 19.606 50.049 19.654 50.085 ;
      RECT 18.08 50.049 18.12 50.085 ;
      RECT 16.718 50.049 16.772 50.085 ;
      RECT 16.346 50.049 16.394 50.085 ;
      RECT 20.37 50.0545 20.442 50.0795 ;
      RECT 18.764 50.0545 18.836 50.0795 ;
      RECT 15.558 50.0545 15.63 50.0795 ;
      RECT 21.978 49.902 22.022 49.938 ;
      RECT 13.978 49.902 14.022 49.938 ;
      RECT 18.764 49.9075 18.836 49.9325 ;
      RECT 19.762 49.755 19.81 49.791 ;
      RECT 17.616 49.755 17.656 49.791 ;
      RECT 16.19 49.755 16.238 49.791 ;
      RECT 35.254 49.526 35.306 49.562 ;
      RECT 34.854 49.526 34.906 49.562 ;
      RECT 34.454 49.526 34.506 49.562 ;
      RECT 34.054 49.526 34.106 49.562 ;
      RECT 33.654 49.526 33.706 49.562 ;
      RECT 33.254 49.526 33.306 49.562 ;
      RECT 32.854 49.526 32.906 49.562 ;
      RECT 32.454 49.526 32.506 49.562 ;
      RECT 32.054 49.526 32.106 49.562 ;
      RECT 31.654 49.526 31.706 49.562 ;
      RECT 31.254 49.526 31.306 49.562 ;
      RECT 30.854 49.526 30.906 49.562 ;
      RECT 30.454 49.526 30.506 49.562 ;
      RECT 30.054 49.526 30.106 49.562 ;
      RECT 29.654 49.526 29.706 49.562 ;
      RECT 29.254 49.526 29.306 49.562 ;
      RECT 28.854 49.526 28.906 49.562 ;
      RECT 28.454 49.526 28.506 49.562 ;
      RECT 28.054 49.526 28.106 49.562 ;
      RECT 27.654 49.526 27.706 49.562 ;
      RECT 27.254 49.526 27.306 49.562 ;
      RECT 26.854 49.526 26.906 49.562 ;
      RECT 26.454 49.526 26.506 49.562 ;
      RECT 26.054 49.526 26.106 49.562 ;
      RECT 25.654 49.526 25.706 49.562 ;
      RECT 25.254 49.526 25.306 49.562 ;
      RECT 24.854 49.526 24.906 49.562 ;
      RECT 24.454 49.526 24.506 49.562 ;
      RECT 24.054 49.526 24.106 49.562 ;
      RECT 23.654 49.526 23.706 49.562 ;
      RECT 23.254 49.526 23.306 49.562 ;
      RECT 22.854 49.526 22.906 49.562 ;
      RECT 22.694 49.526 22.746 49.562 ;
      RECT 21.732 49.526 21.786 49.562 ;
      RECT 14.214 49.526 14.268 49.562 ;
      RECT 13.054 49.526 13.106 49.562 ;
      RECT 12.654 49.526 12.706 49.562 ;
      RECT 12.254 49.526 12.306 49.562 ;
      RECT 11.854 49.526 11.906 49.562 ;
      RECT 11.454 49.526 11.506 49.562 ;
      RECT 11.054 49.526 11.106 49.562 ;
      RECT 10.654 49.526 10.706 49.562 ;
      RECT 10.254 49.526 10.306 49.562 ;
      RECT 9.854 49.526 9.906 49.562 ;
      RECT 9.454 49.526 9.506 49.562 ;
      RECT 9.054 49.526 9.106 49.562 ;
      RECT 8.654 49.526 8.706 49.562 ;
      RECT 8.254 49.526 8.306 49.562 ;
      RECT 7.854 49.526 7.906 49.562 ;
      RECT 7.454 49.526 7.506 49.562 ;
      RECT 7.054 49.526 7.106 49.562 ;
      RECT 6.654 49.526 6.706 49.562 ;
      RECT 6.254 49.526 6.306 49.562 ;
      RECT 5.854 49.526 5.906 49.562 ;
      RECT 5.454 49.526 5.506 49.562 ;
      RECT 5.054 49.526 5.106 49.562 ;
      RECT 4.654 49.526 4.706 49.562 ;
      RECT 4.254 49.526 4.306 49.562 ;
      RECT 3.854 49.526 3.906 49.562 ;
      RECT 3.454 49.526 3.506 49.562 ;
      RECT 3.054 49.526 3.106 49.562 ;
      RECT 2.654 49.526 2.706 49.562 ;
      RECT 2.254 49.526 2.306 49.562 ;
      RECT 1.854 49.526 1.906 49.562 ;
      RECT 1.454 49.526 1.506 49.562 ;
      RECT 1.054 49.526 1.106 49.562 ;
      RECT 0.654 49.526 0.706 49.562 ;
      RECT 21.978 49.302 22.022 49.338 ;
      RECT 21.096 49.302 21.14 49.338 ;
      RECT 14.86 49.302 14.904 49.338 ;
      RECT 13.978 49.302 14.022 49.338 ;
      RECT 35.494 49.078 35.546 49.114 ;
      RECT 35.094 49.078 35.146 49.114 ;
      RECT 34.694 49.078 34.746 49.114 ;
      RECT 34.294 49.078 34.346 49.114 ;
      RECT 33.894 49.078 33.946 49.114 ;
      RECT 33.494 49.078 33.546 49.114 ;
      RECT 33.094 49.078 33.146 49.114 ;
      RECT 32.694 49.078 32.746 49.114 ;
      RECT 32.294 49.078 32.346 49.114 ;
      RECT 31.894 49.078 31.946 49.114 ;
      RECT 31.494 49.078 31.546 49.114 ;
      RECT 31.094 49.078 31.146 49.114 ;
      RECT 30.694 49.078 30.746 49.114 ;
      RECT 30.294 49.078 30.346 49.114 ;
      RECT 29.894 49.078 29.946 49.114 ;
      RECT 29.494 49.078 29.546 49.114 ;
      RECT 29.094 49.078 29.146 49.114 ;
      RECT 28.694 49.078 28.746 49.114 ;
      RECT 28.294 49.078 28.346 49.114 ;
      RECT 27.894 49.078 27.946 49.114 ;
      RECT 27.494 49.078 27.546 49.114 ;
      RECT 27.094 49.078 27.146 49.114 ;
      RECT 26.694 49.078 26.746 49.114 ;
      RECT 26.294 49.078 26.346 49.114 ;
      RECT 25.894 49.078 25.946 49.114 ;
      RECT 25.494 49.078 25.546 49.114 ;
      RECT 25.094 49.078 25.146 49.114 ;
      RECT 24.694 49.078 24.746 49.114 ;
      RECT 24.294 49.078 24.346 49.114 ;
      RECT 23.894 49.078 23.946 49.114 ;
      RECT 23.494 49.078 23.546 49.114 ;
      RECT 23.094 49.078 23.146 49.114 ;
      RECT 21.814 49.078 21.868 49.114 ;
      RECT 19.838 49.078 19.886 49.114 ;
      RECT 19.53 49.078 19.578 49.114 ;
      RECT 16.882 49.078 16.936 49.114 ;
      RECT 16.422 49.078 16.47 49.114 ;
      RECT 16.114 49.078 16.162 49.114 ;
      RECT 14.132 49.078 14.186 49.114 ;
      RECT 13.294 49.078 13.346 49.114 ;
      RECT 12.894 49.078 12.946 49.114 ;
      RECT 12.494 49.078 12.546 49.114 ;
      RECT 12.094 49.078 12.146 49.114 ;
      RECT 11.694 49.078 11.746 49.114 ;
      RECT 11.294 49.078 11.346 49.114 ;
      RECT 10.894 49.078 10.946 49.114 ;
      RECT 10.494 49.078 10.546 49.114 ;
      RECT 10.094 49.078 10.146 49.114 ;
      RECT 9.694 49.078 9.746 49.114 ;
      RECT 9.294 49.078 9.346 49.114 ;
      RECT 8.894 49.078 8.946 49.114 ;
      RECT 8.494 49.078 8.546 49.114 ;
      RECT 8.094 49.078 8.146 49.114 ;
      RECT 7.694 49.078 7.746 49.114 ;
      RECT 7.294 49.078 7.346 49.114 ;
      RECT 6.894 49.078 6.946 49.114 ;
      RECT 6.494 49.078 6.546 49.114 ;
      RECT 6.094 49.078 6.146 49.114 ;
      RECT 5.694 49.078 5.746 49.114 ;
      RECT 5.294 49.078 5.346 49.114 ;
      RECT 4.894 49.078 4.946 49.114 ;
      RECT 4.494 49.078 4.546 49.114 ;
      RECT 4.094 49.078 4.146 49.114 ;
      RECT 3.694 49.078 3.746 49.114 ;
      RECT 3.294 49.078 3.346 49.114 ;
      RECT 2.894 49.078 2.946 49.114 ;
      RECT 2.494 49.078 2.546 49.114 ;
      RECT 2.094 49.078 2.146 49.114 ;
      RECT 1.694 49.078 1.746 49.114 ;
      RECT 1.294 49.078 1.346 49.114 ;
      RECT 0.894 49.078 0.946 49.114 ;
      RECT 21.414 49.002 21.468 49.038 ;
      RECT 14.532 49.002 14.586 49.038 ;
      RECT 19.606 48.849 19.654 48.885 ;
      RECT 18.08 48.849 18.12 48.885 ;
      RECT 16.718 48.849 16.772 48.885 ;
      RECT 16.346 48.849 16.394 48.885 ;
      RECT 20.37 48.8545 20.442 48.8795 ;
      RECT 18.764 48.8545 18.836 48.8795 ;
      RECT 15.558 48.8545 15.63 48.8795 ;
      RECT 21.978 48.702 22.022 48.738 ;
      RECT 13.978 48.702 14.022 48.738 ;
      RECT 18.764 48.7075 18.836 48.7325 ;
      RECT 19.762 48.555 19.81 48.591 ;
      RECT 17.616 48.555 17.656 48.591 ;
      RECT 16.19 48.555 16.238 48.591 ;
      RECT 35.254 48.326 35.306 48.362 ;
      RECT 34.854 48.326 34.906 48.362 ;
      RECT 34.454 48.326 34.506 48.362 ;
      RECT 34.054 48.326 34.106 48.362 ;
      RECT 33.654 48.326 33.706 48.362 ;
      RECT 33.254 48.326 33.306 48.362 ;
      RECT 32.854 48.326 32.906 48.362 ;
      RECT 32.454 48.326 32.506 48.362 ;
      RECT 32.054 48.326 32.106 48.362 ;
      RECT 31.654 48.326 31.706 48.362 ;
      RECT 31.254 48.326 31.306 48.362 ;
      RECT 30.854 48.326 30.906 48.362 ;
      RECT 30.454 48.326 30.506 48.362 ;
      RECT 30.054 48.326 30.106 48.362 ;
      RECT 29.654 48.326 29.706 48.362 ;
      RECT 29.254 48.326 29.306 48.362 ;
      RECT 28.854 48.326 28.906 48.362 ;
      RECT 28.454 48.326 28.506 48.362 ;
      RECT 28.054 48.326 28.106 48.362 ;
      RECT 27.654 48.326 27.706 48.362 ;
      RECT 27.254 48.326 27.306 48.362 ;
      RECT 26.854 48.326 26.906 48.362 ;
      RECT 26.454 48.326 26.506 48.362 ;
      RECT 26.054 48.326 26.106 48.362 ;
      RECT 25.654 48.326 25.706 48.362 ;
      RECT 25.254 48.326 25.306 48.362 ;
      RECT 24.854 48.326 24.906 48.362 ;
      RECT 24.454 48.326 24.506 48.362 ;
      RECT 24.054 48.326 24.106 48.362 ;
      RECT 23.654 48.326 23.706 48.362 ;
      RECT 23.254 48.326 23.306 48.362 ;
      RECT 22.854 48.326 22.906 48.362 ;
      RECT 22.694 48.326 22.746 48.362 ;
      RECT 21.732 48.326 21.786 48.362 ;
      RECT 14.214 48.326 14.268 48.362 ;
      RECT 13.054 48.326 13.106 48.362 ;
      RECT 12.654 48.326 12.706 48.362 ;
      RECT 12.254 48.326 12.306 48.362 ;
      RECT 11.854 48.326 11.906 48.362 ;
      RECT 11.454 48.326 11.506 48.362 ;
      RECT 11.054 48.326 11.106 48.362 ;
      RECT 10.654 48.326 10.706 48.362 ;
      RECT 10.254 48.326 10.306 48.362 ;
      RECT 9.854 48.326 9.906 48.362 ;
      RECT 9.454 48.326 9.506 48.362 ;
      RECT 9.054 48.326 9.106 48.362 ;
      RECT 8.654 48.326 8.706 48.362 ;
      RECT 8.254 48.326 8.306 48.362 ;
      RECT 7.854 48.326 7.906 48.362 ;
      RECT 7.454 48.326 7.506 48.362 ;
      RECT 7.054 48.326 7.106 48.362 ;
      RECT 6.654 48.326 6.706 48.362 ;
      RECT 6.254 48.326 6.306 48.362 ;
      RECT 5.854 48.326 5.906 48.362 ;
      RECT 5.454 48.326 5.506 48.362 ;
      RECT 5.054 48.326 5.106 48.362 ;
      RECT 4.654 48.326 4.706 48.362 ;
      RECT 4.254 48.326 4.306 48.362 ;
      RECT 3.854 48.326 3.906 48.362 ;
      RECT 3.454 48.326 3.506 48.362 ;
      RECT 3.054 48.326 3.106 48.362 ;
      RECT 2.654 48.326 2.706 48.362 ;
      RECT 2.254 48.326 2.306 48.362 ;
      RECT 1.854 48.326 1.906 48.362 ;
      RECT 1.454 48.326 1.506 48.362 ;
      RECT 1.054 48.326 1.106 48.362 ;
      RECT 0.654 48.326 0.706 48.362 ;
      RECT 21.978 48.102 22.022 48.138 ;
      RECT 21.096 48.102 21.14 48.138 ;
      RECT 14.86 48.102 14.904 48.138 ;
      RECT 13.978 48.102 14.022 48.138 ;
      RECT 35.494 47.878 35.546 47.914 ;
      RECT 35.094 47.878 35.146 47.914 ;
      RECT 34.694 47.878 34.746 47.914 ;
      RECT 34.294 47.878 34.346 47.914 ;
      RECT 33.894 47.878 33.946 47.914 ;
      RECT 33.494 47.878 33.546 47.914 ;
      RECT 33.094 47.878 33.146 47.914 ;
      RECT 32.694 47.878 32.746 47.914 ;
      RECT 32.294 47.878 32.346 47.914 ;
      RECT 31.894 47.878 31.946 47.914 ;
      RECT 31.494 47.878 31.546 47.914 ;
      RECT 31.094 47.878 31.146 47.914 ;
      RECT 30.694 47.878 30.746 47.914 ;
      RECT 30.294 47.878 30.346 47.914 ;
      RECT 29.894 47.878 29.946 47.914 ;
      RECT 29.494 47.878 29.546 47.914 ;
      RECT 29.094 47.878 29.146 47.914 ;
      RECT 28.694 47.878 28.746 47.914 ;
      RECT 28.294 47.878 28.346 47.914 ;
      RECT 27.894 47.878 27.946 47.914 ;
      RECT 27.494 47.878 27.546 47.914 ;
      RECT 27.094 47.878 27.146 47.914 ;
      RECT 26.694 47.878 26.746 47.914 ;
      RECT 26.294 47.878 26.346 47.914 ;
      RECT 25.894 47.878 25.946 47.914 ;
      RECT 25.494 47.878 25.546 47.914 ;
      RECT 25.094 47.878 25.146 47.914 ;
      RECT 24.694 47.878 24.746 47.914 ;
      RECT 24.294 47.878 24.346 47.914 ;
      RECT 23.894 47.878 23.946 47.914 ;
      RECT 23.494 47.878 23.546 47.914 ;
      RECT 23.094 47.878 23.146 47.914 ;
      RECT 21.814 47.878 21.868 47.914 ;
      RECT 19.838 47.878 19.886 47.914 ;
      RECT 19.53 47.878 19.578 47.914 ;
      RECT 16.882 47.878 16.936 47.914 ;
      RECT 16.422 47.878 16.47 47.914 ;
      RECT 16.114 47.878 16.162 47.914 ;
      RECT 14.132 47.878 14.186 47.914 ;
      RECT 13.294 47.878 13.346 47.914 ;
      RECT 12.894 47.878 12.946 47.914 ;
      RECT 12.494 47.878 12.546 47.914 ;
      RECT 12.094 47.878 12.146 47.914 ;
      RECT 11.694 47.878 11.746 47.914 ;
      RECT 11.294 47.878 11.346 47.914 ;
      RECT 10.894 47.878 10.946 47.914 ;
      RECT 10.494 47.878 10.546 47.914 ;
      RECT 10.094 47.878 10.146 47.914 ;
      RECT 9.694 47.878 9.746 47.914 ;
      RECT 9.294 47.878 9.346 47.914 ;
      RECT 8.894 47.878 8.946 47.914 ;
      RECT 8.494 47.878 8.546 47.914 ;
      RECT 8.094 47.878 8.146 47.914 ;
      RECT 7.694 47.878 7.746 47.914 ;
      RECT 7.294 47.878 7.346 47.914 ;
      RECT 6.894 47.878 6.946 47.914 ;
      RECT 6.494 47.878 6.546 47.914 ;
      RECT 6.094 47.878 6.146 47.914 ;
      RECT 5.694 47.878 5.746 47.914 ;
      RECT 5.294 47.878 5.346 47.914 ;
      RECT 4.894 47.878 4.946 47.914 ;
      RECT 4.494 47.878 4.546 47.914 ;
      RECT 4.094 47.878 4.146 47.914 ;
      RECT 3.694 47.878 3.746 47.914 ;
      RECT 3.294 47.878 3.346 47.914 ;
      RECT 2.894 47.878 2.946 47.914 ;
      RECT 2.494 47.878 2.546 47.914 ;
      RECT 2.094 47.878 2.146 47.914 ;
      RECT 1.694 47.878 1.746 47.914 ;
      RECT 1.294 47.878 1.346 47.914 ;
      RECT 0.894 47.878 0.946 47.914 ;
      RECT 21.414 47.802 21.468 47.838 ;
      RECT 14.532 47.802 14.586 47.838 ;
      RECT 19.606 47.649 19.654 47.685 ;
      RECT 18.08 47.649 18.12 47.685 ;
      RECT 16.718 47.649 16.772 47.685 ;
      RECT 16.346 47.649 16.394 47.685 ;
      RECT 20.37 47.6545 20.442 47.6795 ;
      RECT 18.764 47.6545 18.836 47.6795 ;
      RECT 15.558 47.6545 15.63 47.6795 ;
      RECT 21.978 47.502 22.022 47.538 ;
      RECT 13.978 47.502 14.022 47.538 ;
      RECT 18.764 47.5075 18.836 47.5325 ;
      RECT 19.762 47.355 19.81 47.391 ;
      RECT 17.616 47.355 17.656 47.391 ;
      RECT 16.19 47.355 16.238 47.391 ;
      RECT 35.254 47.126 35.306 47.162 ;
      RECT 34.854 47.126 34.906 47.162 ;
      RECT 34.454 47.126 34.506 47.162 ;
      RECT 34.054 47.126 34.106 47.162 ;
      RECT 33.654 47.126 33.706 47.162 ;
      RECT 33.254 47.126 33.306 47.162 ;
      RECT 32.854 47.126 32.906 47.162 ;
      RECT 32.454 47.126 32.506 47.162 ;
      RECT 32.054 47.126 32.106 47.162 ;
      RECT 31.654 47.126 31.706 47.162 ;
      RECT 31.254 47.126 31.306 47.162 ;
      RECT 30.854 47.126 30.906 47.162 ;
      RECT 30.454 47.126 30.506 47.162 ;
      RECT 30.054 47.126 30.106 47.162 ;
      RECT 29.654 47.126 29.706 47.162 ;
      RECT 29.254 47.126 29.306 47.162 ;
      RECT 28.854 47.126 28.906 47.162 ;
      RECT 28.454 47.126 28.506 47.162 ;
      RECT 28.054 47.126 28.106 47.162 ;
      RECT 27.654 47.126 27.706 47.162 ;
      RECT 27.254 47.126 27.306 47.162 ;
      RECT 26.854 47.126 26.906 47.162 ;
      RECT 26.454 47.126 26.506 47.162 ;
      RECT 26.054 47.126 26.106 47.162 ;
      RECT 25.654 47.126 25.706 47.162 ;
      RECT 25.254 47.126 25.306 47.162 ;
      RECT 24.854 47.126 24.906 47.162 ;
      RECT 24.454 47.126 24.506 47.162 ;
      RECT 24.054 47.126 24.106 47.162 ;
      RECT 23.654 47.126 23.706 47.162 ;
      RECT 23.254 47.126 23.306 47.162 ;
      RECT 22.854 47.126 22.906 47.162 ;
      RECT 22.694 47.126 22.746 47.162 ;
      RECT 21.732 47.126 21.786 47.162 ;
      RECT 14.214 47.126 14.268 47.162 ;
      RECT 13.054 47.126 13.106 47.162 ;
      RECT 12.654 47.126 12.706 47.162 ;
      RECT 12.254 47.126 12.306 47.162 ;
      RECT 11.854 47.126 11.906 47.162 ;
      RECT 11.454 47.126 11.506 47.162 ;
      RECT 11.054 47.126 11.106 47.162 ;
      RECT 10.654 47.126 10.706 47.162 ;
      RECT 10.254 47.126 10.306 47.162 ;
      RECT 9.854 47.126 9.906 47.162 ;
      RECT 9.454 47.126 9.506 47.162 ;
      RECT 9.054 47.126 9.106 47.162 ;
      RECT 8.654 47.126 8.706 47.162 ;
      RECT 8.254 47.126 8.306 47.162 ;
      RECT 7.854 47.126 7.906 47.162 ;
      RECT 7.454 47.126 7.506 47.162 ;
      RECT 7.054 47.126 7.106 47.162 ;
      RECT 6.654 47.126 6.706 47.162 ;
      RECT 6.254 47.126 6.306 47.162 ;
      RECT 5.854 47.126 5.906 47.162 ;
      RECT 5.454 47.126 5.506 47.162 ;
      RECT 5.054 47.126 5.106 47.162 ;
      RECT 4.654 47.126 4.706 47.162 ;
      RECT 4.254 47.126 4.306 47.162 ;
      RECT 3.854 47.126 3.906 47.162 ;
      RECT 3.454 47.126 3.506 47.162 ;
      RECT 3.054 47.126 3.106 47.162 ;
      RECT 2.654 47.126 2.706 47.162 ;
      RECT 2.254 47.126 2.306 47.162 ;
      RECT 1.854 47.126 1.906 47.162 ;
      RECT 1.454 47.126 1.506 47.162 ;
      RECT 1.054 47.126 1.106 47.162 ;
      RECT 0.654 47.126 0.706 47.162 ;
      RECT 21.978 46.902 22.022 46.938 ;
      RECT 21.096 46.902 21.14 46.938 ;
      RECT 14.86 46.902 14.904 46.938 ;
      RECT 13.978 46.902 14.022 46.938 ;
      RECT 35.494 46.678 35.546 46.714 ;
      RECT 35.094 46.678 35.146 46.714 ;
      RECT 34.694 46.678 34.746 46.714 ;
      RECT 34.294 46.678 34.346 46.714 ;
      RECT 33.894 46.678 33.946 46.714 ;
      RECT 33.494 46.678 33.546 46.714 ;
      RECT 33.094 46.678 33.146 46.714 ;
      RECT 32.694 46.678 32.746 46.714 ;
      RECT 32.294 46.678 32.346 46.714 ;
      RECT 31.894 46.678 31.946 46.714 ;
      RECT 31.494 46.678 31.546 46.714 ;
      RECT 31.094 46.678 31.146 46.714 ;
      RECT 30.694 46.678 30.746 46.714 ;
      RECT 30.294 46.678 30.346 46.714 ;
      RECT 29.894 46.678 29.946 46.714 ;
      RECT 29.494 46.678 29.546 46.714 ;
      RECT 29.094 46.678 29.146 46.714 ;
      RECT 28.694 46.678 28.746 46.714 ;
      RECT 28.294 46.678 28.346 46.714 ;
      RECT 27.894 46.678 27.946 46.714 ;
      RECT 27.494 46.678 27.546 46.714 ;
      RECT 27.094 46.678 27.146 46.714 ;
      RECT 26.694 46.678 26.746 46.714 ;
      RECT 26.294 46.678 26.346 46.714 ;
      RECT 25.894 46.678 25.946 46.714 ;
      RECT 25.494 46.678 25.546 46.714 ;
      RECT 25.094 46.678 25.146 46.714 ;
      RECT 24.694 46.678 24.746 46.714 ;
      RECT 24.294 46.678 24.346 46.714 ;
      RECT 23.894 46.678 23.946 46.714 ;
      RECT 23.494 46.678 23.546 46.714 ;
      RECT 23.094 46.678 23.146 46.714 ;
      RECT 21.814 46.678 21.868 46.714 ;
      RECT 19.838 46.678 19.886 46.714 ;
      RECT 19.53 46.678 19.578 46.714 ;
      RECT 16.882 46.678 16.936 46.714 ;
      RECT 16.422 46.678 16.47 46.714 ;
      RECT 16.114 46.678 16.162 46.714 ;
      RECT 14.132 46.678 14.186 46.714 ;
      RECT 13.294 46.678 13.346 46.714 ;
      RECT 12.894 46.678 12.946 46.714 ;
      RECT 12.494 46.678 12.546 46.714 ;
      RECT 12.094 46.678 12.146 46.714 ;
      RECT 11.694 46.678 11.746 46.714 ;
      RECT 11.294 46.678 11.346 46.714 ;
      RECT 10.894 46.678 10.946 46.714 ;
      RECT 10.494 46.678 10.546 46.714 ;
      RECT 10.094 46.678 10.146 46.714 ;
      RECT 9.694 46.678 9.746 46.714 ;
      RECT 9.294 46.678 9.346 46.714 ;
      RECT 8.894 46.678 8.946 46.714 ;
      RECT 8.494 46.678 8.546 46.714 ;
      RECT 8.094 46.678 8.146 46.714 ;
      RECT 7.694 46.678 7.746 46.714 ;
      RECT 7.294 46.678 7.346 46.714 ;
      RECT 6.894 46.678 6.946 46.714 ;
      RECT 6.494 46.678 6.546 46.714 ;
      RECT 6.094 46.678 6.146 46.714 ;
      RECT 5.694 46.678 5.746 46.714 ;
      RECT 5.294 46.678 5.346 46.714 ;
      RECT 4.894 46.678 4.946 46.714 ;
      RECT 4.494 46.678 4.546 46.714 ;
      RECT 4.094 46.678 4.146 46.714 ;
      RECT 3.694 46.678 3.746 46.714 ;
      RECT 3.294 46.678 3.346 46.714 ;
      RECT 2.894 46.678 2.946 46.714 ;
      RECT 2.494 46.678 2.546 46.714 ;
      RECT 2.094 46.678 2.146 46.714 ;
      RECT 1.694 46.678 1.746 46.714 ;
      RECT 1.294 46.678 1.346 46.714 ;
      RECT 0.894 46.678 0.946 46.714 ;
      RECT 21.414 46.602 21.468 46.638 ;
      RECT 14.532 46.602 14.586 46.638 ;
      RECT 19.606 46.449 19.654 46.485 ;
      RECT 18.08 46.449 18.12 46.485 ;
      RECT 16.718 46.449 16.772 46.485 ;
      RECT 16.346 46.449 16.394 46.485 ;
      RECT 20.37 46.4545 20.442 46.4795 ;
      RECT 18.764 46.4545 18.836 46.4795 ;
      RECT 15.558 46.4545 15.63 46.4795 ;
      RECT 21.978 46.302 22.022 46.338 ;
      RECT 13.978 46.302 14.022 46.338 ;
      RECT 18.764 46.3075 18.836 46.3325 ;
      RECT 19.762 46.155 19.81 46.191 ;
      RECT 17.616 46.155 17.656 46.191 ;
      RECT 16.19 46.155 16.238 46.191 ;
      RECT 35.254 45.926 35.306 45.962 ;
      RECT 34.854 45.926 34.906 45.962 ;
      RECT 34.454 45.926 34.506 45.962 ;
      RECT 34.054 45.926 34.106 45.962 ;
      RECT 33.654 45.926 33.706 45.962 ;
      RECT 33.254 45.926 33.306 45.962 ;
      RECT 32.854 45.926 32.906 45.962 ;
      RECT 32.454 45.926 32.506 45.962 ;
      RECT 32.054 45.926 32.106 45.962 ;
      RECT 31.654 45.926 31.706 45.962 ;
      RECT 31.254 45.926 31.306 45.962 ;
      RECT 30.854 45.926 30.906 45.962 ;
      RECT 30.454 45.926 30.506 45.962 ;
      RECT 30.054 45.926 30.106 45.962 ;
      RECT 29.654 45.926 29.706 45.962 ;
      RECT 29.254 45.926 29.306 45.962 ;
      RECT 28.854 45.926 28.906 45.962 ;
      RECT 28.454 45.926 28.506 45.962 ;
      RECT 28.054 45.926 28.106 45.962 ;
      RECT 27.654 45.926 27.706 45.962 ;
      RECT 27.254 45.926 27.306 45.962 ;
      RECT 26.854 45.926 26.906 45.962 ;
      RECT 26.454 45.926 26.506 45.962 ;
      RECT 26.054 45.926 26.106 45.962 ;
      RECT 25.654 45.926 25.706 45.962 ;
      RECT 25.254 45.926 25.306 45.962 ;
      RECT 24.854 45.926 24.906 45.962 ;
      RECT 24.454 45.926 24.506 45.962 ;
      RECT 24.054 45.926 24.106 45.962 ;
      RECT 23.654 45.926 23.706 45.962 ;
      RECT 23.254 45.926 23.306 45.962 ;
      RECT 22.854 45.926 22.906 45.962 ;
      RECT 22.694 45.926 22.746 45.962 ;
      RECT 21.732 45.926 21.786 45.962 ;
      RECT 14.214 45.926 14.268 45.962 ;
      RECT 13.054 45.926 13.106 45.962 ;
      RECT 12.654 45.926 12.706 45.962 ;
      RECT 12.254 45.926 12.306 45.962 ;
      RECT 11.854 45.926 11.906 45.962 ;
      RECT 11.454 45.926 11.506 45.962 ;
      RECT 11.054 45.926 11.106 45.962 ;
      RECT 10.654 45.926 10.706 45.962 ;
      RECT 10.254 45.926 10.306 45.962 ;
      RECT 9.854 45.926 9.906 45.962 ;
      RECT 9.454 45.926 9.506 45.962 ;
      RECT 9.054 45.926 9.106 45.962 ;
      RECT 8.654 45.926 8.706 45.962 ;
      RECT 8.254 45.926 8.306 45.962 ;
      RECT 7.854 45.926 7.906 45.962 ;
      RECT 7.454 45.926 7.506 45.962 ;
      RECT 7.054 45.926 7.106 45.962 ;
      RECT 6.654 45.926 6.706 45.962 ;
      RECT 6.254 45.926 6.306 45.962 ;
      RECT 5.854 45.926 5.906 45.962 ;
      RECT 5.454 45.926 5.506 45.962 ;
      RECT 5.054 45.926 5.106 45.962 ;
      RECT 4.654 45.926 4.706 45.962 ;
      RECT 4.254 45.926 4.306 45.962 ;
      RECT 3.854 45.926 3.906 45.962 ;
      RECT 3.454 45.926 3.506 45.962 ;
      RECT 3.054 45.926 3.106 45.962 ;
      RECT 2.654 45.926 2.706 45.962 ;
      RECT 2.254 45.926 2.306 45.962 ;
      RECT 1.854 45.926 1.906 45.962 ;
      RECT 1.454 45.926 1.506 45.962 ;
      RECT 1.054 45.926 1.106 45.962 ;
      RECT 0.654 45.926 0.706 45.962 ;
      RECT 21.978 45.702 22.022 45.738 ;
      RECT 21.096 45.702 21.14 45.738 ;
      RECT 14.86 45.702 14.904 45.738 ;
      RECT 13.978 45.702 14.022 45.738 ;
      RECT 35.494 45.478 35.546 45.514 ;
      RECT 35.094 45.478 35.146 45.514 ;
      RECT 34.694 45.478 34.746 45.514 ;
      RECT 34.294 45.478 34.346 45.514 ;
      RECT 33.894 45.478 33.946 45.514 ;
      RECT 33.494 45.478 33.546 45.514 ;
      RECT 33.094 45.478 33.146 45.514 ;
      RECT 32.694 45.478 32.746 45.514 ;
      RECT 32.294 45.478 32.346 45.514 ;
      RECT 31.894 45.478 31.946 45.514 ;
      RECT 31.494 45.478 31.546 45.514 ;
      RECT 31.094 45.478 31.146 45.514 ;
      RECT 30.694 45.478 30.746 45.514 ;
      RECT 30.294 45.478 30.346 45.514 ;
      RECT 29.894 45.478 29.946 45.514 ;
      RECT 29.494 45.478 29.546 45.514 ;
      RECT 29.094 45.478 29.146 45.514 ;
      RECT 28.694 45.478 28.746 45.514 ;
      RECT 28.294 45.478 28.346 45.514 ;
      RECT 27.894 45.478 27.946 45.514 ;
      RECT 27.494 45.478 27.546 45.514 ;
      RECT 27.094 45.478 27.146 45.514 ;
      RECT 26.694 45.478 26.746 45.514 ;
      RECT 26.294 45.478 26.346 45.514 ;
      RECT 25.894 45.478 25.946 45.514 ;
      RECT 25.494 45.478 25.546 45.514 ;
      RECT 25.094 45.478 25.146 45.514 ;
      RECT 24.694 45.478 24.746 45.514 ;
      RECT 24.294 45.478 24.346 45.514 ;
      RECT 23.894 45.478 23.946 45.514 ;
      RECT 23.494 45.478 23.546 45.514 ;
      RECT 23.094 45.478 23.146 45.514 ;
      RECT 21.814 45.478 21.868 45.514 ;
      RECT 19.838 45.478 19.886 45.514 ;
      RECT 19.53 45.478 19.578 45.514 ;
      RECT 16.882 45.478 16.936 45.514 ;
      RECT 16.422 45.478 16.47 45.514 ;
      RECT 16.114 45.478 16.162 45.514 ;
      RECT 14.132 45.478 14.186 45.514 ;
      RECT 13.294 45.478 13.346 45.514 ;
      RECT 12.894 45.478 12.946 45.514 ;
      RECT 12.494 45.478 12.546 45.514 ;
      RECT 12.094 45.478 12.146 45.514 ;
      RECT 11.694 45.478 11.746 45.514 ;
      RECT 11.294 45.478 11.346 45.514 ;
      RECT 10.894 45.478 10.946 45.514 ;
      RECT 10.494 45.478 10.546 45.514 ;
      RECT 10.094 45.478 10.146 45.514 ;
      RECT 9.694 45.478 9.746 45.514 ;
      RECT 9.294 45.478 9.346 45.514 ;
      RECT 8.894 45.478 8.946 45.514 ;
      RECT 8.494 45.478 8.546 45.514 ;
      RECT 8.094 45.478 8.146 45.514 ;
      RECT 7.694 45.478 7.746 45.514 ;
      RECT 7.294 45.478 7.346 45.514 ;
      RECT 6.894 45.478 6.946 45.514 ;
      RECT 6.494 45.478 6.546 45.514 ;
      RECT 6.094 45.478 6.146 45.514 ;
      RECT 5.694 45.478 5.746 45.514 ;
      RECT 5.294 45.478 5.346 45.514 ;
      RECT 4.894 45.478 4.946 45.514 ;
      RECT 4.494 45.478 4.546 45.514 ;
      RECT 4.094 45.478 4.146 45.514 ;
      RECT 3.694 45.478 3.746 45.514 ;
      RECT 3.294 45.478 3.346 45.514 ;
      RECT 2.894 45.478 2.946 45.514 ;
      RECT 2.494 45.478 2.546 45.514 ;
      RECT 2.094 45.478 2.146 45.514 ;
      RECT 1.694 45.478 1.746 45.514 ;
      RECT 1.294 45.478 1.346 45.514 ;
      RECT 0.894 45.478 0.946 45.514 ;
      RECT 21.414 45.402 21.468 45.438 ;
      RECT 14.532 45.402 14.586 45.438 ;
      RECT 19.606 45.249 19.654 45.285 ;
      RECT 18.08 45.249 18.12 45.285 ;
      RECT 16.718 45.249 16.772 45.285 ;
      RECT 16.346 45.249 16.394 45.285 ;
      RECT 20.37 45.2545 20.442 45.2795 ;
      RECT 18.764 45.2545 18.836 45.2795 ;
      RECT 15.558 45.2545 15.63 45.2795 ;
      RECT 21.978 45.102 22.022 45.138 ;
      RECT 13.978 45.102 14.022 45.138 ;
      RECT 18.764 45.1075 18.836 45.1325 ;
      RECT 19.762 44.955 19.81 44.991 ;
      RECT 17.616 44.955 17.656 44.991 ;
      RECT 16.19 44.955 16.238 44.991 ;
      RECT 35.254 44.726 35.306 44.762 ;
      RECT 34.854 44.726 34.906 44.762 ;
      RECT 34.454 44.726 34.506 44.762 ;
      RECT 34.054 44.726 34.106 44.762 ;
      RECT 33.654 44.726 33.706 44.762 ;
      RECT 33.254 44.726 33.306 44.762 ;
      RECT 32.854 44.726 32.906 44.762 ;
      RECT 32.454 44.726 32.506 44.762 ;
      RECT 32.054 44.726 32.106 44.762 ;
      RECT 31.654 44.726 31.706 44.762 ;
      RECT 31.254 44.726 31.306 44.762 ;
      RECT 30.854 44.726 30.906 44.762 ;
      RECT 30.454 44.726 30.506 44.762 ;
      RECT 30.054 44.726 30.106 44.762 ;
      RECT 29.654 44.726 29.706 44.762 ;
      RECT 29.254 44.726 29.306 44.762 ;
      RECT 28.854 44.726 28.906 44.762 ;
      RECT 28.454 44.726 28.506 44.762 ;
      RECT 28.054 44.726 28.106 44.762 ;
      RECT 27.654 44.726 27.706 44.762 ;
      RECT 27.254 44.726 27.306 44.762 ;
      RECT 26.854 44.726 26.906 44.762 ;
      RECT 26.454 44.726 26.506 44.762 ;
      RECT 26.054 44.726 26.106 44.762 ;
      RECT 25.654 44.726 25.706 44.762 ;
      RECT 25.254 44.726 25.306 44.762 ;
      RECT 24.854 44.726 24.906 44.762 ;
      RECT 24.454 44.726 24.506 44.762 ;
      RECT 24.054 44.726 24.106 44.762 ;
      RECT 23.654 44.726 23.706 44.762 ;
      RECT 23.254 44.726 23.306 44.762 ;
      RECT 22.854 44.726 22.906 44.762 ;
      RECT 22.694 44.726 22.746 44.762 ;
      RECT 21.732 44.726 21.786 44.762 ;
      RECT 14.214 44.726 14.268 44.762 ;
      RECT 13.054 44.726 13.106 44.762 ;
      RECT 12.654 44.726 12.706 44.762 ;
      RECT 12.254 44.726 12.306 44.762 ;
      RECT 11.854 44.726 11.906 44.762 ;
      RECT 11.454 44.726 11.506 44.762 ;
      RECT 11.054 44.726 11.106 44.762 ;
      RECT 10.654 44.726 10.706 44.762 ;
      RECT 10.254 44.726 10.306 44.762 ;
      RECT 9.854 44.726 9.906 44.762 ;
      RECT 9.454 44.726 9.506 44.762 ;
      RECT 9.054 44.726 9.106 44.762 ;
      RECT 8.654 44.726 8.706 44.762 ;
      RECT 8.254 44.726 8.306 44.762 ;
      RECT 7.854 44.726 7.906 44.762 ;
      RECT 7.454 44.726 7.506 44.762 ;
      RECT 7.054 44.726 7.106 44.762 ;
      RECT 6.654 44.726 6.706 44.762 ;
      RECT 6.254 44.726 6.306 44.762 ;
      RECT 5.854 44.726 5.906 44.762 ;
      RECT 5.454 44.726 5.506 44.762 ;
      RECT 5.054 44.726 5.106 44.762 ;
      RECT 4.654 44.726 4.706 44.762 ;
      RECT 4.254 44.726 4.306 44.762 ;
      RECT 3.854 44.726 3.906 44.762 ;
      RECT 3.454 44.726 3.506 44.762 ;
      RECT 3.054 44.726 3.106 44.762 ;
      RECT 2.654 44.726 2.706 44.762 ;
      RECT 2.254 44.726 2.306 44.762 ;
      RECT 1.854 44.726 1.906 44.762 ;
      RECT 1.454 44.726 1.506 44.762 ;
      RECT 1.054 44.726 1.106 44.762 ;
      RECT 0.654 44.726 0.706 44.762 ;
      RECT 21.978 44.502 22.022 44.538 ;
      RECT 21.096 44.502 21.14 44.538 ;
      RECT 14.86 44.502 14.904 44.538 ;
      RECT 13.978 44.502 14.022 44.538 ;
      RECT 35.494 44.278 35.546 44.314 ;
      RECT 35.094 44.278 35.146 44.314 ;
      RECT 34.694 44.278 34.746 44.314 ;
      RECT 34.294 44.278 34.346 44.314 ;
      RECT 33.894 44.278 33.946 44.314 ;
      RECT 33.494 44.278 33.546 44.314 ;
      RECT 33.094 44.278 33.146 44.314 ;
      RECT 32.694 44.278 32.746 44.314 ;
      RECT 32.294 44.278 32.346 44.314 ;
      RECT 31.894 44.278 31.946 44.314 ;
      RECT 31.494 44.278 31.546 44.314 ;
      RECT 31.094 44.278 31.146 44.314 ;
      RECT 30.694 44.278 30.746 44.314 ;
      RECT 30.294 44.278 30.346 44.314 ;
      RECT 29.894 44.278 29.946 44.314 ;
      RECT 29.494 44.278 29.546 44.314 ;
      RECT 29.094 44.278 29.146 44.314 ;
      RECT 28.694 44.278 28.746 44.314 ;
      RECT 28.294 44.278 28.346 44.314 ;
      RECT 27.894 44.278 27.946 44.314 ;
      RECT 27.494 44.278 27.546 44.314 ;
      RECT 27.094 44.278 27.146 44.314 ;
      RECT 26.694 44.278 26.746 44.314 ;
      RECT 26.294 44.278 26.346 44.314 ;
      RECT 25.894 44.278 25.946 44.314 ;
      RECT 25.494 44.278 25.546 44.314 ;
      RECT 25.094 44.278 25.146 44.314 ;
      RECT 24.694 44.278 24.746 44.314 ;
      RECT 24.294 44.278 24.346 44.314 ;
      RECT 23.894 44.278 23.946 44.314 ;
      RECT 23.494 44.278 23.546 44.314 ;
      RECT 23.094 44.278 23.146 44.314 ;
      RECT 21.814 44.278 21.868 44.314 ;
      RECT 19.838 44.278 19.886 44.314 ;
      RECT 19.53 44.278 19.578 44.314 ;
      RECT 16.882 44.278 16.936 44.314 ;
      RECT 16.422 44.278 16.47 44.314 ;
      RECT 16.114 44.278 16.162 44.314 ;
      RECT 14.132 44.278 14.186 44.314 ;
      RECT 13.294 44.278 13.346 44.314 ;
      RECT 12.894 44.278 12.946 44.314 ;
      RECT 12.494 44.278 12.546 44.314 ;
      RECT 12.094 44.278 12.146 44.314 ;
      RECT 11.694 44.278 11.746 44.314 ;
      RECT 11.294 44.278 11.346 44.314 ;
      RECT 10.894 44.278 10.946 44.314 ;
      RECT 10.494 44.278 10.546 44.314 ;
      RECT 10.094 44.278 10.146 44.314 ;
      RECT 9.694 44.278 9.746 44.314 ;
      RECT 9.294 44.278 9.346 44.314 ;
      RECT 8.894 44.278 8.946 44.314 ;
      RECT 8.494 44.278 8.546 44.314 ;
      RECT 8.094 44.278 8.146 44.314 ;
      RECT 7.694 44.278 7.746 44.314 ;
      RECT 7.294 44.278 7.346 44.314 ;
      RECT 6.894 44.278 6.946 44.314 ;
      RECT 6.494 44.278 6.546 44.314 ;
      RECT 6.094 44.278 6.146 44.314 ;
      RECT 5.694 44.278 5.746 44.314 ;
      RECT 5.294 44.278 5.346 44.314 ;
      RECT 4.894 44.278 4.946 44.314 ;
      RECT 4.494 44.278 4.546 44.314 ;
      RECT 4.094 44.278 4.146 44.314 ;
      RECT 3.694 44.278 3.746 44.314 ;
      RECT 3.294 44.278 3.346 44.314 ;
      RECT 2.894 44.278 2.946 44.314 ;
      RECT 2.494 44.278 2.546 44.314 ;
      RECT 2.094 44.278 2.146 44.314 ;
      RECT 1.694 44.278 1.746 44.314 ;
      RECT 1.294 44.278 1.346 44.314 ;
      RECT 0.894 44.278 0.946 44.314 ;
      RECT 21.414 44.202 21.468 44.238 ;
      RECT 14.532 44.202 14.586 44.238 ;
      RECT 19.606 44.049 19.654 44.085 ;
      RECT 18.08 44.049 18.12 44.085 ;
      RECT 16.718 44.049 16.772 44.085 ;
      RECT 16.346 44.049 16.394 44.085 ;
      RECT 20.37 44.0545 20.442 44.0795 ;
      RECT 18.764 44.0545 18.836 44.0795 ;
      RECT 15.558 44.0545 15.63 44.0795 ;
      RECT 21.978 43.902 22.022 43.938 ;
      RECT 13.978 43.902 14.022 43.938 ;
      RECT 18.764 43.9075 18.836 43.9325 ;
      RECT 19.762 43.755 19.81 43.791 ;
      RECT 17.616 43.755 17.656 43.791 ;
      RECT 16.19 43.755 16.238 43.791 ;
      RECT 35.254 43.526 35.306 43.562 ;
      RECT 34.854 43.526 34.906 43.562 ;
      RECT 34.454 43.526 34.506 43.562 ;
      RECT 34.054 43.526 34.106 43.562 ;
      RECT 33.654 43.526 33.706 43.562 ;
      RECT 33.254 43.526 33.306 43.562 ;
      RECT 32.854 43.526 32.906 43.562 ;
      RECT 32.454 43.526 32.506 43.562 ;
      RECT 32.054 43.526 32.106 43.562 ;
      RECT 31.654 43.526 31.706 43.562 ;
      RECT 31.254 43.526 31.306 43.562 ;
      RECT 30.854 43.526 30.906 43.562 ;
      RECT 30.454 43.526 30.506 43.562 ;
      RECT 30.054 43.526 30.106 43.562 ;
      RECT 29.654 43.526 29.706 43.562 ;
      RECT 29.254 43.526 29.306 43.562 ;
      RECT 28.854 43.526 28.906 43.562 ;
      RECT 28.454 43.526 28.506 43.562 ;
      RECT 28.054 43.526 28.106 43.562 ;
      RECT 27.654 43.526 27.706 43.562 ;
      RECT 27.254 43.526 27.306 43.562 ;
      RECT 26.854 43.526 26.906 43.562 ;
      RECT 26.454 43.526 26.506 43.562 ;
      RECT 26.054 43.526 26.106 43.562 ;
      RECT 25.654 43.526 25.706 43.562 ;
      RECT 25.254 43.526 25.306 43.562 ;
      RECT 24.854 43.526 24.906 43.562 ;
      RECT 24.454 43.526 24.506 43.562 ;
      RECT 24.054 43.526 24.106 43.562 ;
      RECT 23.654 43.526 23.706 43.562 ;
      RECT 23.254 43.526 23.306 43.562 ;
      RECT 22.854 43.526 22.906 43.562 ;
      RECT 22.694 43.526 22.746 43.562 ;
      RECT 21.732 43.526 21.786 43.562 ;
      RECT 14.214 43.526 14.268 43.562 ;
      RECT 13.054 43.526 13.106 43.562 ;
      RECT 12.654 43.526 12.706 43.562 ;
      RECT 12.254 43.526 12.306 43.562 ;
      RECT 11.854 43.526 11.906 43.562 ;
      RECT 11.454 43.526 11.506 43.562 ;
      RECT 11.054 43.526 11.106 43.562 ;
      RECT 10.654 43.526 10.706 43.562 ;
      RECT 10.254 43.526 10.306 43.562 ;
      RECT 9.854 43.526 9.906 43.562 ;
      RECT 9.454 43.526 9.506 43.562 ;
      RECT 9.054 43.526 9.106 43.562 ;
      RECT 8.654 43.526 8.706 43.562 ;
      RECT 8.254 43.526 8.306 43.562 ;
      RECT 7.854 43.526 7.906 43.562 ;
      RECT 7.454 43.526 7.506 43.562 ;
      RECT 7.054 43.526 7.106 43.562 ;
      RECT 6.654 43.526 6.706 43.562 ;
      RECT 6.254 43.526 6.306 43.562 ;
      RECT 5.854 43.526 5.906 43.562 ;
      RECT 5.454 43.526 5.506 43.562 ;
      RECT 5.054 43.526 5.106 43.562 ;
      RECT 4.654 43.526 4.706 43.562 ;
      RECT 4.254 43.526 4.306 43.562 ;
      RECT 3.854 43.526 3.906 43.562 ;
      RECT 3.454 43.526 3.506 43.562 ;
      RECT 3.054 43.526 3.106 43.562 ;
      RECT 2.654 43.526 2.706 43.562 ;
      RECT 2.254 43.526 2.306 43.562 ;
      RECT 1.854 43.526 1.906 43.562 ;
      RECT 1.454 43.526 1.506 43.562 ;
      RECT 1.054 43.526 1.106 43.562 ;
      RECT 0.654 43.526 0.706 43.562 ;
      RECT 21.978 43.302 22.022 43.338 ;
      RECT 21.096 43.302 21.14 43.338 ;
      RECT 14.86 43.302 14.904 43.338 ;
      RECT 13.978 43.302 14.022 43.338 ;
      RECT 35.494 43.078 35.546 43.114 ;
      RECT 35.094 43.078 35.146 43.114 ;
      RECT 34.694 43.078 34.746 43.114 ;
      RECT 34.294 43.078 34.346 43.114 ;
      RECT 33.894 43.078 33.946 43.114 ;
      RECT 33.494 43.078 33.546 43.114 ;
      RECT 33.094 43.078 33.146 43.114 ;
      RECT 32.694 43.078 32.746 43.114 ;
      RECT 32.294 43.078 32.346 43.114 ;
      RECT 31.894 43.078 31.946 43.114 ;
      RECT 31.494 43.078 31.546 43.114 ;
      RECT 31.094 43.078 31.146 43.114 ;
      RECT 30.694 43.078 30.746 43.114 ;
      RECT 30.294 43.078 30.346 43.114 ;
      RECT 29.894 43.078 29.946 43.114 ;
      RECT 29.494 43.078 29.546 43.114 ;
      RECT 29.094 43.078 29.146 43.114 ;
      RECT 28.694 43.078 28.746 43.114 ;
      RECT 28.294 43.078 28.346 43.114 ;
      RECT 27.894 43.078 27.946 43.114 ;
      RECT 27.494 43.078 27.546 43.114 ;
      RECT 27.094 43.078 27.146 43.114 ;
      RECT 26.694 43.078 26.746 43.114 ;
      RECT 26.294 43.078 26.346 43.114 ;
      RECT 25.894 43.078 25.946 43.114 ;
      RECT 25.494 43.078 25.546 43.114 ;
      RECT 25.094 43.078 25.146 43.114 ;
      RECT 24.694 43.078 24.746 43.114 ;
      RECT 24.294 43.078 24.346 43.114 ;
      RECT 23.894 43.078 23.946 43.114 ;
      RECT 23.494 43.078 23.546 43.114 ;
      RECT 23.094 43.078 23.146 43.114 ;
      RECT 21.814 43.078 21.868 43.114 ;
      RECT 19.838 43.078 19.886 43.114 ;
      RECT 19.53 43.078 19.578 43.114 ;
      RECT 16.882 43.078 16.936 43.114 ;
      RECT 16.422 43.078 16.47 43.114 ;
      RECT 16.114 43.078 16.162 43.114 ;
      RECT 14.132 43.078 14.186 43.114 ;
      RECT 13.294 43.078 13.346 43.114 ;
      RECT 12.894 43.078 12.946 43.114 ;
      RECT 12.494 43.078 12.546 43.114 ;
      RECT 12.094 43.078 12.146 43.114 ;
      RECT 11.694 43.078 11.746 43.114 ;
      RECT 11.294 43.078 11.346 43.114 ;
      RECT 10.894 43.078 10.946 43.114 ;
      RECT 10.494 43.078 10.546 43.114 ;
      RECT 10.094 43.078 10.146 43.114 ;
      RECT 9.694 43.078 9.746 43.114 ;
      RECT 9.294 43.078 9.346 43.114 ;
      RECT 8.894 43.078 8.946 43.114 ;
      RECT 8.494 43.078 8.546 43.114 ;
      RECT 8.094 43.078 8.146 43.114 ;
      RECT 7.694 43.078 7.746 43.114 ;
      RECT 7.294 43.078 7.346 43.114 ;
      RECT 6.894 43.078 6.946 43.114 ;
      RECT 6.494 43.078 6.546 43.114 ;
      RECT 6.094 43.078 6.146 43.114 ;
      RECT 5.694 43.078 5.746 43.114 ;
      RECT 5.294 43.078 5.346 43.114 ;
      RECT 4.894 43.078 4.946 43.114 ;
      RECT 4.494 43.078 4.546 43.114 ;
      RECT 4.094 43.078 4.146 43.114 ;
      RECT 3.694 43.078 3.746 43.114 ;
      RECT 3.294 43.078 3.346 43.114 ;
      RECT 2.894 43.078 2.946 43.114 ;
      RECT 2.494 43.078 2.546 43.114 ;
      RECT 2.094 43.078 2.146 43.114 ;
      RECT 1.694 43.078 1.746 43.114 ;
      RECT 1.294 43.078 1.346 43.114 ;
      RECT 0.894 43.078 0.946 43.114 ;
      RECT 21.414 43.002 21.468 43.038 ;
      RECT 14.532 43.002 14.586 43.038 ;
      RECT 19.606 42.849 19.654 42.885 ;
      RECT 18.08 42.849 18.12 42.885 ;
      RECT 16.718 42.849 16.772 42.885 ;
      RECT 16.346 42.849 16.394 42.885 ;
      RECT 20.37 42.8545 20.442 42.8795 ;
      RECT 18.764 42.8545 18.836 42.8795 ;
      RECT 15.558 42.8545 15.63 42.8795 ;
      RECT 21.978 42.702 22.022 42.738 ;
      RECT 13.978 42.702 14.022 42.738 ;
      RECT 18.764 42.7075 18.836 42.7325 ;
      RECT 19.762 42.555 19.81 42.591 ;
      RECT 17.616 42.555 17.656 42.591 ;
      RECT 16.19 42.555 16.238 42.591 ;
      RECT 35.254 42.326 35.306 42.362 ;
      RECT 34.854 42.326 34.906 42.362 ;
      RECT 34.454 42.326 34.506 42.362 ;
      RECT 34.054 42.326 34.106 42.362 ;
      RECT 33.654 42.326 33.706 42.362 ;
      RECT 33.254 42.326 33.306 42.362 ;
      RECT 32.854 42.326 32.906 42.362 ;
      RECT 32.454 42.326 32.506 42.362 ;
      RECT 32.054 42.326 32.106 42.362 ;
      RECT 31.654 42.326 31.706 42.362 ;
      RECT 31.254 42.326 31.306 42.362 ;
      RECT 30.854 42.326 30.906 42.362 ;
      RECT 30.454 42.326 30.506 42.362 ;
      RECT 30.054 42.326 30.106 42.362 ;
      RECT 29.654 42.326 29.706 42.362 ;
      RECT 29.254 42.326 29.306 42.362 ;
      RECT 28.854 42.326 28.906 42.362 ;
      RECT 28.454 42.326 28.506 42.362 ;
      RECT 28.054 42.326 28.106 42.362 ;
      RECT 27.654 42.326 27.706 42.362 ;
      RECT 27.254 42.326 27.306 42.362 ;
      RECT 26.854 42.326 26.906 42.362 ;
      RECT 26.454 42.326 26.506 42.362 ;
      RECT 26.054 42.326 26.106 42.362 ;
      RECT 25.654 42.326 25.706 42.362 ;
      RECT 25.254 42.326 25.306 42.362 ;
      RECT 24.854 42.326 24.906 42.362 ;
      RECT 24.454 42.326 24.506 42.362 ;
      RECT 24.054 42.326 24.106 42.362 ;
      RECT 23.654 42.326 23.706 42.362 ;
      RECT 23.254 42.326 23.306 42.362 ;
      RECT 22.854 42.326 22.906 42.362 ;
      RECT 22.694 42.326 22.746 42.362 ;
      RECT 21.732 42.326 21.786 42.362 ;
      RECT 14.214 42.326 14.268 42.362 ;
      RECT 13.054 42.326 13.106 42.362 ;
      RECT 12.654 42.326 12.706 42.362 ;
      RECT 12.254 42.326 12.306 42.362 ;
      RECT 11.854 42.326 11.906 42.362 ;
      RECT 11.454 42.326 11.506 42.362 ;
      RECT 11.054 42.326 11.106 42.362 ;
      RECT 10.654 42.326 10.706 42.362 ;
      RECT 10.254 42.326 10.306 42.362 ;
      RECT 9.854 42.326 9.906 42.362 ;
      RECT 9.454 42.326 9.506 42.362 ;
      RECT 9.054 42.326 9.106 42.362 ;
      RECT 8.654 42.326 8.706 42.362 ;
      RECT 8.254 42.326 8.306 42.362 ;
      RECT 7.854 42.326 7.906 42.362 ;
      RECT 7.454 42.326 7.506 42.362 ;
      RECT 7.054 42.326 7.106 42.362 ;
      RECT 6.654 42.326 6.706 42.362 ;
      RECT 6.254 42.326 6.306 42.362 ;
      RECT 5.854 42.326 5.906 42.362 ;
      RECT 5.454 42.326 5.506 42.362 ;
      RECT 5.054 42.326 5.106 42.362 ;
      RECT 4.654 42.326 4.706 42.362 ;
      RECT 4.254 42.326 4.306 42.362 ;
      RECT 3.854 42.326 3.906 42.362 ;
      RECT 3.454 42.326 3.506 42.362 ;
      RECT 3.054 42.326 3.106 42.362 ;
      RECT 2.654 42.326 2.706 42.362 ;
      RECT 2.254 42.326 2.306 42.362 ;
      RECT 1.854 42.326 1.906 42.362 ;
      RECT 1.454 42.326 1.506 42.362 ;
      RECT 1.054 42.326 1.106 42.362 ;
      RECT 0.654 42.326 0.706 42.362 ;
      RECT 21.978 42.102 22.022 42.138 ;
      RECT 21.096 42.102 21.14 42.138 ;
      RECT 14.86 42.102 14.904 42.138 ;
      RECT 13.978 42.102 14.022 42.138 ;
      RECT 35.494 41.878 35.546 41.914 ;
      RECT 35.094 41.878 35.146 41.914 ;
      RECT 34.694 41.878 34.746 41.914 ;
      RECT 34.294 41.878 34.346 41.914 ;
      RECT 33.894 41.878 33.946 41.914 ;
      RECT 33.494 41.878 33.546 41.914 ;
      RECT 33.094 41.878 33.146 41.914 ;
      RECT 32.694 41.878 32.746 41.914 ;
      RECT 32.294 41.878 32.346 41.914 ;
      RECT 31.894 41.878 31.946 41.914 ;
      RECT 31.494 41.878 31.546 41.914 ;
      RECT 31.094 41.878 31.146 41.914 ;
      RECT 30.694 41.878 30.746 41.914 ;
      RECT 30.294 41.878 30.346 41.914 ;
      RECT 29.894 41.878 29.946 41.914 ;
      RECT 29.494 41.878 29.546 41.914 ;
      RECT 29.094 41.878 29.146 41.914 ;
      RECT 28.694 41.878 28.746 41.914 ;
      RECT 28.294 41.878 28.346 41.914 ;
      RECT 27.894 41.878 27.946 41.914 ;
      RECT 27.494 41.878 27.546 41.914 ;
      RECT 27.094 41.878 27.146 41.914 ;
      RECT 26.694 41.878 26.746 41.914 ;
      RECT 26.294 41.878 26.346 41.914 ;
      RECT 25.894 41.878 25.946 41.914 ;
      RECT 25.494 41.878 25.546 41.914 ;
      RECT 25.094 41.878 25.146 41.914 ;
      RECT 24.694 41.878 24.746 41.914 ;
      RECT 24.294 41.878 24.346 41.914 ;
      RECT 23.894 41.878 23.946 41.914 ;
      RECT 23.494 41.878 23.546 41.914 ;
      RECT 23.094 41.878 23.146 41.914 ;
      RECT 21.814 41.878 21.868 41.914 ;
      RECT 19.838 41.878 19.886 41.914 ;
      RECT 19.53 41.878 19.578 41.914 ;
      RECT 16.882 41.878 16.936 41.914 ;
      RECT 16.422 41.878 16.47 41.914 ;
      RECT 16.114 41.878 16.162 41.914 ;
      RECT 14.132 41.878 14.186 41.914 ;
      RECT 13.294 41.878 13.346 41.914 ;
      RECT 12.894 41.878 12.946 41.914 ;
      RECT 12.494 41.878 12.546 41.914 ;
      RECT 12.094 41.878 12.146 41.914 ;
      RECT 11.694 41.878 11.746 41.914 ;
      RECT 11.294 41.878 11.346 41.914 ;
      RECT 10.894 41.878 10.946 41.914 ;
      RECT 10.494 41.878 10.546 41.914 ;
      RECT 10.094 41.878 10.146 41.914 ;
      RECT 9.694 41.878 9.746 41.914 ;
      RECT 9.294 41.878 9.346 41.914 ;
      RECT 8.894 41.878 8.946 41.914 ;
      RECT 8.494 41.878 8.546 41.914 ;
      RECT 8.094 41.878 8.146 41.914 ;
      RECT 7.694 41.878 7.746 41.914 ;
      RECT 7.294 41.878 7.346 41.914 ;
      RECT 6.894 41.878 6.946 41.914 ;
      RECT 6.494 41.878 6.546 41.914 ;
      RECT 6.094 41.878 6.146 41.914 ;
      RECT 5.694 41.878 5.746 41.914 ;
      RECT 5.294 41.878 5.346 41.914 ;
      RECT 4.894 41.878 4.946 41.914 ;
      RECT 4.494 41.878 4.546 41.914 ;
      RECT 4.094 41.878 4.146 41.914 ;
      RECT 3.694 41.878 3.746 41.914 ;
      RECT 3.294 41.878 3.346 41.914 ;
      RECT 2.894 41.878 2.946 41.914 ;
      RECT 2.494 41.878 2.546 41.914 ;
      RECT 2.094 41.878 2.146 41.914 ;
      RECT 1.694 41.878 1.746 41.914 ;
      RECT 1.294 41.878 1.346 41.914 ;
      RECT 0.894 41.878 0.946 41.914 ;
      RECT 21.414 41.802 21.468 41.838 ;
      RECT 14.532 41.802 14.586 41.838 ;
      RECT 19.606 41.649 19.654 41.685 ;
      RECT 18.08 41.649 18.12 41.685 ;
      RECT 16.718 41.649 16.772 41.685 ;
      RECT 16.346 41.649 16.394 41.685 ;
      RECT 20.37 41.6545 20.442 41.6795 ;
      RECT 18.764 41.6545 18.836 41.6795 ;
      RECT 15.558 41.6545 15.63 41.6795 ;
      RECT 21.978 41.502 22.022 41.538 ;
      RECT 13.978 41.502 14.022 41.538 ;
      RECT 18.764 41.5075 18.836 41.5325 ;
      RECT 19.762 41.355 19.81 41.391 ;
      RECT 17.616 41.355 17.656 41.391 ;
      RECT 16.19 41.355 16.238 41.391 ;
      RECT 35.254 41.126 35.306 41.162 ;
      RECT 34.854 41.126 34.906 41.162 ;
      RECT 34.454 41.126 34.506 41.162 ;
      RECT 34.054 41.126 34.106 41.162 ;
      RECT 33.654 41.126 33.706 41.162 ;
      RECT 33.254 41.126 33.306 41.162 ;
      RECT 32.854 41.126 32.906 41.162 ;
      RECT 32.454 41.126 32.506 41.162 ;
      RECT 32.054 41.126 32.106 41.162 ;
      RECT 31.654 41.126 31.706 41.162 ;
      RECT 31.254 41.126 31.306 41.162 ;
      RECT 30.854 41.126 30.906 41.162 ;
      RECT 30.454 41.126 30.506 41.162 ;
      RECT 30.054 41.126 30.106 41.162 ;
      RECT 29.654 41.126 29.706 41.162 ;
      RECT 29.254 41.126 29.306 41.162 ;
      RECT 28.854 41.126 28.906 41.162 ;
      RECT 28.454 41.126 28.506 41.162 ;
      RECT 28.054 41.126 28.106 41.162 ;
      RECT 27.654 41.126 27.706 41.162 ;
      RECT 27.254 41.126 27.306 41.162 ;
      RECT 26.854 41.126 26.906 41.162 ;
      RECT 26.454 41.126 26.506 41.162 ;
      RECT 26.054 41.126 26.106 41.162 ;
      RECT 25.654 41.126 25.706 41.162 ;
      RECT 25.254 41.126 25.306 41.162 ;
      RECT 24.854 41.126 24.906 41.162 ;
      RECT 24.454 41.126 24.506 41.162 ;
      RECT 24.054 41.126 24.106 41.162 ;
      RECT 23.654 41.126 23.706 41.162 ;
      RECT 23.254 41.126 23.306 41.162 ;
      RECT 22.854 41.126 22.906 41.162 ;
      RECT 22.694 41.126 22.746 41.162 ;
      RECT 21.732 41.126 21.786 41.162 ;
      RECT 14.214 41.126 14.268 41.162 ;
      RECT 13.054 41.126 13.106 41.162 ;
      RECT 12.654 41.126 12.706 41.162 ;
      RECT 12.254 41.126 12.306 41.162 ;
      RECT 11.854 41.126 11.906 41.162 ;
      RECT 11.454 41.126 11.506 41.162 ;
      RECT 11.054 41.126 11.106 41.162 ;
      RECT 10.654 41.126 10.706 41.162 ;
      RECT 10.254 41.126 10.306 41.162 ;
      RECT 9.854 41.126 9.906 41.162 ;
      RECT 9.454 41.126 9.506 41.162 ;
      RECT 9.054 41.126 9.106 41.162 ;
      RECT 8.654 41.126 8.706 41.162 ;
      RECT 8.254 41.126 8.306 41.162 ;
      RECT 7.854 41.126 7.906 41.162 ;
      RECT 7.454 41.126 7.506 41.162 ;
      RECT 7.054 41.126 7.106 41.162 ;
      RECT 6.654 41.126 6.706 41.162 ;
      RECT 6.254 41.126 6.306 41.162 ;
      RECT 5.854 41.126 5.906 41.162 ;
      RECT 5.454 41.126 5.506 41.162 ;
      RECT 5.054 41.126 5.106 41.162 ;
      RECT 4.654 41.126 4.706 41.162 ;
      RECT 4.254 41.126 4.306 41.162 ;
      RECT 3.854 41.126 3.906 41.162 ;
      RECT 3.454 41.126 3.506 41.162 ;
      RECT 3.054 41.126 3.106 41.162 ;
      RECT 2.654 41.126 2.706 41.162 ;
      RECT 2.254 41.126 2.306 41.162 ;
      RECT 1.854 41.126 1.906 41.162 ;
      RECT 1.454 41.126 1.506 41.162 ;
      RECT 1.054 41.126 1.106 41.162 ;
      RECT 0.654 41.126 0.706 41.162 ;
      RECT 21.978 40.902 22.022 40.938 ;
      RECT 21.096 40.902 21.14 40.938 ;
      RECT 14.86 40.902 14.904 40.938 ;
      RECT 13.978 40.902 14.022 40.938 ;
      RECT 35.494 40.678 35.546 40.714 ;
      RECT 35.094 40.678 35.146 40.714 ;
      RECT 34.694 40.678 34.746 40.714 ;
      RECT 34.294 40.678 34.346 40.714 ;
      RECT 33.894 40.678 33.946 40.714 ;
      RECT 33.494 40.678 33.546 40.714 ;
      RECT 33.094 40.678 33.146 40.714 ;
      RECT 32.694 40.678 32.746 40.714 ;
      RECT 32.294 40.678 32.346 40.714 ;
      RECT 31.894 40.678 31.946 40.714 ;
      RECT 31.494 40.678 31.546 40.714 ;
      RECT 31.094 40.678 31.146 40.714 ;
      RECT 30.694 40.678 30.746 40.714 ;
      RECT 30.294 40.678 30.346 40.714 ;
      RECT 29.894 40.678 29.946 40.714 ;
      RECT 29.494 40.678 29.546 40.714 ;
      RECT 29.094 40.678 29.146 40.714 ;
      RECT 28.694 40.678 28.746 40.714 ;
      RECT 28.294 40.678 28.346 40.714 ;
      RECT 27.894 40.678 27.946 40.714 ;
      RECT 27.494 40.678 27.546 40.714 ;
      RECT 27.094 40.678 27.146 40.714 ;
      RECT 26.694 40.678 26.746 40.714 ;
      RECT 26.294 40.678 26.346 40.714 ;
      RECT 25.894 40.678 25.946 40.714 ;
      RECT 25.494 40.678 25.546 40.714 ;
      RECT 25.094 40.678 25.146 40.714 ;
      RECT 24.694 40.678 24.746 40.714 ;
      RECT 24.294 40.678 24.346 40.714 ;
      RECT 23.894 40.678 23.946 40.714 ;
      RECT 23.494 40.678 23.546 40.714 ;
      RECT 23.094 40.678 23.146 40.714 ;
      RECT 21.814 40.678 21.868 40.714 ;
      RECT 19.838 40.678 19.886 40.714 ;
      RECT 19.53 40.678 19.578 40.714 ;
      RECT 16.882 40.678 16.936 40.714 ;
      RECT 16.422 40.678 16.47 40.714 ;
      RECT 16.114 40.678 16.162 40.714 ;
      RECT 14.132 40.678 14.186 40.714 ;
      RECT 13.294 40.678 13.346 40.714 ;
      RECT 12.894 40.678 12.946 40.714 ;
      RECT 12.494 40.678 12.546 40.714 ;
      RECT 12.094 40.678 12.146 40.714 ;
      RECT 11.694 40.678 11.746 40.714 ;
      RECT 11.294 40.678 11.346 40.714 ;
      RECT 10.894 40.678 10.946 40.714 ;
      RECT 10.494 40.678 10.546 40.714 ;
      RECT 10.094 40.678 10.146 40.714 ;
      RECT 9.694 40.678 9.746 40.714 ;
      RECT 9.294 40.678 9.346 40.714 ;
      RECT 8.894 40.678 8.946 40.714 ;
      RECT 8.494 40.678 8.546 40.714 ;
      RECT 8.094 40.678 8.146 40.714 ;
      RECT 7.694 40.678 7.746 40.714 ;
      RECT 7.294 40.678 7.346 40.714 ;
      RECT 6.894 40.678 6.946 40.714 ;
      RECT 6.494 40.678 6.546 40.714 ;
      RECT 6.094 40.678 6.146 40.714 ;
      RECT 5.694 40.678 5.746 40.714 ;
      RECT 5.294 40.678 5.346 40.714 ;
      RECT 4.894 40.678 4.946 40.714 ;
      RECT 4.494 40.678 4.546 40.714 ;
      RECT 4.094 40.678 4.146 40.714 ;
      RECT 3.694 40.678 3.746 40.714 ;
      RECT 3.294 40.678 3.346 40.714 ;
      RECT 2.894 40.678 2.946 40.714 ;
      RECT 2.494 40.678 2.546 40.714 ;
      RECT 2.094 40.678 2.146 40.714 ;
      RECT 1.694 40.678 1.746 40.714 ;
      RECT 1.294 40.678 1.346 40.714 ;
      RECT 0.894 40.678 0.946 40.714 ;
      RECT 21.414 40.602 21.468 40.638 ;
      RECT 14.532 40.602 14.586 40.638 ;
      RECT 19.606 40.449 19.654 40.485 ;
      RECT 18.08 40.449 18.12 40.485 ;
      RECT 16.718 40.449 16.772 40.485 ;
      RECT 16.346 40.449 16.394 40.485 ;
      RECT 20.37 40.4545 20.442 40.4795 ;
      RECT 18.764 40.4545 18.836 40.4795 ;
      RECT 15.558 40.4545 15.63 40.4795 ;
      RECT 21.978 40.302 22.022 40.338 ;
      RECT 13.978 40.302 14.022 40.338 ;
      RECT 18.764 40.3075 18.836 40.3325 ;
      RECT 19.762 40.155 19.81 40.191 ;
      RECT 17.616 40.155 17.656 40.191 ;
      RECT 16.19 40.155 16.238 40.191 ;
      RECT 35.254 39.926 35.306 39.962 ;
      RECT 34.854 39.926 34.906 39.962 ;
      RECT 34.454 39.926 34.506 39.962 ;
      RECT 34.054 39.926 34.106 39.962 ;
      RECT 33.654 39.926 33.706 39.962 ;
      RECT 33.254 39.926 33.306 39.962 ;
      RECT 32.854 39.926 32.906 39.962 ;
      RECT 32.454 39.926 32.506 39.962 ;
      RECT 32.054 39.926 32.106 39.962 ;
      RECT 31.654 39.926 31.706 39.962 ;
      RECT 31.254 39.926 31.306 39.962 ;
      RECT 30.854 39.926 30.906 39.962 ;
      RECT 30.454 39.926 30.506 39.962 ;
      RECT 30.054 39.926 30.106 39.962 ;
      RECT 29.654 39.926 29.706 39.962 ;
      RECT 29.254 39.926 29.306 39.962 ;
      RECT 28.854 39.926 28.906 39.962 ;
      RECT 28.454 39.926 28.506 39.962 ;
      RECT 28.054 39.926 28.106 39.962 ;
      RECT 27.654 39.926 27.706 39.962 ;
      RECT 27.254 39.926 27.306 39.962 ;
      RECT 26.854 39.926 26.906 39.962 ;
      RECT 26.454 39.926 26.506 39.962 ;
      RECT 26.054 39.926 26.106 39.962 ;
      RECT 25.654 39.926 25.706 39.962 ;
      RECT 25.254 39.926 25.306 39.962 ;
      RECT 24.854 39.926 24.906 39.962 ;
      RECT 24.454 39.926 24.506 39.962 ;
      RECT 24.054 39.926 24.106 39.962 ;
      RECT 23.654 39.926 23.706 39.962 ;
      RECT 23.254 39.926 23.306 39.962 ;
      RECT 22.854 39.926 22.906 39.962 ;
      RECT 22.694 39.926 22.746 39.962 ;
      RECT 21.732 39.926 21.786 39.962 ;
      RECT 14.214 39.926 14.268 39.962 ;
      RECT 13.054 39.926 13.106 39.962 ;
      RECT 12.654 39.926 12.706 39.962 ;
      RECT 12.254 39.926 12.306 39.962 ;
      RECT 11.854 39.926 11.906 39.962 ;
      RECT 11.454 39.926 11.506 39.962 ;
      RECT 11.054 39.926 11.106 39.962 ;
      RECT 10.654 39.926 10.706 39.962 ;
      RECT 10.254 39.926 10.306 39.962 ;
      RECT 9.854 39.926 9.906 39.962 ;
      RECT 9.454 39.926 9.506 39.962 ;
      RECT 9.054 39.926 9.106 39.962 ;
      RECT 8.654 39.926 8.706 39.962 ;
      RECT 8.254 39.926 8.306 39.962 ;
      RECT 7.854 39.926 7.906 39.962 ;
      RECT 7.454 39.926 7.506 39.962 ;
      RECT 7.054 39.926 7.106 39.962 ;
      RECT 6.654 39.926 6.706 39.962 ;
      RECT 6.254 39.926 6.306 39.962 ;
      RECT 5.854 39.926 5.906 39.962 ;
      RECT 5.454 39.926 5.506 39.962 ;
      RECT 5.054 39.926 5.106 39.962 ;
      RECT 4.654 39.926 4.706 39.962 ;
      RECT 4.254 39.926 4.306 39.962 ;
      RECT 3.854 39.926 3.906 39.962 ;
      RECT 3.454 39.926 3.506 39.962 ;
      RECT 3.054 39.926 3.106 39.962 ;
      RECT 2.654 39.926 2.706 39.962 ;
      RECT 2.254 39.926 2.306 39.962 ;
      RECT 1.854 39.926 1.906 39.962 ;
      RECT 1.454 39.926 1.506 39.962 ;
      RECT 1.054 39.926 1.106 39.962 ;
      RECT 0.654 39.926 0.706 39.962 ;
      RECT 21.978 39.702 22.022 39.738 ;
      RECT 21.096 39.702 21.14 39.738 ;
      RECT 14.86 39.702 14.904 39.738 ;
      RECT 13.978 39.702 14.022 39.738 ;
      RECT 21.978 39.342 22.022 39.378 ;
      RECT 21.096 39.342 21.14 39.378 ;
      RECT 14.86 39.342 14.904 39.378 ;
      RECT 13.978 39.342 14.022 39.378 ;
      RECT 16.882 39.2835 16.936 39.3195 ;
      RECT 16.718 39.2835 16.772 39.3195 ;
      RECT 21.414 39.222 21.468 39.258 ;
      RECT 14.532 39.222 14.586 39.258 ;
      RECT 20.37 39.2275 20.442 39.2525 ;
      RECT 15.558 39.2275 15.63 39.2525 ;
      RECT 21.414 38.982 21.468 39.018 ;
      RECT 19.606 38.982 19.654 39.018 ;
      RECT 18.08 38.982 18.12 39.018 ;
      RECT 17.616 38.982 17.656 39.018 ;
      RECT 16.346 38.982 16.394 39.018 ;
      RECT 14.532 38.982 14.586 39.018 ;
      RECT 19.838 38.9205 19.886 38.9565 ;
      RECT 16.114 38.9205 16.162 38.9565 ;
      RECT 35.254 38.862 35.306 38.898 ;
      RECT 34.854 38.862 34.906 38.898 ;
      RECT 34.454 38.862 34.506 38.898 ;
      RECT 34.054 38.862 34.106 38.898 ;
      RECT 33.654 38.862 33.706 38.898 ;
      RECT 33.254 38.862 33.306 38.898 ;
      RECT 32.854 38.862 32.906 38.898 ;
      RECT 32.454 38.862 32.506 38.898 ;
      RECT 32.054 38.862 32.106 38.898 ;
      RECT 31.654 38.862 31.706 38.898 ;
      RECT 31.254 38.862 31.306 38.898 ;
      RECT 30.854 38.862 30.906 38.898 ;
      RECT 30.454 38.862 30.506 38.898 ;
      RECT 30.054 38.862 30.106 38.898 ;
      RECT 29.654 38.862 29.706 38.898 ;
      RECT 29.254 38.862 29.306 38.898 ;
      RECT 28.854 38.862 28.906 38.898 ;
      RECT 28.454 38.862 28.506 38.898 ;
      RECT 28.054 38.862 28.106 38.898 ;
      RECT 27.654 38.862 27.706 38.898 ;
      RECT 27.254 38.862 27.306 38.898 ;
      RECT 26.854 38.862 26.906 38.898 ;
      RECT 26.454 38.862 26.506 38.898 ;
      RECT 26.054 38.862 26.106 38.898 ;
      RECT 25.654 38.862 25.706 38.898 ;
      RECT 25.254 38.862 25.306 38.898 ;
      RECT 24.854 38.862 24.906 38.898 ;
      RECT 24.454 38.862 24.506 38.898 ;
      RECT 24.054 38.862 24.106 38.898 ;
      RECT 23.654 38.862 23.706 38.898 ;
      RECT 23.254 38.862 23.306 38.898 ;
      RECT 22.854 38.862 22.906 38.898 ;
      RECT 21.978 38.862 22.022 38.898 ;
      RECT 21.096 38.862 21.14 38.898 ;
      RECT 14.86 38.862 14.904 38.898 ;
      RECT 13.978 38.862 14.022 38.898 ;
      RECT 13.054 38.862 13.106 38.898 ;
      RECT 12.654 38.862 12.706 38.898 ;
      RECT 12.254 38.862 12.306 38.898 ;
      RECT 11.854 38.862 11.906 38.898 ;
      RECT 11.454 38.862 11.506 38.898 ;
      RECT 11.054 38.862 11.106 38.898 ;
      RECT 10.654 38.862 10.706 38.898 ;
      RECT 10.254 38.862 10.306 38.898 ;
      RECT 9.854 38.862 9.906 38.898 ;
      RECT 9.454 38.862 9.506 38.898 ;
      RECT 9.054 38.862 9.106 38.898 ;
      RECT 8.654 38.862 8.706 38.898 ;
      RECT 8.254 38.862 8.306 38.898 ;
      RECT 7.854 38.862 7.906 38.898 ;
      RECT 7.454 38.862 7.506 38.898 ;
      RECT 7.054 38.862 7.106 38.898 ;
      RECT 6.654 38.862 6.706 38.898 ;
      RECT 6.254 38.862 6.306 38.898 ;
      RECT 5.854 38.862 5.906 38.898 ;
      RECT 5.454 38.862 5.506 38.898 ;
      RECT 5.054 38.862 5.106 38.898 ;
      RECT 4.654 38.862 4.706 38.898 ;
      RECT 4.254 38.862 4.306 38.898 ;
      RECT 3.854 38.862 3.906 38.898 ;
      RECT 3.454 38.862 3.506 38.898 ;
      RECT 3.054 38.862 3.106 38.898 ;
      RECT 2.654 38.862 2.706 38.898 ;
      RECT 2.254 38.862 2.306 38.898 ;
      RECT 1.854 38.862 1.906 38.898 ;
      RECT 1.454 38.862 1.506 38.898 ;
      RECT 1.054 38.862 1.106 38.898 ;
      RECT 0.654 38.862 0.706 38.898 ;
      RECT 19.762 38.742 19.81 38.778 ;
      RECT 16.19 38.742 16.238 38.778 ;
      RECT 19.53 38.6805 19.578 38.7165 ;
      RECT 16.422 38.6805 16.47 38.7165 ;
      RECT 35.254 38.622 35.306 38.658 ;
      RECT 34.854 38.622 34.906 38.658 ;
      RECT 34.454 38.622 34.506 38.658 ;
      RECT 34.054 38.622 34.106 38.658 ;
      RECT 33.654 38.622 33.706 38.658 ;
      RECT 33.254 38.622 33.306 38.658 ;
      RECT 32.854 38.622 32.906 38.658 ;
      RECT 32.454 38.622 32.506 38.658 ;
      RECT 32.054 38.622 32.106 38.658 ;
      RECT 31.654 38.622 31.706 38.658 ;
      RECT 31.254 38.622 31.306 38.658 ;
      RECT 30.854 38.622 30.906 38.658 ;
      RECT 30.454 38.622 30.506 38.658 ;
      RECT 30.054 38.622 30.106 38.658 ;
      RECT 29.654 38.622 29.706 38.658 ;
      RECT 29.254 38.622 29.306 38.658 ;
      RECT 28.854 38.622 28.906 38.658 ;
      RECT 28.454 38.622 28.506 38.658 ;
      RECT 28.054 38.622 28.106 38.658 ;
      RECT 27.654 38.622 27.706 38.658 ;
      RECT 27.254 38.622 27.306 38.658 ;
      RECT 26.854 38.622 26.906 38.658 ;
      RECT 26.454 38.622 26.506 38.658 ;
      RECT 26.054 38.622 26.106 38.658 ;
      RECT 25.654 38.622 25.706 38.658 ;
      RECT 25.254 38.622 25.306 38.658 ;
      RECT 24.854 38.622 24.906 38.658 ;
      RECT 24.454 38.622 24.506 38.658 ;
      RECT 24.054 38.622 24.106 38.658 ;
      RECT 23.654 38.622 23.706 38.658 ;
      RECT 23.254 38.622 23.306 38.658 ;
      RECT 22.854 38.622 22.906 38.658 ;
      RECT 13.054 38.622 13.106 38.658 ;
      RECT 12.654 38.622 12.706 38.658 ;
      RECT 12.254 38.622 12.306 38.658 ;
      RECT 11.854 38.622 11.906 38.658 ;
      RECT 11.454 38.622 11.506 38.658 ;
      RECT 11.054 38.622 11.106 38.658 ;
      RECT 10.654 38.622 10.706 38.658 ;
      RECT 10.254 38.622 10.306 38.658 ;
      RECT 9.854 38.622 9.906 38.658 ;
      RECT 9.454 38.622 9.506 38.658 ;
      RECT 9.054 38.622 9.106 38.658 ;
      RECT 8.654 38.622 8.706 38.658 ;
      RECT 8.254 38.622 8.306 38.658 ;
      RECT 7.854 38.622 7.906 38.658 ;
      RECT 7.454 38.622 7.506 38.658 ;
      RECT 7.054 38.622 7.106 38.658 ;
      RECT 6.654 38.622 6.706 38.658 ;
      RECT 6.254 38.622 6.306 38.658 ;
      RECT 5.854 38.622 5.906 38.658 ;
      RECT 5.454 38.622 5.506 38.658 ;
      RECT 5.054 38.622 5.106 38.658 ;
      RECT 4.654 38.622 4.706 38.658 ;
      RECT 4.254 38.622 4.306 38.658 ;
      RECT 3.854 38.622 3.906 38.658 ;
      RECT 3.454 38.622 3.506 38.658 ;
      RECT 3.054 38.622 3.106 38.658 ;
      RECT 2.654 38.622 2.706 38.658 ;
      RECT 2.254 38.622 2.306 38.658 ;
      RECT 1.854 38.622 1.906 38.658 ;
      RECT 1.454 38.622 1.506 38.658 ;
      RECT 1.054 38.622 1.106 38.658 ;
      RECT 0.654 38.622 0.706 38.658 ;
      RECT 19.762 38.4405 19.81 38.4765 ;
      RECT 16.19 38.4405 16.238 38.4765 ;
      RECT 21.978 38.382 22.022 38.418 ;
      RECT 21.096 38.382 21.14 38.418 ;
      RECT 14.86 38.382 14.904 38.418 ;
      RECT 13.978 38.382 14.022 38.418 ;
      RECT 20.222 38.262 20.262 38.298 ;
      RECT 19.606 38.262 19.654 38.298 ;
      RECT 16.346 38.262 16.394 38.298 ;
      RECT 15.738 38.262 15.778 38.298 ;
      RECT 35.494 38.142 35.546 38.178 ;
      RECT 35.094 38.142 35.146 38.178 ;
      RECT 34.934 38.142 34.986 38.178 ;
      RECT 34.694 38.142 34.746 38.178 ;
      RECT 34.294 38.142 34.346 38.178 ;
      RECT 34.134 38.142 34.186 38.178 ;
      RECT 33.894 38.142 33.946 38.178 ;
      RECT 33.494 38.142 33.546 38.178 ;
      RECT 33.334 38.142 33.386 38.178 ;
      RECT 33.094 38.142 33.146 38.178 ;
      RECT 32.694 38.142 32.746 38.178 ;
      RECT 32.534 38.142 32.586 38.178 ;
      RECT 32.294 38.142 32.346 38.178 ;
      RECT 31.894 38.142 31.946 38.178 ;
      RECT 31.734 38.142 31.786 38.178 ;
      RECT 31.494 38.142 31.546 38.178 ;
      RECT 31.094 38.142 31.146 38.178 ;
      RECT 30.934 38.142 30.986 38.178 ;
      RECT 30.694 38.142 30.746 38.178 ;
      RECT 30.294 38.142 30.346 38.178 ;
      RECT 30.134 38.142 30.186 38.178 ;
      RECT 29.894 38.142 29.946 38.178 ;
      RECT 29.494 38.142 29.546 38.178 ;
      RECT 29.334 38.142 29.386 38.178 ;
      RECT 29.094 38.142 29.146 38.178 ;
      RECT 28.694 38.142 28.746 38.178 ;
      RECT 28.534 38.142 28.586 38.178 ;
      RECT 28.294 38.142 28.346 38.178 ;
      RECT 27.894 38.142 27.946 38.178 ;
      RECT 27.734 38.142 27.786 38.178 ;
      RECT 27.494 38.142 27.546 38.178 ;
      RECT 27.094 38.142 27.146 38.178 ;
      RECT 26.934 38.142 26.986 38.178 ;
      RECT 26.694 38.142 26.746 38.178 ;
      RECT 26.294 38.142 26.346 38.178 ;
      RECT 26.134 38.142 26.186 38.178 ;
      RECT 25.894 38.142 25.946 38.178 ;
      RECT 25.494 38.142 25.546 38.178 ;
      RECT 25.334 38.142 25.386 38.178 ;
      RECT 25.094 38.142 25.146 38.178 ;
      RECT 24.694 38.142 24.746 38.178 ;
      RECT 24.534 38.142 24.586 38.178 ;
      RECT 24.294 38.142 24.346 38.178 ;
      RECT 23.894 38.142 23.946 38.178 ;
      RECT 23.734 38.142 23.786 38.178 ;
      RECT 23.494 38.142 23.546 38.178 ;
      RECT 23.094 38.142 23.146 38.178 ;
      RECT 22.934 38.142 22.986 38.178 ;
      RECT 22.694 38.142 22.746 38.178 ;
      RECT 13.294 38.142 13.346 38.178 ;
      RECT 12.894 38.142 12.946 38.178 ;
      RECT 12.734 38.142 12.786 38.178 ;
      RECT 12.494 38.142 12.546 38.178 ;
      RECT 12.094 38.142 12.146 38.178 ;
      RECT 11.934 38.142 11.986 38.178 ;
      RECT 11.694 38.142 11.746 38.178 ;
      RECT 11.294 38.142 11.346 38.178 ;
      RECT 11.134 38.142 11.186 38.178 ;
      RECT 10.894 38.142 10.946 38.178 ;
      RECT 10.494 38.142 10.546 38.178 ;
      RECT 10.334 38.142 10.386 38.178 ;
      RECT 10.094 38.142 10.146 38.178 ;
      RECT 9.694 38.142 9.746 38.178 ;
      RECT 9.534 38.142 9.586 38.178 ;
      RECT 9.294 38.142 9.346 38.178 ;
      RECT 8.894 38.142 8.946 38.178 ;
      RECT 8.734 38.142 8.786 38.178 ;
      RECT 8.494 38.142 8.546 38.178 ;
      RECT 8.094 38.142 8.146 38.178 ;
      RECT 7.934 38.142 7.986 38.178 ;
      RECT 7.694 38.142 7.746 38.178 ;
      RECT 7.294 38.142 7.346 38.178 ;
      RECT 7.134 38.142 7.186 38.178 ;
      RECT 6.894 38.142 6.946 38.178 ;
      RECT 6.494 38.142 6.546 38.178 ;
      RECT 6.334 38.142 6.386 38.178 ;
      RECT 6.094 38.142 6.146 38.178 ;
      RECT 5.694 38.142 5.746 38.178 ;
      RECT 5.534 38.142 5.586 38.178 ;
      RECT 5.294 38.142 5.346 38.178 ;
      RECT 4.894 38.142 4.946 38.178 ;
      RECT 4.734 38.142 4.786 38.178 ;
      RECT 4.494 38.142 4.546 38.178 ;
      RECT 4.094 38.142 4.146 38.178 ;
      RECT 3.934 38.142 3.986 38.178 ;
      RECT 3.694 38.142 3.746 38.178 ;
      RECT 3.294 38.142 3.346 38.178 ;
      RECT 3.134 38.142 3.186 38.178 ;
      RECT 2.894 38.142 2.946 38.178 ;
      RECT 2.494 38.142 2.546 38.178 ;
      RECT 2.334 38.142 2.386 38.178 ;
      RECT 2.094 38.142 2.146 38.178 ;
      RECT 1.694 38.142 1.746 38.178 ;
      RECT 1.534 38.142 1.586 38.178 ;
      RECT 1.294 38.142 1.346 38.178 ;
      RECT 0.894 38.142 0.946 38.178 ;
      RECT 0.734 38.142 0.786 38.178 ;
      RECT 35.494 37.902 35.546 37.938 ;
      RECT 35.094 37.902 35.146 37.938 ;
      RECT 34.934 37.902 34.986 37.938 ;
      RECT 34.694 37.902 34.746 37.938 ;
      RECT 34.294 37.902 34.346 37.938 ;
      RECT 34.134 37.902 34.186 37.938 ;
      RECT 33.894 37.902 33.946 37.938 ;
      RECT 33.494 37.902 33.546 37.938 ;
      RECT 33.334 37.902 33.386 37.938 ;
      RECT 33.094 37.902 33.146 37.938 ;
      RECT 32.694 37.902 32.746 37.938 ;
      RECT 32.534 37.902 32.586 37.938 ;
      RECT 32.294 37.902 32.346 37.938 ;
      RECT 31.894 37.902 31.946 37.938 ;
      RECT 31.734 37.902 31.786 37.938 ;
      RECT 31.494 37.902 31.546 37.938 ;
      RECT 31.094 37.902 31.146 37.938 ;
      RECT 30.934 37.902 30.986 37.938 ;
      RECT 30.694 37.902 30.746 37.938 ;
      RECT 30.294 37.902 30.346 37.938 ;
      RECT 30.134 37.902 30.186 37.938 ;
      RECT 29.894 37.902 29.946 37.938 ;
      RECT 29.494 37.902 29.546 37.938 ;
      RECT 29.334 37.902 29.386 37.938 ;
      RECT 29.094 37.902 29.146 37.938 ;
      RECT 28.694 37.902 28.746 37.938 ;
      RECT 28.534 37.902 28.586 37.938 ;
      RECT 28.294 37.902 28.346 37.938 ;
      RECT 27.894 37.902 27.946 37.938 ;
      RECT 27.734 37.902 27.786 37.938 ;
      RECT 27.494 37.902 27.546 37.938 ;
      RECT 27.094 37.902 27.146 37.938 ;
      RECT 26.934 37.902 26.986 37.938 ;
      RECT 26.694 37.902 26.746 37.938 ;
      RECT 26.294 37.902 26.346 37.938 ;
      RECT 26.134 37.902 26.186 37.938 ;
      RECT 25.894 37.902 25.946 37.938 ;
      RECT 25.494 37.902 25.546 37.938 ;
      RECT 25.334 37.902 25.386 37.938 ;
      RECT 25.094 37.902 25.146 37.938 ;
      RECT 24.694 37.902 24.746 37.938 ;
      RECT 24.534 37.902 24.586 37.938 ;
      RECT 24.294 37.902 24.346 37.938 ;
      RECT 23.894 37.902 23.946 37.938 ;
      RECT 23.734 37.902 23.786 37.938 ;
      RECT 23.494 37.902 23.546 37.938 ;
      RECT 23.094 37.902 23.146 37.938 ;
      RECT 22.934 37.902 22.986 37.938 ;
      RECT 22.694 37.902 22.746 37.938 ;
      RECT 21.978 37.902 22.022 37.938 ;
      RECT 21.096 37.902 21.14 37.938 ;
      RECT 14.86 37.902 14.904 37.938 ;
      RECT 13.978 37.902 14.022 37.938 ;
      RECT 13.294 37.902 13.346 37.938 ;
      RECT 12.894 37.902 12.946 37.938 ;
      RECT 12.734 37.902 12.786 37.938 ;
      RECT 12.494 37.902 12.546 37.938 ;
      RECT 12.094 37.902 12.146 37.938 ;
      RECT 11.934 37.902 11.986 37.938 ;
      RECT 11.694 37.902 11.746 37.938 ;
      RECT 11.294 37.902 11.346 37.938 ;
      RECT 11.134 37.902 11.186 37.938 ;
      RECT 10.894 37.902 10.946 37.938 ;
      RECT 10.494 37.902 10.546 37.938 ;
      RECT 10.334 37.902 10.386 37.938 ;
      RECT 10.094 37.902 10.146 37.938 ;
      RECT 9.694 37.902 9.746 37.938 ;
      RECT 9.534 37.902 9.586 37.938 ;
      RECT 9.294 37.902 9.346 37.938 ;
      RECT 8.894 37.902 8.946 37.938 ;
      RECT 8.734 37.902 8.786 37.938 ;
      RECT 8.494 37.902 8.546 37.938 ;
      RECT 8.094 37.902 8.146 37.938 ;
      RECT 7.934 37.902 7.986 37.938 ;
      RECT 7.694 37.902 7.746 37.938 ;
      RECT 7.294 37.902 7.346 37.938 ;
      RECT 7.134 37.902 7.186 37.938 ;
      RECT 6.894 37.902 6.946 37.938 ;
      RECT 6.494 37.902 6.546 37.938 ;
      RECT 6.334 37.902 6.386 37.938 ;
      RECT 6.094 37.902 6.146 37.938 ;
      RECT 5.694 37.902 5.746 37.938 ;
      RECT 5.534 37.902 5.586 37.938 ;
      RECT 5.294 37.902 5.346 37.938 ;
      RECT 4.894 37.902 4.946 37.938 ;
      RECT 4.734 37.902 4.786 37.938 ;
      RECT 4.494 37.902 4.546 37.938 ;
      RECT 4.094 37.902 4.146 37.938 ;
      RECT 3.934 37.902 3.986 37.938 ;
      RECT 3.694 37.902 3.746 37.938 ;
      RECT 3.294 37.902 3.346 37.938 ;
      RECT 3.134 37.902 3.186 37.938 ;
      RECT 2.894 37.902 2.946 37.938 ;
      RECT 2.494 37.902 2.546 37.938 ;
      RECT 2.334 37.902 2.386 37.938 ;
      RECT 2.094 37.902 2.146 37.938 ;
      RECT 1.694 37.902 1.746 37.938 ;
      RECT 1.534 37.902 1.586 37.938 ;
      RECT 1.294 37.902 1.346 37.938 ;
      RECT 0.894 37.902 0.946 37.938 ;
      RECT 0.734 37.902 0.786 37.938 ;
      RECT 20.37 37.7875 20.442 37.8125 ;
      RECT 15.558 37.7875 15.63 37.8125 ;
      RECT 21.414 37.6035 21.468 37.6395 ;
      RECT 14.532 37.6035 14.586 37.6395 ;
      RECT 21.978 37.422 22.022 37.458 ;
      RECT 21.096 37.422 21.14 37.458 ;
      RECT 14.86 37.422 14.904 37.458 ;
      RECT 13.978 37.422 14.022 37.458 ;
      RECT 21.814 37.3635 21.868 37.3995 ;
      RECT 20.932 37.3635 20.986 37.3995 ;
      RECT 15.014 37.3635 15.068 37.3995 ;
      RECT 14.132 37.3635 14.186 37.3995 ;
      RECT 21.578 37.302 21.622 37.338 ;
      RECT 20.154 37.302 20.194 37.338 ;
      RECT 15.806 37.302 15.846 37.338 ;
      RECT 14.378 37.302 14.422 37.338 ;
      RECT 16.19 37.2405 16.238 37.2765 ;
      RECT 35.254 37.182 35.306 37.218 ;
      RECT 34.454 37.182 34.506 37.218 ;
      RECT 33.654 37.182 33.706 37.218 ;
      RECT 32.854 37.182 32.906 37.218 ;
      RECT 32.054 37.182 32.106 37.218 ;
      RECT 31.254 37.182 31.306 37.218 ;
      RECT 30.454 37.182 30.506 37.218 ;
      RECT 29.654 37.182 29.706 37.218 ;
      RECT 28.854 37.182 28.906 37.218 ;
      RECT 28.054 37.182 28.106 37.218 ;
      RECT 27.254 37.182 27.306 37.218 ;
      RECT 26.454 37.182 26.506 37.218 ;
      RECT 25.654 37.182 25.706 37.218 ;
      RECT 24.854 37.182 24.906 37.218 ;
      RECT 24.054 37.182 24.106 37.218 ;
      RECT 23.254 37.182 23.306 37.218 ;
      RECT 13.054 37.182 13.106 37.218 ;
      RECT 12.254 37.182 12.306 37.218 ;
      RECT 11.454 37.182 11.506 37.218 ;
      RECT 10.654 37.182 10.706 37.218 ;
      RECT 9.854 37.182 9.906 37.218 ;
      RECT 9.054 37.182 9.106 37.218 ;
      RECT 8.254 37.182 8.306 37.218 ;
      RECT 7.454 37.182 7.506 37.218 ;
      RECT 6.654 37.182 6.706 37.218 ;
      RECT 5.854 37.182 5.906 37.218 ;
      RECT 5.054 37.182 5.106 37.218 ;
      RECT 4.254 37.182 4.306 37.218 ;
      RECT 3.454 37.182 3.506 37.218 ;
      RECT 2.654 37.182 2.706 37.218 ;
      RECT 1.854 37.182 1.906 37.218 ;
      RECT 1.054 37.182 1.106 37.218 ;
      RECT 19.762 37.1235 19.81 37.1595 ;
      RECT 16.422 37.1235 16.47 37.1595 ;
      RECT 21.732 37.0005 21.786 37.0365 ;
      RECT 19.838 37.0005 19.886 37.0365 ;
      RECT 14.214 37.0005 14.268 37.0365 ;
      RECT 21.978 36.942 22.022 36.978 ;
      RECT 21.096 36.942 21.14 36.978 ;
      RECT 14.86 36.942 14.904 36.978 ;
      RECT 13.978 36.942 14.022 36.978 ;
      RECT 35.254 36.702 35.306 36.738 ;
      RECT 34.454 36.702 34.506 36.738 ;
      RECT 33.654 36.702 33.706 36.738 ;
      RECT 32.854 36.702 32.906 36.738 ;
      RECT 32.054 36.702 32.106 36.738 ;
      RECT 31.254 36.702 31.306 36.738 ;
      RECT 30.454 36.702 30.506 36.738 ;
      RECT 29.654 36.702 29.706 36.738 ;
      RECT 28.854 36.702 28.906 36.738 ;
      RECT 28.054 36.702 28.106 36.738 ;
      RECT 27.254 36.702 27.306 36.738 ;
      RECT 26.454 36.702 26.506 36.738 ;
      RECT 25.654 36.702 25.706 36.738 ;
      RECT 24.854 36.702 24.906 36.738 ;
      RECT 24.054 36.702 24.106 36.738 ;
      RECT 23.254 36.702 23.306 36.738 ;
      RECT 13.054 36.702 13.106 36.738 ;
      RECT 12.254 36.702 12.306 36.738 ;
      RECT 11.454 36.702 11.506 36.738 ;
      RECT 10.654 36.702 10.706 36.738 ;
      RECT 9.854 36.702 9.906 36.738 ;
      RECT 9.054 36.702 9.106 36.738 ;
      RECT 8.254 36.702 8.306 36.738 ;
      RECT 7.454 36.702 7.506 36.738 ;
      RECT 6.654 36.702 6.706 36.738 ;
      RECT 5.854 36.702 5.906 36.738 ;
      RECT 5.054 36.702 5.106 36.738 ;
      RECT 4.254 36.702 4.306 36.738 ;
      RECT 3.454 36.702 3.506 36.738 ;
      RECT 2.654 36.702 2.706 36.738 ;
      RECT 1.854 36.702 1.906 36.738 ;
      RECT 1.054 36.702 1.106 36.738 ;
      RECT 21.978 36.462 22.022 36.498 ;
      RECT 21.096 36.462 21.14 36.498 ;
      RECT 14.86 36.462 14.904 36.498 ;
      RECT 13.978 36.462 14.022 36.498 ;
      RECT 21.578 36.342 21.622 36.378 ;
      RECT 14.378 36.342 14.422 36.378 ;
      RECT 20.55 36.102 20.602 36.138 ;
      RECT 15.398 36.102 15.45 36.138 ;
      RECT 21.978 35.982 22.022 36.018 ;
      RECT 21.096 35.982 21.14 36.018 ;
      RECT 14.86 35.982 14.904 36.018 ;
      RECT 13.978 35.982 14.022 36.018 ;
      RECT 21.814 35.9235 21.868 35.9595 ;
      RECT 14.132 35.9235 14.186 35.9595 ;
      RECT 19.606 35.8005 19.654 35.8365 ;
      RECT 20.222 35.6835 20.262 35.7195 ;
      RECT 15.738 35.6835 15.778 35.7195 ;
      RECT 16.346 35.622 16.394 35.658 ;
      RECT 21.978 35.502 22.022 35.538 ;
      RECT 21.096 35.502 21.14 35.538 ;
      RECT 14.86 35.502 14.904 35.538 ;
      RECT 13.978 35.502 14.022 35.538 ;
      RECT 19.838 35.382 19.886 35.418 ;
      RECT 21.978 35.022 22.022 35.058 ;
      RECT 21.096 35.022 21.14 35.058 ;
      RECT 17.944 35.022 17.984 35.058 ;
      RECT 14.86 35.022 14.904 35.058 ;
      RECT 13.978 35.022 14.022 35.058 ;
      RECT 19.838 34.902 19.886 34.938 ;
      RECT 16.422 34.902 16.47 34.938 ;
      RECT 35.254 34.782 35.306 34.818 ;
      RECT 34.454 34.782 34.506 34.818 ;
      RECT 33.654 34.782 33.706 34.818 ;
      RECT 32.854 34.782 32.906 34.818 ;
      RECT 32.054 34.782 32.106 34.818 ;
      RECT 31.254 34.782 31.306 34.818 ;
      RECT 30.454 34.782 30.506 34.818 ;
      RECT 29.654 34.782 29.706 34.818 ;
      RECT 28.854 34.782 28.906 34.818 ;
      RECT 28.054 34.782 28.106 34.818 ;
      RECT 27.254 34.782 27.306 34.818 ;
      RECT 26.454 34.782 26.506 34.818 ;
      RECT 25.654 34.782 25.706 34.818 ;
      RECT 24.854 34.782 24.906 34.818 ;
      RECT 24.054 34.782 24.106 34.818 ;
      RECT 23.254 34.782 23.306 34.818 ;
      RECT 13.054 34.782 13.106 34.818 ;
      RECT 12.254 34.782 12.306 34.818 ;
      RECT 11.454 34.782 11.506 34.818 ;
      RECT 10.654 34.782 10.706 34.818 ;
      RECT 9.854 34.782 9.906 34.818 ;
      RECT 9.054 34.782 9.106 34.818 ;
      RECT 8.254 34.782 8.306 34.818 ;
      RECT 7.454 34.782 7.506 34.818 ;
      RECT 6.654 34.782 6.706 34.818 ;
      RECT 5.854 34.782 5.906 34.818 ;
      RECT 5.054 34.782 5.106 34.818 ;
      RECT 4.254 34.782 4.306 34.818 ;
      RECT 3.454 34.782 3.506 34.818 ;
      RECT 2.654 34.782 2.706 34.818 ;
      RECT 1.854 34.782 1.906 34.818 ;
      RECT 1.054 34.782 1.106 34.818 ;
      RECT 20.55 34.6005 20.602 34.6365 ;
      RECT 15.398 34.6005 15.45 34.6365 ;
      RECT 21.978 34.542 22.022 34.578 ;
      RECT 21.096 34.542 21.14 34.578 ;
      RECT 17.944 34.542 17.984 34.578 ;
      RECT 14.86 34.542 14.904 34.578 ;
      RECT 13.978 34.542 14.022 34.578 ;
      RECT 20.932 34.4835 20.986 34.5195 ;
      RECT 15.014 34.4835 15.068 34.5195 ;
      RECT 21.578 34.422 21.622 34.458 ;
      RECT 17.944 34.422 17.984 34.458 ;
      RECT 14.378 34.422 14.422 34.458 ;
      RECT 21.814 34.3605 21.868 34.3965 ;
      RECT 14.132 34.3605 14.186 34.3965 ;
      RECT 35.254 34.302 35.306 34.338 ;
      RECT 34.454 34.302 34.506 34.338 ;
      RECT 33.654 34.302 33.706 34.338 ;
      RECT 32.854 34.302 32.906 34.338 ;
      RECT 32.054 34.302 32.106 34.338 ;
      RECT 31.254 34.302 31.306 34.338 ;
      RECT 30.454 34.302 30.506 34.338 ;
      RECT 29.654 34.302 29.706 34.338 ;
      RECT 28.854 34.302 28.906 34.338 ;
      RECT 28.054 34.302 28.106 34.338 ;
      RECT 27.254 34.302 27.306 34.338 ;
      RECT 26.454 34.302 26.506 34.338 ;
      RECT 25.654 34.302 25.706 34.338 ;
      RECT 24.854 34.302 24.906 34.338 ;
      RECT 24.054 34.302 24.106 34.338 ;
      RECT 23.254 34.302 23.306 34.338 ;
      RECT 13.054 34.302 13.106 34.338 ;
      RECT 12.254 34.302 12.306 34.338 ;
      RECT 11.454 34.302 11.506 34.338 ;
      RECT 10.654 34.302 10.706 34.338 ;
      RECT 9.854 34.302 9.906 34.338 ;
      RECT 9.054 34.302 9.106 34.338 ;
      RECT 8.254 34.302 8.306 34.338 ;
      RECT 7.454 34.302 7.506 34.338 ;
      RECT 6.654 34.302 6.706 34.338 ;
      RECT 5.854 34.302 5.906 34.338 ;
      RECT 5.054 34.302 5.106 34.338 ;
      RECT 4.254 34.302 4.306 34.338 ;
      RECT 3.454 34.302 3.506 34.338 ;
      RECT 2.654 34.302 2.706 34.338 ;
      RECT 1.854 34.302 1.906 34.338 ;
      RECT 1.054 34.302 1.106 34.338 ;
      RECT 21.578 34.182 21.622 34.218 ;
      RECT 14.378 34.182 14.422 34.218 ;
      RECT 21.814 34.1205 21.868 34.1565 ;
      RECT 14.132 34.1205 14.186 34.1565 ;
      RECT 21.978 34.062 22.022 34.098 ;
      RECT 21.096 34.062 21.14 34.098 ;
      RECT 17.616 34.062 17.656 34.098 ;
      RECT 14.86 34.062 14.904 34.098 ;
      RECT 13.978 34.062 14.022 34.098 ;
      RECT 21.732 34.0035 21.786 34.0395 ;
      RECT 14.214 34.0035 14.268 34.0395 ;
      RECT 35.494 33.582 35.546 33.618 ;
      RECT 35.094 33.582 35.146 33.618 ;
      RECT 34.934 33.582 34.986 33.618 ;
      RECT 34.694 33.582 34.746 33.618 ;
      RECT 34.294 33.582 34.346 33.618 ;
      RECT 34.134 33.582 34.186 33.618 ;
      RECT 33.894 33.582 33.946 33.618 ;
      RECT 33.494 33.582 33.546 33.618 ;
      RECT 33.334 33.582 33.386 33.618 ;
      RECT 33.094 33.582 33.146 33.618 ;
      RECT 32.694 33.582 32.746 33.618 ;
      RECT 32.534 33.582 32.586 33.618 ;
      RECT 32.294 33.582 32.346 33.618 ;
      RECT 31.894 33.582 31.946 33.618 ;
      RECT 31.734 33.582 31.786 33.618 ;
      RECT 31.494 33.582 31.546 33.618 ;
      RECT 31.094 33.582 31.146 33.618 ;
      RECT 30.934 33.582 30.986 33.618 ;
      RECT 30.694 33.582 30.746 33.618 ;
      RECT 30.294 33.582 30.346 33.618 ;
      RECT 30.134 33.582 30.186 33.618 ;
      RECT 29.894 33.582 29.946 33.618 ;
      RECT 29.494 33.582 29.546 33.618 ;
      RECT 29.334 33.582 29.386 33.618 ;
      RECT 29.094 33.582 29.146 33.618 ;
      RECT 28.694 33.582 28.746 33.618 ;
      RECT 28.534 33.582 28.586 33.618 ;
      RECT 28.294 33.582 28.346 33.618 ;
      RECT 27.894 33.582 27.946 33.618 ;
      RECT 27.734 33.582 27.786 33.618 ;
      RECT 27.494 33.582 27.546 33.618 ;
      RECT 27.094 33.582 27.146 33.618 ;
      RECT 26.934 33.582 26.986 33.618 ;
      RECT 26.694 33.582 26.746 33.618 ;
      RECT 26.294 33.582 26.346 33.618 ;
      RECT 26.134 33.582 26.186 33.618 ;
      RECT 25.894 33.582 25.946 33.618 ;
      RECT 25.494 33.582 25.546 33.618 ;
      RECT 25.334 33.582 25.386 33.618 ;
      RECT 25.094 33.582 25.146 33.618 ;
      RECT 24.694 33.582 24.746 33.618 ;
      RECT 24.534 33.582 24.586 33.618 ;
      RECT 24.294 33.582 24.346 33.618 ;
      RECT 23.894 33.582 23.946 33.618 ;
      RECT 23.734 33.582 23.786 33.618 ;
      RECT 23.494 33.582 23.546 33.618 ;
      RECT 23.094 33.582 23.146 33.618 ;
      RECT 22.934 33.582 22.986 33.618 ;
      RECT 22.694 33.582 22.746 33.618 ;
      RECT 21.978 33.582 22.022 33.618 ;
      RECT 21.096 33.582 21.14 33.618 ;
      RECT 17.616 33.582 17.656 33.618 ;
      RECT 14.86 33.582 14.904 33.618 ;
      RECT 13.978 33.582 14.022 33.618 ;
      RECT 13.294 33.582 13.346 33.618 ;
      RECT 12.894 33.582 12.946 33.618 ;
      RECT 12.734 33.582 12.786 33.618 ;
      RECT 12.494 33.582 12.546 33.618 ;
      RECT 12.094 33.582 12.146 33.618 ;
      RECT 11.934 33.582 11.986 33.618 ;
      RECT 11.694 33.582 11.746 33.618 ;
      RECT 11.294 33.582 11.346 33.618 ;
      RECT 11.134 33.582 11.186 33.618 ;
      RECT 10.894 33.582 10.946 33.618 ;
      RECT 10.494 33.582 10.546 33.618 ;
      RECT 10.334 33.582 10.386 33.618 ;
      RECT 10.094 33.582 10.146 33.618 ;
      RECT 9.694 33.582 9.746 33.618 ;
      RECT 9.534 33.582 9.586 33.618 ;
      RECT 9.294 33.582 9.346 33.618 ;
      RECT 8.894 33.582 8.946 33.618 ;
      RECT 8.734 33.582 8.786 33.618 ;
      RECT 8.494 33.582 8.546 33.618 ;
      RECT 8.094 33.582 8.146 33.618 ;
      RECT 7.934 33.582 7.986 33.618 ;
      RECT 7.694 33.582 7.746 33.618 ;
      RECT 7.294 33.582 7.346 33.618 ;
      RECT 7.134 33.582 7.186 33.618 ;
      RECT 6.894 33.582 6.946 33.618 ;
      RECT 6.494 33.582 6.546 33.618 ;
      RECT 6.334 33.582 6.386 33.618 ;
      RECT 6.094 33.582 6.146 33.618 ;
      RECT 5.694 33.582 5.746 33.618 ;
      RECT 5.534 33.582 5.586 33.618 ;
      RECT 5.294 33.582 5.346 33.618 ;
      RECT 4.894 33.582 4.946 33.618 ;
      RECT 4.734 33.582 4.786 33.618 ;
      RECT 4.494 33.582 4.546 33.618 ;
      RECT 4.094 33.582 4.146 33.618 ;
      RECT 3.934 33.582 3.986 33.618 ;
      RECT 3.694 33.582 3.746 33.618 ;
      RECT 3.294 33.582 3.346 33.618 ;
      RECT 3.134 33.582 3.186 33.618 ;
      RECT 2.894 33.582 2.946 33.618 ;
      RECT 2.494 33.582 2.546 33.618 ;
      RECT 2.334 33.582 2.386 33.618 ;
      RECT 2.094 33.582 2.146 33.618 ;
      RECT 1.694 33.582 1.746 33.618 ;
      RECT 1.534 33.582 1.586 33.618 ;
      RECT 1.294 33.582 1.346 33.618 ;
      RECT 0.894 33.582 0.946 33.618 ;
      RECT 0.734 33.582 0.786 33.618 ;
      RECT 15.558 33.4675 15.63 33.4925 ;
      RECT 17.616 33.4005 17.656 33.4365 ;
      RECT 20.37 33.406 20.442 33.431 ;
      RECT 35.494 33.342 35.546 33.378 ;
      RECT 35.094 33.342 35.146 33.378 ;
      RECT 34.934 33.342 34.986 33.378 ;
      RECT 34.694 33.342 34.746 33.378 ;
      RECT 34.294 33.342 34.346 33.378 ;
      RECT 34.134 33.342 34.186 33.378 ;
      RECT 33.894 33.342 33.946 33.378 ;
      RECT 33.494 33.342 33.546 33.378 ;
      RECT 33.334 33.342 33.386 33.378 ;
      RECT 33.094 33.342 33.146 33.378 ;
      RECT 32.694 33.342 32.746 33.378 ;
      RECT 32.534 33.342 32.586 33.378 ;
      RECT 32.294 33.342 32.346 33.378 ;
      RECT 31.894 33.342 31.946 33.378 ;
      RECT 31.734 33.342 31.786 33.378 ;
      RECT 31.494 33.342 31.546 33.378 ;
      RECT 31.094 33.342 31.146 33.378 ;
      RECT 30.934 33.342 30.986 33.378 ;
      RECT 30.694 33.342 30.746 33.378 ;
      RECT 30.294 33.342 30.346 33.378 ;
      RECT 30.134 33.342 30.186 33.378 ;
      RECT 29.894 33.342 29.946 33.378 ;
      RECT 29.494 33.342 29.546 33.378 ;
      RECT 29.334 33.342 29.386 33.378 ;
      RECT 29.094 33.342 29.146 33.378 ;
      RECT 28.694 33.342 28.746 33.378 ;
      RECT 28.534 33.342 28.586 33.378 ;
      RECT 28.294 33.342 28.346 33.378 ;
      RECT 27.894 33.342 27.946 33.378 ;
      RECT 27.734 33.342 27.786 33.378 ;
      RECT 27.494 33.342 27.546 33.378 ;
      RECT 27.094 33.342 27.146 33.378 ;
      RECT 26.934 33.342 26.986 33.378 ;
      RECT 26.694 33.342 26.746 33.378 ;
      RECT 26.294 33.342 26.346 33.378 ;
      RECT 26.134 33.342 26.186 33.378 ;
      RECT 25.894 33.342 25.946 33.378 ;
      RECT 25.494 33.342 25.546 33.378 ;
      RECT 25.334 33.342 25.386 33.378 ;
      RECT 25.094 33.342 25.146 33.378 ;
      RECT 24.694 33.342 24.746 33.378 ;
      RECT 24.534 33.342 24.586 33.378 ;
      RECT 24.294 33.342 24.346 33.378 ;
      RECT 23.894 33.342 23.946 33.378 ;
      RECT 23.734 33.342 23.786 33.378 ;
      RECT 23.494 33.342 23.546 33.378 ;
      RECT 23.094 33.342 23.146 33.378 ;
      RECT 22.934 33.342 22.986 33.378 ;
      RECT 22.694 33.342 22.746 33.378 ;
      RECT 13.294 33.342 13.346 33.378 ;
      RECT 12.894 33.342 12.946 33.378 ;
      RECT 12.734 33.342 12.786 33.378 ;
      RECT 12.494 33.342 12.546 33.378 ;
      RECT 12.094 33.342 12.146 33.378 ;
      RECT 11.934 33.342 11.986 33.378 ;
      RECT 11.694 33.342 11.746 33.378 ;
      RECT 11.294 33.342 11.346 33.378 ;
      RECT 11.134 33.342 11.186 33.378 ;
      RECT 10.894 33.342 10.946 33.378 ;
      RECT 10.494 33.342 10.546 33.378 ;
      RECT 10.334 33.342 10.386 33.378 ;
      RECT 10.094 33.342 10.146 33.378 ;
      RECT 9.694 33.342 9.746 33.378 ;
      RECT 9.534 33.342 9.586 33.378 ;
      RECT 9.294 33.342 9.346 33.378 ;
      RECT 8.894 33.342 8.946 33.378 ;
      RECT 8.734 33.342 8.786 33.378 ;
      RECT 8.494 33.342 8.546 33.378 ;
      RECT 8.094 33.342 8.146 33.378 ;
      RECT 7.934 33.342 7.986 33.378 ;
      RECT 7.694 33.342 7.746 33.378 ;
      RECT 7.294 33.342 7.346 33.378 ;
      RECT 7.134 33.342 7.186 33.378 ;
      RECT 6.894 33.342 6.946 33.378 ;
      RECT 6.494 33.342 6.546 33.378 ;
      RECT 6.334 33.342 6.386 33.378 ;
      RECT 6.094 33.342 6.146 33.378 ;
      RECT 5.694 33.342 5.746 33.378 ;
      RECT 5.534 33.342 5.586 33.378 ;
      RECT 5.294 33.342 5.346 33.378 ;
      RECT 4.894 33.342 4.946 33.378 ;
      RECT 4.734 33.342 4.786 33.378 ;
      RECT 4.494 33.342 4.546 33.378 ;
      RECT 4.094 33.342 4.146 33.378 ;
      RECT 3.934 33.342 3.986 33.378 ;
      RECT 3.694 33.342 3.746 33.378 ;
      RECT 3.294 33.342 3.346 33.378 ;
      RECT 3.134 33.342 3.186 33.378 ;
      RECT 2.894 33.342 2.946 33.378 ;
      RECT 2.494 33.342 2.546 33.378 ;
      RECT 2.334 33.342 2.386 33.378 ;
      RECT 2.094 33.342 2.146 33.378 ;
      RECT 1.694 33.342 1.746 33.378 ;
      RECT 1.534 33.342 1.586 33.378 ;
      RECT 1.294 33.342 1.346 33.378 ;
      RECT 0.894 33.342 0.946 33.378 ;
      RECT 0.734 33.342 0.786 33.378 ;
      RECT 20.222 33.222 20.262 33.258 ;
      RECT 19.762 33.222 19.81 33.258 ;
      RECT 19.606 33.222 19.654 33.258 ;
      RECT 16.346 33.222 16.394 33.258 ;
      RECT 16.19 33.222 16.238 33.258 ;
      RECT 15.738 33.222 15.778 33.258 ;
      RECT 21.978 33.102 22.022 33.138 ;
      RECT 21.096 33.102 21.14 33.138 ;
      RECT 14.86 33.102 14.904 33.138 ;
      RECT 13.978 33.102 14.022 33.138 ;
      RECT 20.154 32.982 20.194 33.018 ;
      RECT 15.806 32.982 15.846 33.018 ;
      RECT 17.944 32.9205 17.984 32.9565 ;
      RECT 35.254 32.862 35.306 32.898 ;
      RECT 34.854 32.862 34.906 32.898 ;
      RECT 34.454 32.862 34.506 32.898 ;
      RECT 34.054 32.862 34.106 32.898 ;
      RECT 33.654 32.862 33.706 32.898 ;
      RECT 33.254 32.862 33.306 32.898 ;
      RECT 32.854 32.862 32.906 32.898 ;
      RECT 32.454 32.862 32.506 32.898 ;
      RECT 32.054 32.862 32.106 32.898 ;
      RECT 31.654 32.862 31.706 32.898 ;
      RECT 31.254 32.862 31.306 32.898 ;
      RECT 30.854 32.862 30.906 32.898 ;
      RECT 30.454 32.862 30.506 32.898 ;
      RECT 30.054 32.862 30.106 32.898 ;
      RECT 29.654 32.862 29.706 32.898 ;
      RECT 29.254 32.862 29.306 32.898 ;
      RECT 28.854 32.862 28.906 32.898 ;
      RECT 28.454 32.862 28.506 32.898 ;
      RECT 28.054 32.862 28.106 32.898 ;
      RECT 27.654 32.862 27.706 32.898 ;
      RECT 27.254 32.862 27.306 32.898 ;
      RECT 26.854 32.862 26.906 32.898 ;
      RECT 26.454 32.862 26.506 32.898 ;
      RECT 26.054 32.862 26.106 32.898 ;
      RECT 25.654 32.862 25.706 32.898 ;
      RECT 25.254 32.862 25.306 32.898 ;
      RECT 24.854 32.862 24.906 32.898 ;
      RECT 24.454 32.862 24.506 32.898 ;
      RECT 24.054 32.862 24.106 32.898 ;
      RECT 23.654 32.862 23.706 32.898 ;
      RECT 23.254 32.862 23.306 32.898 ;
      RECT 22.854 32.862 22.906 32.898 ;
      RECT 13.054 32.862 13.106 32.898 ;
      RECT 12.654 32.862 12.706 32.898 ;
      RECT 12.254 32.862 12.306 32.898 ;
      RECT 11.854 32.862 11.906 32.898 ;
      RECT 11.454 32.862 11.506 32.898 ;
      RECT 11.054 32.862 11.106 32.898 ;
      RECT 10.654 32.862 10.706 32.898 ;
      RECT 10.254 32.862 10.306 32.898 ;
      RECT 9.854 32.862 9.906 32.898 ;
      RECT 9.454 32.862 9.506 32.898 ;
      RECT 9.054 32.862 9.106 32.898 ;
      RECT 8.654 32.862 8.706 32.898 ;
      RECT 8.254 32.862 8.306 32.898 ;
      RECT 7.854 32.862 7.906 32.898 ;
      RECT 7.454 32.862 7.506 32.898 ;
      RECT 7.054 32.862 7.106 32.898 ;
      RECT 6.654 32.862 6.706 32.898 ;
      RECT 6.254 32.862 6.306 32.898 ;
      RECT 5.854 32.862 5.906 32.898 ;
      RECT 5.454 32.862 5.506 32.898 ;
      RECT 5.054 32.862 5.106 32.898 ;
      RECT 4.654 32.862 4.706 32.898 ;
      RECT 4.254 32.862 4.306 32.898 ;
      RECT 3.854 32.862 3.906 32.898 ;
      RECT 3.454 32.862 3.506 32.898 ;
      RECT 3.054 32.862 3.106 32.898 ;
      RECT 2.654 32.862 2.706 32.898 ;
      RECT 2.254 32.862 2.306 32.898 ;
      RECT 1.854 32.862 1.906 32.898 ;
      RECT 1.454 32.862 1.506 32.898 ;
      RECT 1.054 32.862 1.106 32.898 ;
      RECT 0.654 32.862 0.706 32.898 ;
      RECT 19.606 32.742 19.654 32.778 ;
      RECT 17.136 32.742 17.176 32.778 ;
      RECT 16.114 32.742 16.162 32.778 ;
      RECT 16.346 32.6805 16.394 32.7165 ;
      RECT 35.254 32.622 35.306 32.658 ;
      RECT 34.854 32.622 34.906 32.658 ;
      RECT 34.454 32.622 34.506 32.658 ;
      RECT 34.054 32.622 34.106 32.658 ;
      RECT 33.654 32.622 33.706 32.658 ;
      RECT 33.254 32.622 33.306 32.658 ;
      RECT 32.854 32.622 32.906 32.658 ;
      RECT 32.454 32.622 32.506 32.658 ;
      RECT 32.054 32.622 32.106 32.658 ;
      RECT 31.654 32.622 31.706 32.658 ;
      RECT 31.254 32.622 31.306 32.658 ;
      RECT 30.854 32.622 30.906 32.658 ;
      RECT 30.454 32.622 30.506 32.658 ;
      RECT 30.054 32.622 30.106 32.658 ;
      RECT 29.654 32.622 29.706 32.658 ;
      RECT 29.254 32.622 29.306 32.658 ;
      RECT 28.854 32.622 28.906 32.658 ;
      RECT 28.454 32.622 28.506 32.658 ;
      RECT 28.054 32.622 28.106 32.658 ;
      RECT 27.654 32.622 27.706 32.658 ;
      RECT 27.254 32.622 27.306 32.658 ;
      RECT 26.854 32.622 26.906 32.658 ;
      RECT 26.454 32.622 26.506 32.658 ;
      RECT 26.054 32.622 26.106 32.658 ;
      RECT 25.654 32.622 25.706 32.658 ;
      RECT 25.254 32.622 25.306 32.658 ;
      RECT 24.854 32.622 24.906 32.658 ;
      RECT 24.454 32.622 24.506 32.658 ;
      RECT 24.054 32.622 24.106 32.658 ;
      RECT 23.654 32.622 23.706 32.658 ;
      RECT 23.254 32.622 23.306 32.658 ;
      RECT 22.854 32.622 22.906 32.658 ;
      RECT 21.978 32.622 22.022 32.658 ;
      RECT 21.096 32.622 21.14 32.658 ;
      RECT 17.944 32.622 17.984 32.658 ;
      RECT 17.136 32.622 17.176 32.658 ;
      RECT 14.86 32.622 14.904 32.658 ;
      RECT 13.978 32.622 14.022 32.658 ;
      RECT 13.054 32.622 13.106 32.658 ;
      RECT 12.654 32.622 12.706 32.658 ;
      RECT 12.254 32.622 12.306 32.658 ;
      RECT 11.854 32.622 11.906 32.658 ;
      RECT 11.454 32.622 11.506 32.658 ;
      RECT 11.054 32.622 11.106 32.658 ;
      RECT 10.654 32.622 10.706 32.658 ;
      RECT 10.254 32.622 10.306 32.658 ;
      RECT 9.854 32.622 9.906 32.658 ;
      RECT 9.454 32.622 9.506 32.658 ;
      RECT 9.054 32.622 9.106 32.658 ;
      RECT 8.654 32.622 8.706 32.658 ;
      RECT 8.254 32.622 8.306 32.658 ;
      RECT 7.854 32.622 7.906 32.658 ;
      RECT 7.454 32.622 7.506 32.658 ;
      RECT 7.054 32.622 7.106 32.658 ;
      RECT 6.654 32.622 6.706 32.658 ;
      RECT 6.254 32.622 6.306 32.658 ;
      RECT 5.854 32.622 5.906 32.658 ;
      RECT 5.454 32.622 5.506 32.658 ;
      RECT 5.054 32.622 5.106 32.658 ;
      RECT 4.654 32.622 4.706 32.658 ;
      RECT 4.254 32.622 4.306 32.658 ;
      RECT 3.854 32.622 3.906 32.658 ;
      RECT 3.454 32.622 3.506 32.658 ;
      RECT 3.054 32.622 3.106 32.658 ;
      RECT 2.654 32.622 2.706 32.658 ;
      RECT 2.254 32.622 2.306 32.658 ;
      RECT 1.854 32.622 1.906 32.658 ;
      RECT 1.454 32.622 1.506 32.658 ;
      RECT 1.054 32.622 1.106 32.658 ;
      RECT 0.654 32.622 0.706 32.658 ;
      RECT 19.838 32.502 19.886 32.538 ;
      RECT 18.492 32.502 18.536 32.538 ;
      RECT 17.944 32.502 17.984 32.538 ;
      RECT 16.19 32.502 16.238 32.538 ;
      RECT 21.414 32.4405 21.468 32.4765 ;
      RECT 16.422 32.4405 16.47 32.4765 ;
      RECT 14.532 32.4405 14.586 32.4765 ;
      RECT 21.414 32.3235 21.468 32.3595 ;
      RECT 19.53 32.3235 19.578 32.3595 ;
      RECT 14.532 32.3235 14.586 32.3595 ;
      RECT 19.762 32.262 19.81 32.298 ;
      RECT 20.37 32.2675 20.442 32.2925 ;
      RECT 15.558 32.2675 15.63 32.2925 ;
      RECT 16.882 32.2005 16.936 32.2365 ;
      RECT 16.718 32.2005 16.772 32.2365 ;
      RECT 21.978 32.142 22.022 32.178 ;
      RECT 21.096 32.142 21.14 32.178 ;
      RECT 14.86 32.142 14.904 32.178 ;
      RECT 13.978 32.142 14.022 32.178 ;
      RECT 21.978 31.782 22.022 31.818 ;
      RECT 21.096 31.782 21.14 31.818 ;
      RECT 14.86 31.782 14.904 31.818 ;
      RECT 13.978 31.782 14.022 31.818 ;
      RECT 35.494 31.558 35.546 31.594 ;
      RECT 35.094 31.558 35.146 31.594 ;
      RECT 34.694 31.558 34.746 31.594 ;
      RECT 34.294 31.558 34.346 31.594 ;
      RECT 33.894 31.558 33.946 31.594 ;
      RECT 33.494 31.558 33.546 31.594 ;
      RECT 33.094 31.558 33.146 31.594 ;
      RECT 32.694 31.558 32.746 31.594 ;
      RECT 32.294 31.558 32.346 31.594 ;
      RECT 31.894 31.558 31.946 31.594 ;
      RECT 31.494 31.558 31.546 31.594 ;
      RECT 31.094 31.558 31.146 31.594 ;
      RECT 30.694 31.558 30.746 31.594 ;
      RECT 30.294 31.558 30.346 31.594 ;
      RECT 29.894 31.558 29.946 31.594 ;
      RECT 29.494 31.558 29.546 31.594 ;
      RECT 29.094 31.558 29.146 31.594 ;
      RECT 28.694 31.558 28.746 31.594 ;
      RECT 28.294 31.558 28.346 31.594 ;
      RECT 27.894 31.558 27.946 31.594 ;
      RECT 27.494 31.558 27.546 31.594 ;
      RECT 27.094 31.558 27.146 31.594 ;
      RECT 26.694 31.558 26.746 31.594 ;
      RECT 26.294 31.558 26.346 31.594 ;
      RECT 25.894 31.558 25.946 31.594 ;
      RECT 25.494 31.558 25.546 31.594 ;
      RECT 25.094 31.558 25.146 31.594 ;
      RECT 24.694 31.558 24.746 31.594 ;
      RECT 24.294 31.558 24.346 31.594 ;
      RECT 23.894 31.558 23.946 31.594 ;
      RECT 23.494 31.558 23.546 31.594 ;
      RECT 23.094 31.558 23.146 31.594 ;
      RECT 21.814 31.558 21.868 31.594 ;
      RECT 19.838 31.558 19.886 31.594 ;
      RECT 19.53 31.558 19.578 31.594 ;
      RECT 16.882 31.558 16.936 31.594 ;
      RECT 16.422 31.558 16.47 31.594 ;
      RECT 16.114 31.558 16.162 31.594 ;
      RECT 14.132 31.558 14.186 31.594 ;
      RECT 13.294 31.558 13.346 31.594 ;
      RECT 12.894 31.558 12.946 31.594 ;
      RECT 12.494 31.558 12.546 31.594 ;
      RECT 12.094 31.558 12.146 31.594 ;
      RECT 11.694 31.558 11.746 31.594 ;
      RECT 11.294 31.558 11.346 31.594 ;
      RECT 10.894 31.558 10.946 31.594 ;
      RECT 10.494 31.558 10.546 31.594 ;
      RECT 10.094 31.558 10.146 31.594 ;
      RECT 9.694 31.558 9.746 31.594 ;
      RECT 9.294 31.558 9.346 31.594 ;
      RECT 8.894 31.558 8.946 31.594 ;
      RECT 8.494 31.558 8.546 31.594 ;
      RECT 8.094 31.558 8.146 31.594 ;
      RECT 7.694 31.558 7.746 31.594 ;
      RECT 7.294 31.558 7.346 31.594 ;
      RECT 6.894 31.558 6.946 31.594 ;
      RECT 6.494 31.558 6.546 31.594 ;
      RECT 6.094 31.558 6.146 31.594 ;
      RECT 5.694 31.558 5.746 31.594 ;
      RECT 5.294 31.558 5.346 31.594 ;
      RECT 4.894 31.558 4.946 31.594 ;
      RECT 4.494 31.558 4.546 31.594 ;
      RECT 4.094 31.558 4.146 31.594 ;
      RECT 3.694 31.558 3.746 31.594 ;
      RECT 3.294 31.558 3.346 31.594 ;
      RECT 2.894 31.558 2.946 31.594 ;
      RECT 2.494 31.558 2.546 31.594 ;
      RECT 2.094 31.558 2.146 31.594 ;
      RECT 1.694 31.558 1.746 31.594 ;
      RECT 1.294 31.558 1.346 31.594 ;
      RECT 0.894 31.558 0.946 31.594 ;
      RECT 21.414 31.482 21.468 31.518 ;
      RECT 14.532 31.482 14.586 31.518 ;
      RECT 19.606 31.329 19.654 31.365 ;
      RECT 18.08 31.329 18.12 31.365 ;
      RECT 16.718 31.329 16.772 31.365 ;
      RECT 16.346 31.329 16.394 31.365 ;
      RECT 20.37 31.3345 20.442 31.3595 ;
      RECT 18.764 31.3345 18.836 31.3595 ;
      RECT 15.558 31.3345 15.63 31.3595 ;
      RECT 21.978 31.182 22.022 31.218 ;
      RECT 13.978 31.182 14.022 31.218 ;
      RECT 18.764 31.1875 18.836 31.2125 ;
      RECT 19.762 31.035 19.81 31.071 ;
      RECT 17.616 31.035 17.656 31.071 ;
      RECT 16.19 31.035 16.238 31.071 ;
      RECT 35.254 30.806 35.306 30.842 ;
      RECT 34.854 30.806 34.906 30.842 ;
      RECT 34.454 30.806 34.506 30.842 ;
      RECT 34.054 30.806 34.106 30.842 ;
      RECT 33.654 30.806 33.706 30.842 ;
      RECT 33.254 30.806 33.306 30.842 ;
      RECT 32.854 30.806 32.906 30.842 ;
      RECT 32.454 30.806 32.506 30.842 ;
      RECT 32.054 30.806 32.106 30.842 ;
      RECT 31.654 30.806 31.706 30.842 ;
      RECT 31.254 30.806 31.306 30.842 ;
      RECT 30.854 30.806 30.906 30.842 ;
      RECT 30.454 30.806 30.506 30.842 ;
      RECT 30.054 30.806 30.106 30.842 ;
      RECT 29.654 30.806 29.706 30.842 ;
      RECT 29.254 30.806 29.306 30.842 ;
      RECT 28.854 30.806 28.906 30.842 ;
      RECT 28.454 30.806 28.506 30.842 ;
      RECT 28.054 30.806 28.106 30.842 ;
      RECT 27.654 30.806 27.706 30.842 ;
      RECT 27.254 30.806 27.306 30.842 ;
      RECT 26.854 30.806 26.906 30.842 ;
      RECT 26.454 30.806 26.506 30.842 ;
      RECT 26.054 30.806 26.106 30.842 ;
      RECT 25.654 30.806 25.706 30.842 ;
      RECT 25.254 30.806 25.306 30.842 ;
      RECT 24.854 30.806 24.906 30.842 ;
      RECT 24.454 30.806 24.506 30.842 ;
      RECT 24.054 30.806 24.106 30.842 ;
      RECT 23.654 30.806 23.706 30.842 ;
      RECT 23.254 30.806 23.306 30.842 ;
      RECT 22.854 30.806 22.906 30.842 ;
      RECT 22.694 30.806 22.746 30.842 ;
      RECT 21.732 30.806 21.786 30.842 ;
      RECT 14.214 30.806 14.268 30.842 ;
      RECT 13.054 30.806 13.106 30.842 ;
      RECT 12.654 30.806 12.706 30.842 ;
      RECT 12.254 30.806 12.306 30.842 ;
      RECT 11.854 30.806 11.906 30.842 ;
      RECT 11.454 30.806 11.506 30.842 ;
      RECT 11.054 30.806 11.106 30.842 ;
      RECT 10.654 30.806 10.706 30.842 ;
      RECT 10.254 30.806 10.306 30.842 ;
      RECT 9.854 30.806 9.906 30.842 ;
      RECT 9.454 30.806 9.506 30.842 ;
      RECT 9.054 30.806 9.106 30.842 ;
      RECT 8.654 30.806 8.706 30.842 ;
      RECT 8.254 30.806 8.306 30.842 ;
      RECT 7.854 30.806 7.906 30.842 ;
      RECT 7.454 30.806 7.506 30.842 ;
      RECT 7.054 30.806 7.106 30.842 ;
      RECT 6.654 30.806 6.706 30.842 ;
      RECT 6.254 30.806 6.306 30.842 ;
      RECT 5.854 30.806 5.906 30.842 ;
      RECT 5.454 30.806 5.506 30.842 ;
      RECT 5.054 30.806 5.106 30.842 ;
      RECT 4.654 30.806 4.706 30.842 ;
      RECT 4.254 30.806 4.306 30.842 ;
      RECT 3.854 30.806 3.906 30.842 ;
      RECT 3.454 30.806 3.506 30.842 ;
      RECT 3.054 30.806 3.106 30.842 ;
      RECT 2.654 30.806 2.706 30.842 ;
      RECT 2.254 30.806 2.306 30.842 ;
      RECT 1.854 30.806 1.906 30.842 ;
      RECT 1.454 30.806 1.506 30.842 ;
      RECT 1.054 30.806 1.106 30.842 ;
      RECT 0.654 30.806 0.706 30.842 ;
      RECT 21.978 30.582 22.022 30.618 ;
      RECT 21.096 30.582 21.14 30.618 ;
      RECT 14.86 30.582 14.904 30.618 ;
      RECT 13.978 30.582 14.022 30.618 ;
      RECT 35.494 30.358 35.546 30.394 ;
      RECT 35.094 30.358 35.146 30.394 ;
      RECT 34.694 30.358 34.746 30.394 ;
      RECT 34.294 30.358 34.346 30.394 ;
      RECT 33.894 30.358 33.946 30.394 ;
      RECT 33.494 30.358 33.546 30.394 ;
      RECT 33.094 30.358 33.146 30.394 ;
      RECT 32.694 30.358 32.746 30.394 ;
      RECT 32.294 30.358 32.346 30.394 ;
      RECT 31.894 30.358 31.946 30.394 ;
      RECT 31.494 30.358 31.546 30.394 ;
      RECT 31.094 30.358 31.146 30.394 ;
      RECT 30.694 30.358 30.746 30.394 ;
      RECT 30.294 30.358 30.346 30.394 ;
      RECT 29.894 30.358 29.946 30.394 ;
      RECT 29.494 30.358 29.546 30.394 ;
      RECT 29.094 30.358 29.146 30.394 ;
      RECT 28.694 30.358 28.746 30.394 ;
      RECT 28.294 30.358 28.346 30.394 ;
      RECT 27.894 30.358 27.946 30.394 ;
      RECT 27.494 30.358 27.546 30.394 ;
      RECT 27.094 30.358 27.146 30.394 ;
      RECT 26.694 30.358 26.746 30.394 ;
      RECT 26.294 30.358 26.346 30.394 ;
      RECT 25.894 30.358 25.946 30.394 ;
      RECT 25.494 30.358 25.546 30.394 ;
      RECT 25.094 30.358 25.146 30.394 ;
      RECT 24.694 30.358 24.746 30.394 ;
      RECT 24.294 30.358 24.346 30.394 ;
      RECT 23.894 30.358 23.946 30.394 ;
      RECT 23.494 30.358 23.546 30.394 ;
      RECT 23.094 30.358 23.146 30.394 ;
      RECT 21.814 30.358 21.868 30.394 ;
      RECT 19.838 30.358 19.886 30.394 ;
      RECT 19.53 30.358 19.578 30.394 ;
      RECT 16.882 30.358 16.936 30.394 ;
      RECT 16.422 30.358 16.47 30.394 ;
      RECT 16.114 30.358 16.162 30.394 ;
      RECT 14.132 30.358 14.186 30.394 ;
      RECT 13.294 30.358 13.346 30.394 ;
      RECT 12.894 30.358 12.946 30.394 ;
      RECT 12.494 30.358 12.546 30.394 ;
      RECT 12.094 30.358 12.146 30.394 ;
      RECT 11.694 30.358 11.746 30.394 ;
      RECT 11.294 30.358 11.346 30.394 ;
      RECT 10.894 30.358 10.946 30.394 ;
      RECT 10.494 30.358 10.546 30.394 ;
      RECT 10.094 30.358 10.146 30.394 ;
      RECT 9.694 30.358 9.746 30.394 ;
      RECT 9.294 30.358 9.346 30.394 ;
      RECT 8.894 30.358 8.946 30.394 ;
      RECT 8.494 30.358 8.546 30.394 ;
      RECT 8.094 30.358 8.146 30.394 ;
      RECT 7.694 30.358 7.746 30.394 ;
      RECT 7.294 30.358 7.346 30.394 ;
      RECT 6.894 30.358 6.946 30.394 ;
      RECT 6.494 30.358 6.546 30.394 ;
      RECT 6.094 30.358 6.146 30.394 ;
      RECT 5.694 30.358 5.746 30.394 ;
      RECT 5.294 30.358 5.346 30.394 ;
      RECT 4.894 30.358 4.946 30.394 ;
      RECT 4.494 30.358 4.546 30.394 ;
      RECT 4.094 30.358 4.146 30.394 ;
      RECT 3.694 30.358 3.746 30.394 ;
      RECT 3.294 30.358 3.346 30.394 ;
      RECT 2.894 30.358 2.946 30.394 ;
      RECT 2.494 30.358 2.546 30.394 ;
      RECT 2.094 30.358 2.146 30.394 ;
      RECT 1.694 30.358 1.746 30.394 ;
      RECT 1.294 30.358 1.346 30.394 ;
      RECT 0.894 30.358 0.946 30.394 ;
      RECT 21.414 30.282 21.468 30.318 ;
      RECT 14.532 30.282 14.586 30.318 ;
      RECT 19.606 30.129 19.654 30.165 ;
      RECT 18.08 30.129 18.12 30.165 ;
      RECT 16.718 30.129 16.772 30.165 ;
      RECT 16.346 30.129 16.394 30.165 ;
      RECT 20.37 30.1345 20.442 30.1595 ;
      RECT 18.764 30.1345 18.836 30.1595 ;
      RECT 15.558 30.1345 15.63 30.1595 ;
      RECT 21.978 29.982 22.022 30.018 ;
      RECT 13.978 29.982 14.022 30.018 ;
      RECT 18.764 29.9875 18.836 30.0125 ;
      RECT 19.762 29.835 19.81 29.871 ;
      RECT 17.616 29.835 17.656 29.871 ;
      RECT 16.19 29.835 16.238 29.871 ;
      RECT 35.254 29.606 35.306 29.642 ;
      RECT 34.854 29.606 34.906 29.642 ;
      RECT 34.454 29.606 34.506 29.642 ;
      RECT 34.054 29.606 34.106 29.642 ;
      RECT 33.654 29.606 33.706 29.642 ;
      RECT 33.254 29.606 33.306 29.642 ;
      RECT 32.854 29.606 32.906 29.642 ;
      RECT 32.454 29.606 32.506 29.642 ;
      RECT 32.054 29.606 32.106 29.642 ;
      RECT 31.654 29.606 31.706 29.642 ;
      RECT 31.254 29.606 31.306 29.642 ;
      RECT 30.854 29.606 30.906 29.642 ;
      RECT 30.454 29.606 30.506 29.642 ;
      RECT 30.054 29.606 30.106 29.642 ;
      RECT 29.654 29.606 29.706 29.642 ;
      RECT 29.254 29.606 29.306 29.642 ;
      RECT 28.854 29.606 28.906 29.642 ;
      RECT 28.454 29.606 28.506 29.642 ;
      RECT 28.054 29.606 28.106 29.642 ;
      RECT 27.654 29.606 27.706 29.642 ;
      RECT 27.254 29.606 27.306 29.642 ;
      RECT 26.854 29.606 26.906 29.642 ;
      RECT 26.454 29.606 26.506 29.642 ;
      RECT 26.054 29.606 26.106 29.642 ;
      RECT 25.654 29.606 25.706 29.642 ;
      RECT 25.254 29.606 25.306 29.642 ;
      RECT 24.854 29.606 24.906 29.642 ;
      RECT 24.454 29.606 24.506 29.642 ;
      RECT 24.054 29.606 24.106 29.642 ;
      RECT 23.654 29.606 23.706 29.642 ;
      RECT 23.254 29.606 23.306 29.642 ;
      RECT 22.854 29.606 22.906 29.642 ;
      RECT 22.694 29.606 22.746 29.642 ;
      RECT 21.732 29.606 21.786 29.642 ;
      RECT 14.214 29.606 14.268 29.642 ;
      RECT 13.054 29.606 13.106 29.642 ;
      RECT 12.654 29.606 12.706 29.642 ;
      RECT 12.254 29.606 12.306 29.642 ;
      RECT 11.854 29.606 11.906 29.642 ;
      RECT 11.454 29.606 11.506 29.642 ;
      RECT 11.054 29.606 11.106 29.642 ;
      RECT 10.654 29.606 10.706 29.642 ;
      RECT 10.254 29.606 10.306 29.642 ;
      RECT 9.854 29.606 9.906 29.642 ;
      RECT 9.454 29.606 9.506 29.642 ;
      RECT 9.054 29.606 9.106 29.642 ;
      RECT 8.654 29.606 8.706 29.642 ;
      RECT 8.254 29.606 8.306 29.642 ;
      RECT 7.854 29.606 7.906 29.642 ;
      RECT 7.454 29.606 7.506 29.642 ;
      RECT 7.054 29.606 7.106 29.642 ;
      RECT 6.654 29.606 6.706 29.642 ;
      RECT 6.254 29.606 6.306 29.642 ;
      RECT 5.854 29.606 5.906 29.642 ;
      RECT 5.454 29.606 5.506 29.642 ;
      RECT 5.054 29.606 5.106 29.642 ;
      RECT 4.654 29.606 4.706 29.642 ;
      RECT 4.254 29.606 4.306 29.642 ;
      RECT 3.854 29.606 3.906 29.642 ;
      RECT 3.454 29.606 3.506 29.642 ;
      RECT 3.054 29.606 3.106 29.642 ;
      RECT 2.654 29.606 2.706 29.642 ;
      RECT 2.254 29.606 2.306 29.642 ;
      RECT 1.854 29.606 1.906 29.642 ;
      RECT 1.454 29.606 1.506 29.642 ;
      RECT 1.054 29.606 1.106 29.642 ;
      RECT 0.654 29.606 0.706 29.642 ;
      RECT 21.978 29.382 22.022 29.418 ;
      RECT 21.096 29.382 21.14 29.418 ;
      RECT 14.86 29.382 14.904 29.418 ;
      RECT 13.978 29.382 14.022 29.418 ;
      RECT 35.494 29.158 35.546 29.194 ;
      RECT 35.094 29.158 35.146 29.194 ;
      RECT 34.694 29.158 34.746 29.194 ;
      RECT 34.294 29.158 34.346 29.194 ;
      RECT 33.894 29.158 33.946 29.194 ;
      RECT 33.494 29.158 33.546 29.194 ;
      RECT 33.094 29.158 33.146 29.194 ;
      RECT 32.694 29.158 32.746 29.194 ;
      RECT 32.294 29.158 32.346 29.194 ;
      RECT 31.894 29.158 31.946 29.194 ;
      RECT 31.494 29.158 31.546 29.194 ;
      RECT 31.094 29.158 31.146 29.194 ;
      RECT 30.694 29.158 30.746 29.194 ;
      RECT 30.294 29.158 30.346 29.194 ;
      RECT 29.894 29.158 29.946 29.194 ;
      RECT 29.494 29.158 29.546 29.194 ;
      RECT 29.094 29.158 29.146 29.194 ;
      RECT 28.694 29.158 28.746 29.194 ;
      RECT 28.294 29.158 28.346 29.194 ;
      RECT 27.894 29.158 27.946 29.194 ;
      RECT 27.494 29.158 27.546 29.194 ;
      RECT 27.094 29.158 27.146 29.194 ;
      RECT 26.694 29.158 26.746 29.194 ;
      RECT 26.294 29.158 26.346 29.194 ;
      RECT 25.894 29.158 25.946 29.194 ;
      RECT 25.494 29.158 25.546 29.194 ;
      RECT 25.094 29.158 25.146 29.194 ;
      RECT 24.694 29.158 24.746 29.194 ;
      RECT 24.294 29.158 24.346 29.194 ;
      RECT 23.894 29.158 23.946 29.194 ;
      RECT 23.494 29.158 23.546 29.194 ;
      RECT 23.094 29.158 23.146 29.194 ;
      RECT 21.814 29.158 21.868 29.194 ;
      RECT 19.838 29.158 19.886 29.194 ;
      RECT 19.53 29.158 19.578 29.194 ;
      RECT 16.882 29.158 16.936 29.194 ;
      RECT 16.422 29.158 16.47 29.194 ;
      RECT 16.114 29.158 16.162 29.194 ;
      RECT 14.132 29.158 14.186 29.194 ;
      RECT 13.294 29.158 13.346 29.194 ;
      RECT 12.894 29.158 12.946 29.194 ;
      RECT 12.494 29.158 12.546 29.194 ;
      RECT 12.094 29.158 12.146 29.194 ;
      RECT 11.694 29.158 11.746 29.194 ;
      RECT 11.294 29.158 11.346 29.194 ;
      RECT 10.894 29.158 10.946 29.194 ;
      RECT 10.494 29.158 10.546 29.194 ;
      RECT 10.094 29.158 10.146 29.194 ;
      RECT 9.694 29.158 9.746 29.194 ;
      RECT 9.294 29.158 9.346 29.194 ;
      RECT 8.894 29.158 8.946 29.194 ;
      RECT 8.494 29.158 8.546 29.194 ;
      RECT 8.094 29.158 8.146 29.194 ;
      RECT 7.694 29.158 7.746 29.194 ;
      RECT 7.294 29.158 7.346 29.194 ;
      RECT 6.894 29.158 6.946 29.194 ;
      RECT 6.494 29.158 6.546 29.194 ;
      RECT 6.094 29.158 6.146 29.194 ;
      RECT 5.694 29.158 5.746 29.194 ;
      RECT 5.294 29.158 5.346 29.194 ;
      RECT 4.894 29.158 4.946 29.194 ;
      RECT 4.494 29.158 4.546 29.194 ;
      RECT 4.094 29.158 4.146 29.194 ;
      RECT 3.694 29.158 3.746 29.194 ;
      RECT 3.294 29.158 3.346 29.194 ;
      RECT 2.894 29.158 2.946 29.194 ;
      RECT 2.494 29.158 2.546 29.194 ;
      RECT 2.094 29.158 2.146 29.194 ;
      RECT 1.694 29.158 1.746 29.194 ;
      RECT 1.294 29.158 1.346 29.194 ;
      RECT 0.894 29.158 0.946 29.194 ;
      RECT 21.414 29.082 21.468 29.118 ;
      RECT 14.532 29.082 14.586 29.118 ;
      RECT 19.606 28.929 19.654 28.965 ;
      RECT 18.08 28.929 18.12 28.965 ;
      RECT 16.718 28.929 16.772 28.965 ;
      RECT 16.346 28.929 16.394 28.965 ;
      RECT 20.37 28.9345 20.442 28.9595 ;
      RECT 18.764 28.9345 18.836 28.9595 ;
      RECT 15.558 28.9345 15.63 28.9595 ;
      RECT 21.978 28.782 22.022 28.818 ;
      RECT 13.978 28.782 14.022 28.818 ;
      RECT 18.764 28.7875 18.836 28.8125 ;
      RECT 19.762 28.635 19.81 28.671 ;
      RECT 17.616 28.635 17.656 28.671 ;
      RECT 16.19 28.635 16.238 28.671 ;
      RECT 35.254 28.406 35.306 28.442 ;
      RECT 34.854 28.406 34.906 28.442 ;
      RECT 34.454 28.406 34.506 28.442 ;
      RECT 34.054 28.406 34.106 28.442 ;
      RECT 33.654 28.406 33.706 28.442 ;
      RECT 33.254 28.406 33.306 28.442 ;
      RECT 32.854 28.406 32.906 28.442 ;
      RECT 32.454 28.406 32.506 28.442 ;
      RECT 32.054 28.406 32.106 28.442 ;
      RECT 31.654 28.406 31.706 28.442 ;
      RECT 31.254 28.406 31.306 28.442 ;
      RECT 30.854 28.406 30.906 28.442 ;
      RECT 30.454 28.406 30.506 28.442 ;
      RECT 30.054 28.406 30.106 28.442 ;
      RECT 29.654 28.406 29.706 28.442 ;
      RECT 29.254 28.406 29.306 28.442 ;
      RECT 28.854 28.406 28.906 28.442 ;
      RECT 28.454 28.406 28.506 28.442 ;
      RECT 28.054 28.406 28.106 28.442 ;
      RECT 27.654 28.406 27.706 28.442 ;
      RECT 27.254 28.406 27.306 28.442 ;
      RECT 26.854 28.406 26.906 28.442 ;
      RECT 26.454 28.406 26.506 28.442 ;
      RECT 26.054 28.406 26.106 28.442 ;
      RECT 25.654 28.406 25.706 28.442 ;
      RECT 25.254 28.406 25.306 28.442 ;
      RECT 24.854 28.406 24.906 28.442 ;
      RECT 24.454 28.406 24.506 28.442 ;
      RECT 24.054 28.406 24.106 28.442 ;
      RECT 23.654 28.406 23.706 28.442 ;
      RECT 23.254 28.406 23.306 28.442 ;
      RECT 22.854 28.406 22.906 28.442 ;
      RECT 22.694 28.406 22.746 28.442 ;
      RECT 21.732 28.406 21.786 28.442 ;
      RECT 14.214 28.406 14.268 28.442 ;
      RECT 13.054 28.406 13.106 28.442 ;
      RECT 12.654 28.406 12.706 28.442 ;
      RECT 12.254 28.406 12.306 28.442 ;
      RECT 11.854 28.406 11.906 28.442 ;
      RECT 11.454 28.406 11.506 28.442 ;
      RECT 11.054 28.406 11.106 28.442 ;
      RECT 10.654 28.406 10.706 28.442 ;
      RECT 10.254 28.406 10.306 28.442 ;
      RECT 9.854 28.406 9.906 28.442 ;
      RECT 9.454 28.406 9.506 28.442 ;
      RECT 9.054 28.406 9.106 28.442 ;
      RECT 8.654 28.406 8.706 28.442 ;
      RECT 8.254 28.406 8.306 28.442 ;
      RECT 7.854 28.406 7.906 28.442 ;
      RECT 7.454 28.406 7.506 28.442 ;
      RECT 7.054 28.406 7.106 28.442 ;
      RECT 6.654 28.406 6.706 28.442 ;
      RECT 6.254 28.406 6.306 28.442 ;
      RECT 5.854 28.406 5.906 28.442 ;
      RECT 5.454 28.406 5.506 28.442 ;
      RECT 5.054 28.406 5.106 28.442 ;
      RECT 4.654 28.406 4.706 28.442 ;
      RECT 4.254 28.406 4.306 28.442 ;
      RECT 3.854 28.406 3.906 28.442 ;
      RECT 3.454 28.406 3.506 28.442 ;
      RECT 3.054 28.406 3.106 28.442 ;
      RECT 2.654 28.406 2.706 28.442 ;
      RECT 2.254 28.406 2.306 28.442 ;
      RECT 1.854 28.406 1.906 28.442 ;
      RECT 1.454 28.406 1.506 28.442 ;
      RECT 1.054 28.406 1.106 28.442 ;
      RECT 0.654 28.406 0.706 28.442 ;
      RECT 21.978 28.182 22.022 28.218 ;
      RECT 21.096 28.182 21.14 28.218 ;
      RECT 14.86 28.182 14.904 28.218 ;
      RECT 13.978 28.182 14.022 28.218 ;
      RECT 35.494 27.958 35.546 27.994 ;
      RECT 35.094 27.958 35.146 27.994 ;
      RECT 34.694 27.958 34.746 27.994 ;
      RECT 34.294 27.958 34.346 27.994 ;
      RECT 33.894 27.958 33.946 27.994 ;
      RECT 33.494 27.958 33.546 27.994 ;
      RECT 33.094 27.958 33.146 27.994 ;
      RECT 32.694 27.958 32.746 27.994 ;
      RECT 32.294 27.958 32.346 27.994 ;
      RECT 31.894 27.958 31.946 27.994 ;
      RECT 31.494 27.958 31.546 27.994 ;
      RECT 31.094 27.958 31.146 27.994 ;
      RECT 30.694 27.958 30.746 27.994 ;
      RECT 30.294 27.958 30.346 27.994 ;
      RECT 29.894 27.958 29.946 27.994 ;
      RECT 29.494 27.958 29.546 27.994 ;
      RECT 29.094 27.958 29.146 27.994 ;
      RECT 28.694 27.958 28.746 27.994 ;
      RECT 28.294 27.958 28.346 27.994 ;
      RECT 27.894 27.958 27.946 27.994 ;
      RECT 27.494 27.958 27.546 27.994 ;
      RECT 27.094 27.958 27.146 27.994 ;
      RECT 26.694 27.958 26.746 27.994 ;
      RECT 26.294 27.958 26.346 27.994 ;
      RECT 25.894 27.958 25.946 27.994 ;
      RECT 25.494 27.958 25.546 27.994 ;
      RECT 25.094 27.958 25.146 27.994 ;
      RECT 24.694 27.958 24.746 27.994 ;
      RECT 24.294 27.958 24.346 27.994 ;
      RECT 23.894 27.958 23.946 27.994 ;
      RECT 23.494 27.958 23.546 27.994 ;
      RECT 23.094 27.958 23.146 27.994 ;
      RECT 21.814 27.958 21.868 27.994 ;
      RECT 19.838 27.958 19.886 27.994 ;
      RECT 19.53 27.958 19.578 27.994 ;
      RECT 16.882 27.958 16.936 27.994 ;
      RECT 16.422 27.958 16.47 27.994 ;
      RECT 16.114 27.958 16.162 27.994 ;
      RECT 14.132 27.958 14.186 27.994 ;
      RECT 13.294 27.958 13.346 27.994 ;
      RECT 12.894 27.958 12.946 27.994 ;
      RECT 12.494 27.958 12.546 27.994 ;
      RECT 12.094 27.958 12.146 27.994 ;
      RECT 11.694 27.958 11.746 27.994 ;
      RECT 11.294 27.958 11.346 27.994 ;
      RECT 10.894 27.958 10.946 27.994 ;
      RECT 10.494 27.958 10.546 27.994 ;
      RECT 10.094 27.958 10.146 27.994 ;
      RECT 9.694 27.958 9.746 27.994 ;
      RECT 9.294 27.958 9.346 27.994 ;
      RECT 8.894 27.958 8.946 27.994 ;
      RECT 8.494 27.958 8.546 27.994 ;
      RECT 8.094 27.958 8.146 27.994 ;
      RECT 7.694 27.958 7.746 27.994 ;
      RECT 7.294 27.958 7.346 27.994 ;
      RECT 6.894 27.958 6.946 27.994 ;
      RECT 6.494 27.958 6.546 27.994 ;
      RECT 6.094 27.958 6.146 27.994 ;
      RECT 5.694 27.958 5.746 27.994 ;
      RECT 5.294 27.958 5.346 27.994 ;
      RECT 4.894 27.958 4.946 27.994 ;
      RECT 4.494 27.958 4.546 27.994 ;
      RECT 4.094 27.958 4.146 27.994 ;
      RECT 3.694 27.958 3.746 27.994 ;
      RECT 3.294 27.958 3.346 27.994 ;
      RECT 2.894 27.958 2.946 27.994 ;
      RECT 2.494 27.958 2.546 27.994 ;
      RECT 2.094 27.958 2.146 27.994 ;
      RECT 1.694 27.958 1.746 27.994 ;
      RECT 1.294 27.958 1.346 27.994 ;
      RECT 0.894 27.958 0.946 27.994 ;
      RECT 21.414 27.882 21.468 27.918 ;
      RECT 14.532 27.882 14.586 27.918 ;
      RECT 19.606 27.729 19.654 27.765 ;
      RECT 18.08 27.729 18.12 27.765 ;
      RECT 16.718 27.729 16.772 27.765 ;
      RECT 16.346 27.729 16.394 27.765 ;
      RECT 20.37 27.7345 20.442 27.7595 ;
      RECT 18.764 27.7345 18.836 27.7595 ;
      RECT 15.558 27.7345 15.63 27.7595 ;
      RECT 21.978 27.582 22.022 27.618 ;
      RECT 13.978 27.582 14.022 27.618 ;
      RECT 18.764 27.5875 18.836 27.6125 ;
      RECT 19.762 27.435 19.81 27.471 ;
      RECT 17.616 27.435 17.656 27.471 ;
      RECT 16.19 27.435 16.238 27.471 ;
      RECT 35.254 27.206 35.306 27.242 ;
      RECT 34.854 27.206 34.906 27.242 ;
      RECT 34.454 27.206 34.506 27.242 ;
      RECT 34.054 27.206 34.106 27.242 ;
      RECT 33.654 27.206 33.706 27.242 ;
      RECT 33.254 27.206 33.306 27.242 ;
      RECT 32.854 27.206 32.906 27.242 ;
      RECT 32.454 27.206 32.506 27.242 ;
      RECT 32.054 27.206 32.106 27.242 ;
      RECT 31.654 27.206 31.706 27.242 ;
      RECT 31.254 27.206 31.306 27.242 ;
      RECT 30.854 27.206 30.906 27.242 ;
      RECT 30.454 27.206 30.506 27.242 ;
      RECT 30.054 27.206 30.106 27.242 ;
      RECT 29.654 27.206 29.706 27.242 ;
      RECT 29.254 27.206 29.306 27.242 ;
      RECT 28.854 27.206 28.906 27.242 ;
      RECT 28.454 27.206 28.506 27.242 ;
      RECT 28.054 27.206 28.106 27.242 ;
      RECT 27.654 27.206 27.706 27.242 ;
      RECT 27.254 27.206 27.306 27.242 ;
      RECT 26.854 27.206 26.906 27.242 ;
      RECT 26.454 27.206 26.506 27.242 ;
      RECT 26.054 27.206 26.106 27.242 ;
      RECT 25.654 27.206 25.706 27.242 ;
      RECT 25.254 27.206 25.306 27.242 ;
      RECT 24.854 27.206 24.906 27.242 ;
      RECT 24.454 27.206 24.506 27.242 ;
      RECT 24.054 27.206 24.106 27.242 ;
      RECT 23.654 27.206 23.706 27.242 ;
      RECT 23.254 27.206 23.306 27.242 ;
      RECT 22.854 27.206 22.906 27.242 ;
      RECT 22.694 27.206 22.746 27.242 ;
      RECT 21.732 27.206 21.786 27.242 ;
      RECT 14.214 27.206 14.268 27.242 ;
      RECT 13.054 27.206 13.106 27.242 ;
      RECT 12.654 27.206 12.706 27.242 ;
      RECT 12.254 27.206 12.306 27.242 ;
      RECT 11.854 27.206 11.906 27.242 ;
      RECT 11.454 27.206 11.506 27.242 ;
      RECT 11.054 27.206 11.106 27.242 ;
      RECT 10.654 27.206 10.706 27.242 ;
      RECT 10.254 27.206 10.306 27.242 ;
      RECT 9.854 27.206 9.906 27.242 ;
      RECT 9.454 27.206 9.506 27.242 ;
      RECT 9.054 27.206 9.106 27.242 ;
      RECT 8.654 27.206 8.706 27.242 ;
      RECT 8.254 27.206 8.306 27.242 ;
      RECT 7.854 27.206 7.906 27.242 ;
      RECT 7.454 27.206 7.506 27.242 ;
      RECT 7.054 27.206 7.106 27.242 ;
      RECT 6.654 27.206 6.706 27.242 ;
      RECT 6.254 27.206 6.306 27.242 ;
      RECT 5.854 27.206 5.906 27.242 ;
      RECT 5.454 27.206 5.506 27.242 ;
      RECT 5.054 27.206 5.106 27.242 ;
      RECT 4.654 27.206 4.706 27.242 ;
      RECT 4.254 27.206 4.306 27.242 ;
      RECT 3.854 27.206 3.906 27.242 ;
      RECT 3.454 27.206 3.506 27.242 ;
      RECT 3.054 27.206 3.106 27.242 ;
      RECT 2.654 27.206 2.706 27.242 ;
      RECT 2.254 27.206 2.306 27.242 ;
      RECT 1.854 27.206 1.906 27.242 ;
      RECT 1.454 27.206 1.506 27.242 ;
      RECT 1.054 27.206 1.106 27.242 ;
      RECT 0.654 27.206 0.706 27.242 ;
      RECT 21.978 26.982 22.022 27.018 ;
      RECT 21.096 26.982 21.14 27.018 ;
      RECT 14.86 26.982 14.904 27.018 ;
      RECT 13.978 26.982 14.022 27.018 ;
      RECT 35.494 26.758 35.546 26.794 ;
      RECT 35.094 26.758 35.146 26.794 ;
      RECT 34.694 26.758 34.746 26.794 ;
      RECT 34.294 26.758 34.346 26.794 ;
      RECT 33.894 26.758 33.946 26.794 ;
      RECT 33.494 26.758 33.546 26.794 ;
      RECT 33.094 26.758 33.146 26.794 ;
      RECT 32.694 26.758 32.746 26.794 ;
      RECT 32.294 26.758 32.346 26.794 ;
      RECT 31.894 26.758 31.946 26.794 ;
      RECT 31.494 26.758 31.546 26.794 ;
      RECT 31.094 26.758 31.146 26.794 ;
      RECT 30.694 26.758 30.746 26.794 ;
      RECT 30.294 26.758 30.346 26.794 ;
      RECT 29.894 26.758 29.946 26.794 ;
      RECT 29.494 26.758 29.546 26.794 ;
      RECT 29.094 26.758 29.146 26.794 ;
      RECT 28.694 26.758 28.746 26.794 ;
      RECT 28.294 26.758 28.346 26.794 ;
      RECT 27.894 26.758 27.946 26.794 ;
      RECT 27.494 26.758 27.546 26.794 ;
      RECT 27.094 26.758 27.146 26.794 ;
      RECT 26.694 26.758 26.746 26.794 ;
      RECT 26.294 26.758 26.346 26.794 ;
      RECT 25.894 26.758 25.946 26.794 ;
      RECT 25.494 26.758 25.546 26.794 ;
      RECT 25.094 26.758 25.146 26.794 ;
      RECT 24.694 26.758 24.746 26.794 ;
      RECT 24.294 26.758 24.346 26.794 ;
      RECT 23.894 26.758 23.946 26.794 ;
      RECT 23.494 26.758 23.546 26.794 ;
      RECT 23.094 26.758 23.146 26.794 ;
      RECT 21.814 26.758 21.868 26.794 ;
      RECT 19.838 26.758 19.886 26.794 ;
      RECT 19.53 26.758 19.578 26.794 ;
      RECT 16.882 26.758 16.936 26.794 ;
      RECT 16.422 26.758 16.47 26.794 ;
      RECT 16.114 26.758 16.162 26.794 ;
      RECT 14.132 26.758 14.186 26.794 ;
      RECT 13.294 26.758 13.346 26.794 ;
      RECT 12.894 26.758 12.946 26.794 ;
      RECT 12.494 26.758 12.546 26.794 ;
      RECT 12.094 26.758 12.146 26.794 ;
      RECT 11.694 26.758 11.746 26.794 ;
      RECT 11.294 26.758 11.346 26.794 ;
      RECT 10.894 26.758 10.946 26.794 ;
      RECT 10.494 26.758 10.546 26.794 ;
      RECT 10.094 26.758 10.146 26.794 ;
      RECT 9.694 26.758 9.746 26.794 ;
      RECT 9.294 26.758 9.346 26.794 ;
      RECT 8.894 26.758 8.946 26.794 ;
      RECT 8.494 26.758 8.546 26.794 ;
      RECT 8.094 26.758 8.146 26.794 ;
      RECT 7.694 26.758 7.746 26.794 ;
      RECT 7.294 26.758 7.346 26.794 ;
      RECT 6.894 26.758 6.946 26.794 ;
      RECT 6.494 26.758 6.546 26.794 ;
      RECT 6.094 26.758 6.146 26.794 ;
      RECT 5.694 26.758 5.746 26.794 ;
      RECT 5.294 26.758 5.346 26.794 ;
      RECT 4.894 26.758 4.946 26.794 ;
      RECT 4.494 26.758 4.546 26.794 ;
      RECT 4.094 26.758 4.146 26.794 ;
      RECT 3.694 26.758 3.746 26.794 ;
      RECT 3.294 26.758 3.346 26.794 ;
      RECT 2.894 26.758 2.946 26.794 ;
      RECT 2.494 26.758 2.546 26.794 ;
      RECT 2.094 26.758 2.146 26.794 ;
      RECT 1.694 26.758 1.746 26.794 ;
      RECT 1.294 26.758 1.346 26.794 ;
      RECT 0.894 26.758 0.946 26.794 ;
      RECT 21.414 26.682 21.468 26.718 ;
      RECT 14.532 26.682 14.586 26.718 ;
      RECT 19.606 26.529 19.654 26.565 ;
      RECT 18.08 26.529 18.12 26.565 ;
      RECT 16.718 26.529 16.772 26.565 ;
      RECT 16.346 26.529 16.394 26.565 ;
      RECT 20.37 26.5345 20.442 26.5595 ;
      RECT 18.764 26.5345 18.836 26.5595 ;
      RECT 15.558 26.5345 15.63 26.5595 ;
      RECT 21.978 26.382 22.022 26.418 ;
      RECT 13.978 26.382 14.022 26.418 ;
      RECT 18.764 26.3875 18.836 26.4125 ;
      RECT 19.762 26.235 19.81 26.271 ;
      RECT 17.616 26.235 17.656 26.271 ;
      RECT 16.19 26.235 16.238 26.271 ;
      RECT 35.254 26.006 35.306 26.042 ;
      RECT 34.854 26.006 34.906 26.042 ;
      RECT 34.454 26.006 34.506 26.042 ;
      RECT 34.054 26.006 34.106 26.042 ;
      RECT 33.654 26.006 33.706 26.042 ;
      RECT 33.254 26.006 33.306 26.042 ;
      RECT 32.854 26.006 32.906 26.042 ;
      RECT 32.454 26.006 32.506 26.042 ;
      RECT 32.054 26.006 32.106 26.042 ;
      RECT 31.654 26.006 31.706 26.042 ;
      RECT 31.254 26.006 31.306 26.042 ;
      RECT 30.854 26.006 30.906 26.042 ;
      RECT 30.454 26.006 30.506 26.042 ;
      RECT 30.054 26.006 30.106 26.042 ;
      RECT 29.654 26.006 29.706 26.042 ;
      RECT 29.254 26.006 29.306 26.042 ;
      RECT 28.854 26.006 28.906 26.042 ;
      RECT 28.454 26.006 28.506 26.042 ;
      RECT 28.054 26.006 28.106 26.042 ;
      RECT 27.654 26.006 27.706 26.042 ;
      RECT 27.254 26.006 27.306 26.042 ;
      RECT 26.854 26.006 26.906 26.042 ;
      RECT 26.454 26.006 26.506 26.042 ;
      RECT 26.054 26.006 26.106 26.042 ;
      RECT 25.654 26.006 25.706 26.042 ;
      RECT 25.254 26.006 25.306 26.042 ;
      RECT 24.854 26.006 24.906 26.042 ;
      RECT 24.454 26.006 24.506 26.042 ;
      RECT 24.054 26.006 24.106 26.042 ;
      RECT 23.654 26.006 23.706 26.042 ;
      RECT 23.254 26.006 23.306 26.042 ;
      RECT 22.854 26.006 22.906 26.042 ;
      RECT 22.694 26.006 22.746 26.042 ;
      RECT 21.732 26.006 21.786 26.042 ;
      RECT 14.214 26.006 14.268 26.042 ;
      RECT 13.054 26.006 13.106 26.042 ;
      RECT 12.654 26.006 12.706 26.042 ;
      RECT 12.254 26.006 12.306 26.042 ;
      RECT 11.854 26.006 11.906 26.042 ;
      RECT 11.454 26.006 11.506 26.042 ;
      RECT 11.054 26.006 11.106 26.042 ;
      RECT 10.654 26.006 10.706 26.042 ;
      RECT 10.254 26.006 10.306 26.042 ;
      RECT 9.854 26.006 9.906 26.042 ;
      RECT 9.454 26.006 9.506 26.042 ;
      RECT 9.054 26.006 9.106 26.042 ;
      RECT 8.654 26.006 8.706 26.042 ;
      RECT 8.254 26.006 8.306 26.042 ;
      RECT 7.854 26.006 7.906 26.042 ;
      RECT 7.454 26.006 7.506 26.042 ;
      RECT 7.054 26.006 7.106 26.042 ;
      RECT 6.654 26.006 6.706 26.042 ;
      RECT 6.254 26.006 6.306 26.042 ;
      RECT 5.854 26.006 5.906 26.042 ;
      RECT 5.454 26.006 5.506 26.042 ;
      RECT 5.054 26.006 5.106 26.042 ;
      RECT 4.654 26.006 4.706 26.042 ;
      RECT 4.254 26.006 4.306 26.042 ;
      RECT 3.854 26.006 3.906 26.042 ;
      RECT 3.454 26.006 3.506 26.042 ;
      RECT 3.054 26.006 3.106 26.042 ;
      RECT 2.654 26.006 2.706 26.042 ;
      RECT 2.254 26.006 2.306 26.042 ;
      RECT 1.854 26.006 1.906 26.042 ;
      RECT 1.454 26.006 1.506 26.042 ;
      RECT 1.054 26.006 1.106 26.042 ;
      RECT 0.654 26.006 0.706 26.042 ;
      RECT 21.978 25.782 22.022 25.818 ;
      RECT 21.096 25.782 21.14 25.818 ;
      RECT 14.86 25.782 14.904 25.818 ;
      RECT 13.978 25.782 14.022 25.818 ;
      RECT 35.494 25.558 35.546 25.594 ;
      RECT 35.094 25.558 35.146 25.594 ;
      RECT 34.694 25.558 34.746 25.594 ;
      RECT 34.294 25.558 34.346 25.594 ;
      RECT 33.894 25.558 33.946 25.594 ;
      RECT 33.494 25.558 33.546 25.594 ;
      RECT 33.094 25.558 33.146 25.594 ;
      RECT 32.694 25.558 32.746 25.594 ;
      RECT 32.294 25.558 32.346 25.594 ;
      RECT 31.894 25.558 31.946 25.594 ;
      RECT 31.494 25.558 31.546 25.594 ;
      RECT 31.094 25.558 31.146 25.594 ;
      RECT 30.694 25.558 30.746 25.594 ;
      RECT 30.294 25.558 30.346 25.594 ;
      RECT 29.894 25.558 29.946 25.594 ;
      RECT 29.494 25.558 29.546 25.594 ;
      RECT 29.094 25.558 29.146 25.594 ;
      RECT 28.694 25.558 28.746 25.594 ;
      RECT 28.294 25.558 28.346 25.594 ;
      RECT 27.894 25.558 27.946 25.594 ;
      RECT 27.494 25.558 27.546 25.594 ;
      RECT 27.094 25.558 27.146 25.594 ;
      RECT 26.694 25.558 26.746 25.594 ;
      RECT 26.294 25.558 26.346 25.594 ;
      RECT 25.894 25.558 25.946 25.594 ;
      RECT 25.494 25.558 25.546 25.594 ;
      RECT 25.094 25.558 25.146 25.594 ;
      RECT 24.694 25.558 24.746 25.594 ;
      RECT 24.294 25.558 24.346 25.594 ;
      RECT 23.894 25.558 23.946 25.594 ;
      RECT 23.494 25.558 23.546 25.594 ;
      RECT 23.094 25.558 23.146 25.594 ;
      RECT 21.814 25.558 21.868 25.594 ;
      RECT 19.838 25.558 19.886 25.594 ;
      RECT 19.53 25.558 19.578 25.594 ;
      RECT 16.882 25.558 16.936 25.594 ;
      RECT 16.422 25.558 16.47 25.594 ;
      RECT 16.114 25.558 16.162 25.594 ;
      RECT 14.132 25.558 14.186 25.594 ;
      RECT 13.294 25.558 13.346 25.594 ;
      RECT 12.894 25.558 12.946 25.594 ;
      RECT 12.494 25.558 12.546 25.594 ;
      RECT 12.094 25.558 12.146 25.594 ;
      RECT 11.694 25.558 11.746 25.594 ;
      RECT 11.294 25.558 11.346 25.594 ;
      RECT 10.894 25.558 10.946 25.594 ;
      RECT 10.494 25.558 10.546 25.594 ;
      RECT 10.094 25.558 10.146 25.594 ;
      RECT 9.694 25.558 9.746 25.594 ;
      RECT 9.294 25.558 9.346 25.594 ;
      RECT 8.894 25.558 8.946 25.594 ;
      RECT 8.494 25.558 8.546 25.594 ;
      RECT 8.094 25.558 8.146 25.594 ;
      RECT 7.694 25.558 7.746 25.594 ;
      RECT 7.294 25.558 7.346 25.594 ;
      RECT 6.894 25.558 6.946 25.594 ;
      RECT 6.494 25.558 6.546 25.594 ;
      RECT 6.094 25.558 6.146 25.594 ;
      RECT 5.694 25.558 5.746 25.594 ;
      RECT 5.294 25.558 5.346 25.594 ;
      RECT 4.894 25.558 4.946 25.594 ;
      RECT 4.494 25.558 4.546 25.594 ;
      RECT 4.094 25.558 4.146 25.594 ;
      RECT 3.694 25.558 3.746 25.594 ;
      RECT 3.294 25.558 3.346 25.594 ;
      RECT 2.894 25.558 2.946 25.594 ;
      RECT 2.494 25.558 2.546 25.594 ;
      RECT 2.094 25.558 2.146 25.594 ;
      RECT 1.694 25.558 1.746 25.594 ;
      RECT 1.294 25.558 1.346 25.594 ;
      RECT 0.894 25.558 0.946 25.594 ;
      RECT 21.414 25.482 21.468 25.518 ;
      RECT 14.532 25.482 14.586 25.518 ;
      RECT 19.606 25.329 19.654 25.365 ;
      RECT 18.08 25.329 18.12 25.365 ;
      RECT 16.718 25.329 16.772 25.365 ;
      RECT 16.346 25.329 16.394 25.365 ;
      RECT 20.37 25.3345 20.442 25.3595 ;
      RECT 18.764 25.3345 18.836 25.3595 ;
      RECT 15.558 25.3345 15.63 25.3595 ;
      RECT 21.978 25.182 22.022 25.218 ;
      RECT 13.978 25.182 14.022 25.218 ;
      RECT 18.764 25.1875 18.836 25.2125 ;
      RECT 19.762 25.035 19.81 25.071 ;
      RECT 17.616 25.035 17.656 25.071 ;
      RECT 16.19 25.035 16.238 25.071 ;
      RECT 35.254 24.806 35.306 24.842 ;
      RECT 34.854 24.806 34.906 24.842 ;
      RECT 34.454 24.806 34.506 24.842 ;
      RECT 34.054 24.806 34.106 24.842 ;
      RECT 33.654 24.806 33.706 24.842 ;
      RECT 33.254 24.806 33.306 24.842 ;
      RECT 32.854 24.806 32.906 24.842 ;
      RECT 32.454 24.806 32.506 24.842 ;
      RECT 32.054 24.806 32.106 24.842 ;
      RECT 31.654 24.806 31.706 24.842 ;
      RECT 31.254 24.806 31.306 24.842 ;
      RECT 30.854 24.806 30.906 24.842 ;
      RECT 30.454 24.806 30.506 24.842 ;
      RECT 30.054 24.806 30.106 24.842 ;
      RECT 29.654 24.806 29.706 24.842 ;
      RECT 29.254 24.806 29.306 24.842 ;
      RECT 28.854 24.806 28.906 24.842 ;
      RECT 28.454 24.806 28.506 24.842 ;
      RECT 28.054 24.806 28.106 24.842 ;
      RECT 27.654 24.806 27.706 24.842 ;
      RECT 27.254 24.806 27.306 24.842 ;
      RECT 26.854 24.806 26.906 24.842 ;
      RECT 26.454 24.806 26.506 24.842 ;
      RECT 26.054 24.806 26.106 24.842 ;
      RECT 25.654 24.806 25.706 24.842 ;
      RECT 25.254 24.806 25.306 24.842 ;
      RECT 24.854 24.806 24.906 24.842 ;
      RECT 24.454 24.806 24.506 24.842 ;
      RECT 24.054 24.806 24.106 24.842 ;
      RECT 23.654 24.806 23.706 24.842 ;
      RECT 23.254 24.806 23.306 24.842 ;
      RECT 22.854 24.806 22.906 24.842 ;
      RECT 22.694 24.806 22.746 24.842 ;
      RECT 21.732 24.806 21.786 24.842 ;
      RECT 14.214 24.806 14.268 24.842 ;
      RECT 13.054 24.806 13.106 24.842 ;
      RECT 12.654 24.806 12.706 24.842 ;
      RECT 12.254 24.806 12.306 24.842 ;
      RECT 11.854 24.806 11.906 24.842 ;
      RECT 11.454 24.806 11.506 24.842 ;
      RECT 11.054 24.806 11.106 24.842 ;
      RECT 10.654 24.806 10.706 24.842 ;
      RECT 10.254 24.806 10.306 24.842 ;
      RECT 9.854 24.806 9.906 24.842 ;
      RECT 9.454 24.806 9.506 24.842 ;
      RECT 9.054 24.806 9.106 24.842 ;
      RECT 8.654 24.806 8.706 24.842 ;
      RECT 8.254 24.806 8.306 24.842 ;
      RECT 7.854 24.806 7.906 24.842 ;
      RECT 7.454 24.806 7.506 24.842 ;
      RECT 7.054 24.806 7.106 24.842 ;
      RECT 6.654 24.806 6.706 24.842 ;
      RECT 6.254 24.806 6.306 24.842 ;
      RECT 5.854 24.806 5.906 24.842 ;
      RECT 5.454 24.806 5.506 24.842 ;
      RECT 5.054 24.806 5.106 24.842 ;
      RECT 4.654 24.806 4.706 24.842 ;
      RECT 4.254 24.806 4.306 24.842 ;
      RECT 3.854 24.806 3.906 24.842 ;
      RECT 3.454 24.806 3.506 24.842 ;
      RECT 3.054 24.806 3.106 24.842 ;
      RECT 2.654 24.806 2.706 24.842 ;
      RECT 2.254 24.806 2.306 24.842 ;
      RECT 1.854 24.806 1.906 24.842 ;
      RECT 1.454 24.806 1.506 24.842 ;
      RECT 1.054 24.806 1.106 24.842 ;
      RECT 0.654 24.806 0.706 24.842 ;
      RECT 21.978 24.582 22.022 24.618 ;
      RECT 21.096 24.582 21.14 24.618 ;
      RECT 14.86 24.582 14.904 24.618 ;
      RECT 13.978 24.582 14.022 24.618 ;
      RECT 35.494 24.358 35.546 24.394 ;
      RECT 35.094 24.358 35.146 24.394 ;
      RECT 34.694 24.358 34.746 24.394 ;
      RECT 34.294 24.358 34.346 24.394 ;
      RECT 33.894 24.358 33.946 24.394 ;
      RECT 33.494 24.358 33.546 24.394 ;
      RECT 33.094 24.358 33.146 24.394 ;
      RECT 32.694 24.358 32.746 24.394 ;
      RECT 32.294 24.358 32.346 24.394 ;
      RECT 31.894 24.358 31.946 24.394 ;
      RECT 31.494 24.358 31.546 24.394 ;
      RECT 31.094 24.358 31.146 24.394 ;
      RECT 30.694 24.358 30.746 24.394 ;
      RECT 30.294 24.358 30.346 24.394 ;
      RECT 29.894 24.358 29.946 24.394 ;
      RECT 29.494 24.358 29.546 24.394 ;
      RECT 29.094 24.358 29.146 24.394 ;
      RECT 28.694 24.358 28.746 24.394 ;
      RECT 28.294 24.358 28.346 24.394 ;
      RECT 27.894 24.358 27.946 24.394 ;
      RECT 27.494 24.358 27.546 24.394 ;
      RECT 27.094 24.358 27.146 24.394 ;
      RECT 26.694 24.358 26.746 24.394 ;
      RECT 26.294 24.358 26.346 24.394 ;
      RECT 25.894 24.358 25.946 24.394 ;
      RECT 25.494 24.358 25.546 24.394 ;
      RECT 25.094 24.358 25.146 24.394 ;
      RECT 24.694 24.358 24.746 24.394 ;
      RECT 24.294 24.358 24.346 24.394 ;
      RECT 23.894 24.358 23.946 24.394 ;
      RECT 23.494 24.358 23.546 24.394 ;
      RECT 23.094 24.358 23.146 24.394 ;
      RECT 21.814 24.358 21.868 24.394 ;
      RECT 19.838 24.358 19.886 24.394 ;
      RECT 19.53 24.358 19.578 24.394 ;
      RECT 16.882 24.358 16.936 24.394 ;
      RECT 16.422 24.358 16.47 24.394 ;
      RECT 16.114 24.358 16.162 24.394 ;
      RECT 14.132 24.358 14.186 24.394 ;
      RECT 13.294 24.358 13.346 24.394 ;
      RECT 12.894 24.358 12.946 24.394 ;
      RECT 12.494 24.358 12.546 24.394 ;
      RECT 12.094 24.358 12.146 24.394 ;
      RECT 11.694 24.358 11.746 24.394 ;
      RECT 11.294 24.358 11.346 24.394 ;
      RECT 10.894 24.358 10.946 24.394 ;
      RECT 10.494 24.358 10.546 24.394 ;
      RECT 10.094 24.358 10.146 24.394 ;
      RECT 9.694 24.358 9.746 24.394 ;
      RECT 9.294 24.358 9.346 24.394 ;
      RECT 8.894 24.358 8.946 24.394 ;
      RECT 8.494 24.358 8.546 24.394 ;
      RECT 8.094 24.358 8.146 24.394 ;
      RECT 7.694 24.358 7.746 24.394 ;
      RECT 7.294 24.358 7.346 24.394 ;
      RECT 6.894 24.358 6.946 24.394 ;
      RECT 6.494 24.358 6.546 24.394 ;
      RECT 6.094 24.358 6.146 24.394 ;
      RECT 5.694 24.358 5.746 24.394 ;
      RECT 5.294 24.358 5.346 24.394 ;
      RECT 4.894 24.358 4.946 24.394 ;
      RECT 4.494 24.358 4.546 24.394 ;
      RECT 4.094 24.358 4.146 24.394 ;
      RECT 3.694 24.358 3.746 24.394 ;
      RECT 3.294 24.358 3.346 24.394 ;
      RECT 2.894 24.358 2.946 24.394 ;
      RECT 2.494 24.358 2.546 24.394 ;
      RECT 2.094 24.358 2.146 24.394 ;
      RECT 1.694 24.358 1.746 24.394 ;
      RECT 1.294 24.358 1.346 24.394 ;
      RECT 0.894 24.358 0.946 24.394 ;
      RECT 21.414 24.282 21.468 24.318 ;
      RECT 14.532 24.282 14.586 24.318 ;
      RECT 19.606 24.129 19.654 24.165 ;
      RECT 18.08 24.129 18.12 24.165 ;
      RECT 16.718 24.129 16.772 24.165 ;
      RECT 16.346 24.129 16.394 24.165 ;
      RECT 20.37 24.1345 20.442 24.1595 ;
      RECT 18.764 24.1345 18.836 24.1595 ;
      RECT 15.558 24.1345 15.63 24.1595 ;
      RECT 21.978 23.982 22.022 24.018 ;
      RECT 13.978 23.982 14.022 24.018 ;
      RECT 18.764 23.9875 18.836 24.0125 ;
      RECT 19.762 23.835 19.81 23.871 ;
      RECT 17.616 23.835 17.656 23.871 ;
      RECT 16.19 23.835 16.238 23.871 ;
      RECT 35.254 23.606 35.306 23.642 ;
      RECT 34.854 23.606 34.906 23.642 ;
      RECT 34.454 23.606 34.506 23.642 ;
      RECT 34.054 23.606 34.106 23.642 ;
      RECT 33.654 23.606 33.706 23.642 ;
      RECT 33.254 23.606 33.306 23.642 ;
      RECT 32.854 23.606 32.906 23.642 ;
      RECT 32.454 23.606 32.506 23.642 ;
      RECT 32.054 23.606 32.106 23.642 ;
      RECT 31.654 23.606 31.706 23.642 ;
      RECT 31.254 23.606 31.306 23.642 ;
      RECT 30.854 23.606 30.906 23.642 ;
      RECT 30.454 23.606 30.506 23.642 ;
      RECT 30.054 23.606 30.106 23.642 ;
      RECT 29.654 23.606 29.706 23.642 ;
      RECT 29.254 23.606 29.306 23.642 ;
      RECT 28.854 23.606 28.906 23.642 ;
      RECT 28.454 23.606 28.506 23.642 ;
      RECT 28.054 23.606 28.106 23.642 ;
      RECT 27.654 23.606 27.706 23.642 ;
      RECT 27.254 23.606 27.306 23.642 ;
      RECT 26.854 23.606 26.906 23.642 ;
      RECT 26.454 23.606 26.506 23.642 ;
      RECT 26.054 23.606 26.106 23.642 ;
      RECT 25.654 23.606 25.706 23.642 ;
      RECT 25.254 23.606 25.306 23.642 ;
      RECT 24.854 23.606 24.906 23.642 ;
      RECT 24.454 23.606 24.506 23.642 ;
      RECT 24.054 23.606 24.106 23.642 ;
      RECT 23.654 23.606 23.706 23.642 ;
      RECT 23.254 23.606 23.306 23.642 ;
      RECT 22.854 23.606 22.906 23.642 ;
      RECT 22.694 23.606 22.746 23.642 ;
      RECT 21.732 23.606 21.786 23.642 ;
      RECT 14.214 23.606 14.268 23.642 ;
      RECT 13.054 23.606 13.106 23.642 ;
      RECT 12.654 23.606 12.706 23.642 ;
      RECT 12.254 23.606 12.306 23.642 ;
      RECT 11.854 23.606 11.906 23.642 ;
      RECT 11.454 23.606 11.506 23.642 ;
      RECT 11.054 23.606 11.106 23.642 ;
      RECT 10.654 23.606 10.706 23.642 ;
      RECT 10.254 23.606 10.306 23.642 ;
      RECT 9.854 23.606 9.906 23.642 ;
      RECT 9.454 23.606 9.506 23.642 ;
      RECT 9.054 23.606 9.106 23.642 ;
      RECT 8.654 23.606 8.706 23.642 ;
      RECT 8.254 23.606 8.306 23.642 ;
      RECT 7.854 23.606 7.906 23.642 ;
      RECT 7.454 23.606 7.506 23.642 ;
      RECT 7.054 23.606 7.106 23.642 ;
      RECT 6.654 23.606 6.706 23.642 ;
      RECT 6.254 23.606 6.306 23.642 ;
      RECT 5.854 23.606 5.906 23.642 ;
      RECT 5.454 23.606 5.506 23.642 ;
      RECT 5.054 23.606 5.106 23.642 ;
      RECT 4.654 23.606 4.706 23.642 ;
      RECT 4.254 23.606 4.306 23.642 ;
      RECT 3.854 23.606 3.906 23.642 ;
      RECT 3.454 23.606 3.506 23.642 ;
      RECT 3.054 23.606 3.106 23.642 ;
      RECT 2.654 23.606 2.706 23.642 ;
      RECT 2.254 23.606 2.306 23.642 ;
      RECT 1.854 23.606 1.906 23.642 ;
      RECT 1.454 23.606 1.506 23.642 ;
      RECT 1.054 23.606 1.106 23.642 ;
      RECT 0.654 23.606 0.706 23.642 ;
      RECT 21.978 23.382 22.022 23.418 ;
      RECT 21.096 23.382 21.14 23.418 ;
      RECT 14.86 23.382 14.904 23.418 ;
      RECT 13.978 23.382 14.022 23.418 ;
      RECT 35.494 23.158 35.546 23.194 ;
      RECT 35.094 23.158 35.146 23.194 ;
      RECT 34.694 23.158 34.746 23.194 ;
      RECT 34.294 23.158 34.346 23.194 ;
      RECT 33.894 23.158 33.946 23.194 ;
      RECT 33.494 23.158 33.546 23.194 ;
      RECT 33.094 23.158 33.146 23.194 ;
      RECT 32.694 23.158 32.746 23.194 ;
      RECT 32.294 23.158 32.346 23.194 ;
      RECT 31.894 23.158 31.946 23.194 ;
      RECT 31.494 23.158 31.546 23.194 ;
      RECT 31.094 23.158 31.146 23.194 ;
      RECT 30.694 23.158 30.746 23.194 ;
      RECT 30.294 23.158 30.346 23.194 ;
      RECT 29.894 23.158 29.946 23.194 ;
      RECT 29.494 23.158 29.546 23.194 ;
      RECT 29.094 23.158 29.146 23.194 ;
      RECT 28.694 23.158 28.746 23.194 ;
      RECT 28.294 23.158 28.346 23.194 ;
      RECT 27.894 23.158 27.946 23.194 ;
      RECT 27.494 23.158 27.546 23.194 ;
      RECT 27.094 23.158 27.146 23.194 ;
      RECT 26.694 23.158 26.746 23.194 ;
      RECT 26.294 23.158 26.346 23.194 ;
      RECT 25.894 23.158 25.946 23.194 ;
      RECT 25.494 23.158 25.546 23.194 ;
      RECT 25.094 23.158 25.146 23.194 ;
      RECT 24.694 23.158 24.746 23.194 ;
      RECT 24.294 23.158 24.346 23.194 ;
      RECT 23.894 23.158 23.946 23.194 ;
      RECT 23.494 23.158 23.546 23.194 ;
      RECT 23.094 23.158 23.146 23.194 ;
      RECT 21.814 23.158 21.868 23.194 ;
      RECT 19.838 23.158 19.886 23.194 ;
      RECT 19.53 23.158 19.578 23.194 ;
      RECT 16.882 23.158 16.936 23.194 ;
      RECT 16.422 23.158 16.47 23.194 ;
      RECT 16.114 23.158 16.162 23.194 ;
      RECT 14.132 23.158 14.186 23.194 ;
      RECT 13.294 23.158 13.346 23.194 ;
      RECT 12.894 23.158 12.946 23.194 ;
      RECT 12.494 23.158 12.546 23.194 ;
      RECT 12.094 23.158 12.146 23.194 ;
      RECT 11.694 23.158 11.746 23.194 ;
      RECT 11.294 23.158 11.346 23.194 ;
      RECT 10.894 23.158 10.946 23.194 ;
      RECT 10.494 23.158 10.546 23.194 ;
      RECT 10.094 23.158 10.146 23.194 ;
      RECT 9.694 23.158 9.746 23.194 ;
      RECT 9.294 23.158 9.346 23.194 ;
      RECT 8.894 23.158 8.946 23.194 ;
      RECT 8.494 23.158 8.546 23.194 ;
      RECT 8.094 23.158 8.146 23.194 ;
      RECT 7.694 23.158 7.746 23.194 ;
      RECT 7.294 23.158 7.346 23.194 ;
      RECT 6.894 23.158 6.946 23.194 ;
      RECT 6.494 23.158 6.546 23.194 ;
      RECT 6.094 23.158 6.146 23.194 ;
      RECT 5.694 23.158 5.746 23.194 ;
      RECT 5.294 23.158 5.346 23.194 ;
      RECT 4.894 23.158 4.946 23.194 ;
      RECT 4.494 23.158 4.546 23.194 ;
      RECT 4.094 23.158 4.146 23.194 ;
      RECT 3.694 23.158 3.746 23.194 ;
      RECT 3.294 23.158 3.346 23.194 ;
      RECT 2.894 23.158 2.946 23.194 ;
      RECT 2.494 23.158 2.546 23.194 ;
      RECT 2.094 23.158 2.146 23.194 ;
      RECT 1.694 23.158 1.746 23.194 ;
      RECT 1.294 23.158 1.346 23.194 ;
      RECT 0.894 23.158 0.946 23.194 ;
      RECT 21.414 23.082 21.468 23.118 ;
      RECT 14.532 23.082 14.586 23.118 ;
      RECT 19.606 22.929 19.654 22.965 ;
      RECT 18.08 22.929 18.12 22.965 ;
      RECT 16.718 22.929 16.772 22.965 ;
      RECT 16.346 22.929 16.394 22.965 ;
      RECT 20.37 22.9345 20.442 22.9595 ;
      RECT 18.764 22.9345 18.836 22.9595 ;
      RECT 15.558 22.9345 15.63 22.9595 ;
      RECT 21.978 22.782 22.022 22.818 ;
      RECT 13.978 22.782 14.022 22.818 ;
      RECT 18.764 22.7875 18.836 22.8125 ;
      RECT 19.762 22.635 19.81 22.671 ;
      RECT 17.616 22.635 17.656 22.671 ;
      RECT 16.19 22.635 16.238 22.671 ;
      RECT 35.254 22.406 35.306 22.442 ;
      RECT 34.854 22.406 34.906 22.442 ;
      RECT 34.454 22.406 34.506 22.442 ;
      RECT 34.054 22.406 34.106 22.442 ;
      RECT 33.654 22.406 33.706 22.442 ;
      RECT 33.254 22.406 33.306 22.442 ;
      RECT 32.854 22.406 32.906 22.442 ;
      RECT 32.454 22.406 32.506 22.442 ;
      RECT 32.054 22.406 32.106 22.442 ;
      RECT 31.654 22.406 31.706 22.442 ;
      RECT 31.254 22.406 31.306 22.442 ;
      RECT 30.854 22.406 30.906 22.442 ;
      RECT 30.454 22.406 30.506 22.442 ;
      RECT 30.054 22.406 30.106 22.442 ;
      RECT 29.654 22.406 29.706 22.442 ;
      RECT 29.254 22.406 29.306 22.442 ;
      RECT 28.854 22.406 28.906 22.442 ;
      RECT 28.454 22.406 28.506 22.442 ;
      RECT 28.054 22.406 28.106 22.442 ;
      RECT 27.654 22.406 27.706 22.442 ;
      RECT 27.254 22.406 27.306 22.442 ;
      RECT 26.854 22.406 26.906 22.442 ;
      RECT 26.454 22.406 26.506 22.442 ;
      RECT 26.054 22.406 26.106 22.442 ;
      RECT 25.654 22.406 25.706 22.442 ;
      RECT 25.254 22.406 25.306 22.442 ;
      RECT 24.854 22.406 24.906 22.442 ;
      RECT 24.454 22.406 24.506 22.442 ;
      RECT 24.054 22.406 24.106 22.442 ;
      RECT 23.654 22.406 23.706 22.442 ;
      RECT 23.254 22.406 23.306 22.442 ;
      RECT 22.854 22.406 22.906 22.442 ;
      RECT 22.694 22.406 22.746 22.442 ;
      RECT 21.732 22.406 21.786 22.442 ;
      RECT 14.214 22.406 14.268 22.442 ;
      RECT 13.054 22.406 13.106 22.442 ;
      RECT 12.654 22.406 12.706 22.442 ;
      RECT 12.254 22.406 12.306 22.442 ;
      RECT 11.854 22.406 11.906 22.442 ;
      RECT 11.454 22.406 11.506 22.442 ;
      RECT 11.054 22.406 11.106 22.442 ;
      RECT 10.654 22.406 10.706 22.442 ;
      RECT 10.254 22.406 10.306 22.442 ;
      RECT 9.854 22.406 9.906 22.442 ;
      RECT 9.454 22.406 9.506 22.442 ;
      RECT 9.054 22.406 9.106 22.442 ;
      RECT 8.654 22.406 8.706 22.442 ;
      RECT 8.254 22.406 8.306 22.442 ;
      RECT 7.854 22.406 7.906 22.442 ;
      RECT 7.454 22.406 7.506 22.442 ;
      RECT 7.054 22.406 7.106 22.442 ;
      RECT 6.654 22.406 6.706 22.442 ;
      RECT 6.254 22.406 6.306 22.442 ;
      RECT 5.854 22.406 5.906 22.442 ;
      RECT 5.454 22.406 5.506 22.442 ;
      RECT 5.054 22.406 5.106 22.442 ;
      RECT 4.654 22.406 4.706 22.442 ;
      RECT 4.254 22.406 4.306 22.442 ;
      RECT 3.854 22.406 3.906 22.442 ;
      RECT 3.454 22.406 3.506 22.442 ;
      RECT 3.054 22.406 3.106 22.442 ;
      RECT 2.654 22.406 2.706 22.442 ;
      RECT 2.254 22.406 2.306 22.442 ;
      RECT 1.854 22.406 1.906 22.442 ;
      RECT 1.454 22.406 1.506 22.442 ;
      RECT 1.054 22.406 1.106 22.442 ;
      RECT 0.654 22.406 0.706 22.442 ;
      RECT 21.978 22.182 22.022 22.218 ;
      RECT 21.096 22.182 21.14 22.218 ;
      RECT 14.86 22.182 14.904 22.218 ;
      RECT 13.978 22.182 14.022 22.218 ;
      RECT 35.494 21.958 35.546 21.994 ;
      RECT 35.094 21.958 35.146 21.994 ;
      RECT 34.694 21.958 34.746 21.994 ;
      RECT 34.294 21.958 34.346 21.994 ;
      RECT 33.894 21.958 33.946 21.994 ;
      RECT 33.494 21.958 33.546 21.994 ;
      RECT 33.094 21.958 33.146 21.994 ;
      RECT 32.694 21.958 32.746 21.994 ;
      RECT 32.294 21.958 32.346 21.994 ;
      RECT 31.894 21.958 31.946 21.994 ;
      RECT 31.494 21.958 31.546 21.994 ;
      RECT 31.094 21.958 31.146 21.994 ;
      RECT 30.694 21.958 30.746 21.994 ;
      RECT 30.294 21.958 30.346 21.994 ;
      RECT 29.894 21.958 29.946 21.994 ;
      RECT 29.494 21.958 29.546 21.994 ;
      RECT 29.094 21.958 29.146 21.994 ;
      RECT 28.694 21.958 28.746 21.994 ;
      RECT 28.294 21.958 28.346 21.994 ;
      RECT 27.894 21.958 27.946 21.994 ;
      RECT 27.494 21.958 27.546 21.994 ;
      RECT 27.094 21.958 27.146 21.994 ;
      RECT 26.694 21.958 26.746 21.994 ;
      RECT 26.294 21.958 26.346 21.994 ;
      RECT 25.894 21.958 25.946 21.994 ;
      RECT 25.494 21.958 25.546 21.994 ;
      RECT 25.094 21.958 25.146 21.994 ;
      RECT 24.694 21.958 24.746 21.994 ;
      RECT 24.294 21.958 24.346 21.994 ;
      RECT 23.894 21.958 23.946 21.994 ;
      RECT 23.494 21.958 23.546 21.994 ;
      RECT 23.094 21.958 23.146 21.994 ;
      RECT 21.814 21.958 21.868 21.994 ;
      RECT 19.838 21.958 19.886 21.994 ;
      RECT 19.53 21.958 19.578 21.994 ;
      RECT 16.882 21.958 16.936 21.994 ;
      RECT 16.422 21.958 16.47 21.994 ;
      RECT 16.114 21.958 16.162 21.994 ;
      RECT 14.132 21.958 14.186 21.994 ;
      RECT 13.294 21.958 13.346 21.994 ;
      RECT 12.894 21.958 12.946 21.994 ;
      RECT 12.494 21.958 12.546 21.994 ;
      RECT 12.094 21.958 12.146 21.994 ;
      RECT 11.694 21.958 11.746 21.994 ;
      RECT 11.294 21.958 11.346 21.994 ;
      RECT 10.894 21.958 10.946 21.994 ;
      RECT 10.494 21.958 10.546 21.994 ;
      RECT 10.094 21.958 10.146 21.994 ;
      RECT 9.694 21.958 9.746 21.994 ;
      RECT 9.294 21.958 9.346 21.994 ;
      RECT 8.894 21.958 8.946 21.994 ;
      RECT 8.494 21.958 8.546 21.994 ;
      RECT 8.094 21.958 8.146 21.994 ;
      RECT 7.694 21.958 7.746 21.994 ;
      RECT 7.294 21.958 7.346 21.994 ;
      RECT 6.894 21.958 6.946 21.994 ;
      RECT 6.494 21.958 6.546 21.994 ;
      RECT 6.094 21.958 6.146 21.994 ;
      RECT 5.694 21.958 5.746 21.994 ;
      RECT 5.294 21.958 5.346 21.994 ;
      RECT 4.894 21.958 4.946 21.994 ;
      RECT 4.494 21.958 4.546 21.994 ;
      RECT 4.094 21.958 4.146 21.994 ;
      RECT 3.694 21.958 3.746 21.994 ;
      RECT 3.294 21.958 3.346 21.994 ;
      RECT 2.894 21.958 2.946 21.994 ;
      RECT 2.494 21.958 2.546 21.994 ;
      RECT 2.094 21.958 2.146 21.994 ;
      RECT 1.694 21.958 1.746 21.994 ;
      RECT 1.294 21.958 1.346 21.994 ;
      RECT 0.894 21.958 0.946 21.994 ;
      RECT 21.414 21.882 21.468 21.918 ;
      RECT 14.532 21.882 14.586 21.918 ;
      RECT 19.606 21.729 19.654 21.765 ;
      RECT 18.08 21.729 18.12 21.765 ;
      RECT 16.718 21.729 16.772 21.765 ;
      RECT 16.346 21.729 16.394 21.765 ;
      RECT 20.37 21.7345 20.442 21.7595 ;
      RECT 18.764 21.7345 18.836 21.7595 ;
      RECT 15.558 21.7345 15.63 21.7595 ;
      RECT 21.978 21.582 22.022 21.618 ;
      RECT 13.978 21.582 14.022 21.618 ;
      RECT 18.764 21.5875 18.836 21.6125 ;
      RECT 19.762 21.435 19.81 21.471 ;
      RECT 17.616 21.435 17.656 21.471 ;
      RECT 16.19 21.435 16.238 21.471 ;
      RECT 35.254 21.206 35.306 21.242 ;
      RECT 34.854 21.206 34.906 21.242 ;
      RECT 34.454 21.206 34.506 21.242 ;
      RECT 34.054 21.206 34.106 21.242 ;
      RECT 33.654 21.206 33.706 21.242 ;
      RECT 33.254 21.206 33.306 21.242 ;
      RECT 32.854 21.206 32.906 21.242 ;
      RECT 32.454 21.206 32.506 21.242 ;
      RECT 32.054 21.206 32.106 21.242 ;
      RECT 31.654 21.206 31.706 21.242 ;
      RECT 31.254 21.206 31.306 21.242 ;
      RECT 30.854 21.206 30.906 21.242 ;
      RECT 30.454 21.206 30.506 21.242 ;
      RECT 30.054 21.206 30.106 21.242 ;
      RECT 29.654 21.206 29.706 21.242 ;
      RECT 29.254 21.206 29.306 21.242 ;
      RECT 28.854 21.206 28.906 21.242 ;
      RECT 28.454 21.206 28.506 21.242 ;
      RECT 28.054 21.206 28.106 21.242 ;
      RECT 27.654 21.206 27.706 21.242 ;
      RECT 27.254 21.206 27.306 21.242 ;
      RECT 26.854 21.206 26.906 21.242 ;
      RECT 26.454 21.206 26.506 21.242 ;
      RECT 26.054 21.206 26.106 21.242 ;
      RECT 25.654 21.206 25.706 21.242 ;
      RECT 25.254 21.206 25.306 21.242 ;
      RECT 24.854 21.206 24.906 21.242 ;
      RECT 24.454 21.206 24.506 21.242 ;
      RECT 24.054 21.206 24.106 21.242 ;
      RECT 23.654 21.206 23.706 21.242 ;
      RECT 23.254 21.206 23.306 21.242 ;
      RECT 22.854 21.206 22.906 21.242 ;
      RECT 22.694 21.206 22.746 21.242 ;
      RECT 21.732 21.206 21.786 21.242 ;
      RECT 14.214 21.206 14.268 21.242 ;
      RECT 13.054 21.206 13.106 21.242 ;
      RECT 12.654 21.206 12.706 21.242 ;
      RECT 12.254 21.206 12.306 21.242 ;
      RECT 11.854 21.206 11.906 21.242 ;
      RECT 11.454 21.206 11.506 21.242 ;
      RECT 11.054 21.206 11.106 21.242 ;
      RECT 10.654 21.206 10.706 21.242 ;
      RECT 10.254 21.206 10.306 21.242 ;
      RECT 9.854 21.206 9.906 21.242 ;
      RECT 9.454 21.206 9.506 21.242 ;
      RECT 9.054 21.206 9.106 21.242 ;
      RECT 8.654 21.206 8.706 21.242 ;
      RECT 8.254 21.206 8.306 21.242 ;
      RECT 7.854 21.206 7.906 21.242 ;
      RECT 7.454 21.206 7.506 21.242 ;
      RECT 7.054 21.206 7.106 21.242 ;
      RECT 6.654 21.206 6.706 21.242 ;
      RECT 6.254 21.206 6.306 21.242 ;
      RECT 5.854 21.206 5.906 21.242 ;
      RECT 5.454 21.206 5.506 21.242 ;
      RECT 5.054 21.206 5.106 21.242 ;
      RECT 4.654 21.206 4.706 21.242 ;
      RECT 4.254 21.206 4.306 21.242 ;
      RECT 3.854 21.206 3.906 21.242 ;
      RECT 3.454 21.206 3.506 21.242 ;
      RECT 3.054 21.206 3.106 21.242 ;
      RECT 2.654 21.206 2.706 21.242 ;
      RECT 2.254 21.206 2.306 21.242 ;
      RECT 1.854 21.206 1.906 21.242 ;
      RECT 1.454 21.206 1.506 21.242 ;
      RECT 1.054 21.206 1.106 21.242 ;
      RECT 0.654 21.206 0.706 21.242 ;
      RECT 21.978 20.982 22.022 21.018 ;
      RECT 21.096 20.982 21.14 21.018 ;
      RECT 14.86 20.982 14.904 21.018 ;
      RECT 13.978 20.982 14.022 21.018 ;
      RECT 35.494 20.758 35.546 20.794 ;
      RECT 35.094 20.758 35.146 20.794 ;
      RECT 34.694 20.758 34.746 20.794 ;
      RECT 34.294 20.758 34.346 20.794 ;
      RECT 33.894 20.758 33.946 20.794 ;
      RECT 33.494 20.758 33.546 20.794 ;
      RECT 33.094 20.758 33.146 20.794 ;
      RECT 32.694 20.758 32.746 20.794 ;
      RECT 32.294 20.758 32.346 20.794 ;
      RECT 31.894 20.758 31.946 20.794 ;
      RECT 31.494 20.758 31.546 20.794 ;
      RECT 31.094 20.758 31.146 20.794 ;
      RECT 30.694 20.758 30.746 20.794 ;
      RECT 30.294 20.758 30.346 20.794 ;
      RECT 29.894 20.758 29.946 20.794 ;
      RECT 29.494 20.758 29.546 20.794 ;
      RECT 29.094 20.758 29.146 20.794 ;
      RECT 28.694 20.758 28.746 20.794 ;
      RECT 28.294 20.758 28.346 20.794 ;
      RECT 27.894 20.758 27.946 20.794 ;
      RECT 27.494 20.758 27.546 20.794 ;
      RECT 27.094 20.758 27.146 20.794 ;
      RECT 26.694 20.758 26.746 20.794 ;
      RECT 26.294 20.758 26.346 20.794 ;
      RECT 25.894 20.758 25.946 20.794 ;
      RECT 25.494 20.758 25.546 20.794 ;
      RECT 25.094 20.758 25.146 20.794 ;
      RECT 24.694 20.758 24.746 20.794 ;
      RECT 24.294 20.758 24.346 20.794 ;
      RECT 23.894 20.758 23.946 20.794 ;
      RECT 23.494 20.758 23.546 20.794 ;
      RECT 23.094 20.758 23.146 20.794 ;
      RECT 21.814 20.758 21.868 20.794 ;
      RECT 19.838 20.758 19.886 20.794 ;
      RECT 19.53 20.758 19.578 20.794 ;
      RECT 16.882 20.758 16.936 20.794 ;
      RECT 16.422 20.758 16.47 20.794 ;
      RECT 16.114 20.758 16.162 20.794 ;
      RECT 14.132 20.758 14.186 20.794 ;
      RECT 13.294 20.758 13.346 20.794 ;
      RECT 12.894 20.758 12.946 20.794 ;
      RECT 12.494 20.758 12.546 20.794 ;
      RECT 12.094 20.758 12.146 20.794 ;
      RECT 11.694 20.758 11.746 20.794 ;
      RECT 11.294 20.758 11.346 20.794 ;
      RECT 10.894 20.758 10.946 20.794 ;
      RECT 10.494 20.758 10.546 20.794 ;
      RECT 10.094 20.758 10.146 20.794 ;
      RECT 9.694 20.758 9.746 20.794 ;
      RECT 9.294 20.758 9.346 20.794 ;
      RECT 8.894 20.758 8.946 20.794 ;
      RECT 8.494 20.758 8.546 20.794 ;
      RECT 8.094 20.758 8.146 20.794 ;
      RECT 7.694 20.758 7.746 20.794 ;
      RECT 7.294 20.758 7.346 20.794 ;
      RECT 6.894 20.758 6.946 20.794 ;
      RECT 6.494 20.758 6.546 20.794 ;
      RECT 6.094 20.758 6.146 20.794 ;
      RECT 5.694 20.758 5.746 20.794 ;
      RECT 5.294 20.758 5.346 20.794 ;
      RECT 4.894 20.758 4.946 20.794 ;
      RECT 4.494 20.758 4.546 20.794 ;
      RECT 4.094 20.758 4.146 20.794 ;
      RECT 3.694 20.758 3.746 20.794 ;
      RECT 3.294 20.758 3.346 20.794 ;
      RECT 2.894 20.758 2.946 20.794 ;
      RECT 2.494 20.758 2.546 20.794 ;
      RECT 2.094 20.758 2.146 20.794 ;
      RECT 1.694 20.758 1.746 20.794 ;
      RECT 1.294 20.758 1.346 20.794 ;
      RECT 0.894 20.758 0.946 20.794 ;
      RECT 21.414 20.682 21.468 20.718 ;
      RECT 14.532 20.682 14.586 20.718 ;
      RECT 19.606 20.529 19.654 20.565 ;
      RECT 18.08 20.529 18.12 20.565 ;
      RECT 16.718 20.529 16.772 20.565 ;
      RECT 16.346 20.529 16.394 20.565 ;
      RECT 20.37 20.5345 20.442 20.5595 ;
      RECT 18.764 20.5345 18.836 20.5595 ;
      RECT 15.558 20.5345 15.63 20.5595 ;
      RECT 21.978 20.382 22.022 20.418 ;
      RECT 13.978 20.382 14.022 20.418 ;
      RECT 18.764 20.3875 18.836 20.4125 ;
      RECT 19.762 20.235 19.81 20.271 ;
      RECT 17.616 20.235 17.656 20.271 ;
      RECT 16.19 20.235 16.238 20.271 ;
      RECT 35.254 20.006 35.306 20.042 ;
      RECT 34.854 20.006 34.906 20.042 ;
      RECT 34.454 20.006 34.506 20.042 ;
      RECT 34.054 20.006 34.106 20.042 ;
      RECT 33.654 20.006 33.706 20.042 ;
      RECT 33.254 20.006 33.306 20.042 ;
      RECT 32.854 20.006 32.906 20.042 ;
      RECT 32.454 20.006 32.506 20.042 ;
      RECT 32.054 20.006 32.106 20.042 ;
      RECT 31.654 20.006 31.706 20.042 ;
      RECT 31.254 20.006 31.306 20.042 ;
      RECT 30.854 20.006 30.906 20.042 ;
      RECT 30.454 20.006 30.506 20.042 ;
      RECT 30.054 20.006 30.106 20.042 ;
      RECT 29.654 20.006 29.706 20.042 ;
      RECT 29.254 20.006 29.306 20.042 ;
      RECT 28.854 20.006 28.906 20.042 ;
      RECT 28.454 20.006 28.506 20.042 ;
      RECT 28.054 20.006 28.106 20.042 ;
      RECT 27.654 20.006 27.706 20.042 ;
      RECT 27.254 20.006 27.306 20.042 ;
      RECT 26.854 20.006 26.906 20.042 ;
      RECT 26.454 20.006 26.506 20.042 ;
      RECT 26.054 20.006 26.106 20.042 ;
      RECT 25.654 20.006 25.706 20.042 ;
      RECT 25.254 20.006 25.306 20.042 ;
      RECT 24.854 20.006 24.906 20.042 ;
      RECT 24.454 20.006 24.506 20.042 ;
      RECT 24.054 20.006 24.106 20.042 ;
      RECT 23.654 20.006 23.706 20.042 ;
      RECT 23.254 20.006 23.306 20.042 ;
      RECT 22.854 20.006 22.906 20.042 ;
      RECT 22.694 20.006 22.746 20.042 ;
      RECT 21.732 20.006 21.786 20.042 ;
      RECT 14.214 20.006 14.268 20.042 ;
      RECT 13.054 20.006 13.106 20.042 ;
      RECT 12.654 20.006 12.706 20.042 ;
      RECT 12.254 20.006 12.306 20.042 ;
      RECT 11.854 20.006 11.906 20.042 ;
      RECT 11.454 20.006 11.506 20.042 ;
      RECT 11.054 20.006 11.106 20.042 ;
      RECT 10.654 20.006 10.706 20.042 ;
      RECT 10.254 20.006 10.306 20.042 ;
      RECT 9.854 20.006 9.906 20.042 ;
      RECT 9.454 20.006 9.506 20.042 ;
      RECT 9.054 20.006 9.106 20.042 ;
      RECT 8.654 20.006 8.706 20.042 ;
      RECT 8.254 20.006 8.306 20.042 ;
      RECT 7.854 20.006 7.906 20.042 ;
      RECT 7.454 20.006 7.506 20.042 ;
      RECT 7.054 20.006 7.106 20.042 ;
      RECT 6.654 20.006 6.706 20.042 ;
      RECT 6.254 20.006 6.306 20.042 ;
      RECT 5.854 20.006 5.906 20.042 ;
      RECT 5.454 20.006 5.506 20.042 ;
      RECT 5.054 20.006 5.106 20.042 ;
      RECT 4.654 20.006 4.706 20.042 ;
      RECT 4.254 20.006 4.306 20.042 ;
      RECT 3.854 20.006 3.906 20.042 ;
      RECT 3.454 20.006 3.506 20.042 ;
      RECT 3.054 20.006 3.106 20.042 ;
      RECT 2.654 20.006 2.706 20.042 ;
      RECT 2.254 20.006 2.306 20.042 ;
      RECT 1.854 20.006 1.906 20.042 ;
      RECT 1.454 20.006 1.506 20.042 ;
      RECT 1.054 20.006 1.106 20.042 ;
      RECT 0.654 20.006 0.706 20.042 ;
      RECT 21.978 19.782 22.022 19.818 ;
      RECT 21.096 19.782 21.14 19.818 ;
      RECT 14.86 19.782 14.904 19.818 ;
      RECT 13.978 19.782 14.022 19.818 ;
      RECT 35.494 19.558 35.546 19.594 ;
      RECT 35.094 19.558 35.146 19.594 ;
      RECT 34.694 19.558 34.746 19.594 ;
      RECT 34.294 19.558 34.346 19.594 ;
      RECT 33.894 19.558 33.946 19.594 ;
      RECT 33.494 19.558 33.546 19.594 ;
      RECT 33.094 19.558 33.146 19.594 ;
      RECT 32.694 19.558 32.746 19.594 ;
      RECT 32.294 19.558 32.346 19.594 ;
      RECT 31.894 19.558 31.946 19.594 ;
      RECT 31.494 19.558 31.546 19.594 ;
      RECT 31.094 19.558 31.146 19.594 ;
      RECT 30.694 19.558 30.746 19.594 ;
      RECT 30.294 19.558 30.346 19.594 ;
      RECT 29.894 19.558 29.946 19.594 ;
      RECT 29.494 19.558 29.546 19.594 ;
      RECT 29.094 19.558 29.146 19.594 ;
      RECT 28.694 19.558 28.746 19.594 ;
      RECT 28.294 19.558 28.346 19.594 ;
      RECT 27.894 19.558 27.946 19.594 ;
      RECT 27.494 19.558 27.546 19.594 ;
      RECT 27.094 19.558 27.146 19.594 ;
      RECT 26.694 19.558 26.746 19.594 ;
      RECT 26.294 19.558 26.346 19.594 ;
      RECT 25.894 19.558 25.946 19.594 ;
      RECT 25.494 19.558 25.546 19.594 ;
      RECT 25.094 19.558 25.146 19.594 ;
      RECT 24.694 19.558 24.746 19.594 ;
      RECT 24.294 19.558 24.346 19.594 ;
      RECT 23.894 19.558 23.946 19.594 ;
      RECT 23.494 19.558 23.546 19.594 ;
      RECT 23.094 19.558 23.146 19.594 ;
      RECT 21.814 19.558 21.868 19.594 ;
      RECT 19.838 19.558 19.886 19.594 ;
      RECT 19.53 19.558 19.578 19.594 ;
      RECT 16.882 19.558 16.936 19.594 ;
      RECT 16.422 19.558 16.47 19.594 ;
      RECT 16.114 19.558 16.162 19.594 ;
      RECT 14.132 19.558 14.186 19.594 ;
      RECT 13.294 19.558 13.346 19.594 ;
      RECT 12.894 19.558 12.946 19.594 ;
      RECT 12.494 19.558 12.546 19.594 ;
      RECT 12.094 19.558 12.146 19.594 ;
      RECT 11.694 19.558 11.746 19.594 ;
      RECT 11.294 19.558 11.346 19.594 ;
      RECT 10.894 19.558 10.946 19.594 ;
      RECT 10.494 19.558 10.546 19.594 ;
      RECT 10.094 19.558 10.146 19.594 ;
      RECT 9.694 19.558 9.746 19.594 ;
      RECT 9.294 19.558 9.346 19.594 ;
      RECT 8.894 19.558 8.946 19.594 ;
      RECT 8.494 19.558 8.546 19.594 ;
      RECT 8.094 19.558 8.146 19.594 ;
      RECT 7.694 19.558 7.746 19.594 ;
      RECT 7.294 19.558 7.346 19.594 ;
      RECT 6.894 19.558 6.946 19.594 ;
      RECT 6.494 19.558 6.546 19.594 ;
      RECT 6.094 19.558 6.146 19.594 ;
      RECT 5.694 19.558 5.746 19.594 ;
      RECT 5.294 19.558 5.346 19.594 ;
      RECT 4.894 19.558 4.946 19.594 ;
      RECT 4.494 19.558 4.546 19.594 ;
      RECT 4.094 19.558 4.146 19.594 ;
      RECT 3.694 19.558 3.746 19.594 ;
      RECT 3.294 19.558 3.346 19.594 ;
      RECT 2.894 19.558 2.946 19.594 ;
      RECT 2.494 19.558 2.546 19.594 ;
      RECT 2.094 19.558 2.146 19.594 ;
      RECT 1.694 19.558 1.746 19.594 ;
      RECT 1.294 19.558 1.346 19.594 ;
      RECT 0.894 19.558 0.946 19.594 ;
      RECT 21.414 19.482 21.468 19.518 ;
      RECT 14.532 19.482 14.586 19.518 ;
      RECT 19.606 19.329 19.654 19.365 ;
      RECT 18.08 19.329 18.12 19.365 ;
      RECT 16.718 19.329 16.772 19.365 ;
      RECT 16.346 19.329 16.394 19.365 ;
      RECT 20.37 19.3345 20.442 19.3595 ;
      RECT 18.764 19.3345 18.836 19.3595 ;
      RECT 15.558 19.3345 15.63 19.3595 ;
      RECT 21.978 19.182 22.022 19.218 ;
      RECT 13.978 19.182 14.022 19.218 ;
      RECT 18.764 19.1875 18.836 19.2125 ;
      RECT 19.762 19.035 19.81 19.071 ;
      RECT 17.616 19.035 17.656 19.071 ;
      RECT 16.19 19.035 16.238 19.071 ;
      RECT 35.254 18.806 35.306 18.842 ;
      RECT 34.854 18.806 34.906 18.842 ;
      RECT 34.454 18.806 34.506 18.842 ;
      RECT 34.054 18.806 34.106 18.842 ;
      RECT 33.654 18.806 33.706 18.842 ;
      RECT 33.254 18.806 33.306 18.842 ;
      RECT 32.854 18.806 32.906 18.842 ;
      RECT 32.454 18.806 32.506 18.842 ;
      RECT 32.054 18.806 32.106 18.842 ;
      RECT 31.654 18.806 31.706 18.842 ;
      RECT 31.254 18.806 31.306 18.842 ;
      RECT 30.854 18.806 30.906 18.842 ;
      RECT 30.454 18.806 30.506 18.842 ;
      RECT 30.054 18.806 30.106 18.842 ;
      RECT 29.654 18.806 29.706 18.842 ;
      RECT 29.254 18.806 29.306 18.842 ;
      RECT 28.854 18.806 28.906 18.842 ;
      RECT 28.454 18.806 28.506 18.842 ;
      RECT 28.054 18.806 28.106 18.842 ;
      RECT 27.654 18.806 27.706 18.842 ;
      RECT 27.254 18.806 27.306 18.842 ;
      RECT 26.854 18.806 26.906 18.842 ;
      RECT 26.454 18.806 26.506 18.842 ;
      RECT 26.054 18.806 26.106 18.842 ;
      RECT 25.654 18.806 25.706 18.842 ;
      RECT 25.254 18.806 25.306 18.842 ;
      RECT 24.854 18.806 24.906 18.842 ;
      RECT 24.454 18.806 24.506 18.842 ;
      RECT 24.054 18.806 24.106 18.842 ;
      RECT 23.654 18.806 23.706 18.842 ;
      RECT 23.254 18.806 23.306 18.842 ;
      RECT 22.854 18.806 22.906 18.842 ;
      RECT 22.694 18.806 22.746 18.842 ;
      RECT 21.732 18.806 21.786 18.842 ;
      RECT 14.214 18.806 14.268 18.842 ;
      RECT 13.054 18.806 13.106 18.842 ;
      RECT 12.654 18.806 12.706 18.842 ;
      RECT 12.254 18.806 12.306 18.842 ;
      RECT 11.854 18.806 11.906 18.842 ;
      RECT 11.454 18.806 11.506 18.842 ;
      RECT 11.054 18.806 11.106 18.842 ;
      RECT 10.654 18.806 10.706 18.842 ;
      RECT 10.254 18.806 10.306 18.842 ;
      RECT 9.854 18.806 9.906 18.842 ;
      RECT 9.454 18.806 9.506 18.842 ;
      RECT 9.054 18.806 9.106 18.842 ;
      RECT 8.654 18.806 8.706 18.842 ;
      RECT 8.254 18.806 8.306 18.842 ;
      RECT 7.854 18.806 7.906 18.842 ;
      RECT 7.454 18.806 7.506 18.842 ;
      RECT 7.054 18.806 7.106 18.842 ;
      RECT 6.654 18.806 6.706 18.842 ;
      RECT 6.254 18.806 6.306 18.842 ;
      RECT 5.854 18.806 5.906 18.842 ;
      RECT 5.454 18.806 5.506 18.842 ;
      RECT 5.054 18.806 5.106 18.842 ;
      RECT 4.654 18.806 4.706 18.842 ;
      RECT 4.254 18.806 4.306 18.842 ;
      RECT 3.854 18.806 3.906 18.842 ;
      RECT 3.454 18.806 3.506 18.842 ;
      RECT 3.054 18.806 3.106 18.842 ;
      RECT 2.654 18.806 2.706 18.842 ;
      RECT 2.254 18.806 2.306 18.842 ;
      RECT 1.854 18.806 1.906 18.842 ;
      RECT 1.454 18.806 1.506 18.842 ;
      RECT 1.054 18.806 1.106 18.842 ;
      RECT 0.654 18.806 0.706 18.842 ;
      RECT 21.978 18.582 22.022 18.618 ;
      RECT 21.096 18.582 21.14 18.618 ;
      RECT 14.86 18.582 14.904 18.618 ;
      RECT 13.978 18.582 14.022 18.618 ;
      RECT 35.494 18.358 35.546 18.394 ;
      RECT 35.094 18.358 35.146 18.394 ;
      RECT 34.694 18.358 34.746 18.394 ;
      RECT 34.294 18.358 34.346 18.394 ;
      RECT 33.894 18.358 33.946 18.394 ;
      RECT 33.494 18.358 33.546 18.394 ;
      RECT 33.094 18.358 33.146 18.394 ;
      RECT 32.694 18.358 32.746 18.394 ;
      RECT 32.294 18.358 32.346 18.394 ;
      RECT 31.894 18.358 31.946 18.394 ;
      RECT 31.494 18.358 31.546 18.394 ;
      RECT 31.094 18.358 31.146 18.394 ;
      RECT 30.694 18.358 30.746 18.394 ;
      RECT 30.294 18.358 30.346 18.394 ;
      RECT 29.894 18.358 29.946 18.394 ;
      RECT 29.494 18.358 29.546 18.394 ;
      RECT 29.094 18.358 29.146 18.394 ;
      RECT 28.694 18.358 28.746 18.394 ;
      RECT 28.294 18.358 28.346 18.394 ;
      RECT 27.894 18.358 27.946 18.394 ;
      RECT 27.494 18.358 27.546 18.394 ;
      RECT 27.094 18.358 27.146 18.394 ;
      RECT 26.694 18.358 26.746 18.394 ;
      RECT 26.294 18.358 26.346 18.394 ;
      RECT 25.894 18.358 25.946 18.394 ;
      RECT 25.494 18.358 25.546 18.394 ;
      RECT 25.094 18.358 25.146 18.394 ;
      RECT 24.694 18.358 24.746 18.394 ;
      RECT 24.294 18.358 24.346 18.394 ;
      RECT 23.894 18.358 23.946 18.394 ;
      RECT 23.494 18.358 23.546 18.394 ;
      RECT 23.094 18.358 23.146 18.394 ;
      RECT 21.814 18.358 21.868 18.394 ;
      RECT 19.838 18.358 19.886 18.394 ;
      RECT 19.53 18.358 19.578 18.394 ;
      RECT 16.882 18.358 16.936 18.394 ;
      RECT 16.422 18.358 16.47 18.394 ;
      RECT 16.114 18.358 16.162 18.394 ;
      RECT 14.132 18.358 14.186 18.394 ;
      RECT 13.294 18.358 13.346 18.394 ;
      RECT 12.894 18.358 12.946 18.394 ;
      RECT 12.494 18.358 12.546 18.394 ;
      RECT 12.094 18.358 12.146 18.394 ;
      RECT 11.694 18.358 11.746 18.394 ;
      RECT 11.294 18.358 11.346 18.394 ;
      RECT 10.894 18.358 10.946 18.394 ;
      RECT 10.494 18.358 10.546 18.394 ;
      RECT 10.094 18.358 10.146 18.394 ;
      RECT 9.694 18.358 9.746 18.394 ;
      RECT 9.294 18.358 9.346 18.394 ;
      RECT 8.894 18.358 8.946 18.394 ;
      RECT 8.494 18.358 8.546 18.394 ;
      RECT 8.094 18.358 8.146 18.394 ;
      RECT 7.694 18.358 7.746 18.394 ;
      RECT 7.294 18.358 7.346 18.394 ;
      RECT 6.894 18.358 6.946 18.394 ;
      RECT 6.494 18.358 6.546 18.394 ;
      RECT 6.094 18.358 6.146 18.394 ;
      RECT 5.694 18.358 5.746 18.394 ;
      RECT 5.294 18.358 5.346 18.394 ;
      RECT 4.894 18.358 4.946 18.394 ;
      RECT 4.494 18.358 4.546 18.394 ;
      RECT 4.094 18.358 4.146 18.394 ;
      RECT 3.694 18.358 3.746 18.394 ;
      RECT 3.294 18.358 3.346 18.394 ;
      RECT 2.894 18.358 2.946 18.394 ;
      RECT 2.494 18.358 2.546 18.394 ;
      RECT 2.094 18.358 2.146 18.394 ;
      RECT 1.694 18.358 1.746 18.394 ;
      RECT 1.294 18.358 1.346 18.394 ;
      RECT 0.894 18.358 0.946 18.394 ;
      RECT 21.414 18.282 21.468 18.318 ;
      RECT 14.532 18.282 14.586 18.318 ;
      RECT 19.606 18.129 19.654 18.165 ;
      RECT 18.08 18.129 18.12 18.165 ;
      RECT 16.718 18.129 16.772 18.165 ;
      RECT 16.346 18.129 16.394 18.165 ;
      RECT 20.37 18.1345 20.442 18.1595 ;
      RECT 18.764 18.1345 18.836 18.1595 ;
      RECT 15.558 18.1345 15.63 18.1595 ;
      RECT 21.978 17.982 22.022 18.018 ;
      RECT 13.978 17.982 14.022 18.018 ;
      RECT 18.764 17.9875 18.836 18.0125 ;
      RECT 19.762 17.835 19.81 17.871 ;
      RECT 17.616 17.835 17.656 17.871 ;
      RECT 16.19 17.835 16.238 17.871 ;
      RECT 35.254 17.606 35.306 17.642 ;
      RECT 34.854 17.606 34.906 17.642 ;
      RECT 34.454 17.606 34.506 17.642 ;
      RECT 34.054 17.606 34.106 17.642 ;
      RECT 33.654 17.606 33.706 17.642 ;
      RECT 33.254 17.606 33.306 17.642 ;
      RECT 32.854 17.606 32.906 17.642 ;
      RECT 32.454 17.606 32.506 17.642 ;
      RECT 32.054 17.606 32.106 17.642 ;
      RECT 31.654 17.606 31.706 17.642 ;
      RECT 31.254 17.606 31.306 17.642 ;
      RECT 30.854 17.606 30.906 17.642 ;
      RECT 30.454 17.606 30.506 17.642 ;
      RECT 30.054 17.606 30.106 17.642 ;
      RECT 29.654 17.606 29.706 17.642 ;
      RECT 29.254 17.606 29.306 17.642 ;
      RECT 28.854 17.606 28.906 17.642 ;
      RECT 28.454 17.606 28.506 17.642 ;
      RECT 28.054 17.606 28.106 17.642 ;
      RECT 27.654 17.606 27.706 17.642 ;
      RECT 27.254 17.606 27.306 17.642 ;
      RECT 26.854 17.606 26.906 17.642 ;
      RECT 26.454 17.606 26.506 17.642 ;
      RECT 26.054 17.606 26.106 17.642 ;
      RECT 25.654 17.606 25.706 17.642 ;
      RECT 25.254 17.606 25.306 17.642 ;
      RECT 24.854 17.606 24.906 17.642 ;
      RECT 24.454 17.606 24.506 17.642 ;
      RECT 24.054 17.606 24.106 17.642 ;
      RECT 23.654 17.606 23.706 17.642 ;
      RECT 23.254 17.606 23.306 17.642 ;
      RECT 22.854 17.606 22.906 17.642 ;
      RECT 22.694 17.606 22.746 17.642 ;
      RECT 21.732 17.606 21.786 17.642 ;
      RECT 14.214 17.606 14.268 17.642 ;
      RECT 13.054 17.606 13.106 17.642 ;
      RECT 12.654 17.606 12.706 17.642 ;
      RECT 12.254 17.606 12.306 17.642 ;
      RECT 11.854 17.606 11.906 17.642 ;
      RECT 11.454 17.606 11.506 17.642 ;
      RECT 11.054 17.606 11.106 17.642 ;
      RECT 10.654 17.606 10.706 17.642 ;
      RECT 10.254 17.606 10.306 17.642 ;
      RECT 9.854 17.606 9.906 17.642 ;
      RECT 9.454 17.606 9.506 17.642 ;
      RECT 9.054 17.606 9.106 17.642 ;
      RECT 8.654 17.606 8.706 17.642 ;
      RECT 8.254 17.606 8.306 17.642 ;
      RECT 7.854 17.606 7.906 17.642 ;
      RECT 7.454 17.606 7.506 17.642 ;
      RECT 7.054 17.606 7.106 17.642 ;
      RECT 6.654 17.606 6.706 17.642 ;
      RECT 6.254 17.606 6.306 17.642 ;
      RECT 5.854 17.606 5.906 17.642 ;
      RECT 5.454 17.606 5.506 17.642 ;
      RECT 5.054 17.606 5.106 17.642 ;
      RECT 4.654 17.606 4.706 17.642 ;
      RECT 4.254 17.606 4.306 17.642 ;
      RECT 3.854 17.606 3.906 17.642 ;
      RECT 3.454 17.606 3.506 17.642 ;
      RECT 3.054 17.606 3.106 17.642 ;
      RECT 2.654 17.606 2.706 17.642 ;
      RECT 2.254 17.606 2.306 17.642 ;
      RECT 1.854 17.606 1.906 17.642 ;
      RECT 1.454 17.606 1.506 17.642 ;
      RECT 1.054 17.606 1.106 17.642 ;
      RECT 0.654 17.606 0.706 17.642 ;
      RECT 21.978 17.382 22.022 17.418 ;
      RECT 21.096 17.382 21.14 17.418 ;
      RECT 14.86 17.382 14.904 17.418 ;
      RECT 13.978 17.382 14.022 17.418 ;
      RECT 35.494 17.158 35.546 17.194 ;
      RECT 35.094 17.158 35.146 17.194 ;
      RECT 34.694 17.158 34.746 17.194 ;
      RECT 34.294 17.158 34.346 17.194 ;
      RECT 33.894 17.158 33.946 17.194 ;
      RECT 33.494 17.158 33.546 17.194 ;
      RECT 33.094 17.158 33.146 17.194 ;
      RECT 32.694 17.158 32.746 17.194 ;
      RECT 32.294 17.158 32.346 17.194 ;
      RECT 31.894 17.158 31.946 17.194 ;
      RECT 31.494 17.158 31.546 17.194 ;
      RECT 31.094 17.158 31.146 17.194 ;
      RECT 30.694 17.158 30.746 17.194 ;
      RECT 30.294 17.158 30.346 17.194 ;
      RECT 29.894 17.158 29.946 17.194 ;
      RECT 29.494 17.158 29.546 17.194 ;
      RECT 29.094 17.158 29.146 17.194 ;
      RECT 28.694 17.158 28.746 17.194 ;
      RECT 28.294 17.158 28.346 17.194 ;
      RECT 27.894 17.158 27.946 17.194 ;
      RECT 27.494 17.158 27.546 17.194 ;
      RECT 27.094 17.158 27.146 17.194 ;
      RECT 26.694 17.158 26.746 17.194 ;
      RECT 26.294 17.158 26.346 17.194 ;
      RECT 25.894 17.158 25.946 17.194 ;
      RECT 25.494 17.158 25.546 17.194 ;
      RECT 25.094 17.158 25.146 17.194 ;
      RECT 24.694 17.158 24.746 17.194 ;
      RECT 24.294 17.158 24.346 17.194 ;
      RECT 23.894 17.158 23.946 17.194 ;
      RECT 23.494 17.158 23.546 17.194 ;
      RECT 23.094 17.158 23.146 17.194 ;
      RECT 21.814 17.158 21.868 17.194 ;
      RECT 19.838 17.158 19.886 17.194 ;
      RECT 19.53 17.158 19.578 17.194 ;
      RECT 16.882 17.158 16.936 17.194 ;
      RECT 16.422 17.158 16.47 17.194 ;
      RECT 16.114 17.158 16.162 17.194 ;
      RECT 14.132 17.158 14.186 17.194 ;
      RECT 13.294 17.158 13.346 17.194 ;
      RECT 12.894 17.158 12.946 17.194 ;
      RECT 12.494 17.158 12.546 17.194 ;
      RECT 12.094 17.158 12.146 17.194 ;
      RECT 11.694 17.158 11.746 17.194 ;
      RECT 11.294 17.158 11.346 17.194 ;
      RECT 10.894 17.158 10.946 17.194 ;
      RECT 10.494 17.158 10.546 17.194 ;
      RECT 10.094 17.158 10.146 17.194 ;
      RECT 9.694 17.158 9.746 17.194 ;
      RECT 9.294 17.158 9.346 17.194 ;
      RECT 8.894 17.158 8.946 17.194 ;
      RECT 8.494 17.158 8.546 17.194 ;
      RECT 8.094 17.158 8.146 17.194 ;
      RECT 7.694 17.158 7.746 17.194 ;
      RECT 7.294 17.158 7.346 17.194 ;
      RECT 6.894 17.158 6.946 17.194 ;
      RECT 6.494 17.158 6.546 17.194 ;
      RECT 6.094 17.158 6.146 17.194 ;
      RECT 5.694 17.158 5.746 17.194 ;
      RECT 5.294 17.158 5.346 17.194 ;
      RECT 4.894 17.158 4.946 17.194 ;
      RECT 4.494 17.158 4.546 17.194 ;
      RECT 4.094 17.158 4.146 17.194 ;
      RECT 3.694 17.158 3.746 17.194 ;
      RECT 3.294 17.158 3.346 17.194 ;
      RECT 2.894 17.158 2.946 17.194 ;
      RECT 2.494 17.158 2.546 17.194 ;
      RECT 2.094 17.158 2.146 17.194 ;
      RECT 1.694 17.158 1.746 17.194 ;
      RECT 1.294 17.158 1.346 17.194 ;
      RECT 0.894 17.158 0.946 17.194 ;
      RECT 21.414 17.082 21.468 17.118 ;
      RECT 14.532 17.082 14.586 17.118 ;
      RECT 19.606 16.929 19.654 16.965 ;
      RECT 18.08 16.929 18.12 16.965 ;
      RECT 16.718 16.929 16.772 16.965 ;
      RECT 16.346 16.929 16.394 16.965 ;
      RECT 20.37 16.9345 20.442 16.9595 ;
      RECT 18.764 16.9345 18.836 16.9595 ;
      RECT 15.558 16.9345 15.63 16.9595 ;
      RECT 21.978 16.782 22.022 16.818 ;
      RECT 13.978 16.782 14.022 16.818 ;
      RECT 18.764 16.7875 18.836 16.8125 ;
      RECT 19.762 16.635 19.81 16.671 ;
      RECT 17.616 16.635 17.656 16.671 ;
      RECT 16.19 16.635 16.238 16.671 ;
      RECT 35.254 16.406 35.306 16.442 ;
      RECT 34.854 16.406 34.906 16.442 ;
      RECT 34.454 16.406 34.506 16.442 ;
      RECT 34.054 16.406 34.106 16.442 ;
      RECT 33.654 16.406 33.706 16.442 ;
      RECT 33.254 16.406 33.306 16.442 ;
      RECT 32.854 16.406 32.906 16.442 ;
      RECT 32.454 16.406 32.506 16.442 ;
      RECT 32.054 16.406 32.106 16.442 ;
      RECT 31.654 16.406 31.706 16.442 ;
      RECT 31.254 16.406 31.306 16.442 ;
      RECT 30.854 16.406 30.906 16.442 ;
      RECT 30.454 16.406 30.506 16.442 ;
      RECT 30.054 16.406 30.106 16.442 ;
      RECT 29.654 16.406 29.706 16.442 ;
      RECT 29.254 16.406 29.306 16.442 ;
      RECT 28.854 16.406 28.906 16.442 ;
      RECT 28.454 16.406 28.506 16.442 ;
      RECT 28.054 16.406 28.106 16.442 ;
      RECT 27.654 16.406 27.706 16.442 ;
      RECT 27.254 16.406 27.306 16.442 ;
      RECT 26.854 16.406 26.906 16.442 ;
      RECT 26.454 16.406 26.506 16.442 ;
      RECT 26.054 16.406 26.106 16.442 ;
      RECT 25.654 16.406 25.706 16.442 ;
      RECT 25.254 16.406 25.306 16.442 ;
      RECT 24.854 16.406 24.906 16.442 ;
      RECT 24.454 16.406 24.506 16.442 ;
      RECT 24.054 16.406 24.106 16.442 ;
      RECT 23.654 16.406 23.706 16.442 ;
      RECT 23.254 16.406 23.306 16.442 ;
      RECT 22.854 16.406 22.906 16.442 ;
      RECT 22.694 16.406 22.746 16.442 ;
      RECT 21.732 16.406 21.786 16.442 ;
      RECT 14.214 16.406 14.268 16.442 ;
      RECT 13.054 16.406 13.106 16.442 ;
      RECT 12.654 16.406 12.706 16.442 ;
      RECT 12.254 16.406 12.306 16.442 ;
      RECT 11.854 16.406 11.906 16.442 ;
      RECT 11.454 16.406 11.506 16.442 ;
      RECT 11.054 16.406 11.106 16.442 ;
      RECT 10.654 16.406 10.706 16.442 ;
      RECT 10.254 16.406 10.306 16.442 ;
      RECT 9.854 16.406 9.906 16.442 ;
      RECT 9.454 16.406 9.506 16.442 ;
      RECT 9.054 16.406 9.106 16.442 ;
      RECT 8.654 16.406 8.706 16.442 ;
      RECT 8.254 16.406 8.306 16.442 ;
      RECT 7.854 16.406 7.906 16.442 ;
      RECT 7.454 16.406 7.506 16.442 ;
      RECT 7.054 16.406 7.106 16.442 ;
      RECT 6.654 16.406 6.706 16.442 ;
      RECT 6.254 16.406 6.306 16.442 ;
      RECT 5.854 16.406 5.906 16.442 ;
      RECT 5.454 16.406 5.506 16.442 ;
      RECT 5.054 16.406 5.106 16.442 ;
      RECT 4.654 16.406 4.706 16.442 ;
      RECT 4.254 16.406 4.306 16.442 ;
      RECT 3.854 16.406 3.906 16.442 ;
      RECT 3.454 16.406 3.506 16.442 ;
      RECT 3.054 16.406 3.106 16.442 ;
      RECT 2.654 16.406 2.706 16.442 ;
      RECT 2.254 16.406 2.306 16.442 ;
      RECT 1.854 16.406 1.906 16.442 ;
      RECT 1.454 16.406 1.506 16.442 ;
      RECT 1.054 16.406 1.106 16.442 ;
      RECT 0.654 16.406 0.706 16.442 ;
      RECT 21.978 16.182 22.022 16.218 ;
      RECT 21.096 16.182 21.14 16.218 ;
      RECT 14.86 16.182 14.904 16.218 ;
      RECT 13.978 16.182 14.022 16.218 ;
      RECT 35.494 15.958 35.546 15.994 ;
      RECT 35.094 15.958 35.146 15.994 ;
      RECT 34.694 15.958 34.746 15.994 ;
      RECT 34.294 15.958 34.346 15.994 ;
      RECT 33.894 15.958 33.946 15.994 ;
      RECT 33.494 15.958 33.546 15.994 ;
      RECT 33.094 15.958 33.146 15.994 ;
      RECT 32.694 15.958 32.746 15.994 ;
      RECT 32.294 15.958 32.346 15.994 ;
      RECT 31.894 15.958 31.946 15.994 ;
      RECT 31.494 15.958 31.546 15.994 ;
      RECT 31.094 15.958 31.146 15.994 ;
      RECT 30.694 15.958 30.746 15.994 ;
      RECT 30.294 15.958 30.346 15.994 ;
      RECT 29.894 15.958 29.946 15.994 ;
      RECT 29.494 15.958 29.546 15.994 ;
      RECT 29.094 15.958 29.146 15.994 ;
      RECT 28.694 15.958 28.746 15.994 ;
      RECT 28.294 15.958 28.346 15.994 ;
      RECT 27.894 15.958 27.946 15.994 ;
      RECT 27.494 15.958 27.546 15.994 ;
      RECT 27.094 15.958 27.146 15.994 ;
      RECT 26.694 15.958 26.746 15.994 ;
      RECT 26.294 15.958 26.346 15.994 ;
      RECT 25.894 15.958 25.946 15.994 ;
      RECT 25.494 15.958 25.546 15.994 ;
      RECT 25.094 15.958 25.146 15.994 ;
      RECT 24.694 15.958 24.746 15.994 ;
      RECT 24.294 15.958 24.346 15.994 ;
      RECT 23.894 15.958 23.946 15.994 ;
      RECT 23.494 15.958 23.546 15.994 ;
      RECT 23.094 15.958 23.146 15.994 ;
      RECT 21.814 15.958 21.868 15.994 ;
      RECT 19.838 15.958 19.886 15.994 ;
      RECT 19.53 15.958 19.578 15.994 ;
      RECT 16.882 15.958 16.936 15.994 ;
      RECT 16.422 15.958 16.47 15.994 ;
      RECT 16.114 15.958 16.162 15.994 ;
      RECT 14.132 15.958 14.186 15.994 ;
      RECT 13.294 15.958 13.346 15.994 ;
      RECT 12.894 15.958 12.946 15.994 ;
      RECT 12.494 15.958 12.546 15.994 ;
      RECT 12.094 15.958 12.146 15.994 ;
      RECT 11.694 15.958 11.746 15.994 ;
      RECT 11.294 15.958 11.346 15.994 ;
      RECT 10.894 15.958 10.946 15.994 ;
      RECT 10.494 15.958 10.546 15.994 ;
      RECT 10.094 15.958 10.146 15.994 ;
      RECT 9.694 15.958 9.746 15.994 ;
      RECT 9.294 15.958 9.346 15.994 ;
      RECT 8.894 15.958 8.946 15.994 ;
      RECT 8.494 15.958 8.546 15.994 ;
      RECT 8.094 15.958 8.146 15.994 ;
      RECT 7.694 15.958 7.746 15.994 ;
      RECT 7.294 15.958 7.346 15.994 ;
      RECT 6.894 15.958 6.946 15.994 ;
      RECT 6.494 15.958 6.546 15.994 ;
      RECT 6.094 15.958 6.146 15.994 ;
      RECT 5.694 15.958 5.746 15.994 ;
      RECT 5.294 15.958 5.346 15.994 ;
      RECT 4.894 15.958 4.946 15.994 ;
      RECT 4.494 15.958 4.546 15.994 ;
      RECT 4.094 15.958 4.146 15.994 ;
      RECT 3.694 15.958 3.746 15.994 ;
      RECT 3.294 15.958 3.346 15.994 ;
      RECT 2.894 15.958 2.946 15.994 ;
      RECT 2.494 15.958 2.546 15.994 ;
      RECT 2.094 15.958 2.146 15.994 ;
      RECT 1.694 15.958 1.746 15.994 ;
      RECT 1.294 15.958 1.346 15.994 ;
      RECT 0.894 15.958 0.946 15.994 ;
      RECT 21.414 15.882 21.468 15.918 ;
      RECT 14.532 15.882 14.586 15.918 ;
      RECT 19.606 15.729 19.654 15.765 ;
      RECT 18.08 15.729 18.12 15.765 ;
      RECT 16.718 15.729 16.772 15.765 ;
      RECT 16.346 15.729 16.394 15.765 ;
      RECT 20.37 15.7345 20.442 15.7595 ;
      RECT 18.764 15.7345 18.836 15.7595 ;
      RECT 15.558 15.7345 15.63 15.7595 ;
      RECT 21.978 15.582 22.022 15.618 ;
      RECT 13.978 15.582 14.022 15.618 ;
      RECT 18.764 15.5875 18.836 15.6125 ;
      RECT 19.762 15.435 19.81 15.471 ;
      RECT 17.616 15.435 17.656 15.471 ;
      RECT 16.19 15.435 16.238 15.471 ;
      RECT 35.254 15.206 35.306 15.242 ;
      RECT 34.854 15.206 34.906 15.242 ;
      RECT 34.454 15.206 34.506 15.242 ;
      RECT 34.054 15.206 34.106 15.242 ;
      RECT 33.654 15.206 33.706 15.242 ;
      RECT 33.254 15.206 33.306 15.242 ;
      RECT 32.854 15.206 32.906 15.242 ;
      RECT 32.454 15.206 32.506 15.242 ;
      RECT 32.054 15.206 32.106 15.242 ;
      RECT 31.654 15.206 31.706 15.242 ;
      RECT 31.254 15.206 31.306 15.242 ;
      RECT 30.854 15.206 30.906 15.242 ;
      RECT 30.454 15.206 30.506 15.242 ;
      RECT 30.054 15.206 30.106 15.242 ;
      RECT 29.654 15.206 29.706 15.242 ;
      RECT 29.254 15.206 29.306 15.242 ;
      RECT 28.854 15.206 28.906 15.242 ;
      RECT 28.454 15.206 28.506 15.242 ;
      RECT 28.054 15.206 28.106 15.242 ;
      RECT 27.654 15.206 27.706 15.242 ;
      RECT 27.254 15.206 27.306 15.242 ;
      RECT 26.854 15.206 26.906 15.242 ;
      RECT 26.454 15.206 26.506 15.242 ;
      RECT 26.054 15.206 26.106 15.242 ;
      RECT 25.654 15.206 25.706 15.242 ;
      RECT 25.254 15.206 25.306 15.242 ;
      RECT 24.854 15.206 24.906 15.242 ;
      RECT 24.454 15.206 24.506 15.242 ;
      RECT 24.054 15.206 24.106 15.242 ;
      RECT 23.654 15.206 23.706 15.242 ;
      RECT 23.254 15.206 23.306 15.242 ;
      RECT 22.854 15.206 22.906 15.242 ;
      RECT 22.694 15.206 22.746 15.242 ;
      RECT 21.732 15.206 21.786 15.242 ;
      RECT 14.214 15.206 14.268 15.242 ;
      RECT 13.054 15.206 13.106 15.242 ;
      RECT 12.654 15.206 12.706 15.242 ;
      RECT 12.254 15.206 12.306 15.242 ;
      RECT 11.854 15.206 11.906 15.242 ;
      RECT 11.454 15.206 11.506 15.242 ;
      RECT 11.054 15.206 11.106 15.242 ;
      RECT 10.654 15.206 10.706 15.242 ;
      RECT 10.254 15.206 10.306 15.242 ;
      RECT 9.854 15.206 9.906 15.242 ;
      RECT 9.454 15.206 9.506 15.242 ;
      RECT 9.054 15.206 9.106 15.242 ;
      RECT 8.654 15.206 8.706 15.242 ;
      RECT 8.254 15.206 8.306 15.242 ;
      RECT 7.854 15.206 7.906 15.242 ;
      RECT 7.454 15.206 7.506 15.242 ;
      RECT 7.054 15.206 7.106 15.242 ;
      RECT 6.654 15.206 6.706 15.242 ;
      RECT 6.254 15.206 6.306 15.242 ;
      RECT 5.854 15.206 5.906 15.242 ;
      RECT 5.454 15.206 5.506 15.242 ;
      RECT 5.054 15.206 5.106 15.242 ;
      RECT 4.654 15.206 4.706 15.242 ;
      RECT 4.254 15.206 4.306 15.242 ;
      RECT 3.854 15.206 3.906 15.242 ;
      RECT 3.454 15.206 3.506 15.242 ;
      RECT 3.054 15.206 3.106 15.242 ;
      RECT 2.654 15.206 2.706 15.242 ;
      RECT 2.254 15.206 2.306 15.242 ;
      RECT 1.854 15.206 1.906 15.242 ;
      RECT 1.454 15.206 1.506 15.242 ;
      RECT 1.054 15.206 1.106 15.242 ;
      RECT 0.654 15.206 0.706 15.242 ;
      RECT 21.978 14.982 22.022 15.018 ;
      RECT 21.096 14.982 21.14 15.018 ;
      RECT 14.86 14.982 14.904 15.018 ;
      RECT 13.978 14.982 14.022 15.018 ;
      RECT 35.494 14.758 35.546 14.794 ;
      RECT 35.094 14.758 35.146 14.794 ;
      RECT 34.694 14.758 34.746 14.794 ;
      RECT 34.294 14.758 34.346 14.794 ;
      RECT 33.894 14.758 33.946 14.794 ;
      RECT 33.494 14.758 33.546 14.794 ;
      RECT 33.094 14.758 33.146 14.794 ;
      RECT 32.694 14.758 32.746 14.794 ;
      RECT 32.294 14.758 32.346 14.794 ;
      RECT 31.894 14.758 31.946 14.794 ;
      RECT 31.494 14.758 31.546 14.794 ;
      RECT 31.094 14.758 31.146 14.794 ;
      RECT 30.694 14.758 30.746 14.794 ;
      RECT 30.294 14.758 30.346 14.794 ;
      RECT 29.894 14.758 29.946 14.794 ;
      RECT 29.494 14.758 29.546 14.794 ;
      RECT 29.094 14.758 29.146 14.794 ;
      RECT 28.694 14.758 28.746 14.794 ;
      RECT 28.294 14.758 28.346 14.794 ;
      RECT 27.894 14.758 27.946 14.794 ;
      RECT 27.494 14.758 27.546 14.794 ;
      RECT 27.094 14.758 27.146 14.794 ;
      RECT 26.694 14.758 26.746 14.794 ;
      RECT 26.294 14.758 26.346 14.794 ;
      RECT 25.894 14.758 25.946 14.794 ;
      RECT 25.494 14.758 25.546 14.794 ;
      RECT 25.094 14.758 25.146 14.794 ;
      RECT 24.694 14.758 24.746 14.794 ;
      RECT 24.294 14.758 24.346 14.794 ;
      RECT 23.894 14.758 23.946 14.794 ;
      RECT 23.494 14.758 23.546 14.794 ;
      RECT 23.094 14.758 23.146 14.794 ;
      RECT 21.814 14.758 21.868 14.794 ;
      RECT 19.838 14.758 19.886 14.794 ;
      RECT 19.53 14.758 19.578 14.794 ;
      RECT 16.882 14.758 16.936 14.794 ;
      RECT 16.422 14.758 16.47 14.794 ;
      RECT 16.114 14.758 16.162 14.794 ;
      RECT 14.132 14.758 14.186 14.794 ;
      RECT 13.294 14.758 13.346 14.794 ;
      RECT 12.894 14.758 12.946 14.794 ;
      RECT 12.494 14.758 12.546 14.794 ;
      RECT 12.094 14.758 12.146 14.794 ;
      RECT 11.694 14.758 11.746 14.794 ;
      RECT 11.294 14.758 11.346 14.794 ;
      RECT 10.894 14.758 10.946 14.794 ;
      RECT 10.494 14.758 10.546 14.794 ;
      RECT 10.094 14.758 10.146 14.794 ;
      RECT 9.694 14.758 9.746 14.794 ;
      RECT 9.294 14.758 9.346 14.794 ;
      RECT 8.894 14.758 8.946 14.794 ;
      RECT 8.494 14.758 8.546 14.794 ;
      RECT 8.094 14.758 8.146 14.794 ;
      RECT 7.694 14.758 7.746 14.794 ;
      RECT 7.294 14.758 7.346 14.794 ;
      RECT 6.894 14.758 6.946 14.794 ;
      RECT 6.494 14.758 6.546 14.794 ;
      RECT 6.094 14.758 6.146 14.794 ;
      RECT 5.694 14.758 5.746 14.794 ;
      RECT 5.294 14.758 5.346 14.794 ;
      RECT 4.894 14.758 4.946 14.794 ;
      RECT 4.494 14.758 4.546 14.794 ;
      RECT 4.094 14.758 4.146 14.794 ;
      RECT 3.694 14.758 3.746 14.794 ;
      RECT 3.294 14.758 3.346 14.794 ;
      RECT 2.894 14.758 2.946 14.794 ;
      RECT 2.494 14.758 2.546 14.794 ;
      RECT 2.094 14.758 2.146 14.794 ;
      RECT 1.694 14.758 1.746 14.794 ;
      RECT 1.294 14.758 1.346 14.794 ;
      RECT 0.894 14.758 0.946 14.794 ;
      RECT 21.414 14.682 21.468 14.718 ;
      RECT 14.532 14.682 14.586 14.718 ;
      RECT 19.606 14.529 19.654 14.565 ;
      RECT 18.08 14.529 18.12 14.565 ;
      RECT 16.718 14.529 16.772 14.565 ;
      RECT 16.346 14.529 16.394 14.565 ;
      RECT 20.37 14.5345 20.442 14.5595 ;
      RECT 18.764 14.5345 18.836 14.5595 ;
      RECT 15.558 14.5345 15.63 14.5595 ;
      RECT 21.978 14.382 22.022 14.418 ;
      RECT 13.978 14.382 14.022 14.418 ;
      RECT 18.764 14.3875 18.836 14.4125 ;
      RECT 19.762 14.235 19.81 14.271 ;
      RECT 17.616 14.235 17.656 14.271 ;
      RECT 16.19 14.235 16.238 14.271 ;
      RECT 35.254 14.006 35.306 14.042 ;
      RECT 34.854 14.006 34.906 14.042 ;
      RECT 34.454 14.006 34.506 14.042 ;
      RECT 34.054 14.006 34.106 14.042 ;
      RECT 33.654 14.006 33.706 14.042 ;
      RECT 33.254 14.006 33.306 14.042 ;
      RECT 32.854 14.006 32.906 14.042 ;
      RECT 32.454 14.006 32.506 14.042 ;
      RECT 32.054 14.006 32.106 14.042 ;
      RECT 31.654 14.006 31.706 14.042 ;
      RECT 31.254 14.006 31.306 14.042 ;
      RECT 30.854 14.006 30.906 14.042 ;
      RECT 30.454 14.006 30.506 14.042 ;
      RECT 30.054 14.006 30.106 14.042 ;
      RECT 29.654 14.006 29.706 14.042 ;
      RECT 29.254 14.006 29.306 14.042 ;
      RECT 28.854 14.006 28.906 14.042 ;
      RECT 28.454 14.006 28.506 14.042 ;
      RECT 28.054 14.006 28.106 14.042 ;
      RECT 27.654 14.006 27.706 14.042 ;
      RECT 27.254 14.006 27.306 14.042 ;
      RECT 26.854 14.006 26.906 14.042 ;
      RECT 26.454 14.006 26.506 14.042 ;
      RECT 26.054 14.006 26.106 14.042 ;
      RECT 25.654 14.006 25.706 14.042 ;
      RECT 25.254 14.006 25.306 14.042 ;
      RECT 24.854 14.006 24.906 14.042 ;
      RECT 24.454 14.006 24.506 14.042 ;
      RECT 24.054 14.006 24.106 14.042 ;
      RECT 23.654 14.006 23.706 14.042 ;
      RECT 23.254 14.006 23.306 14.042 ;
      RECT 22.854 14.006 22.906 14.042 ;
      RECT 22.694 14.006 22.746 14.042 ;
      RECT 21.732 14.006 21.786 14.042 ;
      RECT 14.214 14.006 14.268 14.042 ;
      RECT 13.054 14.006 13.106 14.042 ;
      RECT 12.654 14.006 12.706 14.042 ;
      RECT 12.254 14.006 12.306 14.042 ;
      RECT 11.854 14.006 11.906 14.042 ;
      RECT 11.454 14.006 11.506 14.042 ;
      RECT 11.054 14.006 11.106 14.042 ;
      RECT 10.654 14.006 10.706 14.042 ;
      RECT 10.254 14.006 10.306 14.042 ;
      RECT 9.854 14.006 9.906 14.042 ;
      RECT 9.454 14.006 9.506 14.042 ;
      RECT 9.054 14.006 9.106 14.042 ;
      RECT 8.654 14.006 8.706 14.042 ;
      RECT 8.254 14.006 8.306 14.042 ;
      RECT 7.854 14.006 7.906 14.042 ;
      RECT 7.454 14.006 7.506 14.042 ;
      RECT 7.054 14.006 7.106 14.042 ;
      RECT 6.654 14.006 6.706 14.042 ;
      RECT 6.254 14.006 6.306 14.042 ;
      RECT 5.854 14.006 5.906 14.042 ;
      RECT 5.454 14.006 5.506 14.042 ;
      RECT 5.054 14.006 5.106 14.042 ;
      RECT 4.654 14.006 4.706 14.042 ;
      RECT 4.254 14.006 4.306 14.042 ;
      RECT 3.854 14.006 3.906 14.042 ;
      RECT 3.454 14.006 3.506 14.042 ;
      RECT 3.054 14.006 3.106 14.042 ;
      RECT 2.654 14.006 2.706 14.042 ;
      RECT 2.254 14.006 2.306 14.042 ;
      RECT 1.854 14.006 1.906 14.042 ;
      RECT 1.454 14.006 1.506 14.042 ;
      RECT 1.054 14.006 1.106 14.042 ;
      RECT 0.654 14.006 0.706 14.042 ;
      RECT 21.978 13.782 22.022 13.818 ;
      RECT 21.096 13.782 21.14 13.818 ;
      RECT 14.86 13.782 14.904 13.818 ;
      RECT 13.978 13.782 14.022 13.818 ;
      RECT 35.494 13.558 35.546 13.594 ;
      RECT 35.094 13.558 35.146 13.594 ;
      RECT 34.694 13.558 34.746 13.594 ;
      RECT 34.294 13.558 34.346 13.594 ;
      RECT 33.894 13.558 33.946 13.594 ;
      RECT 33.494 13.558 33.546 13.594 ;
      RECT 33.094 13.558 33.146 13.594 ;
      RECT 32.694 13.558 32.746 13.594 ;
      RECT 32.294 13.558 32.346 13.594 ;
      RECT 31.894 13.558 31.946 13.594 ;
      RECT 31.494 13.558 31.546 13.594 ;
      RECT 31.094 13.558 31.146 13.594 ;
      RECT 30.694 13.558 30.746 13.594 ;
      RECT 30.294 13.558 30.346 13.594 ;
      RECT 29.894 13.558 29.946 13.594 ;
      RECT 29.494 13.558 29.546 13.594 ;
      RECT 29.094 13.558 29.146 13.594 ;
      RECT 28.694 13.558 28.746 13.594 ;
      RECT 28.294 13.558 28.346 13.594 ;
      RECT 27.894 13.558 27.946 13.594 ;
      RECT 27.494 13.558 27.546 13.594 ;
      RECT 27.094 13.558 27.146 13.594 ;
      RECT 26.694 13.558 26.746 13.594 ;
      RECT 26.294 13.558 26.346 13.594 ;
      RECT 25.894 13.558 25.946 13.594 ;
      RECT 25.494 13.558 25.546 13.594 ;
      RECT 25.094 13.558 25.146 13.594 ;
      RECT 24.694 13.558 24.746 13.594 ;
      RECT 24.294 13.558 24.346 13.594 ;
      RECT 23.894 13.558 23.946 13.594 ;
      RECT 23.494 13.558 23.546 13.594 ;
      RECT 23.094 13.558 23.146 13.594 ;
      RECT 21.814 13.558 21.868 13.594 ;
      RECT 19.838 13.558 19.886 13.594 ;
      RECT 19.53 13.558 19.578 13.594 ;
      RECT 16.882 13.558 16.936 13.594 ;
      RECT 16.422 13.558 16.47 13.594 ;
      RECT 16.114 13.558 16.162 13.594 ;
      RECT 14.132 13.558 14.186 13.594 ;
      RECT 13.294 13.558 13.346 13.594 ;
      RECT 12.894 13.558 12.946 13.594 ;
      RECT 12.494 13.558 12.546 13.594 ;
      RECT 12.094 13.558 12.146 13.594 ;
      RECT 11.694 13.558 11.746 13.594 ;
      RECT 11.294 13.558 11.346 13.594 ;
      RECT 10.894 13.558 10.946 13.594 ;
      RECT 10.494 13.558 10.546 13.594 ;
      RECT 10.094 13.558 10.146 13.594 ;
      RECT 9.694 13.558 9.746 13.594 ;
      RECT 9.294 13.558 9.346 13.594 ;
      RECT 8.894 13.558 8.946 13.594 ;
      RECT 8.494 13.558 8.546 13.594 ;
      RECT 8.094 13.558 8.146 13.594 ;
      RECT 7.694 13.558 7.746 13.594 ;
      RECT 7.294 13.558 7.346 13.594 ;
      RECT 6.894 13.558 6.946 13.594 ;
      RECT 6.494 13.558 6.546 13.594 ;
      RECT 6.094 13.558 6.146 13.594 ;
      RECT 5.694 13.558 5.746 13.594 ;
      RECT 5.294 13.558 5.346 13.594 ;
      RECT 4.894 13.558 4.946 13.594 ;
      RECT 4.494 13.558 4.546 13.594 ;
      RECT 4.094 13.558 4.146 13.594 ;
      RECT 3.694 13.558 3.746 13.594 ;
      RECT 3.294 13.558 3.346 13.594 ;
      RECT 2.894 13.558 2.946 13.594 ;
      RECT 2.494 13.558 2.546 13.594 ;
      RECT 2.094 13.558 2.146 13.594 ;
      RECT 1.694 13.558 1.746 13.594 ;
      RECT 1.294 13.558 1.346 13.594 ;
      RECT 0.894 13.558 0.946 13.594 ;
      RECT 21.414 13.482 21.468 13.518 ;
      RECT 14.532 13.482 14.586 13.518 ;
      RECT 19.606 13.329 19.654 13.365 ;
      RECT 18.08 13.329 18.12 13.365 ;
      RECT 16.718 13.329 16.772 13.365 ;
      RECT 16.346 13.329 16.394 13.365 ;
      RECT 20.37 13.3345 20.442 13.3595 ;
      RECT 18.764 13.3345 18.836 13.3595 ;
      RECT 15.558 13.3345 15.63 13.3595 ;
      RECT 21.978 13.182 22.022 13.218 ;
      RECT 13.978 13.182 14.022 13.218 ;
      RECT 18.764 13.1875 18.836 13.2125 ;
      RECT 19.762 13.035 19.81 13.071 ;
      RECT 17.616 13.035 17.656 13.071 ;
      RECT 16.19 13.035 16.238 13.071 ;
      RECT 35.254 12.806 35.306 12.842 ;
      RECT 34.854 12.806 34.906 12.842 ;
      RECT 34.454 12.806 34.506 12.842 ;
      RECT 34.054 12.806 34.106 12.842 ;
      RECT 33.654 12.806 33.706 12.842 ;
      RECT 33.254 12.806 33.306 12.842 ;
      RECT 32.854 12.806 32.906 12.842 ;
      RECT 32.454 12.806 32.506 12.842 ;
      RECT 32.054 12.806 32.106 12.842 ;
      RECT 31.654 12.806 31.706 12.842 ;
      RECT 31.254 12.806 31.306 12.842 ;
      RECT 30.854 12.806 30.906 12.842 ;
      RECT 30.454 12.806 30.506 12.842 ;
      RECT 30.054 12.806 30.106 12.842 ;
      RECT 29.654 12.806 29.706 12.842 ;
      RECT 29.254 12.806 29.306 12.842 ;
      RECT 28.854 12.806 28.906 12.842 ;
      RECT 28.454 12.806 28.506 12.842 ;
      RECT 28.054 12.806 28.106 12.842 ;
      RECT 27.654 12.806 27.706 12.842 ;
      RECT 27.254 12.806 27.306 12.842 ;
      RECT 26.854 12.806 26.906 12.842 ;
      RECT 26.454 12.806 26.506 12.842 ;
      RECT 26.054 12.806 26.106 12.842 ;
      RECT 25.654 12.806 25.706 12.842 ;
      RECT 25.254 12.806 25.306 12.842 ;
      RECT 24.854 12.806 24.906 12.842 ;
      RECT 24.454 12.806 24.506 12.842 ;
      RECT 24.054 12.806 24.106 12.842 ;
      RECT 23.654 12.806 23.706 12.842 ;
      RECT 23.254 12.806 23.306 12.842 ;
      RECT 22.854 12.806 22.906 12.842 ;
      RECT 22.694 12.806 22.746 12.842 ;
      RECT 21.732 12.806 21.786 12.842 ;
      RECT 14.214 12.806 14.268 12.842 ;
      RECT 13.054 12.806 13.106 12.842 ;
      RECT 12.654 12.806 12.706 12.842 ;
      RECT 12.254 12.806 12.306 12.842 ;
      RECT 11.854 12.806 11.906 12.842 ;
      RECT 11.454 12.806 11.506 12.842 ;
      RECT 11.054 12.806 11.106 12.842 ;
      RECT 10.654 12.806 10.706 12.842 ;
      RECT 10.254 12.806 10.306 12.842 ;
      RECT 9.854 12.806 9.906 12.842 ;
      RECT 9.454 12.806 9.506 12.842 ;
      RECT 9.054 12.806 9.106 12.842 ;
      RECT 8.654 12.806 8.706 12.842 ;
      RECT 8.254 12.806 8.306 12.842 ;
      RECT 7.854 12.806 7.906 12.842 ;
      RECT 7.454 12.806 7.506 12.842 ;
      RECT 7.054 12.806 7.106 12.842 ;
      RECT 6.654 12.806 6.706 12.842 ;
      RECT 6.254 12.806 6.306 12.842 ;
      RECT 5.854 12.806 5.906 12.842 ;
      RECT 5.454 12.806 5.506 12.842 ;
      RECT 5.054 12.806 5.106 12.842 ;
      RECT 4.654 12.806 4.706 12.842 ;
      RECT 4.254 12.806 4.306 12.842 ;
      RECT 3.854 12.806 3.906 12.842 ;
      RECT 3.454 12.806 3.506 12.842 ;
      RECT 3.054 12.806 3.106 12.842 ;
      RECT 2.654 12.806 2.706 12.842 ;
      RECT 2.254 12.806 2.306 12.842 ;
      RECT 1.854 12.806 1.906 12.842 ;
      RECT 1.454 12.806 1.506 12.842 ;
      RECT 1.054 12.806 1.106 12.842 ;
      RECT 0.654 12.806 0.706 12.842 ;
      RECT 21.978 12.582 22.022 12.618 ;
      RECT 21.096 12.582 21.14 12.618 ;
      RECT 14.86 12.582 14.904 12.618 ;
      RECT 13.978 12.582 14.022 12.618 ;
      RECT 35.494 12.358 35.546 12.394 ;
      RECT 35.094 12.358 35.146 12.394 ;
      RECT 34.694 12.358 34.746 12.394 ;
      RECT 34.294 12.358 34.346 12.394 ;
      RECT 33.894 12.358 33.946 12.394 ;
      RECT 33.494 12.358 33.546 12.394 ;
      RECT 33.094 12.358 33.146 12.394 ;
      RECT 32.694 12.358 32.746 12.394 ;
      RECT 32.294 12.358 32.346 12.394 ;
      RECT 31.894 12.358 31.946 12.394 ;
      RECT 31.494 12.358 31.546 12.394 ;
      RECT 31.094 12.358 31.146 12.394 ;
      RECT 30.694 12.358 30.746 12.394 ;
      RECT 30.294 12.358 30.346 12.394 ;
      RECT 29.894 12.358 29.946 12.394 ;
      RECT 29.494 12.358 29.546 12.394 ;
      RECT 29.094 12.358 29.146 12.394 ;
      RECT 28.694 12.358 28.746 12.394 ;
      RECT 28.294 12.358 28.346 12.394 ;
      RECT 27.894 12.358 27.946 12.394 ;
      RECT 27.494 12.358 27.546 12.394 ;
      RECT 27.094 12.358 27.146 12.394 ;
      RECT 26.694 12.358 26.746 12.394 ;
      RECT 26.294 12.358 26.346 12.394 ;
      RECT 25.894 12.358 25.946 12.394 ;
      RECT 25.494 12.358 25.546 12.394 ;
      RECT 25.094 12.358 25.146 12.394 ;
      RECT 24.694 12.358 24.746 12.394 ;
      RECT 24.294 12.358 24.346 12.394 ;
      RECT 23.894 12.358 23.946 12.394 ;
      RECT 23.494 12.358 23.546 12.394 ;
      RECT 23.094 12.358 23.146 12.394 ;
      RECT 21.814 12.358 21.868 12.394 ;
      RECT 19.838 12.358 19.886 12.394 ;
      RECT 19.53 12.358 19.578 12.394 ;
      RECT 16.882 12.358 16.936 12.394 ;
      RECT 16.422 12.358 16.47 12.394 ;
      RECT 16.114 12.358 16.162 12.394 ;
      RECT 14.132 12.358 14.186 12.394 ;
      RECT 13.294 12.358 13.346 12.394 ;
      RECT 12.894 12.358 12.946 12.394 ;
      RECT 12.494 12.358 12.546 12.394 ;
      RECT 12.094 12.358 12.146 12.394 ;
      RECT 11.694 12.358 11.746 12.394 ;
      RECT 11.294 12.358 11.346 12.394 ;
      RECT 10.894 12.358 10.946 12.394 ;
      RECT 10.494 12.358 10.546 12.394 ;
      RECT 10.094 12.358 10.146 12.394 ;
      RECT 9.694 12.358 9.746 12.394 ;
      RECT 9.294 12.358 9.346 12.394 ;
      RECT 8.894 12.358 8.946 12.394 ;
      RECT 8.494 12.358 8.546 12.394 ;
      RECT 8.094 12.358 8.146 12.394 ;
      RECT 7.694 12.358 7.746 12.394 ;
      RECT 7.294 12.358 7.346 12.394 ;
      RECT 6.894 12.358 6.946 12.394 ;
      RECT 6.494 12.358 6.546 12.394 ;
      RECT 6.094 12.358 6.146 12.394 ;
      RECT 5.694 12.358 5.746 12.394 ;
      RECT 5.294 12.358 5.346 12.394 ;
      RECT 4.894 12.358 4.946 12.394 ;
      RECT 4.494 12.358 4.546 12.394 ;
      RECT 4.094 12.358 4.146 12.394 ;
      RECT 3.694 12.358 3.746 12.394 ;
      RECT 3.294 12.358 3.346 12.394 ;
      RECT 2.894 12.358 2.946 12.394 ;
      RECT 2.494 12.358 2.546 12.394 ;
      RECT 2.094 12.358 2.146 12.394 ;
      RECT 1.694 12.358 1.746 12.394 ;
      RECT 1.294 12.358 1.346 12.394 ;
      RECT 0.894 12.358 0.946 12.394 ;
      RECT 21.414 12.282 21.468 12.318 ;
      RECT 14.532 12.282 14.586 12.318 ;
      RECT 19.606 12.129 19.654 12.165 ;
      RECT 18.08 12.129 18.12 12.165 ;
      RECT 16.718 12.129 16.772 12.165 ;
      RECT 16.346 12.129 16.394 12.165 ;
      RECT 20.37 12.1345 20.442 12.1595 ;
      RECT 18.764 12.1345 18.836 12.1595 ;
      RECT 15.558 12.1345 15.63 12.1595 ;
      RECT 21.978 11.982 22.022 12.018 ;
      RECT 13.978 11.982 14.022 12.018 ;
      RECT 18.764 11.9875 18.836 12.0125 ;
      RECT 19.762 11.835 19.81 11.871 ;
      RECT 17.616 11.835 17.656 11.871 ;
      RECT 16.19 11.835 16.238 11.871 ;
      RECT 35.254 11.606 35.306 11.642 ;
      RECT 34.854 11.606 34.906 11.642 ;
      RECT 34.454 11.606 34.506 11.642 ;
      RECT 34.054 11.606 34.106 11.642 ;
      RECT 33.654 11.606 33.706 11.642 ;
      RECT 33.254 11.606 33.306 11.642 ;
      RECT 32.854 11.606 32.906 11.642 ;
      RECT 32.454 11.606 32.506 11.642 ;
      RECT 32.054 11.606 32.106 11.642 ;
      RECT 31.654 11.606 31.706 11.642 ;
      RECT 31.254 11.606 31.306 11.642 ;
      RECT 30.854 11.606 30.906 11.642 ;
      RECT 30.454 11.606 30.506 11.642 ;
      RECT 30.054 11.606 30.106 11.642 ;
      RECT 29.654 11.606 29.706 11.642 ;
      RECT 29.254 11.606 29.306 11.642 ;
      RECT 28.854 11.606 28.906 11.642 ;
      RECT 28.454 11.606 28.506 11.642 ;
      RECT 28.054 11.606 28.106 11.642 ;
      RECT 27.654 11.606 27.706 11.642 ;
      RECT 27.254 11.606 27.306 11.642 ;
      RECT 26.854 11.606 26.906 11.642 ;
      RECT 26.454 11.606 26.506 11.642 ;
      RECT 26.054 11.606 26.106 11.642 ;
      RECT 25.654 11.606 25.706 11.642 ;
      RECT 25.254 11.606 25.306 11.642 ;
      RECT 24.854 11.606 24.906 11.642 ;
      RECT 24.454 11.606 24.506 11.642 ;
      RECT 24.054 11.606 24.106 11.642 ;
      RECT 23.654 11.606 23.706 11.642 ;
      RECT 23.254 11.606 23.306 11.642 ;
      RECT 22.854 11.606 22.906 11.642 ;
      RECT 22.694 11.606 22.746 11.642 ;
      RECT 21.732 11.606 21.786 11.642 ;
      RECT 14.214 11.606 14.268 11.642 ;
      RECT 13.054 11.606 13.106 11.642 ;
      RECT 12.654 11.606 12.706 11.642 ;
      RECT 12.254 11.606 12.306 11.642 ;
      RECT 11.854 11.606 11.906 11.642 ;
      RECT 11.454 11.606 11.506 11.642 ;
      RECT 11.054 11.606 11.106 11.642 ;
      RECT 10.654 11.606 10.706 11.642 ;
      RECT 10.254 11.606 10.306 11.642 ;
      RECT 9.854 11.606 9.906 11.642 ;
      RECT 9.454 11.606 9.506 11.642 ;
      RECT 9.054 11.606 9.106 11.642 ;
      RECT 8.654 11.606 8.706 11.642 ;
      RECT 8.254 11.606 8.306 11.642 ;
      RECT 7.854 11.606 7.906 11.642 ;
      RECT 7.454 11.606 7.506 11.642 ;
      RECT 7.054 11.606 7.106 11.642 ;
      RECT 6.654 11.606 6.706 11.642 ;
      RECT 6.254 11.606 6.306 11.642 ;
      RECT 5.854 11.606 5.906 11.642 ;
      RECT 5.454 11.606 5.506 11.642 ;
      RECT 5.054 11.606 5.106 11.642 ;
      RECT 4.654 11.606 4.706 11.642 ;
      RECT 4.254 11.606 4.306 11.642 ;
      RECT 3.854 11.606 3.906 11.642 ;
      RECT 3.454 11.606 3.506 11.642 ;
      RECT 3.054 11.606 3.106 11.642 ;
      RECT 2.654 11.606 2.706 11.642 ;
      RECT 2.254 11.606 2.306 11.642 ;
      RECT 1.854 11.606 1.906 11.642 ;
      RECT 1.454 11.606 1.506 11.642 ;
      RECT 1.054 11.606 1.106 11.642 ;
      RECT 0.654 11.606 0.706 11.642 ;
      RECT 21.978 11.382 22.022 11.418 ;
      RECT 21.096 11.382 21.14 11.418 ;
      RECT 14.86 11.382 14.904 11.418 ;
      RECT 13.978 11.382 14.022 11.418 ;
      RECT 35.494 11.158 35.546 11.194 ;
      RECT 35.094 11.158 35.146 11.194 ;
      RECT 34.694 11.158 34.746 11.194 ;
      RECT 34.294 11.158 34.346 11.194 ;
      RECT 33.894 11.158 33.946 11.194 ;
      RECT 33.494 11.158 33.546 11.194 ;
      RECT 33.094 11.158 33.146 11.194 ;
      RECT 32.694 11.158 32.746 11.194 ;
      RECT 32.294 11.158 32.346 11.194 ;
      RECT 31.894 11.158 31.946 11.194 ;
      RECT 31.494 11.158 31.546 11.194 ;
      RECT 31.094 11.158 31.146 11.194 ;
      RECT 30.694 11.158 30.746 11.194 ;
      RECT 30.294 11.158 30.346 11.194 ;
      RECT 29.894 11.158 29.946 11.194 ;
      RECT 29.494 11.158 29.546 11.194 ;
      RECT 29.094 11.158 29.146 11.194 ;
      RECT 28.694 11.158 28.746 11.194 ;
      RECT 28.294 11.158 28.346 11.194 ;
      RECT 27.894 11.158 27.946 11.194 ;
      RECT 27.494 11.158 27.546 11.194 ;
      RECT 27.094 11.158 27.146 11.194 ;
      RECT 26.694 11.158 26.746 11.194 ;
      RECT 26.294 11.158 26.346 11.194 ;
      RECT 25.894 11.158 25.946 11.194 ;
      RECT 25.494 11.158 25.546 11.194 ;
      RECT 25.094 11.158 25.146 11.194 ;
      RECT 24.694 11.158 24.746 11.194 ;
      RECT 24.294 11.158 24.346 11.194 ;
      RECT 23.894 11.158 23.946 11.194 ;
      RECT 23.494 11.158 23.546 11.194 ;
      RECT 23.094 11.158 23.146 11.194 ;
      RECT 21.814 11.158 21.868 11.194 ;
      RECT 19.838 11.158 19.886 11.194 ;
      RECT 19.53 11.158 19.578 11.194 ;
      RECT 16.882 11.158 16.936 11.194 ;
      RECT 16.422 11.158 16.47 11.194 ;
      RECT 16.114 11.158 16.162 11.194 ;
      RECT 14.132 11.158 14.186 11.194 ;
      RECT 13.294 11.158 13.346 11.194 ;
      RECT 12.894 11.158 12.946 11.194 ;
      RECT 12.494 11.158 12.546 11.194 ;
      RECT 12.094 11.158 12.146 11.194 ;
      RECT 11.694 11.158 11.746 11.194 ;
      RECT 11.294 11.158 11.346 11.194 ;
      RECT 10.894 11.158 10.946 11.194 ;
      RECT 10.494 11.158 10.546 11.194 ;
      RECT 10.094 11.158 10.146 11.194 ;
      RECT 9.694 11.158 9.746 11.194 ;
      RECT 9.294 11.158 9.346 11.194 ;
      RECT 8.894 11.158 8.946 11.194 ;
      RECT 8.494 11.158 8.546 11.194 ;
      RECT 8.094 11.158 8.146 11.194 ;
      RECT 7.694 11.158 7.746 11.194 ;
      RECT 7.294 11.158 7.346 11.194 ;
      RECT 6.894 11.158 6.946 11.194 ;
      RECT 6.494 11.158 6.546 11.194 ;
      RECT 6.094 11.158 6.146 11.194 ;
      RECT 5.694 11.158 5.746 11.194 ;
      RECT 5.294 11.158 5.346 11.194 ;
      RECT 4.894 11.158 4.946 11.194 ;
      RECT 4.494 11.158 4.546 11.194 ;
      RECT 4.094 11.158 4.146 11.194 ;
      RECT 3.694 11.158 3.746 11.194 ;
      RECT 3.294 11.158 3.346 11.194 ;
      RECT 2.894 11.158 2.946 11.194 ;
      RECT 2.494 11.158 2.546 11.194 ;
      RECT 2.094 11.158 2.146 11.194 ;
      RECT 1.694 11.158 1.746 11.194 ;
      RECT 1.294 11.158 1.346 11.194 ;
      RECT 0.894 11.158 0.946 11.194 ;
      RECT 21.414 11.082 21.468 11.118 ;
      RECT 14.532 11.082 14.586 11.118 ;
      RECT 19.606 10.929 19.654 10.965 ;
      RECT 18.08 10.929 18.12 10.965 ;
      RECT 16.718 10.929 16.772 10.965 ;
      RECT 16.346 10.929 16.394 10.965 ;
      RECT 20.37 10.9345 20.442 10.9595 ;
      RECT 18.764 10.9345 18.836 10.9595 ;
      RECT 15.558 10.9345 15.63 10.9595 ;
      RECT 21.978 10.782 22.022 10.818 ;
      RECT 13.978 10.782 14.022 10.818 ;
      RECT 18.764 10.7875 18.836 10.8125 ;
      RECT 19.762 10.635 19.81 10.671 ;
      RECT 17.616 10.635 17.656 10.671 ;
      RECT 16.19 10.635 16.238 10.671 ;
      RECT 35.254 10.406 35.306 10.442 ;
      RECT 34.854 10.406 34.906 10.442 ;
      RECT 34.454 10.406 34.506 10.442 ;
      RECT 34.054 10.406 34.106 10.442 ;
      RECT 33.654 10.406 33.706 10.442 ;
      RECT 33.254 10.406 33.306 10.442 ;
      RECT 32.854 10.406 32.906 10.442 ;
      RECT 32.454 10.406 32.506 10.442 ;
      RECT 32.054 10.406 32.106 10.442 ;
      RECT 31.654 10.406 31.706 10.442 ;
      RECT 31.254 10.406 31.306 10.442 ;
      RECT 30.854 10.406 30.906 10.442 ;
      RECT 30.454 10.406 30.506 10.442 ;
      RECT 30.054 10.406 30.106 10.442 ;
      RECT 29.654 10.406 29.706 10.442 ;
      RECT 29.254 10.406 29.306 10.442 ;
      RECT 28.854 10.406 28.906 10.442 ;
      RECT 28.454 10.406 28.506 10.442 ;
      RECT 28.054 10.406 28.106 10.442 ;
      RECT 27.654 10.406 27.706 10.442 ;
      RECT 27.254 10.406 27.306 10.442 ;
      RECT 26.854 10.406 26.906 10.442 ;
      RECT 26.454 10.406 26.506 10.442 ;
      RECT 26.054 10.406 26.106 10.442 ;
      RECT 25.654 10.406 25.706 10.442 ;
      RECT 25.254 10.406 25.306 10.442 ;
      RECT 24.854 10.406 24.906 10.442 ;
      RECT 24.454 10.406 24.506 10.442 ;
      RECT 24.054 10.406 24.106 10.442 ;
      RECT 23.654 10.406 23.706 10.442 ;
      RECT 23.254 10.406 23.306 10.442 ;
      RECT 22.854 10.406 22.906 10.442 ;
      RECT 22.694 10.406 22.746 10.442 ;
      RECT 21.732 10.406 21.786 10.442 ;
      RECT 14.214 10.406 14.268 10.442 ;
      RECT 13.054 10.406 13.106 10.442 ;
      RECT 12.654 10.406 12.706 10.442 ;
      RECT 12.254 10.406 12.306 10.442 ;
      RECT 11.854 10.406 11.906 10.442 ;
      RECT 11.454 10.406 11.506 10.442 ;
      RECT 11.054 10.406 11.106 10.442 ;
      RECT 10.654 10.406 10.706 10.442 ;
      RECT 10.254 10.406 10.306 10.442 ;
      RECT 9.854 10.406 9.906 10.442 ;
      RECT 9.454 10.406 9.506 10.442 ;
      RECT 9.054 10.406 9.106 10.442 ;
      RECT 8.654 10.406 8.706 10.442 ;
      RECT 8.254 10.406 8.306 10.442 ;
      RECT 7.854 10.406 7.906 10.442 ;
      RECT 7.454 10.406 7.506 10.442 ;
      RECT 7.054 10.406 7.106 10.442 ;
      RECT 6.654 10.406 6.706 10.442 ;
      RECT 6.254 10.406 6.306 10.442 ;
      RECT 5.854 10.406 5.906 10.442 ;
      RECT 5.454 10.406 5.506 10.442 ;
      RECT 5.054 10.406 5.106 10.442 ;
      RECT 4.654 10.406 4.706 10.442 ;
      RECT 4.254 10.406 4.306 10.442 ;
      RECT 3.854 10.406 3.906 10.442 ;
      RECT 3.454 10.406 3.506 10.442 ;
      RECT 3.054 10.406 3.106 10.442 ;
      RECT 2.654 10.406 2.706 10.442 ;
      RECT 2.254 10.406 2.306 10.442 ;
      RECT 1.854 10.406 1.906 10.442 ;
      RECT 1.454 10.406 1.506 10.442 ;
      RECT 1.054 10.406 1.106 10.442 ;
      RECT 0.654 10.406 0.706 10.442 ;
      RECT 21.978 10.182 22.022 10.218 ;
      RECT 21.096 10.182 21.14 10.218 ;
      RECT 14.86 10.182 14.904 10.218 ;
      RECT 13.978 10.182 14.022 10.218 ;
      RECT 35.494 9.958 35.546 9.994 ;
      RECT 35.094 9.958 35.146 9.994 ;
      RECT 34.694 9.958 34.746 9.994 ;
      RECT 34.294 9.958 34.346 9.994 ;
      RECT 33.894 9.958 33.946 9.994 ;
      RECT 33.494 9.958 33.546 9.994 ;
      RECT 33.094 9.958 33.146 9.994 ;
      RECT 32.694 9.958 32.746 9.994 ;
      RECT 32.294 9.958 32.346 9.994 ;
      RECT 31.894 9.958 31.946 9.994 ;
      RECT 31.494 9.958 31.546 9.994 ;
      RECT 31.094 9.958 31.146 9.994 ;
      RECT 30.694 9.958 30.746 9.994 ;
      RECT 30.294 9.958 30.346 9.994 ;
      RECT 29.894 9.958 29.946 9.994 ;
      RECT 29.494 9.958 29.546 9.994 ;
      RECT 29.094 9.958 29.146 9.994 ;
      RECT 28.694 9.958 28.746 9.994 ;
      RECT 28.294 9.958 28.346 9.994 ;
      RECT 27.894 9.958 27.946 9.994 ;
      RECT 27.494 9.958 27.546 9.994 ;
      RECT 27.094 9.958 27.146 9.994 ;
      RECT 26.694 9.958 26.746 9.994 ;
      RECT 26.294 9.958 26.346 9.994 ;
      RECT 25.894 9.958 25.946 9.994 ;
      RECT 25.494 9.958 25.546 9.994 ;
      RECT 25.094 9.958 25.146 9.994 ;
      RECT 24.694 9.958 24.746 9.994 ;
      RECT 24.294 9.958 24.346 9.994 ;
      RECT 23.894 9.958 23.946 9.994 ;
      RECT 23.494 9.958 23.546 9.994 ;
      RECT 23.094 9.958 23.146 9.994 ;
      RECT 21.814 9.958 21.868 9.994 ;
      RECT 19.838 9.958 19.886 9.994 ;
      RECT 19.53 9.958 19.578 9.994 ;
      RECT 16.882 9.958 16.936 9.994 ;
      RECT 16.422 9.958 16.47 9.994 ;
      RECT 16.114 9.958 16.162 9.994 ;
      RECT 14.132 9.958 14.186 9.994 ;
      RECT 13.294 9.958 13.346 9.994 ;
      RECT 12.894 9.958 12.946 9.994 ;
      RECT 12.494 9.958 12.546 9.994 ;
      RECT 12.094 9.958 12.146 9.994 ;
      RECT 11.694 9.958 11.746 9.994 ;
      RECT 11.294 9.958 11.346 9.994 ;
      RECT 10.894 9.958 10.946 9.994 ;
      RECT 10.494 9.958 10.546 9.994 ;
      RECT 10.094 9.958 10.146 9.994 ;
      RECT 9.694 9.958 9.746 9.994 ;
      RECT 9.294 9.958 9.346 9.994 ;
      RECT 8.894 9.958 8.946 9.994 ;
      RECT 8.494 9.958 8.546 9.994 ;
      RECT 8.094 9.958 8.146 9.994 ;
      RECT 7.694 9.958 7.746 9.994 ;
      RECT 7.294 9.958 7.346 9.994 ;
      RECT 6.894 9.958 6.946 9.994 ;
      RECT 6.494 9.958 6.546 9.994 ;
      RECT 6.094 9.958 6.146 9.994 ;
      RECT 5.694 9.958 5.746 9.994 ;
      RECT 5.294 9.958 5.346 9.994 ;
      RECT 4.894 9.958 4.946 9.994 ;
      RECT 4.494 9.958 4.546 9.994 ;
      RECT 4.094 9.958 4.146 9.994 ;
      RECT 3.694 9.958 3.746 9.994 ;
      RECT 3.294 9.958 3.346 9.994 ;
      RECT 2.894 9.958 2.946 9.994 ;
      RECT 2.494 9.958 2.546 9.994 ;
      RECT 2.094 9.958 2.146 9.994 ;
      RECT 1.694 9.958 1.746 9.994 ;
      RECT 1.294 9.958 1.346 9.994 ;
      RECT 0.894 9.958 0.946 9.994 ;
      RECT 21.414 9.882 21.468 9.918 ;
      RECT 14.532 9.882 14.586 9.918 ;
      RECT 19.606 9.729 19.654 9.765 ;
      RECT 18.08 9.729 18.12 9.765 ;
      RECT 16.718 9.729 16.772 9.765 ;
      RECT 16.346 9.729 16.394 9.765 ;
      RECT 20.37 9.7345 20.442 9.7595 ;
      RECT 18.764 9.7345 18.836 9.7595 ;
      RECT 15.558 9.7345 15.63 9.7595 ;
      RECT 21.978 9.582 22.022 9.618 ;
      RECT 13.978 9.582 14.022 9.618 ;
      RECT 18.764 9.5875 18.836 9.6125 ;
      RECT 19.762 9.435 19.81 9.471 ;
      RECT 17.616 9.435 17.656 9.471 ;
      RECT 16.19 9.435 16.238 9.471 ;
      RECT 35.254 9.206 35.306 9.242 ;
      RECT 34.854 9.206 34.906 9.242 ;
      RECT 34.454 9.206 34.506 9.242 ;
      RECT 34.054 9.206 34.106 9.242 ;
      RECT 33.654 9.206 33.706 9.242 ;
      RECT 33.254 9.206 33.306 9.242 ;
      RECT 32.854 9.206 32.906 9.242 ;
      RECT 32.454 9.206 32.506 9.242 ;
      RECT 32.054 9.206 32.106 9.242 ;
      RECT 31.654 9.206 31.706 9.242 ;
      RECT 31.254 9.206 31.306 9.242 ;
      RECT 30.854 9.206 30.906 9.242 ;
      RECT 30.454 9.206 30.506 9.242 ;
      RECT 30.054 9.206 30.106 9.242 ;
      RECT 29.654 9.206 29.706 9.242 ;
      RECT 29.254 9.206 29.306 9.242 ;
      RECT 28.854 9.206 28.906 9.242 ;
      RECT 28.454 9.206 28.506 9.242 ;
      RECT 28.054 9.206 28.106 9.242 ;
      RECT 27.654 9.206 27.706 9.242 ;
      RECT 27.254 9.206 27.306 9.242 ;
      RECT 26.854 9.206 26.906 9.242 ;
      RECT 26.454 9.206 26.506 9.242 ;
      RECT 26.054 9.206 26.106 9.242 ;
      RECT 25.654 9.206 25.706 9.242 ;
      RECT 25.254 9.206 25.306 9.242 ;
      RECT 24.854 9.206 24.906 9.242 ;
      RECT 24.454 9.206 24.506 9.242 ;
      RECT 24.054 9.206 24.106 9.242 ;
      RECT 23.654 9.206 23.706 9.242 ;
      RECT 23.254 9.206 23.306 9.242 ;
      RECT 22.854 9.206 22.906 9.242 ;
      RECT 22.694 9.206 22.746 9.242 ;
      RECT 21.732 9.206 21.786 9.242 ;
      RECT 14.214 9.206 14.268 9.242 ;
      RECT 13.054 9.206 13.106 9.242 ;
      RECT 12.654 9.206 12.706 9.242 ;
      RECT 12.254 9.206 12.306 9.242 ;
      RECT 11.854 9.206 11.906 9.242 ;
      RECT 11.454 9.206 11.506 9.242 ;
      RECT 11.054 9.206 11.106 9.242 ;
      RECT 10.654 9.206 10.706 9.242 ;
      RECT 10.254 9.206 10.306 9.242 ;
      RECT 9.854 9.206 9.906 9.242 ;
      RECT 9.454 9.206 9.506 9.242 ;
      RECT 9.054 9.206 9.106 9.242 ;
      RECT 8.654 9.206 8.706 9.242 ;
      RECT 8.254 9.206 8.306 9.242 ;
      RECT 7.854 9.206 7.906 9.242 ;
      RECT 7.454 9.206 7.506 9.242 ;
      RECT 7.054 9.206 7.106 9.242 ;
      RECT 6.654 9.206 6.706 9.242 ;
      RECT 6.254 9.206 6.306 9.242 ;
      RECT 5.854 9.206 5.906 9.242 ;
      RECT 5.454 9.206 5.506 9.242 ;
      RECT 5.054 9.206 5.106 9.242 ;
      RECT 4.654 9.206 4.706 9.242 ;
      RECT 4.254 9.206 4.306 9.242 ;
      RECT 3.854 9.206 3.906 9.242 ;
      RECT 3.454 9.206 3.506 9.242 ;
      RECT 3.054 9.206 3.106 9.242 ;
      RECT 2.654 9.206 2.706 9.242 ;
      RECT 2.254 9.206 2.306 9.242 ;
      RECT 1.854 9.206 1.906 9.242 ;
      RECT 1.454 9.206 1.506 9.242 ;
      RECT 1.054 9.206 1.106 9.242 ;
      RECT 0.654 9.206 0.706 9.242 ;
      RECT 21.978 8.982 22.022 9.018 ;
      RECT 21.096 8.982 21.14 9.018 ;
      RECT 14.86 8.982 14.904 9.018 ;
      RECT 13.978 8.982 14.022 9.018 ;
      RECT 35.494 8.758 35.546 8.794 ;
      RECT 35.094 8.758 35.146 8.794 ;
      RECT 34.694 8.758 34.746 8.794 ;
      RECT 34.294 8.758 34.346 8.794 ;
      RECT 33.894 8.758 33.946 8.794 ;
      RECT 33.494 8.758 33.546 8.794 ;
      RECT 33.094 8.758 33.146 8.794 ;
      RECT 32.694 8.758 32.746 8.794 ;
      RECT 32.294 8.758 32.346 8.794 ;
      RECT 31.894 8.758 31.946 8.794 ;
      RECT 31.494 8.758 31.546 8.794 ;
      RECT 31.094 8.758 31.146 8.794 ;
      RECT 30.694 8.758 30.746 8.794 ;
      RECT 30.294 8.758 30.346 8.794 ;
      RECT 29.894 8.758 29.946 8.794 ;
      RECT 29.494 8.758 29.546 8.794 ;
      RECT 29.094 8.758 29.146 8.794 ;
      RECT 28.694 8.758 28.746 8.794 ;
      RECT 28.294 8.758 28.346 8.794 ;
      RECT 27.894 8.758 27.946 8.794 ;
      RECT 27.494 8.758 27.546 8.794 ;
      RECT 27.094 8.758 27.146 8.794 ;
      RECT 26.694 8.758 26.746 8.794 ;
      RECT 26.294 8.758 26.346 8.794 ;
      RECT 25.894 8.758 25.946 8.794 ;
      RECT 25.494 8.758 25.546 8.794 ;
      RECT 25.094 8.758 25.146 8.794 ;
      RECT 24.694 8.758 24.746 8.794 ;
      RECT 24.294 8.758 24.346 8.794 ;
      RECT 23.894 8.758 23.946 8.794 ;
      RECT 23.494 8.758 23.546 8.794 ;
      RECT 23.094 8.758 23.146 8.794 ;
      RECT 21.814 8.758 21.868 8.794 ;
      RECT 19.838 8.758 19.886 8.794 ;
      RECT 19.53 8.758 19.578 8.794 ;
      RECT 16.882 8.758 16.936 8.794 ;
      RECT 16.422 8.758 16.47 8.794 ;
      RECT 16.114 8.758 16.162 8.794 ;
      RECT 14.132 8.758 14.186 8.794 ;
      RECT 13.294 8.758 13.346 8.794 ;
      RECT 12.894 8.758 12.946 8.794 ;
      RECT 12.494 8.758 12.546 8.794 ;
      RECT 12.094 8.758 12.146 8.794 ;
      RECT 11.694 8.758 11.746 8.794 ;
      RECT 11.294 8.758 11.346 8.794 ;
      RECT 10.894 8.758 10.946 8.794 ;
      RECT 10.494 8.758 10.546 8.794 ;
      RECT 10.094 8.758 10.146 8.794 ;
      RECT 9.694 8.758 9.746 8.794 ;
      RECT 9.294 8.758 9.346 8.794 ;
      RECT 8.894 8.758 8.946 8.794 ;
      RECT 8.494 8.758 8.546 8.794 ;
      RECT 8.094 8.758 8.146 8.794 ;
      RECT 7.694 8.758 7.746 8.794 ;
      RECT 7.294 8.758 7.346 8.794 ;
      RECT 6.894 8.758 6.946 8.794 ;
      RECT 6.494 8.758 6.546 8.794 ;
      RECT 6.094 8.758 6.146 8.794 ;
      RECT 5.694 8.758 5.746 8.794 ;
      RECT 5.294 8.758 5.346 8.794 ;
      RECT 4.894 8.758 4.946 8.794 ;
      RECT 4.494 8.758 4.546 8.794 ;
      RECT 4.094 8.758 4.146 8.794 ;
      RECT 3.694 8.758 3.746 8.794 ;
      RECT 3.294 8.758 3.346 8.794 ;
      RECT 2.894 8.758 2.946 8.794 ;
      RECT 2.494 8.758 2.546 8.794 ;
      RECT 2.094 8.758 2.146 8.794 ;
      RECT 1.694 8.758 1.746 8.794 ;
      RECT 1.294 8.758 1.346 8.794 ;
      RECT 0.894 8.758 0.946 8.794 ;
      RECT 21.414 8.682 21.468 8.718 ;
      RECT 14.532 8.682 14.586 8.718 ;
      RECT 19.606 8.529 19.654 8.565 ;
      RECT 18.08 8.529 18.12 8.565 ;
      RECT 16.718 8.529 16.772 8.565 ;
      RECT 16.346 8.529 16.394 8.565 ;
      RECT 20.37 8.5345 20.442 8.5595 ;
      RECT 18.764 8.5345 18.836 8.5595 ;
      RECT 15.558 8.5345 15.63 8.5595 ;
      RECT 21.978 8.382 22.022 8.418 ;
      RECT 13.978 8.382 14.022 8.418 ;
      RECT 18.764 8.3875 18.836 8.4125 ;
      RECT 19.762 8.235 19.81 8.271 ;
      RECT 17.616 8.235 17.656 8.271 ;
      RECT 16.19 8.235 16.238 8.271 ;
      RECT 35.254 8.006 35.306 8.042 ;
      RECT 34.854 8.006 34.906 8.042 ;
      RECT 34.454 8.006 34.506 8.042 ;
      RECT 34.054 8.006 34.106 8.042 ;
      RECT 33.654 8.006 33.706 8.042 ;
      RECT 33.254 8.006 33.306 8.042 ;
      RECT 32.854 8.006 32.906 8.042 ;
      RECT 32.454 8.006 32.506 8.042 ;
      RECT 32.054 8.006 32.106 8.042 ;
      RECT 31.654 8.006 31.706 8.042 ;
      RECT 31.254 8.006 31.306 8.042 ;
      RECT 30.854 8.006 30.906 8.042 ;
      RECT 30.454 8.006 30.506 8.042 ;
      RECT 30.054 8.006 30.106 8.042 ;
      RECT 29.654 8.006 29.706 8.042 ;
      RECT 29.254 8.006 29.306 8.042 ;
      RECT 28.854 8.006 28.906 8.042 ;
      RECT 28.454 8.006 28.506 8.042 ;
      RECT 28.054 8.006 28.106 8.042 ;
      RECT 27.654 8.006 27.706 8.042 ;
      RECT 27.254 8.006 27.306 8.042 ;
      RECT 26.854 8.006 26.906 8.042 ;
      RECT 26.454 8.006 26.506 8.042 ;
      RECT 26.054 8.006 26.106 8.042 ;
      RECT 25.654 8.006 25.706 8.042 ;
      RECT 25.254 8.006 25.306 8.042 ;
      RECT 24.854 8.006 24.906 8.042 ;
      RECT 24.454 8.006 24.506 8.042 ;
      RECT 24.054 8.006 24.106 8.042 ;
      RECT 23.654 8.006 23.706 8.042 ;
      RECT 23.254 8.006 23.306 8.042 ;
      RECT 22.854 8.006 22.906 8.042 ;
      RECT 22.694 8.006 22.746 8.042 ;
      RECT 21.732 8.006 21.786 8.042 ;
      RECT 14.214 8.006 14.268 8.042 ;
      RECT 13.054 8.006 13.106 8.042 ;
      RECT 12.654 8.006 12.706 8.042 ;
      RECT 12.254 8.006 12.306 8.042 ;
      RECT 11.854 8.006 11.906 8.042 ;
      RECT 11.454 8.006 11.506 8.042 ;
      RECT 11.054 8.006 11.106 8.042 ;
      RECT 10.654 8.006 10.706 8.042 ;
      RECT 10.254 8.006 10.306 8.042 ;
      RECT 9.854 8.006 9.906 8.042 ;
      RECT 9.454 8.006 9.506 8.042 ;
      RECT 9.054 8.006 9.106 8.042 ;
      RECT 8.654 8.006 8.706 8.042 ;
      RECT 8.254 8.006 8.306 8.042 ;
      RECT 7.854 8.006 7.906 8.042 ;
      RECT 7.454 8.006 7.506 8.042 ;
      RECT 7.054 8.006 7.106 8.042 ;
      RECT 6.654 8.006 6.706 8.042 ;
      RECT 6.254 8.006 6.306 8.042 ;
      RECT 5.854 8.006 5.906 8.042 ;
      RECT 5.454 8.006 5.506 8.042 ;
      RECT 5.054 8.006 5.106 8.042 ;
      RECT 4.654 8.006 4.706 8.042 ;
      RECT 4.254 8.006 4.306 8.042 ;
      RECT 3.854 8.006 3.906 8.042 ;
      RECT 3.454 8.006 3.506 8.042 ;
      RECT 3.054 8.006 3.106 8.042 ;
      RECT 2.654 8.006 2.706 8.042 ;
      RECT 2.254 8.006 2.306 8.042 ;
      RECT 1.854 8.006 1.906 8.042 ;
      RECT 1.454 8.006 1.506 8.042 ;
      RECT 1.054 8.006 1.106 8.042 ;
      RECT 0.654 8.006 0.706 8.042 ;
      RECT 21.978 7.782 22.022 7.818 ;
      RECT 21.096 7.782 21.14 7.818 ;
      RECT 14.86 7.782 14.904 7.818 ;
      RECT 13.978 7.782 14.022 7.818 ;
      RECT 35.494 7.558 35.546 7.594 ;
      RECT 35.094 7.558 35.146 7.594 ;
      RECT 34.694 7.558 34.746 7.594 ;
      RECT 34.294 7.558 34.346 7.594 ;
      RECT 33.894 7.558 33.946 7.594 ;
      RECT 33.494 7.558 33.546 7.594 ;
      RECT 33.094 7.558 33.146 7.594 ;
      RECT 32.694 7.558 32.746 7.594 ;
      RECT 32.294 7.558 32.346 7.594 ;
      RECT 31.894 7.558 31.946 7.594 ;
      RECT 31.494 7.558 31.546 7.594 ;
      RECT 31.094 7.558 31.146 7.594 ;
      RECT 30.694 7.558 30.746 7.594 ;
      RECT 30.294 7.558 30.346 7.594 ;
      RECT 29.894 7.558 29.946 7.594 ;
      RECT 29.494 7.558 29.546 7.594 ;
      RECT 29.094 7.558 29.146 7.594 ;
      RECT 28.694 7.558 28.746 7.594 ;
      RECT 28.294 7.558 28.346 7.594 ;
      RECT 27.894 7.558 27.946 7.594 ;
      RECT 27.494 7.558 27.546 7.594 ;
      RECT 27.094 7.558 27.146 7.594 ;
      RECT 26.694 7.558 26.746 7.594 ;
      RECT 26.294 7.558 26.346 7.594 ;
      RECT 25.894 7.558 25.946 7.594 ;
      RECT 25.494 7.558 25.546 7.594 ;
      RECT 25.094 7.558 25.146 7.594 ;
      RECT 24.694 7.558 24.746 7.594 ;
      RECT 24.294 7.558 24.346 7.594 ;
      RECT 23.894 7.558 23.946 7.594 ;
      RECT 23.494 7.558 23.546 7.594 ;
      RECT 23.094 7.558 23.146 7.594 ;
      RECT 21.814 7.558 21.868 7.594 ;
      RECT 19.838 7.558 19.886 7.594 ;
      RECT 19.53 7.558 19.578 7.594 ;
      RECT 16.882 7.558 16.936 7.594 ;
      RECT 16.422 7.558 16.47 7.594 ;
      RECT 16.114 7.558 16.162 7.594 ;
      RECT 14.132 7.558 14.186 7.594 ;
      RECT 13.294 7.558 13.346 7.594 ;
      RECT 12.894 7.558 12.946 7.594 ;
      RECT 12.494 7.558 12.546 7.594 ;
      RECT 12.094 7.558 12.146 7.594 ;
      RECT 11.694 7.558 11.746 7.594 ;
      RECT 11.294 7.558 11.346 7.594 ;
      RECT 10.894 7.558 10.946 7.594 ;
      RECT 10.494 7.558 10.546 7.594 ;
      RECT 10.094 7.558 10.146 7.594 ;
      RECT 9.694 7.558 9.746 7.594 ;
      RECT 9.294 7.558 9.346 7.594 ;
      RECT 8.894 7.558 8.946 7.594 ;
      RECT 8.494 7.558 8.546 7.594 ;
      RECT 8.094 7.558 8.146 7.594 ;
      RECT 7.694 7.558 7.746 7.594 ;
      RECT 7.294 7.558 7.346 7.594 ;
      RECT 6.894 7.558 6.946 7.594 ;
      RECT 6.494 7.558 6.546 7.594 ;
      RECT 6.094 7.558 6.146 7.594 ;
      RECT 5.694 7.558 5.746 7.594 ;
      RECT 5.294 7.558 5.346 7.594 ;
      RECT 4.894 7.558 4.946 7.594 ;
      RECT 4.494 7.558 4.546 7.594 ;
      RECT 4.094 7.558 4.146 7.594 ;
      RECT 3.694 7.558 3.746 7.594 ;
      RECT 3.294 7.558 3.346 7.594 ;
      RECT 2.894 7.558 2.946 7.594 ;
      RECT 2.494 7.558 2.546 7.594 ;
      RECT 2.094 7.558 2.146 7.594 ;
      RECT 1.694 7.558 1.746 7.594 ;
      RECT 1.294 7.558 1.346 7.594 ;
      RECT 0.894 7.558 0.946 7.594 ;
      RECT 21.414 7.482 21.468 7.518 ;
      RECT 14.532 7.482 14.586 7.518 ;
      RECT 19.606 7.329 19.654 7.365 ;
      RECT 18.08 7.329 18.12 7.365 ;
      RECT 16.718 7.329 16.772 7.365 ;
      RECT 16.346 7.329 16.394 7.365 ;
      RECT 20.37 7.3345 20.442 7.3595 ;
      RECT 18.764 7.3345 18.836 7.3595 ;
      RECT 15.558 7.3345 15.63 7.3595 ;
      RECT 21.978 7.182 22.022 7.218 ;
      RECT 13.978 7.182 14.022 7.218 ;
      RECT 18.764 7.1875 18.836 7.2125 ;
      RECT 19.762 7.035 19.81 7.071 ;
      RECT 17.616 7.035 17.656 7.071 ;
      RECT 16.19 7.035 16.238 7.071 ;
      RECT 35.254 6.806 35.306 6.842 ;
      RECT 34.854 6.806 34.906 6.842 ;
      RECT 34.454 6.806 34.506 6.842 ;
      RECT 34.054 6.806 34.106 6.842 ;
      RECT 33.654 6.806 33.706 6.842 ;
      RECT 33.254 6.806 33.306 6.842 ;
      RECT 32.854 6.806 32.906 6.842 ;
      RECT 32.454 6.806 32.506 6.842 ;
      RECT 32.054 6.806 32.106 6.842 ;
      RECT 31.654 6.806 31.706 6.842 ;
      RECT 31.254 6.806 31.306 6.842 ;
      RECT 30.854 6.806 30.906 6.842 ;
      RECT 30.454 6.806 30.506 6.842 ;
      RECT 30.054 6.806 30.106 6.842 ;
      RECT 29.654 6.806 29.706 6.842 ;
      RECT 29.254 6.806 29.306 6.842 ;
      RECT 28.854 6.806 28.906 6.842 ;
      RECT 28.454 6.806 28.506 6.842 ;
      RECT 28.054 6.806 28.106 6.842 ;
      RECT 27.654 6.806 27.706 6.842 ;
      RECT 27.254 6.806 27.306 6.842 ;
      RECT 26.854 6.806 26.906 6.842 ;
      RECT 26.454 6.806 26.506 6.842 ;
      RECT 26.054 6.806 26.106 6.842 ;
      RECT 25.654 6.806 25.706 6.842 ;
      RECT 25.254 6.806 25.306 6.842 ;
      RECT 24.854 6.806 24.906 6.842 ;
      RECT 24.454 6.806 24.506 6.842 ;
      RECT 24.054 6.806 24.106 6.842 ;
      RECT 23.654 6.806 23.706 6.842 ;
      RECT 23.254 6.806 23.306 6.842 ;
      RECT 22.854 6.806 22.906 6.842 ;
      RECT 22.694 6.806 22.746 6.842 ;
      RECT 21.732 6.806 21.786 6.842 ;
      RECT 14.214 6.806 14.268 6.842 ;
      RECT 13.054 6.806 13.106 6.842 ;
      RECT 12.654 6.806 12.706 6.842 ;
      RECT 12.254 6.806 12.306 6.842 ;
      RECT 11.854 6.806 11.906 6.842 ;
      RECT 11.454 6.806 11.506 6.842 ;
      RECT 11.054 6.806 11.106 6.842 ;
      RECT 10.654 6.806 10.706 6.842 ;
      RECT 10.254 6.806 10.306 6.842 ;
      RECT 9.854 6.806 9.906 6.842 ;
      RECT 9.454 6.806 9.506 6.842 ;
      RECT 9.054 6.806 9.106 6.842 ;
      RECT 8.654 6.806 8.706 6.842 ;
      RECT 8.254 6.806 8.306 6.842 ;
      RECT 7.854 6.806 7.906 6.842 ;
      RECT 7.454 6.806 7.506 6.842 ;
      RECT 7.054 6.806 7.106 6.842 ;
      RECT 6.654 6.806 6.706 6.842 ;
      RECT 6.254 6.806 6.306 6.842 ;
      RECT 5.854 6.806 5.906 6.842 ;
      RECT 5.454 6.806 5.506 6.842 ;
      RECT 5.054 6.806 5.106 6.842 ;
      RECT 4.654 6.806 4.706 6.842 ;
      RECT 4.254 6.806 4.306 6.842 ;
      RECT 3.854 6.806 3.906 6.842 ;
      RECT 3.454 6.806 3.506 6.842 ;
      RECT 3.054 6.806 3.106 6.842 ;
      RECT 2.654 6.806 2.706 6.842 ;
      RECT 2.254 6.806 2.306 6.842 ;
      RECT 1.854 6.806 1.906 6.842 ;
      RECT 1.454 6.806 1.506 6.842 ;
      RECT 1.054 6.806 1.106 6.842 ;
      RECT 0.654 6.806 0.706 6.842 ;
      RECT 21.978 6.582 22.022 6.618 ;
      RECT 21.096 6.582 21.14 6.618 ;
      RECT 14.86 6.582 14.904 6.618 ;
      RECT 13.978 6.582 14.022 6.618 ;
      RECT 35.494 6.358 35.546 6.394 ;
      RECT 35.094 6.358 35.146 6.394 ;
      RECT 34.694 6.358 34.746 6.394 ;
      RECT 34.294 6.358 34.346 6.394 ;
      RECT 33.894 6.358 33.946 6.394 ;
      RECT 33.494 6.358 33.546 6.394 ;
      RECT 33.094 6.358 33.146 6.394 ;
      RECT 32.694 6.358 32.746 6.394 ;
      RECT 32.294 6.358 32.346 6.394 ;
      RECT 31.894 6.358 31.946 6.394 ;
      RECT 31.494 6.358 31.546 6.394 ;
      RECT 31.094 6.358 31.146 6.394 ;
      RECT 30.694 6.358 30.746 6.394 ;
      RECT 30.294 6.358 30.346 6.394 ;
      RECT 29.894 6.358 29.946 6.394 ;
      RECT 29.494 6.358 29.546 6.394 ;
      RECT 29.094 6.358 29.146 6.394 ;
      RECT 28.694 6.358 28.746 6.394 ;
      RECT 28.294 6.358 28.346 6.394 ;
      RECT 27.894 6.358 27.946 6.394 ;
      RECT 27.494 6.358 27.546 6.394 ;
      RECT 27.094 6.358 27.146 6.394 ;
      RECT 26.694 6.358 26.746 6.394 ;
      RECT 26.294 6.358 26.346 6.394 ;
      RECT 25.894 6.358 25.946 6.394 ;
      RECT 25.494 6.358 25.546 6.394 ;
      RECT 25.094 6.358 25.146 6.394 ;
      RECT 24.694 6.358 24.746 6.394 ;
      RECT 24.294 6.358 24.346 6.394 ;
      RECT 23.894 6.358 23.946 6.394 ;
      RECT 23.494 6.358 23.546 6.394 ;
      RECT 23.094 6.358 23.146 6.394 ;
      RECT 21.814 6.358 21.868 6.394 ;
      RECT 19.838 6.358 19.886 6.394 ;
      RECT 19.53 6.358 19.578 6.394 ;
      RECT 16.882 6.358 16.936 6.394 ;
      RECT 16.422 6.358 16.47 6.394 ;
      RECT 16.114 6.358 16.162 6.394 ;
      RECT 14.132 6.358 14.186 6.394 ;
      RECT 13.294 6.358 13.346 6.394 ;
      RECT 12.894 6.358 12.946 6.394 ;
      RECT 12.494 6.358 12.546 6.394 ;
      RECT 12.094 6.358 12.146 6.394 ;
      RECT 11.694 6.358 11.746 6.394 ;
      RECT 11.294 6.358 11.346 6.394 ;
      RECT 10.894 6.358 10.946 6.394 ;
      RECT 10.494 6.358 10.546 6.394 ;
      RECT 10.094 6.358 10.146 6.394 ;
      RECT 9.694 6.358 9.746 6.394 ;
      RECT 9.294 6.358 9.346 6.394 ;
      RECT 8.894 6.358 8.946 6.394 ;
      RECT 8.494 6.358 8.546 6.394 ;
      RECT 8.094 6.358 8.146 6.394 ;
      RECT 7.694 6.358 7.746 6.394 ;
      RECT 7.294 6.358 7.346 6.394 ;
      RECT 6.894 6.358 6.946 6.394 ;
      RECT 6.494 6.358 6.546 6.394 ;
      RECT 6.094 6.358 6.146 6.394 ;
      RECT 5.694 6.358 5.746 6.394 ;
      RECT 5.294 6.358 5.346 6.394 ;
      RECT 4.894 6.358 4.946 6.394 ;
      RECT 4.494 6.358 4.546 6.394 ;
      RECT 4.094 6.358 4.146 6.394 ;
      RECT 3.694 6.358 3.746 6.394 ;
      RECT 3.294 6.358 3.346 6.394 ;
      RECT 2.894 6.358 2.946 6.394 ;
      RECT 2.494 6.358 2.546 6.394 ;
      RECT 2.094 6.358 2.146 6.394 ;
      RECT 1.694 6.358 1.746 6.394 ;
      RECT 1.294 6.358 1.346 6.394 ;
      RECT 0.894 6.358 0.946 6.394 ;
      RECT 21.414 6.282 21.468 6.318 ;
      RECT 14.532 6.282 14.586 6.318 ;
      RECT 19.606 6.129 19.654 6.165 ;
      RECT 18.08 6.129 18.12 6.165 ;
      RECT 16.718 6.129 16.772 6.165 ;
      RECT 16.346 6.129 16.394 6.165 ;
      RECT 20.37 6.1345 20.442 6.1595 ;
      RECT 18.764 6.1345 18.836 6.1595 ;
      RECT 15.558 6.1345 15.63 6.1595 ;
      RECT 21.978 5.982 22.022 6.018 ;
      RECT 13.978 5.982 14.022 6.018 ;
      RECT 18.764 5.9875 18.836 6.0125 ;
      RECT 19.762 5.835 19.81 5.871 ;
      RECT 17.616 5.835 17.656 5.871 ;
      RECT 16.19 5.835 16.238 5.871 ;
      RECT 35.254 5.606 35.306 5.642 ;
      RECT 34.854 5.606 34.906 5.642 ;
      RECT 34.454 5.606 34.506 5.642 ;
      RECT 34.054 5.606 34.106 5.642 ;
      RECT 33.654 5.606 33.706 5.642 ;
      RECT 33.254 5.606 33.306 5.642 ;
      RECT 32.854 5.606 32.906 5.642 ;
      RECT 32.454 5.606 32.506 5.642 ;
      RECT 32.054 5.606 32.106 5.642 ;
      RECT 31.654 5.606 31.706 5.642 ;
      RECT 31.254 5.606 31.306 5.642 ;
      RECT 30.854 5.606 30.906 5.642 ;
      RECT 30.454 5.606 30.506 5.642 ;
      RECT 30.054 5.606 30.106 5.642 ;
      RECT 29.654 5.606 29.706 5.642 ;
      RECT 29.254 5.606 29.306 5.642 ;
      RECT 28.854 5.606 28.906 5.642 ;
      RECT 28.454 5.606 28.506 5.642 ;
      RECT 28.054 5.606 28.106 5.642 ;
      RECT 27.654 5.606 27.706 5.642 ;
      RECT 27.254 5.606 27.306 5.642 ;
      RECT 26.854 5.606 26.906 5.642 ;
      RECT 26.454 5.606 26.506 5.642 ;
      RECT 26.054 5.606 26.106 5.642 ;
      RECT 25.654 5.606 25.706 5.642 ;
      RECT 25.254 5.606 25.306 5.642 ;
      RECT 24.854 5.606 24.906 5.642 ;
      RECT 24.454 5.606 24.506 5.642 ;
      RECT 24.054 5.606 24.106 5.642 ;
      RECT 23.654 5.606 23.706 5.642 ;
      RECT 23.254 5.606 23.306 5.642 ;
      RECT 22.854 5.606 22.906 5.642 ;
      RECT 22.694 5.606 22.746 5.642 ;
      RECT 21.732 5.606 21.786 5.642 ;
      RECT 14.214 5.606 14.268 5.642 ;
      RECT 13.054 5.606 13.106 5.642 ;
      RECT 12.654 5.606 12.706 5.642 ;
      RECT 12.254 5.606 12.306 5.642 ;
      RECT 11.854 5.606 11.906 5.642 ;
      RECT 11.454 5.606 11.506 5.642 ;
      RECT 11.054 5.606 11.106 5.642 ;
      RECT 10.654 5.606 10.706 5.642 ;
      RECT 10.254 5.606 10.306 5.642 ;
      RECT 9.854 5.606 9.906 5.642 ;
      RECT 9.454 5.606 9.506 5.642 ;
      RECT 9.054 5.606 9.106 5.642 ;
      RECT 8.654 5.606 8.706 5.642 ;
      RECT 8.254 5.606 8.306 5.642 ;
      RECT 7.854 5.606 7.906 5.642 ;
      RECT 7.454 5.606 7.506 5.642 ;
      RECT 7.054 5.606 7.106 5.642 ;
      RECT 6.654 5.606 6.706 5.642 ;
      RECT 6.254 5.606 6.306 5.642 ;
      RECT 5.854 5.606 5.906 5.642 ;
      RECT 5.454 5.606 5.506 5.642 ;
      RECT 5.054 5.606 5.106 5.642 ;
      RECT 4.654 5.606 4.706 5.642 ;
      RECT 4.254 5.606 4.306 5.642 ;
      RECT 3.854 5.606 3.906 5.642 ;
      RECT 3.454 5.606 3.506 5.642 ;
      RECT 3.054 5.606 3.106 5.642 ;
      RECT 2.654 5.606 2.706 5.642 ;
      RECT 2.254 5.606 2.306 5.642 ;
      RECT 1.854 5.606 1.906 5.642 ;
      RECT 1.454 5.606 1.506 5.642 ;
      RECT 1.054 5.606 1.106 5.642 ;
      RECT 0.654 5.606 0.706 5.642 ;
      RECT 21.978 5.382 22.022 5.418 ;
      RECT 21.096 5.382 21.14 5.418 ;
      RECT 14.86 5.382 14.904 5.418 ;
      RECT 13.978 5.382 14.022 5.418 ;
      RECT 35.494 5.158 35.546 5.194 ;
      RECT 35.094 5.158 35.146 5.194 ;
      RECT 34.694 5.158 34.746 5.194 ;
      RECT 34.294 5.158 34.346 5.194 ;
      RECT 33.894 5.158 33.946 5.194 ;
      RECT 33.494 5.158 33.546 5.194 ;
      RECT 33.094 5.158 33.146 5.194 ;
      RECT 32.694 5.158 32.746 5.194 ;
      RECT 32.294 5.158 32.346 5.194 ;
      RECT 31.894 5.158 31.946 5.194 ;
      RECT 31.494 5.158 31.546 5.194 ;
      RECT 31.094 5.158 31.146 5.194 ;
      RECT 30.694 5.158 30.746 5.194 ;
      RECT 30.294 5.158 30.346 5.194 ;
      RECT 29.894 5.158 29.946 5.194 ;
      RECT 29.494 5.158 29.546 5.194 ;
      RECT 29.094 5.158 29.146 5.194 ;
      RECT 28.694 5.158 28.746 5.194 ;
      RECT 28.294 5.158 28.346 5.194 ;
      RECT 27.894 5.158 27.946 5.194 ;
      RECT 27.494 5.158 27.546 5.194 ;
      RECT 27.094 5.158 27.146 5.194 ;
      RECT 26.694 5.158 26.746 5.194 ;
      RECT 26.294 5.158 26.346 5.194 ;
      RECT 25.894 5.158 25.946 5.194 ;
      RECT 25.494 5.158 25.546 5.194 ;
      RECT 25.094 5.158 25.146 5.194 ;
      RECT 24.694 5.158 24.746 5.194 ;
      RECT 24.294 5.158 24.346 5.194 ;
      RECT 23.894 5.158 23.946 5.194 ;
      RECT 23.494 5.158 23.546 5.194 ;
      RECT 23.094 5.158 23.146 5.194 ;
      RECT 21.814 5.158 21.868 5.194 ;
      RECT 19.838 5.158 19.886 5.194 ;
      RECT 19.53 5.158 19.578 5.194 ;
      RECT 16.882 5.158 16.936 5.194 ;
      RECT 16.422 5.158 16.47 5.194 ;
      RECT 16.114 5.158 16.162 5.194 ;
      RECT 14.132 5.158 14.186 5.194 ;
      RECT 13.294 5.158 13.346 5.194 ;
      RECT 12.894 5.158 12.946 5.194 ;
      RECT 12.494 5.158 12.546 5.194 ;
      RECT 12.094 5.158 12.146 5.194 ;
      RECT 11.694 5.158 11.746 5.194 ;
      RECT 11.294 5.158 11.346 5.194 ;
      RECT 10.894 5.158 10.946 5.194 ;
      RECT 10.494 5.158 10.546 5.194 ;
      RECT 10.094 5.158 10.146 5.194 ;
      RECT 9.694 5.158 9.746 5.194 ;
      RECT 9.294 5.158 9.346 5.194 ;
      RECT 8.894 5.158 8.946 5.194 ;
      RECT 8.494 5.158 8.546 5.194 ;
      RECT 8.094 5.158 8.146 5.194 ;
      RECT 7.694 5.158 7.746 5.194 ;
      RECT 7.294 5.158 7.346 5.194 ;
      RECT 6.894 5.158 6.946 5.194 ;
      RECT 6.494 5.158 6.546 5.194 ;
      RECT 6.094 5.158 6.146 5.194 ;
      RECT 5.694 5.158 5.746 5.194 ;
      RECT 5.294 5.158 5.346 5.194 ;
      RECT 4.894 5.158 4.946 5.194 ;
      RECT 4.494 5.158 4.546 5.194 ;
      RECT 4.094 5.158 4.146 5.194 ;
      RECT 3.694 5.158 3.746 5.194 ;
      RECT 3.294 5.158 3.346 5.194 ;
      RECT 2.894 5.158 2.946 5.194 ;
      RECT 2.494 5.158 2.546 5.194 ;
      RECT 2.094 5.158 2.146 5.194 ;
      RECT 1.694 5.158 1.746 5.194 ;
      RECT 1.294 5.158 1.346 5.194 ;
      RECT 0.894 5.158 0.946 5.194 ;
      RECT 21.414 5.082 21.468 5.118 ;
      RECT 14.532 5.082 14.586 5.118 ;
      RECT 19.606 4.929 19.654 4.965 ;
      RECT 18.08 4.929 18.12 4.965 ;
      RECT 16.718 4.929 16.772 4.965 ;
      RECT 16.346 4.929 16.394 4.965 ;
      RECT 20.37 4.9345 20.442 4.9595 ;
      RECT 18.764 4.9345 18.836 4.9595 ;
      RECT 15.558 4.9345 15.63 4.9595 ;
      RECT 21.978 4.782 22.022 4.818 ;
      RECT 13.978 4.782 14.022 4.818 ;
      RECT 18.764 4.7875 18.836 4.8125 ;
      RECT 19.762 4.635 19.81 4.671 ;
      RECT 17.616 4.635 17.656 4.671 ;
      RECT 16.19 4.635 16.238 4.671 ;
      RECT 35.254 4.406 35.306 4.442 ;
      RECT 34.854 4.406 34.906 4.442 ;
      RECT 34.454 4.406 34.506 4.442 ;
      RECT 34.054 4.406 34.106 4.442 ;
      RECT 33.654 4.406 33.706 4.442 ;
      RECT 33.254 4.406 33.306 4.442 ;
      RECT 32.854 4.406 32.906 4.442 ;
      RECT 32.454 4.406 32.506 4.442 ;
      RECT 32.054 4.406 32.106 4.442 ;
      RECT 31.654 4.406 31.706 4.442 ;
      RECT 31.254 4.406 31.306 4.442 ;
      RECT 30.854 4.406 30.906 4.442 ;
      RECT 30.454 4.406 30.506 4.442 ;
      RECT 30.054 4.406 30.106 4.442 ;
      RECT 29.654 4.406 29.706 4.442 ;
      RECT 29.254 4.406 29.306 4.442 ;
      RECT 28.854 4.406 28.906 4.442 ;
      RECT 28.454 4.406 28.506 4.442 ;
      RECT 28.054 4.406 28.106 4.442 ;
      RECT 27.654 4.406 27.706 4.442 ;
      RECT 27.254 4.406 27.306 4.442 ;
      RECT 26.854 4.406 26.906 4.442 ;
      RECT 26.454 4.406 26.506 4.442 ;
      RECT 26.054 4.406 26.106 4.442 ;
      RECT 25.654 4.406 25.706 4.442 ;
      RECT 25.254 4.406 25.306 4.442 ;
      RECT 24.854 4.406 24.906 4.442 ;
      RECT 24.454 4.406 24.506 4.442 ;
      RECT 24.054 4.406 24.106 4.442 ;
      RECT 23.654 4.406 23.706 4.442 ;
      RECT 23.254 4.406 23.306 4.442 ;
      RECT 22.854 4.406 22.906 4.442 ;
      RECT 22.694 4.406 22.746 4.442 ;
      RECT 21.732 4.406 21.786 4.442 ;
      RECT 14.214 4.406 14.268 4.442 ;
      RECT 13.054 4.406 13.106 4.442 ;
      RECT 12.654 4.406 12.706 4.442 ;
      RECT 12.254 4.406 12.306 4.442 ;
      RECT 11.854 4.406 11.906 4.442 ;
      RECT 11.454 4.406 11.506 4.442 ;
      RECT 11.054 4.406 11.106 4.442 ;
      RECT 10.654 4.406 10.706 4.442 ;
      RECT 10.254 4.406 10.306 4.442 ;
      RECT 9.854 4.406 9.906 4.442 ;
      RECT 9.454 4.406 9.506 4.442 ;
      RECT 9.054 4.406 9.106 4.442 ;
      RECT 8.654 4.406 8.706 4.442 ;
      RECT 8.254 4.406 8.306 4.442 ;
      RECT 7.854 4.406 7.906 4.442 ;
      RECT 7.454 4.406 7.506 4.442 ;
      RECT 7.054 4.406 7.106 4.442 ;
      RECT 6.654 4.406 6.706 4.442 ;
      RECT 6.254 4.406 6.306 4.442 ;
      RECT 5.854 4.406 5.906 4.442 ;
      RECT 5.454 4.406 5.506 4.442 ;
      RECT 5.054 4.406 5.106 4.442 ;
      RECT 4.654 4.406 4.706 4.442 ;
      RECT 4.254 4.406 4.306 4.442 ;
      RECT 3.854 4.406 3.906 4.442 ;
      RECT 3.454 4.406 3.506 4.442 ;
      RECT 3.054 4.406 3.106 4.442 ;
      RECT 2.654 4.406 2.706 4.442 ;
      RECT 2.254 4.406 2.306 4.442 ;
      RECT 1.854 4.406 1.906 4.442 ;
      RECT 1.454 4.406 1.506 4.442 ;
      RECT 1.054 4.406 1.106 4.442 ;
      RECT 0.654 4.406 0.706 4.442 ;
      RECT 21.978 4.182 22.022 4.218 ;
      RECT 21.096 4.182 21.14 4.218 ;
      RECT 14.86 4.182 14.904 4.218 ;
      RECT 13.978 4.182 14.022 4.218 ;
      RECT 35.494 3.958 35.546 3.994 ;
      RECT 35.094 3.958 35.146 3.994 ;
      RECT 34.694 3.958 34.746 3.994 ;
      RECT 34.294 3.958 34.346 3.994 ;
      RECT 33.894 3.958 33.946 3.994 ;
      RECT 33.494 3.958 33.546 3.994 ;
      RECT 33.094 3.958 33.146 3.994 ;
      RECT 32.694 3.958 32.746 3.994 ;
      RECT 32.294 3.958 32.346 3.994 ;
      RECT 31.894 3.958 31.946 3.994 ;
      RECT 31.494 3.958 31.546 3.994 ;
      RECT 31.094 3.958 31.146 3.994 ;
      RECT 30.694 3.958 30.746 3.994 ;
      RECT 30.294 3.958 30.346 3.994 ;
      RECT 29.894 3.958 29.946 3.994 ;
      RECT 29.494 3.958 29.546 3.994 ;
      RECT 29.094 3.958 29.146 3.994 ;
      RECT 28.694 3.958 28.746 3.994 ;
      RECT 28.294 3.958 28.346 3.994 ;
      RECT 27.894 3.958 27.946 3.994 ;
      RECT 27.494 3.958 27.546 3.994 ;
      RECT 27.094 3.958 27.146 3.994 ;
      RECT 26.694 3.958 26.746 3.994 ;
      RECT 26.294 3.958 26.346 3.994 ;
      RECT 25.894 3.958 25.946 3.994 ;
      RECT 25.494 3.958 25.546 3.994 ;
      RECT 25.094 3.958 25.146 3.994 ;
      RECT 24.694 3.958 24.746 3.994 ;
      RECT 24.294 3.958 24.346 3.994 ;
      RECT 23.894 3.958 23.946 3.994 ;
      RECT 23.494 3.958 23.546 3.994 ;
      RECT 23.094 3.958 23.146 3.994 ;
      RECT 21.814 3.958 21.868 3.994 ;
      RECT 19.838 3.958 19.886 3.994 ;
      RECT 19.53 3.958 19.578 3.994 ;
      RECT 16.882 3.958 16.936 3.994 ;
      RECT 16.422 3.958 16.47 3.994 ;
      RECT 16.114 3.958 16.162 3.994 ;
      RECT 14.132 3.958 14.186 3.994 ;
      RECT 13.294 3.958 13.346 3.994 ;
      RECT 12.894 3.958 12.946 3.994 ;
      RECT 12.494 3.958 12.546 3.994 ;
      RECT 12.094 3.958 12.146 3.994 ;
      RECT 11.694 3.958 11.746 3.994 ;
      RECT 11.294 3.958 11.346 3.994 ;
      RECT 10.894 3.958 10.946 3.994 ;
      RECT 10.494 3.958 10.546 3.994 ;
      RECT 10.094 3.958 10.146 3.994 ;
      RECT 9.694 3.958 9.746 3.994 ;
      RECT 9.294 3.958 9.346 3.994 ;
      RECT 8.894 3.958 8.946 3.994 ;
      RECT 8.494 3.958 8.546 3.994 ;
      RECT 8.094 3.958 8.146 3.994 ;
      RECT 7.694 3.958 7.746 3.994 ;
      RECT 7.294 3.958 7.346 3.994 ;
      RECT 6.894 3.958 6.946 3.994 ;
      RECT 6.494 3.958 6.546 3.994 ;
      RECT 6.094 3.958 6.146 3.994 ;
      RECT 5.694 3.958 5.746 3.994 ;
      RECT 5.294 3.958 5.346 3.994 ;
      RECT 4.894 3.958 4.946 3.994 ;
      RECT 4.494 3.958 4.546 3.994 ;
      RECT 4.094 3.958 4.146 3.994 ;
      RECT 3.694 3.958 3.746 3.994 ;
      RECT 3.294 3.958 3.346 3.994 ;
      RECT 2.894 3.958 2.946 3.994 ;
      RECT 2.494 3.958 2.546 3.994 ;
      RECT 2.094 3.958 2.146 3.994 ;
      RECT 1.694 3.958 1.746 3.994 ;
      RECT 1.294 3.958 1.346 3.994 ;
      RECT 0.894 3.958 0.946 3.994 ;
      RECT 21.414 3.882 21.468 3.918 ;
      RECT 14.532 3.882 14.586 3.918 ;
      RECT 19.606 3.729 19.654 3.765 ;
      RECT 18.08 3.729 18.12 3.765 ;
      RECT 16.718 3.729 16.772 3.765 ;
      RECT 16.346 3.729 16.394 3.765 ;
      RECT 20.37 3.7345 20.442 3.7595 ;
      RECT 18.764 3.7345 18.836 3.7595 ;
      RECT 15.558 3.7345 15.63 3.7595 ;
      RECT 21.978 3.582 22.022 3.618 ;
      RECT 13.978 3.582 14.022 3.618 ;
      RECT 18.764 3.5875 18.836 3.6125 ;
      RECT 19.762 3.435 19.81 3.471 ;
      RECT 17.616 3.435 17.656 3.471 ;
      RECT 16.19 3.435 16.238 3.471 ;
      RECT 35.254 3.206 35.306 3.242 ;
      RECT 34.854 3.206 34.906 3.242 ;
      RECT 34.454 3.206 34.506 3.242 ;
      RECT 34.054 3.206 34.106 3.242 ;
      RECT 33.654 3.206 33.706 3.242 ;
      RECT 33.254 3.206 33.306 3.242 ;
      RECT 32.854 3.206 32.906 3.242 ;
      RECT 32.454 3.206 32.506 3.242 ;
      RECT 32.054 3.206 32.106 3.242 ;
      RECT 31.654 3.206 31.706 3.242 ;
      RECT 31.254 3.206 31.306 3.242 ;
      RECT 30.854 3.206 30.906 3.242 ;
      RECT 30.454 3.206 30.506 3.242 ;
      RECT 30.054 3.206 30.106 3.242 ;
      RECT 29.654 3.206 29.706 3.242 ;
      RECT 29.254 3.206 29.306 3.242 ;
      RECT 28.854 3.206 28.906 3.242 ;
      RECT 28.454 3.206 28.506 3.242 ;
      RECT 28.054 3.206 28.106 3.242 ;
      RECT 27.654 3.206 27.706 3.242 ;
      RECT 27.254 3.206 27.306 3.242 ;
      RECT 26.854 3.206 26.906 3.242 ;
      RECT 26.454 3.206 26.506 3.242 ;
      RECT 26.054 3.206 26.106 3.242 ;
      RECT 25.654 3.206 25.706 3.242 ;
      RECT 25.254 3.206 25.306 3.242 ;
      RECT 24.854 3.206 24.906 3.242 ;
      RECT 24.454 3.206 24.506 3.242 ;
      RECT 24.054 3.206 24.106 3.242 ;
      RECT 23.654 3.206 23.706 3.242 ;
      RECT 23.254 3.206 23.306 3.242 ;
      RECT 22.854 3.206 22.906 3.242 ;
      RECT 22.694 3.206 22.746 3.242 ;
      RECT 21.732 3.206 21.786 3.242 ;
      RECT 14.214 3.206 14.268 3.242 ;
      RECT 13.054 3.206 13.106 3.242 ;
      RECT 12.654 3.206 12.706 3.242 ;
      RECT 12.254 3.206 12.306 3.242 ;
      RECT 11.854 3.206 11.906 3.242 ;
      RECT 11.454 3.206 11.506 3.242 ;
      RECT 11.054 3.206 11.106 3.242 ;
      RECT 10.654 3.206 10.706 3.242 ;
      RECT 10.254 3.206 10.306 3.242 ;
      RECT 9.854 3.206 9.906 3.242 ;
      RECT 9.454 3.206 9.506 3.242 ;
      RECT 9.054 3.206 9.106 3.242 ;
      RECT 8.654 3.206 8.706 3.242 ;
      RECT 8.254 3.206 8.306 3.242 ;
      RECT 7.854 3.206 7.906 3.242 ;
      RECT 7.454 3.206 7.506 3.242 ;
      RECT 7.054 3.206 7.106 3.242 ;
      RECT 6.654 3.206 6.706 3.242 ;
      RECT 6.254 3.206 6.306 3.242 ;
      RECT 5.854 3.206 5.906 3.242 ;
      RECT 5.454 3.206 5.506 3.242 ;
      RECT 5.054 3.206 5.106 3.242 ;
      RECT 4.654 3.206 4.706 3.242 ;
      RECT 4.254 3.206 4.306 3.242 ;
      RECT 3.854 3.206 3.906 3.242 ;
      RECT 3.454 3.206 3.506 3.242 ;
      RECT 3.054 3.206 3.106 3.242 ;
      RECT 2.654 3.206 2.706 3.242 ;
      RECT 2.254 3.206 2.306 3.242 ;
      RECT 1.854 3.206 1.906 3.242 ;
      RECT 1.454 3.206 1.506 3.242 ;
      RECT 1.054 3.206 1.106 3.242 ;
      RECT 0.654 3.206 0.706 3.242 ;
      RECT 21.978 2.982 22.022 3.018 ;
      RECT 21.096 2.982 21.14 3.018 ;
      RECT 14.86 2.982 14.904 3.018 ;
      RECT 13.978 2.982 14.022 3.018 ;
      RECT 35.494 2.758 35.546 2.794 ;
      RECT 35.094 2.758 35.146 2.794 ;
      RECT 34.694 2.758 34.746 2.794 ;
      RECT 34.294 2.758 34.346 2.794 ;
      RECT 33.894 2.758 33.946 2.794 ;
      RECT 33.494 2.758 33.546 2.794 ;
      RECT 33.094 2.758 33.146 2.794 ;
      RECT 32.694 2.758 32.746 2.794 ;
      RECT 32.294 2.758 32.346 2.794 ;
      RECT 31.894 2.758 31.946 2.794 ;
      RECT 31.494 2.758 31.546 2.794 ;
      RECT 31.094 2.758 31.146 2.794 ;
      RECT 30.694 2.758 30.746 2.794 ;
      RECT 30.294 2.758 30.346 2.794 ;
      RECT 29.894 2.758 29.946 2.794 ;
      RECT 29.494 2.758 29.546 2.794 ;
      RECT 29.094 2.758 29.146 2.794 ;
      RECT 28.694 2.758 28.746 2.794 ;
      RECT 28.294 2.758 28.346 2.794 ;
      RECT 27.894 2.758 27.946 2.794 ;
      RECT 27.494 2.758 27.546 2.794 ;
      RECT 27.094 2.758 27.146 2.794 ;
      RECT 26.694 2.758 26.746 2.794 ;
      RECT 26.294 2.758 26.346 2.794 ;
      RECT 25.894 2.758 25.946 2.794 ;
      RECT 25.494 2.758 25.546 2.794 ;
      RECT 25.094 2.758 25.146 2.794 ;
      RECT 24.694 2.758 24.746 2.794 ;
      RECT 24.294 2.758 24.346 2.794 ;
      RECT 23.894 2.758 23.946 2.794 ;
      RECT 23.494 2.758 23.546 2.794 ;
      RECT 23.094 2.758 23.146 2.794 ;
      RECT 21.814 2.758 21.868 2.794 ;
      RECT 19.838 2.758 19.886 2.794 ;
      RECT 19.53 2.758 19.578 2.794 ;
      RECT 16.882 2.758 16.936 2.794 ;
      RECT 16.422 2.758 16.47 2.794 ;
      RECT 16.114 2.758 16.162 2.794 ;
      RECT 14.132 2.758 14.186 2.794 ;
      RECT 13.294 2.758 13.346 2.794 ;
      RECT 12.894 2.758 12.946 2.794 ;
      RECT 12.494 2.758 12.546 2.794 ;
      RECT 12.094 2.758 12.146 2.794 ;
      RECT 11.694 2.758 11.746 2.794 ;
      RECT 11.294 2.758 11.346 2.794 ;
      RECT 10.894 2.758 10.946 2.794 ;
      RECT 10.494 2.758 10.546 2.794 ;
      RECT 10.094 2.758 10.146 2.794 ;
      RECT 9.694 2.758 9.746 2.794 ;
      RECT 9.294 2.758 9.346 2.794 ;
      RECT 8.894 2.758 8.946 2.794 ;
      RECT 8.494 2.758 8.546 2.794 ;
      RECT 8.094 2.758 8.146 2.794 ;
      RECT 7.694 2.758 7.746 2.794 ;
      RECT 7.294 2.758 7.346 2.794 ;
      RECT 6.894 2.758 6.946 2.794 ;
      RECT 6.494 2.758 6.546 2.794 ;
      RECT 6.094 2.758 6.146 2.794 ;
      RECT 5.694 2.758 5.746 2.794 ;
      RECT 5.294 2.758 5.346 2.794 ;
      RECT 4.894 2.758 4.946 2.794 ;
      RECT 4.494 2.758 4.546 2.794 ;
      RECT 4.094 2.758 4.146 2.794 ;
      RECT 3.694 2.758 3.746 2.794 ;
      RECT 3.294 2.758 3.346 2.794 ;
      RECT 2.894 2.758 2.946 2.794 ;
      RECT 2.494 2.758 2.546 2.794 ;
      RECT 2.094 2.758 2.146 2.794 ;
      RECT 1.694 2.758 1.746 2.794 ;
      RECT 1.294 2.758 1.346 2.794 ;
      RECT 0.894 2.758 0.946 2.794 ;
      RECT 21.414 2.682 21.468 2.718 ;
      RECT 14.532 2.682 14.586 2.718 ;
      RECT 19.606 2.529 19.654 2.565 ;
      RECT 18.08 2.529 18.12 2.565 ;
      RECT 16.718 2.529 16.772 2.565 ;
      RECT 16.346 2.529 16.394 2.565 ;
      RECT 20.37 2.5345 20.442 2.5595 ;
      RECT 18.764 2.5345 18.836 2.5595 ;
      RECT 15.558 2.5345 15.63 2.5595 ;
      RECT 21.978 2.382 22.022 2.418 ;
      RECT 13.978 2.382 14.022 2.418 ;
      RECT 18.764 2.3875 18.836 2.4125 ;
      RECT 19.762 2.235 19.81 2.271 ;
      RECT 17.616 2.235 17.656 2.271 ;
      RECT 16.19 2.235 16.238 2.271 ;
      RECT 35.254 2.006 35.306 2.042 ;
      RECT 34.854 2.006 34.906 2.042 ;
      RECT 34.454 2.006 34.506 2.042 ;
      RECT 34.054 2.006 34.106 2.042 ;
      RECT 33.654 2.006 33.706 2.042 ;
      RECT 33.254 2.006 33.306 2.042 ;
      RECT 32.854 2.006 32.906 2.042 ;
      RECT 32.454 2.006 32.506 2.042 ;
      RECT 32.054 2.006 32.106 2.042 ;
      RECT 31.654 2.006 31.706 2.042 ;
      RECT 31.254 2.006 31.306 2.042 ;
      RECT 30.854 2.006 30.906 2.042 ;
      RECT 30.454 2.006 30.506 2.042 ;
      RECT 30.054 2.006 30.106 2.042 ;
      RECT 29.654 2.006 29.706 2.042 ;
      RECT 29.254 2.006 29.306 2.042 ;
      RECT 28.854 2.006 28.906 2.042 ;
      RECT 28.454 2.006 28.506 2.042 ;
      RECT 28.054 2.006 28.106 2.042 ;
      RECT 27.654 2.006 27.706 2.042 ;
      RECT 27.254 2.006 27.306 2.042 ;
      RECT 26.854 2.006 26.906 2.042 ;
      RECT 26.454 2.006 26.506 2.042 ;
      RECT 26.054 2.006 26.106 2.042 ;
      RECT 25.654 2.006 25.706 2.042 ;
      RECT 25.254 2.006 25.306 2.042 ;
      RECT 24.854 2.006 24.906 2.042 ;
      RECT 24.454 2.006 24.506 2.042 ;
      RECT 24.054 2.006 24.106 2.042 ;
      RECT 23.654 2.006 23.706 2.042 ;
      RECT 23.254 2.006 23.306 2.042 ;
      RECT 22.854 2.006 22.906 2.042 ;
      RECT 22.694 2.006 22.746 2.042 ;
      RECT 21.732 2.006 21.786 2.042 ;
      RECT 14.214 2.006 14.268 2.042 ;
      RECT 13.054 2.006 13.106 2.042 ;
      RECT 12.654 2.006 12.706 2.042 ;
      RECT 12.254 2.006 12.306 2.042 ;
      RECT 11.854 2.006 11.906 2.042 ;
      RECT 11.454 2.006 11.506 2.042 ;
      RECT 11.054 2.006 11.106 2.042 ;
      RECT 10.654 2.006 10.706 2.042 ;
      RECT 10.254 2.006 10.306 2.042 ;
      RECT 9.854 2.006 9.906 2.042 ;
      RECT 9.454 2.006 9.506 2.042 ;
      RECT 9.054 2.006 9.106 2.042 ;
      RECT 8.654 2.006 8.706 2.042 ;
      RECT 8.254 2.006 8.306 2.042 ;
      RECT 7.854 2.006 7.906 2.042 ;
      RECT 7.454 2.006 7.506 2.042 ;
      RECT 7.054 2.006 7.106 2.042 ;
      RECT 6.654 2.006 6.706 2.042 ;
      RECT 6.254 2.006 6.306 2.042 ;
      RECT 5.854 2.006 5.906 2.042 ;
      RECT 5.454 2.006 5.506 2.042 ;
      RECT 5.054 2.006 5.106 2.042 ;
      RECT 4.654 2.006 4.706 2.042 ;
      RECT 4.254 2.006 4.306 2.042 ;
      RECT 3.854 2.006 3.906 2.042 ;
      RECT 3.454 2.006 3.506 2.042 ;
      RECT 3.054 2.006 3.106 2.042 ;
      RECT 2.654 2.006 2.706 2.042 ;
      RECT 2.254 2.006 2.306 2.042 ;
      RECT 1.854 2.006 1.906 2.042 ;
      RECT 1.454 2.006 1.506 2.042 ;
      RECT 1.054 2.006 1.106 2.042 ;
      RECT 0.654 2.006 0.706 2.042 ;
      RECT 21.978 1.782 22.022 1.818 ;
      RECT 21.096 1.782 21.14 1.818 ;
      RECT 14.86 1.782 14.904 1.818 ;
      RECT 13.978 1.782 14.022 1.818 ;
      RECT 35.494 1.558 35.546 1.594 ;
      RECT 35.094 1.558 35.146 1.594 ;
      RECT 34.694 1.558 34.746 1.594 ;
      RECT 34.294 1.558 34.346 1.594 ;
      RECT 33.894 1.558 33.946 1.594 ;
      RECT 33.494 1.558 33.546 1.594 ;
      RECT 33.094 1.558 33.146 1.594 ;
      RECT 32.694 1.558 32.746 1.594 ;
      RECT 32.294 1.558 32.346 1.594 ;
      RECT 31.894 1.558 31.946 1.594 ;
      RECT 31.494 1.558 31.546 1.594 ;
      RECT 31.094 1.558 31.146 1.594 ;
      RECT 30.694 1.558 30.746 1.594 ;
      RECT 30.294 1.558 30.346 1.594 ;
      RECT 29.894 1.558 29.946 1.594 ;
      RECT 29.494 1.558 29.546 1.594 ;
      RECT 29.094 1.558 29.146 1.594 ;
      RECT 28.694 1.558 28.746 1.594 ;
      RECT 28.294 1.558 28.346 1.594 ;
      RECT 27.894 1.558 27.946 1.594 ;
      RECT 27.494 1.558 27.546 1.594 ;
      RECT 27.094 1.558 27.146 1.594 ;
      RECT 26.694 1.558 26.746 1.594 ;
      RECT 26.294 1.558 26.346 1.594 ;
      RECT 25.894 1.558 25.946 1.594 ;
      RECT 25.494 1.558 25.546 1.594 ;
      RECT 25.094 1.558 25.146 1.594 ;
      RECT 24.694 1.558 24.746 1.594 ;
      RECT 24.294 1.558 24.346 1.594 ;
      RECT 23.894 1.558 23.946 1.594 ;
      RECT 23.494 1.558 23.546 1.594 ;
      RECT 23.094 1.558 23.146 1.594 ;
      RECT 21.814 1.558 21.868 1.594 ;
      RECT 19.838 1.558 19.886 1.594 ;
      RECT 19.53 1.558 19.578 1.594 ;
      RECT 16.882 1.558 16.936 1.594 ;
      RECT 16.422 1.558 16.47 1.594 ;
      RECT 16.114 1.558 16.162 1.594 ;
      RECT 14.132 1.558 14.186 1.594 ;
      RECT 13.294 1.558 13.346 1.594 ;
      RECT 12.894 1.558 12.946 1.594 ;
      RECT 12.494 1.558 12.546 1.594 ;
      RECT 12.094 1.558 12.146 1.594 ;
      RECT 11.694 1.558 11.746 1.594 ;
      RECT 11.294 1.558 11.346 1.594 ;
      RECT 10.894 1.558 10.946 1.594 ;
      RECT 10.494 1.558 10.546 1.594 ;
      RECT 10.094 1.558 10.146 1.594 ;
      RECT 9.694 1.558 9.746 1.594 ;
      RECT 9.294 1.558 9.346 1.594 ;
      RECT 8.894 1.558 8.946 1.594 ;
      RECT 8.494 1.558 8.546 1.594 ;
      RECT 8.094 1.558 8.146 1.594 ;
      RECT 7.694 1.558 7.746 1.594 ;
      RECT 7.294 1.558 7.346 1.594 ;
      RECT 6.894 1.558 6.946 1.594 ;
      RECT 6.494 1.558 6.546 1.594 ;
      RECT 6.094 1.558 6.146 1.594 ;
      RECT 5.694 1.558 5.746 1.594 ;
      RECT 5.294 1.558 5.346 1.594 ;
      RECT 4.894 1.558 4.946 1.594 ;
      RECT 4.494 1.558 4.546 1.594 ;
      RECT 4.094 1.558 4.146 1.594 ;
      RECT 3.694 1.558 3.746 1.594 ;
      RECT 3.294 1.558 3.346 1.594 ;
      RECT 2.894 1.558 2.946 1.594 ;
      RECT 2.494 1.558 2.546 1.594 ;
      RECT 2.094 1.558 2.146 1.594 ;
      RECT 1.694 1.558 1.746 1.594 ;
      RECT 1.294 1.558 1.346 1.594 ;
      RECT 0.894 1.558 0.946 1.594 ;
      RECT 21.414 1.482 21.468 1.518 ;
      RECT 14.532 1.482 14.586 1.518 ;
      RECT 19.606 1.329 19.654 1.365 ;
      RECT 18.08 1.329 18.12 1.365 ;
      RECT 16.718 1.329 16.772 1.365 ;
      RECT 16.346 1.329 16.394 1.365 ;
      RECT 20.37 1.3345 20.442 1.3595 ;
      RECT 18.764 1.3345 18.836 1.3595 ;
      RECT 15.558 1.3345 15.63 1.3595 ;
      RECT 21.978 1.182 22.022 1.218 ;
      RECT 13.978 1.182 14.022 1.218 ;
      RECT 18.764 1.1875 18.836 1.2125 ;
      RECT 19.762 1.035 19.81 1.071 ;
      RECT 17.616 1.035 17.656 1.071 ;
      RECT 16.19 1.035 16.238 1.071 ;
      RECT 35.254 0.806 35.306 0.842 ;
      RECT 34.854 0.806 34.906 0.842 ;
      RECT 34.454 0.806 34.506 0.842 ;
      RECT 34.054 0.806 34.106 0.842 ;
      RECT 33.654 0.806 33.706 0.842 ;
      RECT 33.254 0.806 33.306 0.842 ;
      RECT 32.854 0.806 32.906 0.842 ;
      RECT 32.454 0.806 32.506 0.842 ;
      RECT 32.054 0.806 32.106 0.842 ;
      RECT 31.654 0.806 31.706 0.842 ;
      RECT 31.254 0.806 31.306 0.842 ;
      RECT 30.854 0.806 30.906 0.842 ;
      RECT 30.454 0.806 30.506 0.842 ;
      RECT 30.054 0.806 30.106 0.842 ;
      RECT 29.654 0.806 29.706 0.842 ;
      RECT 29.254 0.806 29.306 0.842 ;
      RECT 28.854 0.806 28.906 0.842 ;
      RECT 28.454 0.806 28.506 0.842 ;
      RECT 28.054 0.806 28.106 0.842 ;
      RECT 27.654 0.806 27.706 0.842 ;
      RECT 27.254 0.806 27.306 0.842 ;
      RECT 26.854 0.806 26.906 0.842 ;
      RECT 26.454 0.806 26.506 0.842 ;
      RECT 26.054 0.806 26.106 0.842 ;
      RECT 25.654 0.806 25.706 0.842 ;
      RECT 25.254 0.806 25.306 0.842 ;
      RECT 24.854 0.806 24.906 0.842 ;
      RECT 24.454 0.806 24.506 0.842 ;
      RECT 24.054 0.806 24.106 0.842 ;
      RECT 23.654 0.806 23.706 0.842 ;
      RECT 23.254 0.806 23.306 0.842 ;
      RECT 22.854 0.806 22.906 0.842 ;
      RECT 22.694 0.806 22.746 0.842 ;
      RECT 21.732 0.806 21.786 0.842 ;
      RECT 14.214 0.806 14.268 0.842 ;
      RECT 13.054 0.806 13.106 0.842 ;
      RECT 12.654 0.806 12.706 0.842 ;
      RECT 12.254 0.806 12.306 0.842 ;
      RECT 11.854 0.806 11.906 0.842 ;
      RECT 11.454 0.806 11.506 0.842 ;
      RECT 11.054 0.806 11.106 0.842 ;
      RECT 10.654 0.806 10.706 0.842 ;
      RECT 10.254 0.806 10.306 0.842 ;
      RECT 9.854 0.806 9.906 0.842 ;
      RECT 9.454 0.806 9.506 0.842 ;
      RECT 9.054 0.806 9.106 0.842 ;
      RECT 8.654 0.806 8.706 0.842 ;
      RECT 8.254 0.806 8.306 0.842 ;
      RECT 7.854 0.806 7.906 0.842 ;
      RECT 7.454 0.806 7.506 0.842 ;
      RECT 7.054 0.806 7.106 0.842 ;
      RECT 6.654 0.806 6.706 0.842 ;
      RECT 6.254 0.806 6.306 0.842 ;
      RECT 5.854 0.806 5.906 0.842 ;
      RECT 5.454 0.806 5.506 0.842 ;
      RECT 5.054 0.806 5.106 0.842 ;
      RECT 4.654 0.806 4.706 0.842 ;
      RECT 4.254 0.806 4.306 0.842 ;
      RECT 3.854 0.806 3.906 0.842 ;
      RECT 3.454 0.806 3.506 0.842 ;
      RECT 3.054 0.806 3.106 0.842 ;
      RECT 2.654 0.806 2.706 0.842 ;
      RECT 2.254 0.806 2.306 0.842 ;
      RECT 1.854 0.806 1.906 0.842 ;
      RECT 1.454 0.806 1.506 0.842 ;
      RECT 1.054 0.806 1.106 0.842 ;
      RECT 0.654 0.806 0.706 0.842 ;
      RECT 21.978 0.582 22.022 0.618 ;
      RECT 21.096 0.582 21.14 0.618 ;
      RECT 14.86 0.582 14.904 0.618 ;
      RECT 13.978 0.582 14.022 0.618 ;
      RECT 0.574 0.281 0.626 0.317 ;
      RECT 0.574 72.403 0.626 72.439 ;
      RECT 0.654 0.806 0.706 0.842 ;
      RECT 0.654 2.006 0.706 2.042 ;
      RECT 0.654 3.206 0.706 3.242 ;
      RECT 0.654 4.406 0.706 4.442 ;
      RECT 0.654 5.606 0.706 5.642 ;
      RECT 0.654 6.806 0.706 6.842 ;
      RECT 0.654 8.006 0.706 8.042 ;
      RECT 0.654 9.206 0.706 9.242 ;
      RECT 0.654 10.406 0.706 10.442 ;
      RECT 0.654 11.606 0.706 11.642 ;
      RECT 0.654 12.806 0.706 12.842 ;
      RECT 0.654 14.006 0.706 14.042 ;
      RECT 0.654 15.206 0.706 15.242 ;
      RECT 0.654 16.406 0.706 16.442 ;
      RECT 0.654 17.606 0.706 17.642 ;
      RECT 0.654 18.806 0.706 18.842 ;
      RECT 0.654 20.006 0.706 20.042 ;
      RECT 0.654 21.206 0.706 21.242 ;
      RECT 0.654 22.406 0.706 22.442 ;
      RECT 0.654 23.606 0.706 23.642 ;
      RECT 0.654 24.806 0.706 24.842 ;
      RECT 0.654 26.006 0.706 26.042 ;
      RECT 0.654 27.206 0.706 27.242 ;
      RECT 0.654 28.406 0.706 28.442 ;
      RECT 0.654 29.606 0.706 29.642 ;
      RECT 0.654 30.806 0.706 30.842 ;
      RECT 0.654 32.622 0.706 32.658 ;
      RECT 0.654 32.862 0.706 32.898 ;
      RECT 0.654 38.622 0.706 38.658 ;
      RECT 0.654 38.862 0.706 38.898 ;
      RECT 0.654 39.926 0.706 39.962 ;
      RECT 0.654 41.126 0.706 41.162 ;
      RECT 0.654 42.326 0.706 42.362 ;
      RECT 0.654 43.526 0.706 43.562 ;
      RECT 0.654 44.726 0.706 44.762 ;
      RECT 0.654 45.926 0.706 45.962 ;
      RECT 0.654 47.126 0.706 47.162 ;
      RECT 0.654 48.326 0.706 48.362 ;
      RECT 0.654 49.526 0.706 49.562 ;
      RECT 0.654 50.726 0.706 50.762 ;
      RECT 0.654 51.926 0.706 51.962 ;
      RECT 0.654 53.126 0.706 53.162 ;
      RECT 0.654 54.326 0.706 54.362 ;
      RECT 0.654 55.526 0.706 55.562 ;
      RECT 0.654 56.726 0.706 56.762 ;
      RECT 0.654 57.926 0.706 57.962 ;
      RECT 0.654 59.126 0.706 59.162 ;
      RECT 0.654 60.326 0.706 60.362 ;
      RECT 0.654 61.526 0.706 61.562 ;
      RECT 0.654 62.726 0.706 62.762 ;
      RECT 0.654 63.926 0.706 63.962 ;
      RECT 0.654 65.126 0.706 65.162 ;
      RECT 0.654 66.326 0.706 66.362 ;
      RECT 0.654 67.526 0.706 67.562 ;
      RECT 0.654 68.726 0.706 68.762 ;
      RECT 0.654 69.926 0.706 69.962 ;
      RECT 0.654 71.126 0.706 71.162 ;
      RECT 0.734 1.558 0.786 1.594 ;
      RECT 0.734 2.758 0.786 2.794 ;
      RECT 0.734 3.958 0.786 3.994 ;
      RECT 0.734 5.158 0.786 5.194 ;
      RECT 0.734 6.358 0.786 6.394 ;
      RECT 0.734 7.558 0.786 7.594 ;
      RECT 0.734 8.758 0.786 8.794 ;
      RECT 0.734 9.958 0.786 9.994 ;
      RECT 0.734 11.158 0.786 11.194 ;
      RECT 0.734 12.358 0.786 12.394 ;
      RECT 0.734 13.558 0.786 13.594 ;
      RECT 0.734 14.758 0.786 14.794 ;
      RECT 0.734 15.958 0.786 15.994 ;
      RECT 0.734 17.158 0.786 17.194 ;
      RECT 0.734 18.358 0.786 18.394 ;
      RECT 0.734 19.558 0.786 19.594 ;
      RECT 0.734 20.758 0.786 20.794 ;
      RECT 0.734 21.958 0.786 21.994 ;
      RECT 0.734 23.158 0.786 23.194 ;
      RECT 0.734 24.358 0.786 24.394 ;
      RECT 0.734 25.558 0.786 25.594 ;
      RECT 0.734 26.758 0.786 26.794 ;
      RECT 0.734 27.958 0.786 27.994 ;
      RECT 0.734 29.158 0.786 29.194 ;
      RECT 0.734 30.358 0.786 30.394 ;
      RECT 0.734 31.558 0.786 31.594 ;
      RECT 0.734 33.342 0.786 33.378 ;
      RECT 0.734 33.582 0.786 33.618 ;
      RECT 0.734 37.902 0.786 37.938 ;
      RECT 0.734 38.142 0.786 38.178 ;
      RECT 0.734 40.678 0.786 40.714 ;
      RECT 0.734 41.878 0.786 41.914 ;
      RECT 0.734 43.078 0.786 43.114 ;
      RECT 0.734 44.278 0.786 44.314 ;
      RECT 0.734 45.478 0.786 45.514 ;
      RECT 0.734 46.678 0.786 46.714 ;
      RECT 0.734 47.878 0.786 47.914 ;
      RECT 0.734 49.078 0.786 49.114 ;
      RECT 0.734 50.278 0.786 50.314 ;
      RECT 0.734 51.478 0.786 51.514 ;
      RECT 0.734 52.678 0.786 52.714 ;
      RECT 0.734 53.878 0.786 53.914 ;
      RECT 0.734 55.078 0.786 55.114 ;
      RECT 0.734 56.278 0.786 56.314 ;
      RECT 0.734 57.478 0.786 57.514 ;
      RECT 0.734 58.678 0.786 58.714 ;
      RECT 0.734 59.878 0.786 59.914 ;
      RECT 0.734 61.078 0.786 61.114 ;
      RECT 0.734 62.278 0.786 62.314 ;
      RECT 0.734 63.478 0.786 63.514 ;
      RECT 0.734 64.678 0.786 64.714 ;
      RECT 0.734 65.878 0.786 65.914 ;
      RECT 0.734 67.078 0.786 67.114 ;
      RECT 0.734 68.278 0.786 68.314 ;
      RECT 0.734 69.478 0.786 69.514 ;
      RECT 0.734 70.678 0.786 70.714 ;
      RECT 0.734 71.878 0.786 71.914 ;
      RECT 0.814 0.806 0.866 0.842 ;
      RECT 0.814 2.006 0.866 2.042 ;
      RECT 0.814 3.206 0.866 3.242 ;
      RECT 0.814 4.406 0.866 4.442 ;
      RECT 0.814 5.606 0.866 5.642 ;
      RECT 0.814 6.806 0.866 6.842 ;
      RECT 0.814 8.006 0.866 8.042 ;
      RECT 0.814 9.206 0.866 9.242 ;
      RECT 0.814 10.406 0.866 10.442 ;
      RECT 0.814 11.606 0.866 11.642 ;
      RECT 0.814 12.806 0.866 12.842 ;
      RECT 0.814 14.006 0.866 14.042 ;
      RECT 0.814 15.206 0.866 15.242 ;
      RECT 0.814 16.406 0.866 16.442 ;
      RECT 0.814 17.606 0.866 17.642 ;
      RECT 0.814 18.806 0.866 18.842 ;
      RECT 0.814 20.006 0.866 20.042 ;
      RECT 0.814 21.206 0.866 21.242 ;
      RECT 0.814 22.406 0.866 22.442 ;
      RECT 0.814 23.606 0.866 23.642 ;
      RECT 0.814 24.806 0.866 24.842 ;
      RECT 0.814 26.006 0.866 26.042 ;
      RECT 0.814 27.206 0.866 27.242 ;
      RECT 0.814 28.406 0.866 28.442 ;
      RECT 0.814 29.606 0.866 29.642 ;
      RECT 0.814 30.806 0.866 30.842 ;
      RECT 0.814 32.622 0.866 32.658 ;
      RECT 0.814 32.862 0.866 32.898 ;
      RECT 0.814 38.622 0.866 38.658 ;
      RECT 0.814 38.862 0.866 38.898 ;
      RECT 0.814 39.926 0.866 39.962 ;
      RECT 0.814 41.126 0.866 41.162 ;
      RECT 0.814 42.326 0.866 42.362 ;
      RECT 0.814 43.526 0.866 43.562 ;
      RECT 0.814 44.726 0.866 44.762 ;
      RECT 0.814 45.926 0.866 45.962 ;
      RECT 0.814 47.126 0.866 47.162 ;
      RECT 0.814 48.326 0.866 48.362 ;
      RECT 0.814 49.526 0.866 49.562 ;
      RECT 0.814 50.726 0.866 50.762 ;
      RECT 0.814 51.926 0.866 51.962 ;
      RECT 0.814 53.126 0.866 53.162 ;
      RECT 0.814 54.326 0.866 54.362 ;
      RECT 0.814 55.526 0.866 55.562 ;
      RECT 0.814 56.726 0.866 56.762 ;
      RECT 0.814 57.926 0.866 57.962 ;
      RECT 0.814 59.126 0.866 59.162 ;
      RECT 0.814 60.326 0.866 60.362 ;
      RECT 0.814 61.526 0.866 61.562 ;
      RECT 0.814 62.726 0.866 62.762 ;
      RECT 0.814 63.926 0.866 63.962 ;
      RECT 0.814 65.126 0.866 65.162 ;
      RECT 0.814 66.326 0.866 66.362 ;
      RECT 0.814 67.526 0.866 67.562 ;
      RECT 0.814 68.726 0.866 68.762 ;
      RECT 0.814 69.926 0.866 69.962 ;
      RECT 0.814 71.126 0.866 71.162 ;
      RECT 0.894 1.558 0.946 1.594 ;
      RECT 0.894 2.758 0.946 2.794 ;
      RECT 0.894 3.958 0.946 3.994 ;
      RECT 0.894 5.158 0.946 5.194 ;
      RECT 0.894 6.358 0.946 6.394 ;
      RECT 0.894 7.558 0.946 7.594 ;
      RECT 0.894 8.758 0.946 8.794 ;
      RECT 0.894 9.958 0.946 9.994 ;
      RECT 0.894 11.158 0.946 11.194 ;
      RECT 0.894 12.358 0.946 12.394 ;
      RECT 0.894 13.558 0.946 13.594 ;
      RECT 0.894 14.758 0.946 14.794 ;
      RECT 0.894 15.958 0.946 15.994 ;
      RECT 0.894 17.158 0.946 17.194 ;
      RECT 0.894 18.358 0.946 18.394 ;
      RECT 0.894 19.558 0.946 19.594 ;
      RECT 0.894 20.758 0.946 20.794 ;
      RECT 0.894 21.958 0.946 21.994 ;
      RECT 0.894 23.158 0.946 23.194 ;
      RECT 0.894 24.358 0.946 24.394 ;
      RECT 0.894 25.558 0.946 25.594 ;
      RECT 0.894 26.758 0.946 26.794 ;
      RECT 0.894 27.958 0.946 27.994 ;
      RECT 0.894 29.158 0.946 29.194 ;
      RECT 0.894 30.358 0.946 30.394 ;
      RECT 0.894 31.558 0.946 31.594 ;
      RECT 0.894 33.342 0.946 33.378 ;
      RECT 0.894 33.582 0.946 33.618 ;
      RECT 0.894 37.902 0.946 37.938 ;
      RECT 0.894 38.142 0.946 38.178 ;
      RECT 0.894 40.678 0.946 40.714 ;
      RECT 0.894 41.878 0.946 41.914 ;
      RECT 0.894 43.078 0.946 43.114 ;
      RECT 0.894 44.278 0.946 44.314 ;
      RECT 0.894 45.478 0.946 45.514 ;
      RECT 0.894 46.678 0.946 46.714 ;
      RECT 0.894 47.878 0.946 47.914 ;
      RECT 0.894 49.078 0.946 49.114 ;
      RECT 0.894 50.278 0.946 50.314 ;
      RECT 0.894 51.478 0.946 51.514 ;
      RECT 0.894 52.678 0.946 52.714 ;
      RECT 0.894 53.878 0.946 53.914 ;
      RECT 0.894 55.078 0.946 55.114 ;
      RECT 0.894 56.278 0.946 56.314 ;
      RECT 0.894 57.478 0.946 57.514 ;
      RECT 0.894 58.678 0.946 58.714 ;
      RECT 0.894 59.878 0.946 59.914 ;
      RECT 0.894 61.078 0.946 61.114 ;
      RECT 0.894 62.278 0.946 62.314 ;
      RECT 0.894 63.478 0.946 63.514 ;
      RECT 0.894 64.678 0.946 64.714 ;
      RECT 0.894 65.878 0.946 65.914 ;
      RECT 0.894 67.078 0.946 67.114 ;
      RECT 0.894 68.278 0.946 68.314 ;
      RECT 0.894 69.478 0.946 69.514 ;
      RECT 0.894 70.678 0.946 70.714 ;
      RECT 0.894 71.878 0.946 71.914 ;
      RECT 0.974 0.281 1.026 0.317 ;
      RECT 0.974 72.403 1.026 72.439 ;
      RECT 1.054 0.806 1.106 0.842 ;
      RECT 1.054 2.006 1.106 2.042 ;
      RECT 1.054 3.206 1.106 3.242 ;
      RECT 1.054 4.406 1.106 4.442 ;
      RECT 1.054 5.606 1.106 5.642 ;
      RECT 1.054 6.806 1.106 6.842 ;
      RECT 1.054 8.006 1.106 8.042 ;
      RECT 1.054 9.206 1.106 9.242 ;
      RECT 1.054 10.406 1.106 10.442 ;
      RECT 1.054 11.606 1.106 11.642 ;
      RECT 1.054 12.806 1.106 12.842 ;
      RECT 1.054 14.006 1.106 14.042 ;
      RECT 1.054 15.206 1.106 15.242 ;
      RECT 1.054 16.406 1.106 16.442 ;
      RECT 1.054 17.606 1.106 17.642 ;
      RECT 1.054 18.806 1.106 18.842 ;
      RECT 1.054 20.006 1.106 20.042 ;
      RECT 1.054 21.206 1.106 21.242 ;
      RECT 1.054 22.406 1.106 22.442 ;
      RECT 1.054 23.606 1.106 23.642 ;
      RECT 1.054 24.806 1.106 24.842 ;
      RECT 1.054 26.006 1.106 26.042 ;
      RECT 1.054 27.206 1.106 27.242 ;
      RECT 1.054 28.406 1.106 28.442 ;
      RECT 1.054 29.606 1.106 29.642 ;
      RECT 1.054 30.806 1.106 30.842 ;
      RECT 1.054 32.622 1.106 32.658 ;
      RECT 1.054 32.862 1.106 32.898 ;
      RECT 1.054 34.302 1.106 34.338 ;
      RECT 1.054 34.782 1.106 34.818 ;
      RECT 1.054 36.702 1.106 36.738 ;
      RECT 1.054 37.182 1.106 37.218 ;
      RECT 1.054 38.622 1.106 38.658 ;
      RECT 1.054 38.862 1.106 38.898 ;
      RECT 1.054 39.926 1.106 39.962 ;
      RECT 1.054 41.126 1.106 41.162 ;
      RECT 1.054 42.326 1.106 42.362 ;
      RECT 1.054 43.526 1.106 43.562 ;
      RECT 1.054 44.726 1.106 44.762 ;
      RECT 1.054 45.926 1.106 45.962 ;
      RECT 1.054 47.126 1.106 47.162 ;
      RECT 1.054 48.326 1.106 48.362 ;
      RECT 1.054 49.526 1.106 49.562 ;
      RECT 1.054 50.726 1.106 50.762 ;
      RECT 1.054 51.926 1.106 51.962 ;
      RECT 1.054 53.126 1.106 53.162 ;
      RECT 1.054 54.326 1.106 54.362 ;
      RECT 1.054 55.526 1.106 55.562 ;
      RECT 1.054 56.726 1.106 56.762 ;
      RECT 1.054 57.926 1.106 57.962 ;
      RECT 1.054 59.126 1.106 59.162 ;
      RECT 1.054 60.326 1.106 60.362 ;
      RECT 1.054 61.526 1.106 61.562 ;
      RECT 1.054 62.726 1.106 62.762 ;
      RECT 1.054 63.926 1.106 63.962 ;
      RECT 1.054 65.126 1.106 65.162 ;
      RECT 1.054 66.326 1.106 66.362 ;
      RECT 1.054 67.526 1.106 67.562 ;
      RECT 1.054 68.726 1.106 68.762 ;
      RECT 1.054 69.926 1.106 69.962 ;
      RECT 1.054 71.126 1.106 71.162 ;
      RECT 1.134 1.558 1.186 1.594 ;
      RECT 1.134 2.758 1.186 2.794 ;
      RECT 1.134 3.958 1.186 3.994 ;
      RECT 1.134 5.158 1.186 5.194 ;
      RECT 1.134 6.358 1.186 6.394 ;
      RECT 1.134 7.558 1.186 7.594 ;
      RECT 1.134 8.758 1.186 8.794 ;
      RECT 1.134 9.958 1.186 9.994 ;
      RECT 1.134 11.158 1.186 11.194 ;
      RECT 1.134 12.358 1.186 12.394 ;
      RECT 1.134 13.558 1.186 13.594 ;
      RECT 1.134 14.758 1.186 14.794 ;
      RECT 1.134 15.958 1.186 15.994 ;
      RECT 1.134 17.158 1.186 17.194 ;
      RECT 1.134 18.358 1.186 18.394 ;
      RECT 1.134 19.558 1.186 19.594 ;
      RECT 1.134 20.758 1.186 20.794 ;
      RECT 1.134 21.958 1.186 21.994 ;
      RECT 1.134 23.158 1.186 23.194 ;
      RECT 1.134 24.358 1.186 24.394 ;
      RECT 1.134 25.558 1.186 25.594 ;
      RECT 1.134 26.758 1.186 26.794 ;
      RECT 1.134 27.958 1.186 27.994 ;
      RECT 1.134 29.158 1.186 29.194 ;
      RECT 1.134 30.358 1.186 30.394 ;
      RECT 1.134 31.558 1.186 31.594 ;
      RECT 1.134 33.342 1.186 33.378 ;
      RECT 1.134 33.582 1.186 33.618 ;
      RECT 1.134 37.902 1.186 37.938 ;
      RECT 1.134 38.142 1.186 38.178 ;
      RECT 1.134 40.678 1.186 40.714 ;
      RECT 1.134 41.878 1.186 41.914 ;
      RECT 1.134 43.078 1.186 43.114 ;
      RECT 1.134 44.278 1.186 44.314 ;
      RECT 1.134 45.478 1.186 45.514 ;
      RECT 1.134 46.678 1.186 46.714 ;
      RECT 1.134 47.878 1.186 47.914 ;
      RECT 1.134 49.078 1.186 49.114 ;
      RECT 1.134 50.278 1.186 50.314 ;
      RECT 1.134 51.478 1.186 51.514 ;
      RECT 1.134 52.678 1.186 52.714 ;
      RECT 1.134 53.878 1.186 53.914 ;
      RECT 1.134 55.078 1.186 55.114 ;
      RECT 1.134 56.278 1.186 56.314 ;
      RECT 1.134 57.478 1.186 57.514 ;
      RECT 1.134 58.678 1.186 58.714 ;
      RECT 1.134 59.878 1.186 59.914 ;
      RECT 1.134 61.078 1.186 61.114 ;
      RECT 1.134 62.278 1.186 62.314 ;
      RECT 1.134 63.478 1.186 63.514 ;
      RECT 1.134 64.678 1.186 64.714 ;
      RECT 1.134 65.878 1.186 65.914 ;
      RECT 1.134 67.078 1.186 67.114 ;
      RECT 1.134 68.278 1.186 68.314 ;
      RECT 1.134 69.478 1.186 69.514 ;
      RECT 1.134 70.678 1.186 70.714 ;
      RECT 1.134 71.878 1.186 71.914 ;
      RECT 1.214 0.806 1.266 0.842 ;
      RECT 1.214 2.006 1.266 2.042 ;
      RECT 1.214 3.206 1.266 3.242 ;
      RECT 1.214 4.406 1.266 4.442 ;
      RECT 1.214 5.606 1.266 5.642 ;
      RECT 1.214 6.806 1.266 6.842 ;
      RECT 1.214 8.006 1.266 8.042 ;
      RECT 1.214 9.206 1.266 9.242 ;
      RECT 1.214 10.406 1.266 10.442 ;
      RECT 1.214 11.606 1.266 11.642 ;
      RECT 1.214 12.806 1.266 12.842 ;
      RECT 1.214 14.006 1.266 14.042 ;
      RECT 1.214 15.206 1.266 15.242 ;
      RECT 1.214 16.406 1.266 16.442 ;
      RECT 1.214 17.606 1.266 17.642 ;
      RECT 1.214 18.806 1.266 18.842 ;
      RECT 1.214 20.006 1.266 20.042 ;
      RECT 1.214 21.206 1.266 21.242 ;
      RECT 1.214 22.406 1.266 22.442 ;
      RECT 1.214 23.606 1.266 23.642 ;
      RECT 1.214 24.806 1.266 24.842 ;
      RECT 1.214 26.006 1.266 26.042 ;
      RECT 1.214 27.206 1.266 27.242 ;
      RECT 1.214 28.406 1.266 28.442 ;
      RECT 1.214 29.606 1.266 29.642 ;
      RECT 1.214 30.806 1.266 30.842 ;
      RECT 1.214 32.622 1.266 32.658 ;
      RECT 1.214 32.862 1.266 32.898 ;
      RECT 1.214 38.622 1.266 38.658 ;
      RECT 1.214 38.862 1.266 38.898 ;
      RECT 1.214 39.926 1.266 39.962 ;
      RECT 1.214 41.126 1.266 41.162 ;
      RECT 1.214 42.326 1.266 42.362 ;
      RECT 1.214 43.526 1.266 43.562 ;
      RECT 1.214 44.726 1.266 44.762 ;
      RECT 1.214 45.926 1.266 45.962 ;
      RECT 1.214 47.126 1.266 47.162 ;
      RECT 1.214 48.326 1.266 48.362 ;
      RECT 1.214 49.526 1.266 49.562 ;
      RECT 1.214 50.726 1.266 50.762 ;
      RECT 1.214 51.926 1.266 51.962 ;
      RECT 1.214 53.126 1.266 53.162 ;
      RECT 1.214 54.326 1.266 54.362 ;
      RECT 1.214 55.526 1.266 55.562 ;
      RECT 1.214 56.726 1.266 56.762 ;
      RECT 1.214 57.926 1.266 57.962 ;
      RECT 1.214 59.126 1.266 59.162 ;
      RECT 1.214 60.326 1.266 60.362 ;
      RECT 1.214 61.526 1.266 61.562 ;
      RECT 1.214 62.726 1.266 62.762 ;
      RECT 1.214 63.926 1.266 63.962 ;
      RECT 1.214 65.126 1.266 65.162 ;
      RECT 1.214 66.326 1.266 66.362 ;
      RECT 1.214 67.526 1.266 67.562 ;
      RECT 1.214 68.726 1.266 68.762 ;
      RECT 1.214 69.926 1.266 69.962 ;
      RECT 1.214 71.126 1.266 71.162 ;
      RECT 1.294 1.558 1.346 1.594 ;
      RECT 1.294 2.758 1.346 2.794 ;
      RECT 1.294 3.958 1.346 3.994 ;
      RECT 1.294 5.158 1.346 5.194 ;
      RECT 1.294 6.358 1.346 6.394 ;
      RECT 1.294 7.558 1.346 7.594 ;
      RECT 1.294 8.758 1.346 8.794 ;
      RECT 1.294 9.958 1.346 9.994 ;
      RECT 1.294 11.158 1.346 11.194 ;
      RECT 1.294 12.358 1.346 12.394 ;
      RECT 1.294 13.558 1.346 13.594 ;
      RECT 1.294 14.758 1.346 14.794 ;
      RECT 1.294 15.958 1.346 15.994 ;
      RECT 1.294 17.158 1.346 17.194 ;
      RECT 1.294 18.358 1.346 18.394 ;
      RECT 1.294 19.558 1.346 19.594 ;
      RECT 1.294 20.758 1.346 20.794 ;
      RECT 1.294 21.958 1.346 21.994 ;
      RECT 1.294 23.158 1.346 23.194 ;
      RECT 1.294 24.358 1.346 24.394 ;
      RECT 1.294 25.558 1.346 25.594 ;
      RECT 1.294 26.758 1.346 26.794 ;
      RECT 1.294 27.958 1.346 27.994 ;
      RECT 1.294 29.158 1.346 29.194 ;
      RECT 1.294 30.358 1.346 30.394 ;
      RECT 1.294 31.558 1.346 31.594 ;
      RECT 1.294 33.342 1.346 33.378 ;
      RECT 1.294 33.582 1.346 33.618 ;
      RECT 1.294 37.902 1.346 37.938 ;
      RECT 1.294 38.142 1.346 38.178 ;
      RECT 1.294 40.678 1.346 40.714 ;
      RECT 1.294 41.878 1.346 41.914 ;
      RECT 1.294 43.078 1.346 43.114 ;
      RECT 1.294 44.278 1.346 44.314 ;
      RECT 1.294 45.478 1.346 45.514 ;
      RECT 1.294 46.678 1.346 46.714 ;
      RECT 1.294 47.878 1.346 47.914 ;
      RECT 1.294 49.078 1.346 49.114 ;
      RECT 1.294 50.278 1.346 50.314 ;
      RECT 1.294 51.478 1.346 51.514 ;
      RECT 1.294 52.678 1.346 52.714 ;
      RECT 1.294 53.878 1.346 53.914 ;
      RECT 1.294 55.078 1.346 55.114 ;
      RECT 1.294 56.278 1.346 56.314 ;
      RECT 1.294 57.478 1.346 57.514 ;
      RECT 1.294 58.678 1.346 58.714 ;
      RECT 1.294 59.878 1.346 59.914 ;
      RECT 1.294 61.078 1.346 61.114 ;
      RECT 1.294 62.278 1.346 62.314 ;
      RECT 1.294 63.478 1.346 63.514 ;
      RECT 1.294 64.678 1.346 64.714 ;
      RECT 1.294 65.878 1.346 65.914 ;
      RECT 1.294 67.078 1.346 67.114 ;
      RECT 1.294 68.278 1.346 68.314 ;
      RECT 1.294 69.478 1.346 69.514 ;
      RECT 1.294 70.678 1.346 70.714 ;
      RECT 1.294 71.878 1.346 71.914 ;
      RECT 1.374 0.281 1.426 0.317 ;
      RECT 1.374 72.403 1.426 72.439 ;
      RECT 1.454 0.806 1.506 0.842 ;
      RECT 1.454 2.006 1.506 2.042 ;
      RECT 1.454 3.206 1.506 3.242 ;
      RECT 1.454 4.406 1.506 4.442 ;
      RECT 1.454 5.606 1.506 5.642 ;
      RECT 1.454 6.806 1.506 6.842 ;
      RECT 1.454 8.006 1.506 8.042 ;
      RECT 1.454 9.206 1.506 9.242 ;
      RECT 1.454 10.406 1.506 10.442 ;
      RECT 1.454 11.606 1.506 11.642 ;
      RECT 1.454 12.806 1.506 12.842 ;
      RECT 1.454 14.006 1.506 14.042 ;
      RECT 1.454 15.206 1.506 15.242 ;
      RECT 1.454 16.406 1.506 16.442 ;
      RECT 1.454 17.606 1.506 17.642 ;
      RECT 1.454 18.806 1.506 18.842 ;
      RECT 1.454 20.006 1.506 20.042 ;
      RECT 1.454 21.206 1.506 21.242 ;
      RECT 1.454 22.406 1.506 22.442 ;
      RECT 1.454 23.606 1.506 23.642 ;
      RECT 1.454 24.806 1.506 24.842 ;
      RECT 1.454 26.006 1.506 26.042 ;
      RECT 1.454 27.206 1.506 27.242 ;
      RECT 1.454 28.406 1.506 28.442 ;
      RECT 1.454 29.606 1.506 29.642 ;
      RECT 1.454 30.806 1.506 30.842 ;
      RECT 1.454 32.622 1.506 32.658 ;
      RECT 1.454 32.862 1.506 32.898 ;
      RECT 1.454 38.622 1.506 38.658 ;
      RECT 1.454 38.862 1.506 38.898 ;
      RECT 1.454 39.926 1.506 39.962 ;
      RECT 1.454 41.126 1.506 41.162 ;
      RECT 1.454 42.326 1.506 42.362 ;
      RECT 1.454 43.526 1.506 43.562 ;
      RECT 1.454 44.726 1.506 44.762 ;
      RECT 1.454 45.926 1.506 45.962 ;
      RECT 1.454 47.126 1.506 47.162 ;
      RECT 1.454 48.326 1.506 48.362 ;
      RECT 1.454 49.526 1.506 49.562 ;
      RECT 1.454 50.726 1.506 50.762 ;
      RECT 1.454 51.926 1.506 51.962 ;
      RECT 1.454 53.126 1.506 53.162 ;
      RECT 1.454 54.326 1.506 54.362 ;
      RECT 1.454 55.526 1.506 55.562 ;
      RECT 1.454 56.726 1.506 56.762 ;
      RECT 1.454 57.926 1.506 57.962 ;
      RECT 1.454 59.126 1.506 59.162 ;
      RECT 1.454 60.326 1.506 60.362 ;
      RECT 1.454 61.526 1.506 61.562 ;
      RECT 1.454 62.726 1.506 62.762 ;
      RECT 1.454 63.926 1.506 63.962 ;
      RECT 1.454 65.126 1.506 65.162 ;
      RECT 1.454 66.326 1.506 66.362 ;
      RECT 1.454 67.526 1.506 67.562 ;
      RECT 1.454 68.726 1.506 68.762 ;
      RECT 1.454 69.926 1.506 69.962 ;
      RECT 1.454 71.126 1.506 71.162 ;
      RECT 1.534 1.558 1.586 1.594 ;
      RECT 1.534 2.758 1.586 2.794 ;
      RECT 1.534 3.958 1.586 3.994 ;
      RECT 1.534 5.158 1.586 5.194 ;
      RECT 1.534 6.358 1.586 6.394 ;
      RECT 1.534 7.558 1.586 7.594 ;
      RECT 1.534 8.758 1.586 8.794 ;
      RECT 1.534 9.958 1.586 9.994 ;
      RECT 1.534 11.158 1.586 11.194 ;
      RECT 1.534 12.358 1.586 12.394 ;
      RECT 1.534 13.558 1.586 13.594 ;
      RECT 1.534 14.758 1.586 14.794 ;
      RECT 1.534 15.958 1.586 15.994 ;
      RECT 1.534 17.158 1.586 17.194 ;
      RECT 1.534 18.358 1.586 18.394 ;
      RECT 1.534 19.558 1.586 19.594 ;
      RECT 1.534 20.758 1.586 20.794 ;
      RECT 1.534 21.958 1.586 21.994 ;
      RECT 1.534 23.158 1.586 23.194 ;
      RECT 1.534 24.358 1.586 24.394 ;
      RECT 1.534 25.558 1.586 25.594 ;
      RECT 1.534 26.758 1.586 26.794 ;
      RECT 1.534 27.958 1.586 27.994 ;
      RECT 1.534 29.158 1.586 29.194 ;
      RECT 1.534 30.358 1.586 30.394 ;
      RECT 1.534 31.558 1.586 31.594 ;
      RECT 1.534 33.342 1.586 33.378 ;
      RECT 1.534 33.582 1.586 33.618 ;
      RECT 1.534 37.902 1.586 37.938 ;
      RECT 1.534 38.142 1.586 38.178 ;
      RECT 1.534 40.678 1.586 40.714 ;
      RECT 1.534 41.878 1.586 41.914 ;
      RECT 1.534 43.078 1.586 43.114 ;
      RECT 1.534 44.278 1.586 44.314 ;
      RECT 1.534 45.478 1.586 45.514 ;
      RECT 1.534 46.678 1.586 46.714 ;
      RECT 1.534 47.878 1.586 47.914 ;
      RECT 1.534 49.078 1.586 49.114 ;
      RECT 1.534 50.278 1.586 50.314 ;
      RECT 1.534 51.478 1.586 51.514 ;
      RECT 1.534 52.678 1.586 52.714 ;
      RECT 1.534 53.878 1.586 53.914 ;
      RECT 1.534 55.078 1.586 55.114 ;
      RECT 1.534 56.278 1.586 56.314 ;
      RECT 1.534 57.478 1.586 57.514 ;
      RECT 1.534 58.678 1.586 58.714 ;
      RECT 1.534 59.878 1.586 59.914 ;
      RECT 1.534 61.078 1.586 61.114 ;
      RECT 1.534 62.278 1.586 62.314 ;
      RECT 1.534 63.478 1.586 63.514 ;
      RECT 1.534 64.678 1.586 64.714 ;
      RECT 1.534 65.878 1.586 65.914 ;
      RECT 1.534 67.078 1.586 67.114 ;
      RECT 1.534 68.278 1.586 68.314 ;
      RECT 1.534 69.478 1.586 69.514 ;
      RECT 1.534 70.678 1.586 70.714 ;
      RECT 1.534 71.878 1.586 71.914 ;
      RECT 1.614 0.806 1.666 0.842 ;
      RECT 1.614 2.006 1.666 2.042 ;
      RECT 1.614 3.206 1.666 3.242 ;
      RECT 1.614 4.406 1.666 4.442 ;
      RECT 1.614 5.606 1.666 5.642 ;
      RECT 1.614 6.806 1.666 6.842 ;
      RECT 1.614 8.006 1.666 8.042 ;
      RECT 1.614 9.206 1.666 9.242 ;
      RECT 1.614 10.406 1.666 10.442 ;
      RECT 1.614 11.606 1.666 11.642 ;
      RECT 1.614 12.806 1.666 12.842 ;
      RECT 1.614 14.006 1.666 14.042 ;
      RECT 1.614 15.206 1.666 15.242 ;
      RECT 1.614 16.406 1.666 16.442 ;
      RECT 1.614 17.606 1.666 17.642 ;
      RECT 1.614 18.806 1.666 18.842 ;
      RECT 1.614 20.006 1.666 20.042 ;
      RECT 1.614 21.206 1.666 21.242 ;
      RECT 1.614 22.406 1.666 22.442 ;
      RECT 1.614 23.606 1.666 23.642 ;
      RECT 1.614 24.806 1.666 24.842 ;
      RECT 1.614 26.006 1.666 26.042 ;
      RECT 1.614 27.206 1.666 27.242 ;
      RECT 1.614 28.406 1.666 28.442 ;
      RECT 1.614 29.606 1.666 29.642 ;
      RECT 1.614 30.806 1.666 30.842 ;
      RECT 1.614 32.622 1.666 32.658 ;
      RECT 1.614 32.862 1.666 32.898 ;
      RECT 1.614 38.622 1.666 38.658 ;
      RECT 1.614 38.862 1.666 38.898 ;
      RECT 1.614 39.926 1.666 39.962 ;
      RECT 1.614 41.126 1.666 41.162 ;
      RECT 1.614 42.326 1.666 42.362 ;
      RECT 1.614 43.526 1.666 43.562 ;
      RECT 1.614 44.726 1.666 44.762 ;
      RECT 1.614 45.926 1.666 45.962 ;
      RECT 1.614 47.126 1.666 47.162 ;
      RECT 1.614 48.326 1.666 48.362 ;
      RECT 1.614 49.526 1.666 49.562 ;
      RECT 1.614 50.726 1.666 50.762 ;
      RECT 1.614 51.926 1.666 51.962 ;
      RECT 1.614 53.126 1.666 53.162 ;
      RECT 1.614 54.326 1.666 54.362 ;
      RECT 1.614 55.526 1.666 55.562 ;
      RECT 1.614 56.726 1.666 56.762 ;
      RECT 1.614 57.926 1.666 57.962 ;
      RECT 1.614 59.126 1.666 59.162 ;
      RECT 1.614 60.326 1.666 60.362 ;
      RECT 1.614 61.526 1.666 61.562 ;
      RECT 1.614 62.726 1.666 62.762 ;
      RECT 1.614 63.926 1.666 63.962 ;
      RECT 1.614 65.126 1.666 65.162 ;
      RECT 1.614 66.326 1.666 66.362 ;
      RECT 1.614 67.526 1.666 67.562 ;
      RECT 1.614 68.726 1.666 68.762 ;
      RECT 1.614 69.926 1.666 69.962 ;
      RECT 1.614 71.126 1.666 71.162 ;
      RECT 1.694 1.558 1.746 1.594 ;
      RECT 1.694 2.758 1.746 2.794 ;
      RECT 1.694 3.958 1.746 3.994 ;
      RECT 1.694 5.158 1.746 5.194 ;
      RECT 1.694 6.358 1.746 6.394 ;
      RECT 1.694 7.558 1.746 7.594 ;
      RECT 1.694 8.758 1.746 8.794 ;
      RECT 1.694 9.958 1.746 9.994 ;
      RECT 1.694 11.158 1.746 11.194 ;
      RECT 1.694 12.358 1.746 12.394 ;
      RECT 1.694 13.558 1.746 13.594 ;
      RECT 1.694 14.758 1.746 14.794 ;
      RECT 1.694 15.958 1.746 15.994 ;
      RECT 1.694 17.158 1.746 17.194 ;
      RECT 1.694 18.358 1.746 18.394 ;
      RECT 1.694 19.558 1.746 19.594 ;
      RECT 1.694 20.758 1.746 20.794 ;
      RECT 1.694 21.958 1.746 21.994 ;
      RECT 1.694 23.158 1.746 23.194 ;
      RECT 1.694 24.358 1.746 24.394 ;
      RECT 1.694 25.558 1.746 25.594 ;
      RECT 1.694 26.758 1.746 26.794 ;
      RECT 1.694 27.958 1.746 27.994 ;
      RECT 1.694 29.158 1.746 29.194 ;
      RECT 1.694 30.358 1.746 30.394 ;
      RECT 1.694 31.558 1.746 31.594 ;
      RECT 1.694 33.342 1.746 33.378 ;
      RECT 1.694 33.582 1.746 33.618 ;
      RECT 1.694 37.902 1.746 37.938 ;
      RECT 1.694 38.142 1.746 38.178 ;
      RECT 1.694 40.678 1.746 40.714 ;
      RECT 1.694 41.878 1.746 41.914 ;
      RECT 1.694 43.078 1.746 43.114 ;
      RECT 1.694 44.278 1.746 44.314 ;
      RECT 1.694 45.478 1.746 45.514 ;
      RECT 1.694 46.678 1.746 46.714 ;
      RECT 1.694 47.878 1.746 47.914 ;
      RECT 1.694 49.078 1.746 49.114 ;
      RECT 1.694 50.278 1.746 50.314 ;
      RECT 1.694 51.478 1.746 51.514 ;
      RECT 1.694 52.678 1.746 52.714 ;
      RECT 1.694 53.878 1.746 53.914 ;
      RECT 1.694 55.078 1.746 55.114 ;
      RECT 1.694 56.278 1.746 56.314 ;
      RECT 1.694 57.478 1.746 57.514 ;
      RECT 1.694 58.678 1.746 58.714 ;
      RECT 1.694 59.878 1.746 59.914 ;
      RECT 1.694 61.078 1.746 61.114 ;
      RECT 1.694 62.278 1.746 62.314 ;
      RECT 1.694 63.478 1.746 63.514 ;
      RECT 1.694 64.678 1.746 64.714 ;
      RECT 1.694 65.878 1.746 65.914 ;
      RECT 1.694 67.078 1.746 67.114 ;
      RECT 1.694 68.278 1.746 68.314 ;
      RECT 1.694 69.478 1.746 69.514 ;
      RECT 1.694 70.678 1.746 70.714 ;
      RECT 1.694 71.878 1.746 71.914 ;
      RECT 1.774 0.281 1.826 0.317 ;
      RECT 1.774 72.403 1.826 72.439 ;
      RECT 1.854 0.806 1.906 0.842 ;
      RECT 1.854 2.006 1.906 2.042 ;
      RECT 1.854 3.206 1.906 3.242 ;
      RECT 1.854 4.406 1.906 4.442 ;
      RECT 1.854 5.606 1.906 5.642 ;
      RECT 1.854 6.806 1.906 6.842 ;
      RECT 1.854 8.006 1.906 8.042 ;
      RECT 1.854 9.206 1.906 9.242 ;
      RECT 1.854 10.406 1.906 10.442 ;
      RECT 1.854 11.606 1.906 11.642 ;
      RECT 1.854 12.806 1.906 12.842 ;
      RECT 1.854 14.006 1.906 14.042 ;
      RECT 1.854 15.206 1.906 15.242 ;
      RECT 1.854 16.406 1.906 16.442 ;
      RECT 1.854 17.606 1.906 17.642 ;
      RECT 1.854 18.806 1.906 18.842 ;
      RECT 1.854 20.006 1.906 20.042 ;
      RECT 1.854 21.206 1.906 21.242 ;
      RECT 1.854 22.406 1.906 22.442 ;
      RECT 1.854 23.606 1.906 23.642 ;
      RECT 1.854 24.806 1.906 24.842 ;
      RECT 1.854 26.006 1.906 26.042 ;
      RECT 1.854 27.206 1.906 27.242 ;
      RECT 1.854 28.406 1.906 28.442 ;
      RECT 1.854 29.606 1.906 29.642 ;
      RECT 1.854 30.806 1.906 30.842 ;
      RECT 1.854 32.622 1.906 32.658 ;
      RECT 1.854 32.862 1.906 32.898 ;
      RECT 1.854 34.302 1.906 34.338 ;
      RECT 1.854 34.782 1.906 34.818 ;
      RECT 1.854 36.702 1.906 36.738 ;
      RECT 1.854 37.182 1.906 37.218 ;
      RECT 1.854 38.622 1.906 38.658 ;
      RECT 1.854 38.862 1.906 38.898 ;
      RECT 1.854 39.926 1.906 39.962 ;
      RECT 1.854 41.126 1.906 41.162 ;
      RECT 1.854 42.326 1.906 42.362 ;
      RECT 1.854 43.526 1.906 43.562 ;
      RECT 1.854 44.726 1.906 44.762 ;
      RECT 1.854 45.926 1.906 45.962 ;
      RECT 1.854 47.126 1.906 47.162 ;
      RECT 1.854 48.326 1.906 48.362 ;
      RECT 1.854 49.526 1.906 49.562 ;
      RECT 1.854 50.726 1.906 50.762 ;
      RECT 1.854 51.926 1.906 51.962 ;
      RECT 1.854 53.126 1.906 53.162 ;
      RECT 1.854 54.326 1.906 54.362 ;
      RECT 1.854 55.526 1.906 55.562 ;
      RECT 1.854 56.726 1.906 56.762 ;
      RECT 1.854 57.926 1.906 57.962 ;
      RECT 1.854 59.126 1.906 59.162 ;
      RECT 1.854 60.326 1.906 60.362 ;
      RECT 1.854 61.526 1.906 61.562 ;
      RECT 1.854 62.726 1.906 62.762 ;
      RECT 1.854 63.926 1.906 63.962 ;
      RECT 1.854 65.126 1.906 65.162 ;
      RECT 1.854 66.326 1.906 66.362 ;
      RECT 1.854 67.526 1.906 67.562 ;
      RECT 1.854 68.726 1.906 68.762 ;
      RECT 1.854 69.926 1.906 69.962 ;
      RECT 1.854 71.126 1.906 71.162 ;
      RECT 1.934 1.558 1.986 1.594 ;
      RECT 1.934 2.758 1.986 2.794 ;
      RECT 1.934 3.958 1.986 3.994 ;
      RECT 1.934 5.158 1.986 5.194 ;
      RECT 1.934 6.358 1.986 6.394 ;
      RECT 1.934 7.558 1.986 7.594 ;
      RECT 1.934 8.758 1.986 8.794 ;
      RECT 1.934 9.958 1.986 9.994 ;
      RECT 1.934 11.158 1.986 11.194 ;
      RECT 1.934 12.358 1.986 12.394 ;
      RECT 1.934 13.558 1.986 13.594 ;
      RECT 1.934 14.758 1.986 14.794 ;
      RECT 1.934 15.958 1.986 15.994 ;
      RECT 1.934 17.158 1.986 17.194 ;
      RECT 1.934 18.358 1.986 18.394 ;
      RECT 1.934 19.558 1.986 19.594 ;
      RECT 1.934 20.758 1.986 20.794 ;
      RECT 1.934 21.958 1.986 21.994 ;
      RECT 1.934 23.158 1.986 23.194 ;
      RECT 1.934 24.358 1.986 24.394 ;
      RECT 1.934 25.558 1.986 25.594 ;
      RECT 1.934 26.758 1.986 26.794 ;
      RECT 1.934 27.958 1.986 27.994 ;
      RECT 1.934 29.158 1.986 29.194 ;
      RECT 1.934 30.358 1.986 30.394 ;
      RECT 1.934 31.558 1.986 31.594 ;
      RECT 1.934 33.342 1.986 33.378 ;
      RECT 1.934 33.582 1.986 33.618 ;
      RECT 1.934 37.902 1.986 37.938 ;
      RECT 1.934 38.142 1.986 38.178 ;
      RECT 1.934 40.678 1.986 40.714 ;
      RECT 1.934 41.878 1.986 41.914 ;
      RECT 1.934 43.078 1.986 43.114 ;
      RECT 1.934 44.278 1.986 44.314 ;
      RECT 1.934 45.478 1.986 45.514 ;
      RECT 1.934 46.678 1.986 46.714 ;
      RECT 1.934 47.878 1.986 47.914 ;
      RECT 1.934 49.078 1.986 49.114 ;
      RECT 1.934 50.278 1.986 50.314 ;
      RECT 1.934 51.478 1.986 51.514 ;
      RECT 1.934 52.678 1.986 52.714 ;
      RECT 1.934 53.878 1.986 53.914 ;
      RECT 1.934 55.078 1.986 55.114 ;
      RECT 1.934 56.278 1.986 56.314 ;
      RECT 1.934 57.478 1.986 57.514 ;
      RECT 1.934 58.678 1.986 58.714 ;
      RECT 1.934 59.878 1.986 59.914 ;
      RECT 1.934 61.078 1.986 61.114 ;
      RECT 1.934 62.278 1.986 62.314 ;
      RECT 1.934 63.478 1.986 63.514 ;
      RECT 1.934 64.678 1.986 64.714 ;
      RECT 1.934 65.878 1.986 65.914 ;
      RECT 1.934 67.078 1.986 67.114 ;
      RECT 1.934 68.278 1.986 68.314 ;
      RECT 1.934 69.478 1.986 69.514 ;
      RECT 1.934 70.678 1.986 70.714 ;
      RECT 1.934 71.878 1.986 71.914 ;
      RECT 2.014 0.806 2.066 0.842 ;
      RECT 2.014 2.006 2.066 2.042 ;
      RECT 2.014 3.206 2.066 3.242 ;
      RECT 2.014 4.406 2.066 4.442 ;
      RECT 2.014 5.606 2.066 5.642 ;
      RECT 2.014 6.806 2.066 6.842 ;
      RECT 2.014 8.006 2.066 8.042 ;
      RECT 2.014 9.206 2.066 9.242 ;
      RECT 2.014 10.406 2.066 10.442 ;
      RECT 2.014 11.606 2.066 11.642 ;
      RECT 2.014 12.806 2.066 12.842 ;
      RECT 2.014 14.006 2.066 14.042 ;
      RECT 2.014 15.206 2.066 15.242 ;
      RECT 2.014 16.406 2.066 16.442 ;
      RECT 2.014 17.606 2.066 17.642 ;
      RECT 2.014 18.806 2.066 18.842 ;
      RECT 2.014 20.006 2.066 20.042 ;
      RECT 2.014 21.206 2.066 21.242 ;
      RECT 2.014 22.406 2.066 22.442 ;
      RECT 2.014 23.606 2.066 23.642 ;
      RECT 2.014 24.806 2.066 24.842 ;
      RECT 2.014 26.006 2.066 26.042 ;
      RECT 2.014 27.206 2.066 27.242 ;
      RECT 2.014 28.406 2.066 28.442 ;
      RECT 2.014 29.606 2.066 29.642 ;
      RECT 2.014 30.806 2.066 30.842 ;
      RECT 2.014 32.622 2.066 32.658 ;
      RECT 2.014 32.862 2.066 32.898 ;
      RECT 2.014 38.622 2.066 38.658 ;
      RECT 2.014 38.862 2.066 38.898 ;
      RECT 2.014 39.926 2.066 39.962 ;
      RECT 2.014 41.126 2.066 41.162 ;
      RECT 2.014 42.326 2.066 42.362 ;
      RECT 2.014 43.526 2.066 43.562 ;
      RECT 2.014 44.726 2.066 44.762 ;
      RECT 2.014 45.926 2.066 45.962 ;
      RECT 2.014 47.126 2.066 47.162 ;
      RECT 2.014 48.326 2.066 48.362 ;
      RECT 2.014 49.526 2.066 49.562 ;
      RECT 2.014 50.726 2.066 50.762 ;
      RECT 2.014 51.926 2.066 51.962 ;
      RECT 2.014 53.126 2.066 53.162 ;
      RECT 2.014 54.326 2.066 54.362 ;
      RECT 2.014 55.526 2.066 55.562 ;
      RECT 2.014 56.726 2.066 56.762 ;
      RECT 2.014 57.926 2.066 57.962 ;
      RECT 2.014 59.126 2.066 59.162 ;
      RECT 2.014 60.326 2.066 60.362 ;
      RECT 2.014 61.526 2.066 61.562 ;
      RECT 2.014 62.726 2.066 62.762 ;
      RECT 2.014 63.926 2.066 63.962 ;
      RECT 2.014 65.126 2.066 65.162 ;
      RECT 2.014 66.326 2.066 66.362 ;
      RECT 2.014 67.526 2.066 67.562 ;
      RECT 2.014 68.726 2.066 68.762 ;
      RECT 2.014 69.926 2.066 69.962 ;
      RECT 2.014 71.126 2.066 71.162 ;
      RECT 2.094 1.558 2.146 1.594 ;
      RECT 2.094 2.758 2.146 2.794 ;
      RECT 2.094 3.958 2.146 3.994 ;
      RECT 2.094 5.158 2.146 5.194 ;
      RECT 2.094 6.358 2.146 6.394 ;
      RECT 2.094 7.558 2.146 7.594 ;
      RECT 2.094 8.758 2.146 8.794 ;
      RECT 2.094 9.958 2.146 9.994 ;
      RECT 2.094 11.158 2.146 11.194 ;
      RECT 2.094 12.358 2.146 12.394 ;
      RECT 2.094 13.558 2.146 13.594 ;
      RECT 2.094 14.758 2.146 14.794 ;
      RECT 2.094 15.958 2.146 15.994 ;
      RECT 2.094 17.158 2.146 17.194 ;
      RECT 2.094 18.358 2.146 18.394 ;
      RECT 2.094 19.558 2.146 19.594 ;
      RECT 2.094 20.758 2.146 20.794 ;
      RECT 2.094 21.958 2.146 21.994 ;
      RECT 2.094 23.158 2.146 23.194 ;
      RECT 2.094 24.358 2.146 24.394 ;
      RECT 2.094 25.558 2.146 25.594 ;
      RECT 2.094 26.758 2.146 26.794 ;
      RECT 2.094 27.958 2.146 27.994 ;
      RECT 2.094 29.158 2.146 29.194 ;
      RECT 2.094 30.358 2.146 30.394 ;
      RECT 2.094 31.558 2.146 31.594 ;
      RECT 2.094 33.342 2.146 33.378 ;
      RECT 2.094 33.582 2.146 33.618 ;
      RECT 2.094 37.902 2.146 37.938 ;
      RECT 2.094 38.142 2.146 38.178 ;
      RECT 2.094 40.678 2.146 40.714 ;
      RECT 2.094 41.878 2.146 41.914 ;
      RECT 2.094 43.078 2.146 43.114 ;
      RECT 2.094 44.278 2.146 44.314 ;
      RECT 2.094 45.478 2.146 45.514 ;
      RECT 2.094 46.678 2.146 46.714 ;
      RECT 2.094 47.878 2.146 47.914 ;
      RECT 2.094 49.078 2.146 49.114 ;
      RECT 2.094 50.278 2.146 50.314 ;
      RECT 2.094 51.478 2.146 51.514 ;
      RECT 2.094 52.678 2.146 52.714 ;
      RECT 2.094 53.878 2.146 53.914 ;
      RECT 2.094 55.078 2.146 55.114 ;
      RECT 2.094 56.278 2.146 56.314 ;
      RECT 2.094 57.478 2.146 57.514 ;
      RECT 2.094 58.678 2.146 58.714 ;
      RECT 2.094 59.878 2.146 59.914 ;
      RECT 2.094 61.078 2.146 61.114 ;
      RECT 2.094 62.278 2.146 62.314 ;
      RECT 2.094 63.478 2.146 63.514 ;
      RECT 2.094 64.678 2.146 64.714 ;
      RECT 2.094 65.878 2.146 65.914 ;
      RECT 2.094 67.078 2.146 67.114 ;
      RECT 2.094 68.278 2.146 68.314 ;
      RECT 2.094 69.478 2.146 69.514 ;
      RECT 2.094 70.678 2.146 70.714 ;
      RECT 2.094 71.878 2.146 71.914 ;
      RECT 2.174 0.281 2.226 0.317 ;
      RECT 2.174 72.403 2.226 72.439 ;
      RECT 2.254 0.806 2.306 0.842 ;
      RECT 2.254 2.006 2.306 2.042 ;
      RECT 2.254 3.206 2.306 3.242 ;
      RECT 2.254 4.406 2.306 4.442 ;
      RECT 2.254 5.606 2.306 5.642 ;
      RECT 2.254 6.806 2.306 6.842 ;
      RECT 2.254 8.006 2.306 8.042 ;
      RECT 2.254 9.206 2.306 9.242 ;
      RECT 2.254 10.406 2.306 10.442 ;
      RECT 2.254 11.606 2.306 11.642 ;
      RECT 2.254 12.806 2.306 12.842 ;
      RECT 2.254 14.006 2.306 14.042 ;
      RECT 2.254 15.206 2.306 15.242 ;
      RECT 2.254 16.406 2.306 16.442 ;
      RECT 2.254 17.606 2.306 17.642 ;
      RECT 2.254 18.806 2.306 18.842 ;
      RECT 2.254 20.006 2.306 20.042 ;
      RECT 2.254 21.206 2.306 21.242 ;
      RECT 2.254 22.406 2.306 22.442 ;
      RECT 2.254 23.606 2.306 23.642 ;
      RECT 2.254 24.806 2.306 24.842 ;
      RECT 2.254 26.006 2.306 26.042 ;
      RECT 2.254 27.206 2.306 27.242 ;
      RECT 2.254 28.406 2.306 28.442 ;
      RECT 2.254 29.606 2.306 29.642 ;
      RECT 2.254 30.806 2.306 30.842 ;
      RECT 2.254 32.622 2.306 32.658 ;
      RECT 2.254 32.862 2.306 32.898 ;
      RECT 2.254 38.622 2.306 38.658 ;
      RECT 2.254 38.862 2.306 38.898 ;
      RECT 2.254 39.926 2.306 39.962 ;
      RECT 2.254 41.126 2.306 41.162 ;
      RECT 2.254 42.326 2.306 42.362 ;
      RECT 2.254 43.526 2.306 43.562 ;
      RECT 2.254 44.726 2.306 44.762 ;
      RECT 2.254 45.926 2.306 45.962 ;
      RECT 2.254 47.126 2.306 47.162 ;
      RECT 2.254 48.326 2.306 48.362 ;
      RECT 2.254 49.526 2.306 49.562 ;
      RECT 2.254 50.726 2.306 50.762 ;
      RECT 2.254 51.926 2.306 51.962 ;
      RECT 2.254 53.126 2.306 53.162 ;
      RECT 2.254 54.326 2.306 54.362 ;
      RECT 2.254 55.526 2.306 55.562 ;
      RECT 2.254 56.726 2.306 56.762 ;
      RECT 2.254 57.926 2.306 57.962 ;
      RECT 2.254 59.126 2.306 59.162 ;
      RECT 2.254 60.326 2.306 60.362 ;
      RECT 2.254 61.526 2.306 61.562 ;
      RECT 2.254 62.726 2.306 62.762 ;
      RECT 2.254 63.926 2.306 63.962 ;
      RECT 2.254 65.126 2.306 65.162 ;
      RECT 2.254 66.326 2.306 66.362 ;
      RECT 2.254 67.526 2.306 67.562 ;
      RECT 2.254 68.726 2.306 68.762 ;
      RECT 2.254 69.926 2.306 69.962 ;
      RECT 2.254 71.126 2.306 71.162 ;
      RECT 2.334 1.558 2.386 1.594 ;
      RECT 2.334 2.758 2.386 2.794 ;
      RECT 2.334 3.958 2.386 3.994 ;
      RECT 2.334 5.158 2.386 5.194 ;
      RECT 2.334 6.358 2.386 6.394 ;
      RECT 2.334 7.558 2.386 7.594 ;
      RECT 2.334 8.758 2.386 8.794 ;
      RECT 2.334 9.958 2.386 9.994 ;
      RECT 2.334 11.158 2.386 11.194 ;
      RECT 2.334 12.358 2.386 12.394 ;
      RECT 2.334 13.558 2.386 13.594 ;
      RECT 2.334 14.758 2.386 14.794 ;
      RECT 2.334 15.958 2.386 15.994 ;
      RECT 2.334 17.158 2.386 17.194 ;
      RECT 2.334 18.358 2.386 18.394 ;
      RECT 2.334 19.558 2.386 19.594 ;
      RECT 2.334 20.758 2.386 20.794 ;
      RECT 2.334 21.958 2.386 21.994 ;
      RECT 2.334 23.158 2.386 23.194 ;
      RECT 2.334 24.358 2.386 24.394 ;
      RECT 2.334 25.558 2.386 25.594 ;
      RECT 2.334 26.758 2.386 26.794 ;
      RECT 2.334 27.958 2.386 27.994 ;
      RECT 2.334 29.158 2.386 29.194 ;
      RECT 2.334 30.358 2.386 30.394 ;
      RECT 2.334 31.558 2.386 31.594 ;
      RECT 2.334 33.342 2.386 33.378 ;
      RECT 2.334 33.582 2.386 33.618 ;
      RECT 2.334 37.902 2.386 37.938 ;
      RECT 2.334 38.142 2.386 38.178 ;
      RECT 2.334 40.678 2.386 40.714 ;
      RECT 2.334 41.878 2.386 41.914 ;
      RECT 2.334 43.078 2.386 43.114 ;
      RECT 2.334 44.278 2.386 44.314 ;
      RECT 2.334 45.478 2.386 45.514 ;
      RECT 2.334 46.678 2.386 46.714 ;
      RECT 2.334 47.878 2.386 47.914 ;
      RECT 2.334 49.078 2.386 49.114 ;
      RECT 2.334 50.278 2.386 50.314 ;
      RECT 2.334 51.478 2.386 51.514 ;
      RECT 2.334 52.678 2.386 52.714 ;
      RECT 2.334 53.878 2.386 53.914 ;
      RECT 2.334 55.078 2.386 55.114 ;
      RECT 2.334 56.278 2.386 56.314 ;
      RECT 2.334 57.478 2.386 57.514 ;
      RECT 2.334 58.678 2.386 58.714 ;
      RECT 2.334 59.878 2.386 59.914 ;
      RECT 2.334 61.078 2.386 61.114 ;
      RECT 2.334 62.278 2.386 62.314 ;
      RECT 2.334 63.478 2.386 63.514 ;
      RECT 2.334 64.678 2.386 64.714 ;
      RECT 2.334 65.878 2.386 65.914 ;
      RECT 2.334 67.078 2.386 67.114 ;
      RECT 2.334 68.278 2.386 68.314 ;
      RECT 2.334 69.478 2.386 69.514 ;
      RECT 2.334 70.678 2.386 70.714 ;
      RECT 2.334 71.878 2.386 71.914 ;
      RECT 2.414 0.806 2.466 0.842 ;
      RECT 2.414 2.006 2.466 2.042 ;
      RECT 2.414 3.206 2.466 3.242 ;
      RECT 2.414 4.406 2.466 4.442 ;
      RECT 2.414 5.606 2.466 5.642 ;
      RECT 2.414 6.806 2.466 6.842 ;
      RECT 2.414 8.006 2.466 8.042 ;
      RECT 2.414 9.206 2.466 9.242 ;
      RECT 2.414 10.406 2.466 10.442 ;
      RECT 2.414 11.606 2.466 11.642 ;
      RECT 2.414 12.806 2.466 12.842 ;
      RECT 2.414 14.006 2.466 14.042 ;
      RECT 2.414 15.206 2.466 15.242 ;
      RECT 2.414 16.406 2.466 16.442 ;
      RECT 2.414 17.606 2.466 17.642 ;
      RECT 2.414 18.806 2.466 18.842 ;
      RECT 2.414 20.006 2.466 20.042 ;
      RECT 2.414 21.206 2.466 21.242 ;
      RECT 2.414 22.406 2.466 22.442 ;
      RECT 2.414 23.606 2.466 23.642 ;
      RECT 2.414 24.806 2.466 24.842 ;
      RECT 2.414 26.006 2.466 26.042 ;
      RECT 2.414 27.206 2.466 27.242 ;
      RECT 2.414 28.406 2.466 28.442 ;
      RECT 2.414 29.606 2.466 29.642 ;
      RECT 2.414 30.806 2.466 30.842 ;
      RECT 2.414 32.622 2.466 32.658 ;
      RECT 2.414 32.862 2.466 32.898 ;
      RECT 2.414 38.622 2.466 38.658 ;
      RECT 2.414 38.862 2.466 38.898 ;
      RECT 2.414 39.926 2.466 39.962 ;
      RECT 2.414 41.126 2.466 41.162 ;
      RECT 2.414 42.326 2.466 42.362 ;
      RECT 2.414 43.526 2.466 43.562 ;
      RECT 2.414 44.726 2.466 44.762 ;
      RECT 2.414 45.926 2.466 45.962 ;
      RECT 2.414 47.126 2.466 47.162 ;
      RECT 2.414 48.326 2.466 48.362 ;
      RECT 2.414 49.526 2.466 49.562 ;
      RECT 2.414 50.726 2.466 50.762 ;
      RECT 2.414 51.926 2.466 51.962 ;
      RECT 2.414 53.126 2.466 53.162 ;
      RECT 2.414 54.326 2.466 54.362 ;
      RECT 2.414 55.526 2.466 55.562 ;
      RECT 2.414 56.726 2.466 56.762 ;
      RECT 2.414 57.926 2.466 57.962 ;
      RECT 2.414 59.126 2.466 59.162 ;
      RECT 2.414 60.326 2.466 60.362 ;
      RECT 2.414 61.526 2.466 61.562 ;
      RECT 2.414 62.726 2.466 62.762 ;
      RECT 2.414 63.926 2.466 63.962 ;
      RECT 2.414 65.126 2.466 65.162 ;
      RECT 2.414 66.326 2.466 66.362 ;
      RECT 2.414 67.526 2.466 67.562 ;
      RECT 2.414 68.726 2.466 68.762 ;
      RECT 2.414 69.926 2.466 69.962 ;
      RECT 2.414 71.126 2.466 71.162 ;
      RECT 2.494 1.558 2.546 1.594 ;
      RECT 2.494 2.758 2.546 2.794 ;
      RECT 2.494 3.958 2.546 3.994 ;
      RECT 2.494 5.158 2.546 5.194 ;
      RECT 2.494 6.358 2.546 6.394 ;
      RECT 2.494 7.558 2.546 7.594 ;
      RECT 2.494 8.758 2.546 8.794 ;
      RECT 2.494 9.958 2.546 9.994 ;
      RECT 2.494 11.158 2.546 11.194 ;
      RECT 2.494 12.358 2.546 12.394 ;
      RECT 2.494 13.558 2.546 13.594 ;
      RECT 2.494 14.758 2.546 14.794 ;
      RECT 2.494 15.958 2.546 15.994 ;
      RECT 2.494 17.158 2.546 17.194 ;
      RECT 2.494 18.358 2.546 18.394 ;
      RECT 2.494 19.558 2.546 19.594 ;
      RECT 2.494 20.758 2.546 20.794 ;
      RECT 2.494 21.958 2.546 21.994 ;
      RECT 2.494 23.158 2.546 23.194 ;
      RECT 2.494 24.358 2.546 24.394 ;
      RECT 2.494 25.558 2.546 25.594 ;
      RECT 2.494 26.758 2.546 26.794 ;
      RECT 2.494 27.958 2.546 27.994 ;
      RECT 2.494 29.158 2.546 29.194 ;
      RECT 2.494 30.358 2.546 30.394 ;
      RECT 2.494 31.558 2.546 31.594 ;
      RECT 2.494 33.342 2.546 33.378 ;
      RECT 2.494 33.582 2.546 33.618 ;
      RECT 2.494 37.902 2.546 37.938 ;
      RECT 2.494 38.142 2.546 38.178 ;
      RECT 2.494 40.678 2.546 40.714 ;
      RECT 2.494 41.878 2.546 41.914 ;
      RECT 2.494 43.078 2.546 43.114 ;
      RECT 2.494 44.278 2.546 44.314 ;
      RECT 2.494 45.478 2.546 45.514 ;
      RECT 2.494 46.678 2.546 46.714 ;
      RECT 2.494 47.878 2.546 47.914 ;
      RECT 2.494 49.078 2.546 49.114 ;
      RECT 2.494 50.278 2.546 50.314 ;
      RECT 2.494 51.478 2.546 51.514 ;
      RECT 2.494 52.678 2.546 52.714 ;
      RECT 2.494 53.878 2.546 53.914 ;
      RECT 2.494 55.078 2.546 55.114 ;
      RECT 2.494 56.278 2.546 56.314 ;
      RECT 2.494 57.478 2.546 57.514 ;
      RECT 2.494 58.678 2.546 58.714 ;
      RECT 2.494 59.878 2.546 59.914 ;
      RECT 2.494 61.078 2.546 61.114 ;
      RECT 2.494 62.278 2.546 62.314 ;
      RECT 2.494 63.478 2.546 63.514 ;
      RECT 2.494 64.678 2.546 64.714 ;
      RECT 2.494 65.878 2.546 65.914 ;
      RECT 2.494 67.078 2.546 67.114 ;
      RECT 2.494 68.278 2.546 68.314 ;
      RECT 2.494 69.478 2.546 69.514 ;
      RECT 2.494 70.678 2.546 70.714 ;
      RECT 2.494 71.878 2.546 71.914 ;
      RECT 2.574 0.281 2.626 0.317 ;
      RECT 2.574 72.403 2.626 72.439 ;
      RECT 2.654 0.806 2.706 0.842 ;
      RECT 2.654 2.006 2.706 2.042 ;
      RECT 2.654 3.206 2.706 3.242 ;
      RECT 2.654 4.406 2.706 4.442 ;
      RECT 2.654 5.606 2.706 5.642 ;
      RECT 2.654 6.806 2.706 6.842 ;
      RECT 2.654 8.006 2.706 8.042 ;
      RECT 2.654 9.206 2.706 9.242 ;
      RECT 2.654 10.406 2.706 10.442 ;
      RECT 2.654 11.606 2.706 11.642 ;
      RECT 2.654 12.806 2.706 12.842 ;
      RECT 2.654 14.006 2.706 14.042 ;
      RECT 2.654 15.206 2.706 15.242 ;
      RECT 2.654 16.406 2.706 16.442 ;
      RECT 2.654 17.606 2.706 17.642 ;
      RECT 2.654 18.806 2.706 18.842 ;
      RECT 2.654 20.006 2.706 20.042 ;
      RECT 2.654 21.206 2.706 21.242 ;
      RECT 2.654 22.406 2.706 22.442 ;
      RECT 2.654 23.606 2.706 23.642 ;
      RECT 2.654 24.806 2.706 24.842 ;
      RECT 2.654 26.006 2.706 26.042 ;
      RECT 2.654 27.206 2.706 27.242 ;
      RECT 2.654 28.406 2.706 28.442 ;
      RECT 2.654 29.606 2.706 29.642 ;
      RECT 2.654 30.806 2.706 30.842 ;
      RECT 2.654 32.622 2.706 32.658 ;
      RECT 2.654 32.862 2.706 32.898 ;
      RECT 2.654 34.302 2.706 34.338 ;
      RECT 2.654 34.782 2.706 34.818 ;
      RECT 2.654 36.702 2.706 36.738 ;
      RECT 2.654 37.182 2.706 37.218 ;
      RECT 2.654 38.622 2.706 38.658 ;
      RECT 2.654 38.862 2.706 38.898 ;
      RECT 2.654 39.926 2.706 39.962 ;
      RECT 2.654 41.126 2.706 41.162 ;
      RECT 2.654 42.326 2.706 42.362 ;
      RECT 2.654 43.526 2.706 43.562 ;
      RECT 2.654 44.726 2.706 44.762 ;
      RECT 2.654 45.926 2.706 45.962 ;
      RECT 2.654 47.126 2.706 47.162 ;
      RECT 2.654 48.326 2.706 48.362 ;
      RECT 2.654 49.526 2.706 49.562 ;
      RECT 2.654 50.726 2.706 50.762 ;
      RECT 2.654 51.926 2.706 51.962 ;
      RECT 2.654 53.126 2.706 53.162 ;
      RECT 2.654 54.326 2.706 54.362 ;
      RECT 2.654 55.526 2.706 55.562 ;
      RECT 2.654 56.726 2.706 56.762 ;
      RECT 2.654 57.926 2.706 57.962 ;
      RECT 2.654 59.126 2.706 59.162 ;
      RECT 2.654 60.326 2.706 60.362 ;
      RECT 2.654 61.526 2.706 61.562 ;
      RECT 2.654 62.726 2.706 62.762 ;
      RECT 2.654 63.926 2.706 63.962 ;
      RECT 2.654 65.126 2.706 65.162 ;
      RECT 2.654 66.326 2.706 66.362 ;
      RECT 2.654 67.526 2.706 67.562 ;
      RECT 2.654 68.726 2.706 68.762 ;
      RECT 2.654 69.926 2.706 69.962 ;
      RECT 2.654 71.126 2.706 71.162 ;
      RECT 2.734 1.558 2.786 1.594 ;
      RECT 2.734 2.758 2.786 2.794 ;
      RECT 2.734 3.958 2.786 3.994 ;
      RECT 2.734 5.158 2.786 5.194 ;
      RECT 2.734 6.358 2.786 6.394 ;
      RECT 2.734 7.558 2.786 7.594 ;
      RECT 2.734 8.758 2.786 8.794 ;
      RECT 2.734 9.958 2.786 9.994 ;
      RECT 2.734 11.158 2.786 11.194 ;
      RECT 2.734 12.358 2.786 12.394 ;
      RECT 2.734 13.558 2.786 13.594 ;
      RECT 2.734 14.758 2.786 14.794 ;
      RECT 2.734 15.958 2.786 15.994 ;
      RECT 2.734 17.158 2.786 17.194 ;
      RECT 2.734 18.358 2.786 18.394 ;
      RECT 2.734 19.558 2.786 19.594 ;
      RECT 2.734 20.758 2.786 20.794 ;
      RECT 2.734 21.958 2.786 21.994 ;
      RECT 2.734 23.158 2.786 23.194 ;
      RECT 2.734 24.358 2.786 24.394 ;
      RECT 2.734 25.558 2.786 25.594 ;
      RECT 2.734 26.758 2.786 26.794 ;
      RECT 2.734 27.958 2.786 27.994 ;
      RECT 2.734 29.158 2.786 29.194 ;
      RECT 2.734 30.358 2.786 30.394 ;
      RECT 2.734 31.558 2.786 31.594 ;
      RECT 2.734 33.342 2.786 33.378 ;
      RECT 2.734 33.582 2.786 33.618 ;
      RECT 2.734 37.902 2.786 37.938 ;
      RECT 2.734 38.142 2.786 38.178 ;
      RECT 2.734 40.678 2.786 40.714 ;
      RECT 2.734 41.878 2.786 41.914 ;
      RECT 2.734 43.078 2.786 43.114 ;
      RECT 2.734 44.278 2.786 44.314 ;
      RECT 2.734 45.478 2.786 45.514 ;
      RECT 2.734 46.678 2.786 46.714 ;
      RECT 2.734 47.878 2.786 47.914 ;
      RECT 2.734 49.078 2.786 49.114 ;
      RECT 2.734 50.278 2.786 50.314 ;
      RECT 2.734 51.478 2.786 51.514 ;
      RECT 2.734 52.678 2.786 52.714 ;
      RECT 2.734 53.878 2.786 53.914 ;
      RECT 2.734 55.078 2.786 55.114 ;
      RECT 2.734 56.278 2.786 56.314 ;
      RECT 2.734 57.478 2.786 57.514 ;
      RECT 2.734 58.678 2.786 58.714 ;
      RECT 2.734 59.878 2.786 59.914 ;
      RECT 2.734 61.078 2.786 61.114 ;
      RECT 2.734 62.278 2.786 62.314 ;
      RECT 2.734 63.478 2.786 63.514 ;
      RECT 2.734 64.678 2.786 64.714 ;
      RECT 2.734 65.878 2.786 65.914 ;
      RECT 2.734 67.078 2.786 67.114 ;
      RECT 2.734 68.278 2.786 68.314 ;
      RECT 2.734 69.478 2.786 69.514 ;
      RECT 2.734 70.678 2.786 70.714 ;
      RECT 2.734 71.878 2.786 71.914 ;
      RECT 2.814 0.806 2.866 0.842 ;
      RECT 2.814 2.006 2.866 2.042 ;
      RECT 2.814 3.206 2.866 3.242 ;
      RECT 2.814 4.406 2.866 4.442 ;
      RECT 2.814 5.606 2.866 5.642 ;
      RECT 2.814 6.806 2.866 6.842 ;
      RECT 2.814 8.006 2.866 8.042 ;
      RECT 2.814 9.206 2.866 9.242 ;
      RECT 2.814 10.406 2.866 10.442 ;
      RECT 2.814 11.606 2.866 11.642 ;
      RECT 2.814 12.806 2.866 12.842 ;
      RECT 2.814 14.006 2.866 14.042 ;
      RECT 2.814 15.206 2.866 15.242 ;
      RECT 2.814 16.406 2.866 16.442 ;
      RECT 2.814 17.606 2.866 17.642 ;
      RECT 2.814 18.806 2.866 18.842 ;
      RECT 2.814 20.006 2.866 20.042 ;
      RECT 2.814 21.206 2.866 21.242 ;
      RECT 2.814 22.406 2.866 22.442 ;
      RECT 2.814 23.606 2.866 23.642 ;
      RECT 2.814 24.806 2.866 24.842 ;
      RECT 2.814 26.006 2.866 26.042 ;
      RECT 2.814 27.206 2.866 27.242 ;
      RECT 2.814 28.406 2.866 28.442 ;
      RECT 2.814 29.606 2.866 29.642 ;
      RECT 2.814 30.806 2.866 30.842 ;
      RECT 2.814 32.622 2.866 32.658 ;
      RECT 2.814 32.862 2.866 32.898 ;
      RECT 2.814 38.622 2.866 38.658 ;
      RECT 2.814 38.862 2.866 38.898 ;
      RECT 2.814 39.926 2.866 39.962 ;
      RECT 2.814 41.126 2.866 41.162 ;
      RECT 2.814 42.326 2.866 42.362 ;
      RECT 2.814 43.526 2.866 43.562 ;
      RECT 2.814 44.726 2.866 44.762 ;
      RECT 2.814 45.926 2.866 45.962 ;
      RECT 2.814 47.126 2.866 47.162 ;
      RECT 2.814 48.326 2.866 48.362 ;
      RECT 2.814 49.526 2.866 49.562 ;
      RECT 2.814 50.726 2.866 50.762 ;
      RECT 2.814 51.926 2.866 51.962 ;
      RECT 2.814 53.126 2.866 53.162 ;
      RECT 2.814 54.326 2.866 54.362 ;
      RECT 2.814 55.526 2.866 55.562 ;
      RECT 2.814 56.726 2.866 56.762 ;
      RECT 2.814 57.926 2.866 57.962 ;
      RECT 2.814 59.126 2.866 59.162 ;
      RECT 2.814 60.326 2.866 60.362 ;
      RECT 2.814 61.526 2.866 61.562 ;
      RECT 2.814 62.726 2.866 62.762 ;
      RECT 2.814 63.926 2.866 63.962 ;
      RECT 2.814 65.126 2.866 65.162 ;
      RECT 2.814 66.326 2.866 66.362 ;
      RECT 2.814 67.526 2.866 67.562 ;
      RECT 2.814 68.726 2.866 68.762 ;
      RECT 2.814 69.926 2.866 69.962 ;
      RECT 2.814 71.126 2.866 71.162 ;
      RECT 2.894 1.558 2.946 1.594 ;
      RECT 2.894 2.758 2.946 2.794 ;
      RECT 2.894 3.958 2.946 3.994 ;
      RECT 2.894 5.158 2.946 5.194 ;
      RECT 2.894 6.358 2.946 6.394 ;
      RECT 2.894 7.558 2.946 7.594 ;
      RECT 2.894 8.758 2.946 8.794 ;
      RECT 2.894 9.958 2.946 9.994 ;
      RECT 2.894 11.158 2.946 11.194 ;
      RECT 2.894 12.358 2.946 12.394 ;
      RECT 2.894 13.558 2.946 13.594 ;
      RECT 2.894 14.758 2.946 14.794 ;
      RECT 2.894 15.958 2.946 15.994 ;
      RECT 2.894 17.158 2.946 17.194 ;
      RECT 2.894 18.358 2.946 18.394 ;
      RECT 2.894 19.558 2.946 19.594 ;
      RECT 2.894 20.758 2.946 20.794 ;
      RECT 2.894 21.958 2.946 21.994 ;
      RECT 2.894 23.158 2.946 23.194 ;
      RECT 2.894 24.358 2.946 24.394 ;
      RECT 2.894 25.558 2.946 25.594 ;
      RECT 2.894 26.758 2.946 26.794 ;
      RECT 2.894 27.958 2.946 27.994 ;
      RECT 2.894 29.158 2.946 29.194 ;
      RECT 2.894 30.358 2.946 30.394 ;
      RECT 2.894 31.558 2.946 31.594 ;
      RECT 2.894 33.342 2.946 33.378 ;
      RECT 2.894 33.582 2.946 33.618 ;
      RECT 2.894 37.902 2.946 37.938 ;
      RECT 2.894 38.142 2.946 38.178 ;
      RECT 2.894 40.678 2.946 40.714 ;
      RECT 2.894 41.878 2.946 41.914 ;
      RECT 2.894 43.078 2.946 43.114 ;
      RECT 2.894 44.278 2.946 44.314 ;
      RECT 2.894 45.478 2.946 45.514 ;
      RECT 2.894 46.678 2.946 46.714 ;
      RECT 2.894 47.878 2.946 47.914 ;
      RECT 2.894 49.078 2.946 49.114 ;
      RECT 2.894 50.278 2.946 50.314 ;
      RECT 2.894 51.478 2.946 51.514 ;
      RECT 2.894 52.678 2.946 52.714 ;
      RECT 2.894 53.878 2.946 53.914 ;
      RECT 2.894 55.078 2.946 55.114 ;
      RECT 2.894 56.278 2.946 56.314 ;
      RECT 2.894 57.478 2.946 57.514 ;
      RECT 2.894 58.678 2.946 58.714 ;
      RECT 2.894 59.878 2.946 59.914 ;
      RECT 2.894 61.078 2.946 61.114 ;
      RECT 2.894 62.278 2.946 62.314 ;
      RECT 2.894 63.478 2.946 63.514 ;
      RECT 2.894 64.678 2.946 64.714 ;
      RECT 2.894 65.878 2.946 65.914 ;
      RECT 2.894 67.078 2.946 67.114 ;
      RECT 2.894 68.278 2.946 68.314 ;
      RECT 2.894 69.478 2.946 69.514 ;
      RECT 2.894 70.678 2.946 70.714 ;
      RECT 2.894 71.878 2.946 71.914 ;
      RECT 2.974 0.281 3.026 0.317 ;
      RECT 2.974 72.403 3.026 72.439 ;
      RECT 3.054 0.806 3.106 0.842 ;
      RECT 3.054 2.006 3.106 2.042 ;
      RECT 3.054 3.206 3.106 3.242 ;
      RECT 3.054 4.406 3.106 4.442 ;
      RECT 3.054 5.606 3.106 5.642 ;
      RECT 3.054 6.806 3.106 6.842 ;
      RECT 3.054 8.006 3.106 8.042 ;
      RECT 3.054 9.206 3.106 9.242 ;
      RECT 3.054 10.406 3.106 10.442 ;
      RECT 3.054 11.606 3.106 11.642 ;
      RECT 3.054 12.806 3.106 12.842 ;
      RECT 3.054 14.006 3.106 14.042 ;
      RECT 3.054 15.206 3.106 15.242 ;
      RECT 3.054 16.406 3.106 16.442 ;
      RECT 3.054 17.606 3.106 17.642 ;
      RECT 3.054 18.806 3.106 18.842 ;
      RECT 3.054 20.006 3.106 20.042 ;
      RECT 3.054 21.206 3.106 21.242 ;
      RECT 3.054 22.406 3.106 22.442 ;
      RECT 3.054 23.606 3.106 23.642 ;
      RECT 3.054 24.806 3.106 24.842 ;
      RECT 3.054 26.006 3.106 26.042 ;
      RECT 3.054 27.206 3.106 27.242 ;
      RECT 3.054 28.406 3.106 28.442 ;
      RECT 3.054 29.606 3.106 29.642 ;
      RECT 3.054 30.806 3.106 30.842 ;
      RECT 3.054 32.622 3.106 32.658 ;
      RECT 3.054 32.862 3.106 32.898 ;
      RECT 3.054 38.622 3.106 38.658 ;
      RECT 3.054 38.862 3.106 38.898 ;
      RECT 3.054 39.926 3.106 39.962 ;
      RECT 3.054 41.126 3.106 41.162 ;
      RECT 3.054 42.326 3.106 42.362 ;
      RECT 3.054 43.526 3.106 43.562 ;
      RECT 3.054 44.726 3.106 44.762 ;
      RECT 3.054 45.926 3.106 45.962 ;
      RECT 3.054 47.126 3.106 47.162 ;
      RECT 3.054 48.326 3.106 48.362 ;
      RECT 3.054 49.526 3.106 49.562 ;
      RECT 3.054 50.726 3.106 50.762 ;
      RECT 3.054 51.926 3.106 51.962 ;
      RECT 3.054 53.126 3.106 53.162 ;
      RECT 3.054 54.326 3.106 54.362 ;
      RECT 3.054 55.526 3.106 55.562 ;
      RECT 3.054 56.726 3.106 56.762 ;
      RECT 3.054 57.926 3.106 57.962 ;
      RECT 3.054 59.126 3.106 59.162 ;
      RECT 3.054 60.326 3.106 60.362 ;
      RECT 3.054 61.526 3.106 61.562 ;
      RECT 3.054 62.726 3.106 62.762 ;
      RECT 3.054 63.926 3.106 63.962 ;
      RECT 3.054 65.126 3.106 65.162 ;
      RECT 3.054 66.326 3.106 66.362 ;
      RECT 3.054 67.526 3.106 67.562 ;
      RECT 3.054 68.726 3.106 68.762 ;
      RECT 3.054 69.926 3.106 69.962 ;
      RECT 3.054 71.126 3.106 71.162 ;
      RECT 3.134 1.558 3.186 1.594 ;
      RECT 3.134 2.758 3.186 2.794 ;
      RECT 3.134 3.958 3.186 3.994 ;
      RECT 3.134 5.158 3.186 5.194 ;
      RECT 3.134 6.358 3.186 6.394 ;
      RECT 3.134 7.558 3.186 7.594 ;
      RECT 3.134 8.758 3.186 8.794 ;
      RECT 3.134 9.958 3.186 9.994 ;
      RECT 3.134 11.158 3.186 11.194 ;
      RECT 3.134 12.358 3.186 12.394 ;
      RECT 3.134 13.558 3.186 13.594 ;
      RECT 3.134 14.758 3.186 14.794 ;
      RECT 3.134 15.958 3.186 15.994 ;
      RECT 3.134 17.158 3.186 17.194 ;
      RECT 3.134 18.358 3.186 18.394 ;
      RECT 3.134 19.558 3.186 19.594 ;
      RECT 3.134 20.758 3.186 20.794 ;
      RECT 3.134 21.958 3.186 21.994 ;
      RECT 3.134 23.158 3.186 23.194 ;
      RECT 3.134 24.358 3.186 24.394 ;
      RECT 3.134 25.558 3.186 25.594 ;
      RECT 3.134 26.758 3.186 26.794 ;
      RECT 3.134 27.958 3.186 27.994 ;
      RECT 3.134 29.158 3.186 29.194 ;
      RECT 3.134 30.358 3.186 30.394 ;
      RECT 3.134 31.558 3.186 31.594 ;
      RECT 3.134 33.342 3.186 33.378 ;
      RECT 3.134 33.582 3.186 33.618 ;
      RECT 3.134 37.902 3.186 37.938 ;
      RECT 3.134 38.142 3.186 38.178 ;
      RECT 3.134 40.678 3.186 40.714 ;
      RECT 3.134 41.878 3.186 41.914 ;
      RECT 3.134 43.078 3.186 43.114 ;
      RECT 3.134 44.278 3.186 44.314 ;
      RECT 3.134 45.478 3.186 45.514 ;
      RECT 3.134 46.678 3.186 46.714 ;
      RECT 3.134 47.878 3.186 47.914 ;
      RECT 3.134 49.078 3.186 49.114 ;
      RECT 3.134 50.278 3.186 50.314 ;
      RECT 3.134 51.478 3.186 51.514 ;
      RECT 3.134 52.678 3.186 52.714 ;
      RECT 3.134 53.878 3.186 53.914 ;
      RECT 3.134 55.078 3.186 55.114 ;
      RECT 3.134 56.278 3.186 56.314 ;
      RECT 3.134 57.478 3.186 57.514 ;
      RECT 3.134 58.678 3.186 58.714 ;
      RECT 3.134 59.878 3.186 59.914 ;
      RECT 3.134 61.078 3.186 61.114 ;
      RECT 3.134 62.278 3.186 62.314 ;
      RECT 3.134 63.478 3.186 63.514 ;
      RECT 3.134 64.678 3.186 64.714 ;
      RECT 3.134 65.878 3.186 65.914 ;
      RECT 3.134 67.078 3.186 67.114 ;
      RECT 3.134 68.278 3.186 68.314 ;
      RECT 3.134 69.478 3.186 69.514 ;
      RECT 3.134 70.678 3.186 70.714 ;
      RECT 3.134 71.878 3.186 71.914 ;
      RECT 3.214 0.806 3.266 0.842 ;
      RECT 3.214 2.006 3.266 2.042 ;
      RECT 3.214 3.206 3.266 3.242 ;
      RECT 3.214 4.406 3.266 4.442 ;
      RECT 3.214 5.606 3.266 5.642 ;
      RECT 3.214 6.806 3.266 6.842 ;
      RECT 3.214 8.006 3.266 8.042 ;
      RECT 3.214 9.206 3.266 9.242 ;
      RECT 3.214 10.406 3.266 10.442 ;
      RECT 3.214 11.606 3.266 11.642 ;
      RECT 3.214 12.806 3.266 12.842 ;
      RECT 3.214 14.006 3.266 14.042 ;
      RECT 3.214 15.206 3.266 15.242 ;
      RECT 3.214 16.406 3.266 16.442 ;
      RECT 3.214 17.606 3.266 17.642 ;
      RECT 3.214 18.806 3.266 18.842 ;
      RECT 3.214 20.006 3.266 20.042 ;
      RECT 3.214 21.206 3.266 21.242 ;
      RECT 3.214 22.406 3.266 22.442 ;
      RECT 3.214 23.606 3.266 23.642 ;
      RECT 3.214 24.806 3.266 24.842 ;
      RECT 3.214 26.006 3.266 26.042 ;
      RECT 3.214 27.206 3.266 27.242 ;
      RECT 3.214 28.406 3.266 28.442 ;
      RECT 3.214 29.606 3.266 29.642 ;
      RECT 3.214 30.806 3.266 30.842 ;
      RECT 3.214 32.622 3.266 32.658 ;
      RECT 3.214 32.862 3.266 32.898 ;
      RECT 3.214 38.622 3.266 38.658 ;
      RECT 3.214 38.862 3.266 38.898 ;
      RECT 3.214 39.926 3.266 39.962 ;
      RECT 3.214 41.126 3.266 41.162 ;
      RECT 3.214 42.326 3.266 42.362 ;
      RECT 3.214 43.526 3.266 43.562 ;
      RECT 3.214 44.726 3.266 44.762 ;
      RECT 3.214 45.926 3.266 45.962 ;
      RECT 3.214 47.126 3.266 47.162 ;
      RECT 3.214 48.326 3.266 48.362 ;
      RECT 3.214 49.526 3.266 49.562 ;
      RECT 3.214 50.726 3.266 50.762 ;
      RECT 3.214 51.926 3.266 51.962 ;
      RECT 3.214 53.126 3.266 53.162 ;
      RECT 3.214 54.326 3.266 54.362 ;
      RECT 3.214 55.526 3.266 55.562 ;
      RECT 3.214 56.726 3.266 56.762 ;
      RECT 3.214 57.926 3.266 57.962 ;
      RECT 3.214 59.126 3.266 59.162 ;
      RECT 3.214 60.326 3.266 60.362 ;
      RECT 3.214 61.526 3.266 61.562 ;
      RECT 3.214 62.726 3.266 62.762 ;
      RECT 3.214 63.926 3.266 63.962 ;
      RECT 3.214 65.126 3.266 65.162 ;
      RECT 3.214 66.326 3.266 66.362 ;
      RECT 3.214 67.526 3.266 67.562 ;
      RECT 3.214 68.726 3.266 68.762 ;
      RECT 3.214 69.926 3.266 69.962 ;
      RECT 3.214 71.126 3.266 71.162 ;
      RECT 3.294 1.558 3.346 1.594 ;
      RECT 3.294 2.758 3.346 2.794 ;
      RECT 3.294 3.958 3.346 3.994 ;
      RECT 3.294 5.158 3.346 5.194 ;
      RECT 3.294 6.358 3.346 6.394 ;
      RECT 3.294 7.558 3.346 7.594 ;
      RECT 3.294 8.758 3.346 8.794 ;
      RECT 3.294 9.958 3.346 9.994 ;
      RECT 3.294 11.158 3.346 11.194 ;
      RECT 3.294 12.358 3.346 12.394 ;
      RECT 3.294 13.558 3.346 13.594 ;
      RECT 3.294 14.758 3.346 14.794 ;
      RECT 3.294 15.958 3.346 15.994 ;
      RECT 3.294 17.158 3.346 17.194 ;
      RECT 3.294 18.358 3.346 18.394 ;
      RECT 3.294 19.558 3.346 19.594 ;
      RECT 3.294 20.758 3.346 20.794 ;
      RECT 3.294 21.958 3.346 21.994 ;
      RECT 3.294 23.158 3.346 23.194 ;
      RECT 3.294 24.358 3.346 24.394 ;
      RECT 3.294 25.558 3.346 25.594 ;
      RECT 3.294 26.758 3.346 26.794 ;
      RECT 3.294 27.958 3.346 27.994 ;
      RECT 3.294 29.158 3.346 29.194 ;
      RECT 3.294 30.358 3.346 30.394 ;
      RECT 3.294 31.558 3.346 31.594 ;
      RECT 3.294 33.342 3.346 33.378 ;
      RECT 3.294 33.582 3.346 33.618 ;
      RECT 3.294 37.902 3.346 37.938 ;
      RECT 3.294 38.142 3.346 38.178 ;
      RECT 3.294 40.678 3.346 40.714 ;
      RECT 3.294 41.878 3.346 41.914 ;
      RECT 3.294 43.078 3.346 43.114 ;
      RECT 3.294 44.278 3.346 44.314 ;
      RECT 3.294 45.478 3.346 45.514 ;
      RECT 3.294 46.678 3.346 46.714 ;
      RECT 3.294 47.878 3.346 47.914 ;
      RECT 3.294 49.078 3.346 49.114 ;
      RECT 3.294 50.278 3.346 50.314 ;
      RECT 3.294 51.478 3.346 51.514 ;
      RECT 3.294 52.678 3.346 52.714 ;
      RECT 3.294 53.878 3.346 53.914 ;
      RECT 3.294 55.078 3.346 55.114 ;
      RECT 3.294 56.278 3.346 56.314 ;
      RECT 3.294 57.478 3.346 57.514 ;
      RECT 3.294 58.678 3.346 58.714 ;
      RECT 3.294 59.878 3.346 59.914 ;
      RECT 3.294 61.078 3.346 61.114 ;
      RECT 3.294 62.278 3.346 62.314 ;
      RECT 3.294 63.478 3.346 63.514 ;
      RECT 3.294 64.678 3.346 64.714 ;
      RECT 3.294 65.878 3.346 65.914 ;
      RECT 3.294 67.078 3.346 67.114 ;
      RECT 3.294 68.278 3.346 68.314 ;
      RECT 3.294 69.478 3.346 69.514 ;
      RECT 3.294 70.678 3.346 70.714 ;
      RECT 3.294 71.878 3.346 71.914 ;
      RECT 3.374 0.281 3.426 0.317 ;
      RECT 3.374 72.403 3.426 72.439 ;
      RECT 3.454 0.806 3.506 0.842 ;
      RECT 3.454 2.006 3.506 2.042 ;
      RECT 3.454 3.206 3.506 3.242 ;
      RECT 3.454 4.406 3.506 4.442 ;
      RECT 3.454 5.606 3.506 5.642 ;
      RECT 3.454 6.806 3.506 6.842 ;
      RECT 3.454 8.006 3.506 8.042 ;
      RECT 3.454 9.206 3.506 9.242 ;
      RECT 3.454 10.406 3.506 10.442 ;
      RECT 3.454 11.606 3.506 11.642 ;
      RECT 3.454 12.806 3.506 12.842 ;
      RECT 3.454 14.006 3.506 14.042 ;
      RECT 3.454 15.206 3.506 15.242 ;
      RECT 3.454 16.406 3.506 16.442 ;
      RECT 3.454 17.606 3.506 17.642 ;
      RECT 3.454 18.806 3.506 18.842 ;
      RECT 3.454 20.006 3.506 20.042 ;
      RECT 3.454 21.206 3.506 21.242 ;
      RECT 3.454 22.406 3.506 22.442 ;
      RECT 3.454 23.606 3.506 23.642 ;
      RECT 3.454 24.806 3.506 24.842 ;
      RECT 3.454 26.006 3.506 26.042 ;
      RECT 3.454 27.206 3.506 27.242 ;
      RECT 3.454 28.406 3.506 28.442 ;
      RECT 3.454 29.606 3.506 29.642 ;
      RECT 3.454 30.806 3.506 30.842 ;
      RECT 3.454 32.622 3.506 32.658 ;
      RECT 3.454 32.862 3.506 32.898 ;
      RECT 3.454 34.302 3.506 34.338 ;
      RECT 3.454 34.782 3.506 34.818 ;
      RECT 3.454 36.702 3.506 36.738 ;
      RECT 3.454 37.182 3.506 37.218 ;
      RECT 3.454 38.622 3.506 38.658 ;
      RECT 3.454 38.862 3.506 38.898 ;
      RECT 3.454 39.926 3.506 39.962 ;
      RECT 3.454 41.126 3.506 41.162 ;
      RECT 3.454 42.326 3.506 42.362 ;
      RECT 3.454 43.526 3.506 43.562 ;
      RECT 3.454 44.726 3.506 44.762 ;
      RECT 3.454 45.926 3.506 45.962 ;
      RECT 3.454 47.126 3.506 47.162 ;
      RECT 3.454 48.326 3.506 48.362 ;
      RECT 3.454 49.526 3.506 49.562 ;
      RECT 3.454 50.726 3.506 50.762 ;
      RECT 3.454 51.926 3.506 51.962 ;
      RECT 3.454 53.126 3.506 53.162 ;
      RECT 3.454 54.326 3.506 54.362 ;
      RECT 3.454 55.526 3.506 55.562 ;
      RECT 3.454 56.726 3.506 56.762 ;
      RECT 3.454 57.926 3.506 57.962 ;
      RECT 3.454 59.126 3.506 59.162 ;
      RECT 3.454 60.326 3.506 60.362 ;
      RECT 3.454 61.526 3.506 61.562 ;
      RECT 3.454 62.726 3.506 62.762 ;
      RECT 3.454 63.926 3.506 63.962 ;
      RECT 3.454 65.126 3.506 65.162 ;
      RECT 3.454 66.326 3.506 66.362 ;
      RECT 3.454 67.526 3.506 67.562 ;
      RECT 3.454 68.726 3.506 68.762 ;
      RECT 3.454 69.926 3.506 69.962 ;
      RECT 3.454 71.126 3.506 71.162 ;
      RECT 3.534 1.558 3.586 1.594 ;
      RECT 3.534 2.758 3.586 2.794 ;
      RECT 3.534 3.958 3.586 3.994 ;
      RECT 3.534 5.158 3.586 5.194 ;
      RECT 3.534 6.358 3.586 6.394 ;
      RECT 3.534 7.558 3.586 7.594 ;
      RECT 3.534 8.758 3.586 8.794 ;
      RECT 3.534 9.958 3.586 9.994 ;
      RECT 3.534 11.158 3.586 11.194 ;
      RECT 3.534 12.358 3.586 12.394 ;
      RECT 3.534 13.558 3.586 13.594 ;
      RECT 3.534 14.758 3.586 14.794 ;
      RECT 3.534 15.958 3.586 15.994 ;
      RECT 3.534 17.158 3.586 17.194 ;
      RECT 3.534 18.358 3.586 18.394 ;
      RECT 3.534 19.558 3.586 19.594 ;
      RECT 3.534 20.758 3.586 20.794 ;
      RECT 3.534 21.958 3.586 21.994 ;
      RECT 3.534 23.158 3.586 23.194 ;
      RECT 3.534 24.358 3.586 24.394 ;
      RECT 3.534 25.558 3.586 25.594 ;
      RECT 3.534 26.758 3.586 26.794 ;
      RECT 3.534 27.958 3.586 27.994 ;
      RECT 3.534 29.158 3.586 29.194 ;
      RECT 3.534 30.358 3.586 30.394 ;
      RECT 3.534 31.558 3.586 31.594 ;
      RECT 3.534 33.342 3.586 33.378 ;
      RECT 3.534 33.582 3.586 33.618 ;
      RECT 3.534 37.902 3.586 37.938 ;
      RECT 3.534 38.142 3.586 38.178 ;
      RECT 3.534 40.678 3.586 40.714 ;
      RECT 3.534 41.878 3.586 41.914 ;
      RECT 3.534 43.078 3.586 43.114 ;
      RECT 3.534 44.278 3.586 44.314 ;
      RECT 3.534 45.478 3.586 45.514 ;
      RECT 3.534 46.678 3.586 46.714 ;
      RECT 3.534 47.878 3.586 47.914 ;
      RECT 3.534 49.078 3.586 49.114 ;
      RECT 3.534 50.278 3.586 50.314 ;
      RECT 3.534 51.478 3.586 51.514 ;
      RECT 3.534 52.678 3.586 52.714 ;
      RECT 3.534 53.878 3.586 53.914 ;
      RECT 3.534 55.078 3.586 55.114 ;
      RECT 3.534 56.278 3.586 56.314 ;
      RECT 3.534 57.478 3.586 57.514 ;
      RECT 3.534 58.678 3.586 58.714 ;
      RECT 3.534 59.878 3.586 59.914 ;
      RECT 3.534 61.078 3.586 61.114 ;
      RECT 3.534 62.278 3.586 62.314 ;
      RECT 3.534 63.478 3.586 63.514 ;
      RECT 3.534 64.678 3.586 64.714 ;
      RECT 3.534 65.878 3.586 65.914 ;
      RECT 3.534 67.078 3.586 67.114 ;
      RECT 3.534 68.278 3.586 68.314 ;
      RECT 3.534 69.478 3.586 69.514 ;
      RECT 3.534 70.678 3.586 70.714 ;
      RECT 3.534 71.878 3.586 71.914 ;
      RECT 3.614 0.806 3.666 0.842 ;
      RECT 3.614 2.006 3.666 2.042 ;
      RECT 3.614 3.206 3.666 3.242 ;
      RECT 3.614 4.406 3.666 4.442 ;
      RECT 3.614 5.606 3.666 5.642 ;
      RECT 3.614 6.806 3.666 6.842 ;
      RECT 3.614 8.006 3.666 8.042 ;
      RECT 3.614 9.206 3.666 9.242 ;
      RECT 3.614 10.406 3.666 10.442 ;
      RECT 3.614 11.606 3.666 11.642 ;
      RECT 3.614 12.806 3.666 12.842 ;
      RECT 3.614 14.006 3.666 14.042 ;
      RECT 3.614 15.206 3.666 15.242 ;
      RECT 3.614 16.406 3.666 16.442 ;
      RECT 3.614 17.606 3.666 17.642 ;
      RECT 3.614 18.806 3.666 18.842 ;
      RECT 3.614 20.006 3.666 20.042 ;
      RECT 3.614 21.206 3.666 21.242 ;
      RECT 3.614 22.406 3.666 22.442 ;
      RECT 3.614 23.606 3.666 23.642 ;
      RECT 3.614 24.806 3.666 24.842 ;
      RECT 3.614 26.006 3.666 26.042 ;
      RECT 3.614 27.206 3.666 27.242 ;
      RECT 3.614 28.406 3.666 28.442 ;
      RECT 3.614 29.606 3.666 29.642 ;
      RECT 3.614 30.806 3.666 30.842 ;
      RECT 3.614 32.622 3.666 32.658 ;
      RECT 3.614 32.862 3.666 32.898 ;
      RECT 3.614 38.622 3.666 38.658 ;
      RECT 3.614 38.862 3.666 38.898 ;
      RECT 3.614 39.926 3.666 39.962 ;
      RECT 3.614 41.126 3.666 41.162 ;
      RECT 3.614 42.326 3.666 42.362 ;
      RECT 3.614 43.526 3.666 43.562 ;
      RECT 3.614 44.726 3.666 44.762 ;
      RECT 3.614 45.926 3.666 45.962 ;
      RECT 3.614 47.126 3.666 47.162 ;
      RECT 3.614 48.326 3.666 48.362 ;
      RECT 3.614 49.526 3.666 49.562 ;
      RECT 3.614 50.726 3.666 50.762 ;
      RECT 3.614 51.926 3.666 51.962 ;
      RECT 3.614 53.126 3.666 53.162 ;
      RECT 3.614 54.326 3.666 54.362 ;
      RECT 3.614 55.526 3.666 55.562 ;
      RECT 3.614 56.726 3.666 56.762 ;
      RECT 3.614 57.926 3.666 57.962 ;
      RECT 3.614 59.126 3.666 59.162 ;
      RECT 3.614 60.326 3.666 60.362 ;
      RECT 3.614 61.526 3.666 61.562 ;
      RECT 3.614 62.726 3.666 62.762 ;
      RECT 3.614 63.926 3.666 63.962 ;
      RECT 3.614 65.126 3.666 65.162 ;
      RECT 3.614 66.326 3.666 66.362 ;
      RECT 3.614 67.526 3.666 67.562 ;
      RECT 3.614 68.726 3.666 68.762 ;
      RECT 3.614 69.926 3.666 69.962 ;
      RECT 3.614 71.126 3.666 71.162 ;
      RECT 3.694 1.558 3.746 1.594 ;
      RECT 3.694 2.758 3.746 2.794 ;
      RECT 3.694 3.958 3.746 3.994 ;
      RECT 3.694 5.158 3.746 5.194 ;
      RECT 3.694 6.358 3.746 6.394 ;
      RECT 3.694 7.558 3.746 7.594 ;
      RECT 3.694 8.758 3.746 8.794 ;
      RECT 3.694 9.958 3.746 9.994 ;
      RECT 3.694 11.158 3.746 11.194 ;
      RECT 3.694 12.358 3.746 12.394 ;
      RECT 3.694 13.558 3.746 13.594 ;
      RECT 3.694 14.758 3.746 14.794 ;
      RECT 3.694 15.958 3.746 15.994 ;
      RECT 3.694 17.158 3.746 17.194 ;
      RECT 3.694 18.358 3.746 18.394 ;
      RECT 3.694 19.558 3.746 19.594 ;
      RECT 3.694 20.758 3.746 20.794 ;
      RECT 3.694 21.958 3.746 21.994 ;
      RECT 3.694 23.158 3.746 23.194 ;
      RECT 3.694 24.358 3.746 24.394 ;
      RECT 3.694 25.558 3.746 25.594 ;
      RECT 3.694 26.758 3.746 26.794 ;
      RECT 3.694 27.958 3.746 27.994 ;
      RECT 3.694 29.158 3.746 29.194 ;
      RECT 3.694 30.358 3.746 30.394 ;
      RECT 3.694 31.558 3.746 31.594 ;
      RECT 3.694 33.342 3.746 33.378 ;
      RECT 3.694 33.582 3.746 33.618 ;
      RECT 3.694 37.902 3.746 37.938 ;
      RECT 3.694 38.142 3.746 38.178 ;
      RECT 3.694 40.678 3.746 40.714 ;
      RECT 3.694 41.878 3.746 41.914 ;
      RECT 3.694 43.078 3.746 43.114 ;
      RECT 3.694 44.278 3.746 44.314 ;
      RECT 3.694 45.478 3.746 45.514 ;
      RECT 3.694 46.678 3.746 46.714 ;
      RECT 3.694 47.878 3.746 47.914 ;
      RECT 3.694 49.078 3.746 49.114 ;
      RECT 3.694 50.278 3.746 50.314 ;
      RECT 3.694 51.478 3.746 51.514 ;
      RECT 3.694 52.678 3.746 52.714 ;
      RECT 3.694 53.878 3.746 53.914 ;
      RECT 3.694 55.078 3.746 55.114 ;
      RECT 3.694 56.278 3.746 56.314 ;
      RECT 3.694 57.478 3.746 57.514 ;
      RECT 3.694 58.678 3.746 58.714 ;
      RECT 3.694 59.878 3.746 59.914 ;
      RECT 3.694 61.078 3.746 61.114 ;
      RECT 3.694 62.278 3.746 62.314 ;
      RECT 3.694 63.478 3.746 63.514 ;
      RECT 3.694 64.678 3.746 64.714 ;
      RECT 3.694 65.878 3.746 65.914 ;
      RECT 3.694 67.078 3.746 67.114 ;
      RECT 3.694 68.278 3.746 68.314 ;
      RECT 3.694 69.478 3.746 69.514 ;
      RECT 3.694 70.678 3.746 70.714 ;
      RECT 3.694 71.878 3.746 71.914 ;
      RECT 3.774 0.281 3.826 0.317 ;
      RECT 3.774 72.403 3.826 72.439 ;
      RECT 3.854 0.806 3.906 0.842 ;
      RECT 3.854 2.006 3.906 2.042 ;
      RECT 3.854 3.206 3.906 3.242 ;
      RECT 3.854 4.406 3.906 4.442 ;
      RECT 3.854 5.606 3.906 5.642 ;
      RECT 3.854 6.806 3.906 6.842 ;
      RECT 3.854 8.006 3.906 8.042 ;
      RECT 3.854 9.206 3.906 9.242 ;
      RECT 3.854 10.406 3.906 10.442 ;
      RECT 3.854 11.606 3.906 11.642 ;
      RECT 3.854 12.806 3.906 12.842 ;
      RECT 3.854 14.006 3.906 14.042 ;
      RECT 3.854 15.206 3.906 15.242 ;
      RECT 3.854 16.406 3.906 16.442 ;
      RECT 3.854 17.606 3.906 17.642 ;
      RECT 3.854 18.806 3.906 18.842 ;
      RECT 3.854 20.006 3.906 20.042 ;
      RECT 3.854 21.206 3.906 21.242 ;
      RECT 3.854 22.406 3.906 22.442 ;
      RECT 3.854 23.606 3.906 23.642 ;
      RECT 3.854 24.806 3.906 24.842 ;
      RECT 3.854 26.006 3.906 26.042 ;
      RECT 3.854 27.206 3.906 27.242 ;
      RECT 3.854 28.406 3.906 28.442 ;
      RECT 3.854 29.606 3.906 29.642 ;
      RECT 3.854 30.806 3.906 30.842 ;
      RECT 3.854 32.622 3.906 32.658 ;
      RECT 3.854 32.862 3.906 32.898 ;
      RECT 3.854 38.622 3.906 38.658 ;
      RECT 3.854 38.862 3.906 38.898 ;
      RECT 3.854 39.926 3.906 39.962 ;
      RECT 3.854 41.126 3.906 41.162 ;
      RECT 3.854 42.326 3.906 42.362 ;
      RECT 3.854 43.526 3.906 43.562 ;
      RECT 3.854 44.726 3.906 44.762 ;
      RECT 3.854 45.926 3.906 45.962 ;
      RECT 3.854 47.126 3.906 47.162 ;
      RECT 3.854 48.326 3.906 48.362 ;
      RECT 3.854 49.526 3.906 49.562 ;
      RECT 3.854 50.726 3.906 50.762 ;
      RECT 3.854 51.926 3.906 51.962 ;
      RECT 3.854 53.126 3.906 53.162 ;
      RECT 3.854 54.326 3.906 54.362 ;
      RECT 3.854 55.526 3.906 55.562 ;
      RECT 3.854 56.726 3.906 56.762 ;
      RECT 3.854 57.926 3.906 57.962 ;
      RECT 3.854 59.126 3.906 59.162 ;
      RECT 3.854 60.326 3.906 60.362 ;
      RECT 3.854 61.526 3.906 61.562 ;
      RECT 3.854 62.726 3.906 62.762 ;
      RECT 3.854 63.926 3.906 63.962 ;
      RECT 3.854 65.126 3.906 65.162 ;
      RECT 3.854 66.326 3.906 66.362 ;
      RECT 3.854 67.526 3.906 67.562 ;
      RECT 3.854 68.726 3.906 68.762 ;
      RECT 3.854 69.926 3.906 69.962 ;
      RECT 3.854 71.126 3.906 71.162 ;
      RECT 3.934 1.558 3.986 1.594 ;
      RECT 3.934 2.758 3.986 2.794 ;
      RECT 3.934 3.958 3.986 3.994 ;
      RECT 3.934 5.158 3.986 5.194 ;
      RECT 3.934 6.358 3.986 6.394 ;
      RECT 3.934 7.558 3.986 7.594 ;
      RECT 3.934 8.758 3.986 8.794 ;
      RECT 3.934 9.958 3.986 9.994 ;
      RECT 3.934 11.158 3.986 11.194 ;
      RECT 3.934 12.358 3.986 12.394 ;
      RECT 3.934 13.558 3.986 13.594 ;
      RECT 3.934 14.758 3.986 14.794 ;
      RECT 3.934 15.958 3.986 15.994 ;
      RECT 3.934 17.158 3.986 17.194 ;
      RECT 3.934 18.358 3.986 18.394 ;
      RECT 3.934 19.558 3.986 19.594 ;
      RECT 3.934 20.758 3.986 20.794 ;
      RECT 3.934 21.958 3.986 21.994 ;
      RECT 3.934 23.158 3.986 23.194 ;
      RECT 3.934 24.358 3.986 24.394 ;
      RECT 3.934 25.558 3.986 25.594 ;
      RECT 3.934 26.758 3.986 26.794 ;
      RECT 3.934 27.958 3.986 27.994 ;
      RECT 3.934 29.158 3.986 29.194 ;
      RECT 3.934 30.358 3.986 30.394 ;
      RECT 3.934 31.558 3.986 31.594 ;
      RECT 3.934 33.342 3.986 33.378 ;
      RECT 3.934 33.582 3.986 33.618 ;
      RECT 3.934 37.902 3.986 37.938 ;
      RECT 3.934 38.142 3.986 38.178 ;
      RECT 3.934 40.678 3.986 40.714 ;
      RECT 3.934 41.878 3.986 41.914 ;
      RECT 3.934 43.078 3.986 43.114 ;
      RECT 3.934 44.278 3.986 44.314 ;
      RECT 3.934 45.478 3.986 45.514 ;
      RECT 3.934 46.678 3.986 46.714 ;
      RECT 3.934 47.878 3.986 47.914 ;
      RECT 3.934 49.078 3.986 49.114 ;
      RECT 3.934 50.278 3.986 50.314 ;
      RECT 3.934 51.478 3.986 51.514 ;
      RECT 3.934 52.678 3.986 52.714 ;
      RECT 3.934 53.878 3.986 53.914 ;
      RECT 3.934 55.078 3.986 55.114 ;
      RECT 3.934 56.278 3.986 56.314 ;
      RECT 3.934 57.478 3.986 57.514 ;
      RECT 3.934 58.678 3.986 58.714 ;
      RECT 3.934 59.878 3.986 59.914 ;
      RECT 3.934 61.078 3.986 61.114 ;
      RECT 3.934 62.278 3.986 62.314 ;
      RECT 3.934 63.478 3.986 63.514 ;
      RECT 3.934 64.678 3.986 64.714 ;
      RECT 3.934 65.878 3.986 65.914 ;
      RECT 3.934 67.078 3.986 67.114 ;
      RECT 3.934 68.278 3.986 68.314 ;
      RECT 3.934 69.478 3.986 69.514 ;
      RECT 3.934 70.678 3.986 70.714 ;
      RECT 3.934 71.878 3.986 71.914 ;
      RECT 4.014 0.806 4.066 0.842 ;
      RECT 4.014 2.006 4.066 2.042 ;
      RECT 4.014 3.206 4.066 3.242 ;
      RECT 4.014 4.406 4.066 4.442 ;
      RECT 4.014 5.606 4.066 5.642 ;
      RECT 4.014 6.806 4.066 6.842 ;
      RECT 4.014 8.006 4.066 8.042 ;
      RECT 4.014 9.206 4.066 9.242 ;
      RECT 4.014 10.406 4.066 10.442 ;
      RECT 4.014 11.606 4.066 11.642 ;
      RECT 4.014 12.806 4.066 12.842 ;
      RECT 4.014 14.006 4.066 14.042 ;
      RECT 4.014 15.206 4.066 15.242 ;
      RECT 4.014 16.406 4.066 16.442 ;
      RECT 4.014 17.606 4.066 17.642 ;
      RECT 4.014 18.806 4.066 18.842 ;
      RECT 4.014 20.006 4.066 20.042 ;
      RECT 4.014 21.206 4.066 21.242 ;
      RECT 4.014 22.406 4.066 22.442 ;
      RECT 4.014 23.606 4.066 23.642 ;
      RECT 4.014 24.806 4.066 24.842 ;
      RECT 4.014 26.006 4.066 26.042 ;
      RECT 4.014 27.206 4.066 27.242 ;
      RECT 4.014 28.406 4.066 28.442 ;
      RECT 4.014 29.606 4.066 29.642 ;
      RECT 4.014 30.806 4.066 30.842 ;
      RECT 4.014 32.622 4.066 32.658 ;
      RECT 4.014 32.862 4.066 32.898 ;
      RECT 4.014 38.622 4.066 38.658 ;
      RECT 4.014 38.862 4.066 38.898 ;
      RECT 4.014 39.926 4.066 39.962 ;
      RECT 4.014 41.126 4.066 41.162 ;
      RECT 4.014 42.326 4.066 42.362 ;
      RECT 4.014 43.526 4.066 43.562 ;
      RECT 4.014 44.726 4.066 44.762 ;
      RECT 4.014 45.926 4.066 45.962 ;
      RECT 4.014 47.126 4.066 47.162 ;
      RECT 4.014 48.326 4.066 48.362 ;
      RECT 4.014 49.526 4.066 49.562 ;
      RECT 4.014 50.726 4.066 50.762 ;
      RECT 4.014 51.926 4.066 51.962 ;
      RECT 4.014 53.126 4.066 53.162 ;
      RECT 4.014 54.326 4.066 54.362 ;
      RECT 4.014 55.526 4.066 55.562 ;
      RECT 4.014 56.726 4.066 56.762 ;
      RECT 4.014 57.926 4.066 57.962 ;
      RECT 4.014 59.126 4.066 59.162 ;
      RECT 4.014 60.326 4.066 60.362 ;
      RECT 4.014 61.526 4.066 61.562 ;
      RECT 4.014 62.726 4.066 62.762 ;
      RECT 4.014 63.926 4.066 63.962 ;
      RECT 4.014 65.126 4.066 65.162 ;
      RECT 4.014 66.326 4.066 66.362 ;
      RECT 4.014 67.526 4.066 67.562 ;
      RECT 4.014 68.726 4.066 68.762 ;
      RECT 4.014 69.926 4.066 69.962 ;
      RECT 4.014 71.126 4.066 71.162 ;
      RECT 4.094 1.558 4.146 1.594 ;
      RECT 4.094 2.758 4.146 2.794 ;
      RECT 4.094 3.958 4.146 3.994 ;
      RECT 4.094 5.158 4.146 5.194 ;
      RECT 4.094 6.358 4.146 6.394 ;
      RECT 4.094 7.558 4.146 7.594 ;
      RECT 4.094 8.758 4.146 8.794 ;
      RECT 4.094 9.958 4.146 9.994 ;
      RECT 4.094 11.158 4.146 11.194 ;
      RECT 4.094 12.358 4.146 12.394 ;
      RECT 4.094 13.558 4.146 13.594 ;
      RECT 4.094 14.758 4.146 14.794 ;
      RECT 4.094 15.958 4.146 15.994 ;
      RECT 4.094 17.158 4.146 17.194 ;
      RECT 4.094 18.358 4.146 18.394 ;
      RECT 4.094 19.558 4.146 19.594 ;
      RECT 4.094 20.758 4.146 20.794 ;
      RECT 4.094 21.958 4.146 21.994 ;
      RECT 4.094 23.158 4.146 23.194 ;
      RECT 4.094 24.358 4.146 24.394 ;
      RECT 4.094 25.558 4.146 25.594 ;
      RECT 4.094 26.758 4.146 26.794 ;
      RECT 4.094 27.958 4.146 27.994 ;
      RECT 4.094 29.158 4.146 29.194 ;
      RECT 4.094 30.358 4.146 30.394 ;
      RECT 4.094 31.558 4.146 31.594 ;
      RECT 4.094 33.342 4.146 33.378 ;
      RECT 4.094 33.582 4.146 33.618 ;
      RECT 4.094 37.902 4.146 37.938 ;
      RECT 4.094 38.142 4.146 38.178 ;
      RECT 4.094 40.678 4.146 40.714 ;
      RECT 4.094 41.878 4.146 41.914 ;
      RECT 4.094 43.078 4.146 43.114 ;
      RECT 4.094 44.278 4.146 44.314 ;
      RECT 4.094 45.478 4.146 45.514 ;
      RECT 4.094 46.678 4.146 46.714 ;
      RECT 4.094 47.878 4.146 47.914 ;
      RECT 4.094 49.078 4.146 49.114 ;
      RECT 4.094 50.278 4.146 50.314 ;
      RECT 4.094 51.478 4.146 51.514 ;
      RECT 4.094 52.678 4.146 52.714 ;
      RECT 4.094 53.878 4.146 53.914 ;
      RECT 4.094 55.078 4.146 55.114 ;
      RECT 4.094 56.278 4.146 56.314 ;
      RECT 4.094 57.478 4.146 57.514 ;
      RECT 4.094 58.678 4.146 58.714 ;
      RECT 4.094 59.878 4.146 59.914 ;
      RECT 4.094 61.078 4.146 61.114 ;
      RECT 4.094 62.278 4.146 62.314 ;
      RECT 4.094 63.478 4.146 63.514 ;
      RECT 4.094 64.678 4.146 64.714 ;
      RECT 4.094 65.878 4.146 65.914 ;
      RECT 4.094 67.078 4.146 67.114 ;
      RECT 4.094 68.278 4.146 68.314 ;
      RECT 4.094 69.478 4.146 69.514 ;
      RECT 4.094 70.678 4.146 70.714 ;
      RECT 4.094 71.878 4.146 71.914 ;
      RECT 4.174 0.281 4.226 0.317 ;
      RECT 4.174 72.403 4.226 72.439 ;
      RECT 4.254 0.806 4.306 0.842 ;
      RECT 4.254 2.006 4.306 2.042 ;
      RECT 4.254 3.206 4.306 3.242 ;
      RECT 4.254 4.406 4.306 4.442 ;
      RECT 4.254 5.606 4.306 5.642 ;
      RECT 4.254 6.806 4.306 6.842 ;
      RECT 4.254 8.006 4.306 8.042 ;
      RECT 4.254 9.206 4.306 9.242 ;
      RECT 4.254 10.406 4.306 10.442 ;
      RECT 4.254 11.606 4.306 11.642 ;
      RECT 4.254 12.806 4.306 12.842 ;
      RECT 4.254 14.006 4.306 14.042 ;
      RECT 4.254 15.206 4.306 15.242 ;
      RECT 4.254 16.406 4.306 16.442 ;
      RECT 4.254 17.606 4.306 17.642 ;
      RECT 4.254 18.806 4.306 18.842 ;
      RECT 4.254 20.006 4.306 20.042 ;
      RECT 4.254 21.206 4.306 21.242 ;
      RECT 4.254 22.406 4.306 22.442 ;
      RECT 4.254 23.606 4.306 23.642 ;
      RECT 4.254 24.806 4.306 24.842 ;
      RECT 4.254 26.006 4.306 26.042 ;
      RECT 4.254 27.206 4.306 27.242 ;
      RECT 4.254 28.406 4.306 28.442 ;
      RECT 4.254 29.606 4.306 29.642 ;
      RECT 4.254 30.806 4.306 30.842 ;
      RECT 4.254 32.622 4.306 32.658 ;
      RECT 4.254 32.862 4.306 32.898 ;
      RECT 4.254 34.302 4.306 34.338 ;
      RECT 4.254 34.782 4.306 34.818 ;
      RECT 4.254 36.702 4.306 36.738 ;
      RECT 4.254 37.182 4.306 37.218 ;
      RECT 4.254 38.622 4.306 38.658 ;
      RECT 4.254 38.862 4.306 38.898 ;
      RECT 4.254 39.926 4.306 39.962 ;
      RECT 4.254 41.126 4.306 41.162 ;
      RECT 4.254 42.326 4.306 42.362 ;
      RECT 4.254 43.526 4.306 43.562 ;
      RECT 4.254 44.726 4.306 44.762 ;
      RECT 4.254 45.926 4.306 45.962 ;
      RECT 4.254 47.126 4.306 47.162 ;
      RECT 4.254 48.326 4.306 48.362 ;
      RECT 4.254 49.526 4.306 49.562 ;
      RECT 4.254 50.726 4.306 50.762 ;
      RECT 4.254 51.926 4.306 51.962 ;
      RECT 4.254 53.126 4.306 53.162 ;
      RECT 4.254 54.326 4.306 54.362 ;
      RECT 4.254 55.526 4.306 55.562 ;
      RECT 4.254 56.726 4.306 56.762 ;
      RECT 4.254 57.926 4.306 57.962 ;
      RECT 4.254 59.126 4.306 59.162 ;
      RECT 4.254 60.326 4.306 60.362 ;
      RECT 4.254 61.526 4.306 61.562 ;
      RECT 4.254 62.726 4.306 62.762 ;
      RECT 4.254 63.926 4.306 63.962 ;
      RECT 4.254 65.126 4.306 65.162 ;
      RECT 4.254 66.326 4.306 66.362 ;
      RECT 4.254 67.526 4.306 67.562 ;
      RECT 4.254 68.726 4.306 68.762 ;
      RECT 4.254 69.926 4.306 69.962 ;
      RECT 4.254 71.126 4.306 71.162 ;
      RECT 4.334 1.558 4.386 1.594 ;
      RECT 4.334 2.758 4.386 2.794 ;
      RECT 4.334 3.958 4.386 3.994 ;
      RECT 4.334 5.158 4.386 5.194 ;
      RECT 4.334 6.358 4.386 6.394 ;
      RECT 4.334 7.558 4.386 7.594 ;
      RECT 4.334 8.758 4.386 8.794 ;
      RECT 4.334 9.958 4.386 9.994 ;
      RECT 4.334 11.158 4.386 11.194 ;
      RECT 4.334 12.358 4.386 12.394 ;
      RECT 4.334 13.558 4.386 13.594 ;
      RECT 4.334 14.758 4.386 14.794 ;
      RECT 4.334 15.958 4.386 15.994 ;
      RECT 4.334 17.158 4.386 17.194 ;
      RECT 4.334 18.358 4.386 18.394 ;
      RECT 4.334 19.558 4.386 19.594 ;
      RECT 4.334 20.758 4.386 20.794 ;
      RECT 4.334 21.958 4.386 21.994 ;
      RECT 4.334 23.158 4.386 23.194 ;
      RECT 4.334 24.358 4.386 24.394 ;
      RECT 4.334 25.558 4.386 25.594 ;
      RECT 4.334 26.758 4.386 26.794 ;
      RECT 4.334 27.958 4.386 27.994 ;
      RECT 4.334 29.158 4.386 29.194 ;
      RECT 4.334 30.358 4.386 30.394 ;
      RECT 4.334 31.558 4.386 31.594 ;
      RECT 4.334 33.342 4.386 33.378 ;
      RECT 4.334 33.582 4.386 33.618 ;
      RECT 4.334 37.902 4.386 37.938 ;
      RECT 4.334 38.142 4.386 38.178 ;
      RECT 4.334 40.678 4.386 40.714 ;
      RECT 4.334 41.878 4.386 41.914 ;
      RECT 4.334 43.078 4.386 43.114 ;
      RECT 4.334 44.278 4.386 44.314 ;
      RECT 4.334 45.478 4.386 45.514 ;
      RECT 4.334 46.678 4.386 46.714 ;
      RECT 4.334 47.878 4.386 47.914 ;
      RECT 4.334 49.078 4.386 49.114 ;
      RECT 4.334 50.278 4.386 50.314 ;
      RECT 4.334 51.478 4.386 51.514 ;
      RECT 4.334 52.678 4.386 52.714 ;
      RECT 4.334 53.878 4.386 53.914 ;
      RECT 4.334 55.078 4.386 55.114 ;
      RECT 4.334 56.278 4.386 56.314 ;
      RECT 4.334 57.478 4.386 57.514 ;
      RECT 4.334 58.678 4.386 58.714 ;
      RECT 4.334 59.878 4.386 59.914 ;
      RECT 4.334 61.078 4.386 61.114 ;
      RECT 4.334 62.278 4.386 62.314 ;
      RECT 4.334 63.478 4.386 63.514 ;
      RECT 4.334 64.678 4.386 64.714 ;
      RECT 4.334 65.878 4.386 65.914 ;
      RECT 4.334 67.078 4.386 67.114 ;
      RECT 4.334 68.278 4.386 68.314 ;
      RECT 4.334 69.478 4.386 69.514 ;
      RECT 4.334 70.678 4.386 70.714 ;
      RECT 4.334 71.878 4.386 71.914 ;
      RECT 4.414 0.806 4.466 0.842 ;
      RECT 4.414 2.006 4.466 2.042 ;
      RECT 4.414 3.206 4.466 3.242 ;
      RECT 4.414 4.406 4.466 4.442 ;
      RECT 4.414 5.606 4.466 5.642 ;
      RECT 4.414 6.806 4.466 6.842 ;
      RECT 4.414 8.006 4.466 8.042 ;
      RECT 4.414 9.206 4.466 9.242 ;
      RECT 4.414 10.406 4.466 10.442 ;
      RECT 4.414 11.606 4.466 11.642 ;
      RECT 4.414 12.806 4.466 12.842 ;
      RECT 4.414 14.006 4.466 14.042 ;
      RECT 4.414 15.206 4.466 15.242 ;
      RECT 4.414 16.406 4.466 16.442 ;
      RECT 4.414 17.606 4.466 17.642 ;
      RECT 4.414 18.806 4.466 18.842 ;
      RECT 4.414 20.006 4.466 20.042 ;
      RECT 4.414 21.206 4.466 21.242 ;
      RECT 4.414 22.406 4.466 22.442 ;
      RECT 4.414 23.606 4.466 23.642 ;
      RECT 4.414 24.806 4.466 24.842 ;
      RECT 4.414 26.006 4.466 26.042 ;
      RECT 4.414 27.206 4.466 27.242 ;
      RECT 4.414 28.406 4.466 28.442 ;
      RECT 4.414 29.606 4.466 29.642 ;
      RECT 4.414 30.806 4.466 30.842 ;
      RECT 4.414 32.622 4.466 32.658 ;
      RECT 4.414 32.862 4.466 32.898 ;
      RECT 4.414 38.622 4.466 38.658 ;
      RECT 4.414 38.862 4.466 38.898 ;
      RECT 4.414 39.926 4.466 39.962 ;
      RECT 4.414 41.126 4.466 41.162 ;
      RECT 4.414 42.326 4.466 42.362 ;
      RECT 4.414 43.526 4.466 43.562 ;
      RECT 4.414 44.726 4.466 44.762 ;
      RECT 4.414 45.926 4.466 45.962 ;
      RECT 4.414 47.126 4.466 47.162 ;
      RECT 4.414 48.326 4.466 48.362 ;
      RECT 4.414 49.526 4.466 49.562 ;
      RECT 4.414 50.726 4.466 50.762 ;
      RECT 4.414 51.926 4.466 51.962 ;
      RECT 4.414 53.126 4.466 53.162 ;
      RECT 4.414 54.326 4.466 54.362 ;
      RECT 4.414 55.526 4.466 55.562 ;
      RECT 4.414 56.726 4.466 56.762 ;
      RECT 4.414 57.926 4.466 57.962 ;
      RECT 4.414 59.126 4.466 59.162 ;
      RECT 4.414 60.326 4.466 60.362 ;
      RECT 4.414 61.526 4.466 61.562 ;
      RECT 4.414 62.726 4.466 62.762 ;
      RECT 4.414 63.926 4.466 63.962 ;
      RECT 4.414 65.126 4.466 65.162 ;
      RECT 4.414 66.326 4.466 66.362 ;
      RECT 4.414 67.526 4.466 67.562 ;
      RECT 4.414 68.726 4.466 68.762 ;
      RECT 4.414 69.926 4.466 69.962 ;
      RECT 4.414 71.126 4.466 71.162 ;
      RECT 4.494 1.558 4.546 1.594 ;
      RECT 4.494 2.758 4.546 2.794 ;
      RECT 4.494 3.958 4.546 3.994 ;
      RECT 4.494 5.158 4.546 5.194 ;
      RECT 4.494 6.358 4.546 6.394 ;
      RECT 4.494 7.558 4.546 7.594 ;
      RECT 4.494 8.758 4.546 8.794 ;
      RECT 4.494 9.958 4.546 9.994 ;
      RECT 4.494 11.158 4.546 11.194 ;
      RECT 4.494 12.358 4.546 12.394 ;
      RECT 4.494 13.558 4.546 13.594 ;
      RECT 4.494 14.758 4.546 14.794 ;
      RECT 4.494 15.958 4.546 15.994 ;
      RECT 4.494 17.158 4.546 17.194 ;
      RECT 4.494 18.358 4.546 18.394 ;
      RECT 4.494 19.558 4.546 19.594 ;
      RECT 4.494 20.758 4.546 20.794 ;
      RECT 4.494 21.958 4.546 21.994 ;
      RECT 4.494 23.158 4.546 23.194 ;
      RECT 4.494 24.358 4.546 24.394 ;
      RECT 4.494 25.558 4.546 25.594 ;
      RECT 4.494 26.758 4.546 26.794 ;
      RECT 4.494 27.958 4.546 27.994 ;
      RECT 4.494 29.158 4.546 29.194 ;
      RECT 4.494 30.358 4.546 30.394 ;
      RECT 4.494 31.558 4.546 31.594 ;
      RECT 4.494 33.342 4.546 33.378 ;
      RECT 4.494 33.582 4.546 33.618 ;
      RECT 4.494 37.902 4.546 37.938 ;
      RECT 4.494 38.142 4.546 38.178 ;
      RECT 4.494 40.678 4.546 40.714 ;
      RECT 4.494 41.878 4.546 41.914 ;
      RECT 4.494 43.078 4.546 43.114 ;
      RECT 4.494 44.278 4.546 44.314 ;
      RECT 4.494 45.478 4.546 45.514 ;
      RECT 4.494 46.678 4.546 46.714 ;
      RECT 4.494 47.878 4.546 47.914 ;
      RECT 4.494 49.078 4.546 49.114 ;
      RECT 4.494 50.278 4.546 50.314 ;
      RECT 4.494 51.478 4.546 51.514 ;
      RECT 4.494 52.678 4.546 52.714 ;
      RECT 4.494 53.878 4.546 53.914 ;
      RECT 4.494 55.078 4.546 55.114 ;
      RECT 4.494 56.278 4.546 56.314 ;
      RECT 4.494 57.478 4.546 57.514 ;
      RECT 4.494 58.678 4.546 58.714 ;
      RECT 4.494 59.878 4.546 59.914 ;
      RECT 4.494 61.078 4.546 61.114 ;
      RECT 4.494 62.278 4.546 62.314 ;
      RECT 4.494 63.478 4.546 63.514 ;
      RECT 4.494 64.678 4.546 64.714 ;
      RECT 4.494 65.878 4.546 65.914 ;
      RECT 4.494 67.078 4.546 67.114 ;
      RECT 4.494 68.278 4.546 68.314 ;
      RECT 4.494 69.478 4.546 69.514 ;
      RECT 4.494 70.678 4.546 70.714 ;
      RECT 4.494 71.878 4.546 71.914 ;
      RECT 4.574 0.281 4.626 0.317 ;
      RECT 4.574 72.403 4.626 72.439 ;
      RECT 4.654 0.806 4.706 0.842 ;
      RECT 4.654 2.006 4.706 2.042 ;
      RECT 4.654 3.206 4.706 3.242 ;
      RECT 4.654 4.406 4.706 4.442 ;
      RECT 4.654 5.606 4.706 5.642 ;
      RECT 4.654 6.806 4.706 6.842 ;
      RECT 4.654 8.006 4.706 8.042 ;
      RECT 4.654 9.206 4.706 9.242 ;
      RECT 4.654 10.406 4.706 10.442 ;
      RECT 4.654 11.606 4.706 11.642 ;
      RECT 4.654 12.806 4.706 12.842 ;
      RECT 4.654 14.006 4.706 14.042 ;
      RECT 4.654 15.206 4.706 15.242 ;
      RECT 4.654 16.406 4.706 16.442 ;
      RECT 4.654 17.606 4.706 17.642 ;
      RECT 4.654 18.806 4.706 18.842 ;
      RECT 4.654 20.006 4.706 20.042 ;
      RECT 4.654 21.206 4.706 21.242 ;
      RECT 4.654 22.406 4.706 22.442 ;
      RECT 4.654 23.606 4.706 23.642 ;
      RECT 4.654 24.806 4.706 24.842 ;
      RECT 4.654 26.006 4.706 26.042 ;
      RECT 4.654 27.206 4.706 27.242 ;
      RECT 4.654 28.406 4.706 28.442 ;
      RECT 4.654 29.606 4.706 29.642 ;
      RECT 4.654 30.806 4.706 30.842 ;
      RECT 4.654 32.622 4.706 32.658 ;
      RECT 4.654 32.862 4.706 32.898 ;
      RECT 4.654 38.622 4.706 38.658 ;
      RECT 4.654 38.862 4.706 38.898 ;
      RECT 4.654 39.926 4.706 39.962 ;
      RECT 4.654 41.126 4.706 41.162 ;
      RECT 4.654 42.326 4.706 42.362 ;
      RECT 4.654 43.526 4.706 43.562 ;
      RECT 4.654 44.726 4.706 44.762 ;
      RECT 4.654 45.926 4.706 45.962 ;
      RECT 4.654 47.126 4.706 47.162 ;
      RECT 4.654 48.326 4.706 48.362 ;
      RECT 4.654 49.526 4.706 49.562 ;
      RECT 4.654 50.726 4.706 50.762 ;
      RECT 4.654 51.926 4.706 51.962 ;
      RECT 4.654 53.126 4.706 53.162 ;
      RECT 4.654 54.326 4.706 54.362 ;
      RECT 4.654 55.526 4.706 55.562 ;
      RECT 4.654 56.726 4.706 56.762 ;
      RECT 4.654 57.926 4.706 57.962 ;
      RECT 4.654 59.126 4.706 59.162 ;
      RECT 4.654 60.326 4.706 60.362 ;
      RECT 4.654 61.526 4.706 61.562 ;
      RECT 4.654 62.726 4.706 62.762 ;
      RECT 4.654 63.926 4.706 63.962 ;
      RECT 4.654 65.126 4.706 65.162 ;
      RECT 4.654 66.326 4.706 66.362 ;
      RECT 4.654 67.526 4.706 67.562 ;
      RECT 4.654 68.726 4.706 68.762 ;
      RECT 4.654 69.926 4.706 69.962 ;
      RECT 4.654 71.126 4.706 71.162 ;
      RECT 4.734 1.558 4.786 1.594 ;
      RECT 4.734 2.758 4.786 2.794 ;
      RECT 4.734 3.958 4.786 3.994 ;
      RECT 4.734 5.158 4.786 5.194 ;
      RECT 4.734 6.358 4.786 6.394 ;
      RECT 4.734 7.558 4.786 7.594 ;
      RECT 4.734 8.758 4.786 8.794 ;
      RECT 4.734 9.958 4.786 9.994 ;
      RECT 4.734 11.158 4.786 11.194 ;
      RECT 4.734 12.358 4.786 12.394 ;
      RECT 4.734 13.558 4.786 13.594 ;
      RECT 4.734 14.758 4.786 14.794 ;
      RECT 4.734 15.958 4.786 15.994 ;
      RECT 4.734 17.158 4.786 17.194 ;
      RECT 4.734 18.358 4.786 18.394 ;
      RECT 4.734 19.558 4.786 19.594 ;
      RECT 4.734 20.758 4.786 20.794 ;
      RECT 4.734 21.958 4.786 21.994 ;
      RECT 4.734 23.158 4.786 23.194 ;
      RECT 4.734 24.358 4.786 24.394 ;
      RECT 4.734 25.558 4.786 25.594 ;
      RECT 4.734 26.758 4.786 26.794 ;
      RECT 4.734 27.958 4.786 27.994 ;
      RECT 4.734 29.158 4.786 29.194 ;
      RECT 4.734 30.358 4.786 30.394 ;
      RECT 4.734 31.558 4.786 31.594 ;
      RECT 4.734 33.342 4.786 33.378 ;
      RECT 4.734 33.582 4.786 33.618 ;
      RECT 4.734 37.902 4.786 37.938 ;
      RECT 4.734 38.142 4.786 38.178 ;
      RECT 4.734 40.678 4.786 40.714 ;
      RECT 4.734 41.878 4.786 41.914 ;
      RECT 4.734 43.078 4.786 43.114 ;
      RECT 4.734 44.278 4.786 44.314 ;
      RECT 4.734 45.478 4.786 45.514 ;
      RECT 4.734 46.678 4.786 46.714 ;
      RECT 4.734 47.878 4.786 47.914 ;
      RECT 4.734 49.078 4.786 49.114 ;
      RECT 4.734 50.278 4.786 50.314 ;
      RECT 4.734 51.478 4.786 51.514 ;
      RECT 4.734 52.678 4.786 52.714 ;
      RECT 4.734 53.878 4.786 53.914 ;
      RECT 4.734 55.078 4.786 55.114 ;
      RECT 4.734 56.278 4.786 56.314 ;
      RECT 4.734 57.478 4.786 57.514 ;
      RECT 4.734 58.678 4.786 58.714 ;
      RECT 4.734 59.878 4.786 59.914 ;
      RECT 4.734 61.078 4.786 61.114 ;
      RECT 4.734 62.278 4.786 62.314 ;
      RECT 4.734 63.478 4.786 63.514 ;
      RECT 4.734 64.678 4.786 64.714 ;
      RECT 4.734 65.878 4.786 65.914 ;
      RECT 4.734 67.078 4.786 67.114 ;
      RECT 4.734 68.278 4.786 68.314 ;
      RECT 4.734 69.478 4.786 69.514 ;
      RECT 4.734 70.678 4.786 70.714 ;
      RECT 4.734 71.878 4.786 71.914 ;
      RECT 4.814 0.806 4.866 0.842 ;
      RECT 4.814 2.006 4.866 2.042 ;
      RECT 4.814 3.206 4.866 3.242 ;
      RECT 4.814 4.406 4.866 4.442 ;
      RECT 4.814 5.606 4.866 5.642 ;
      RECT 4.814 6.806 4.866 6.842 ;
      RECT 4.814 8.006 4.866 8.042 ;
      RECT 4.814 9.206 4.866 9.242 ;
      RECT 4.814 10.406 4.866 10.442 ;
      RECT 4.814 11.606 4.866 11.642 ;
      RECT 4.814 12.806 4.866 12.842 ;
      RECT 4.814 14.006 4.866 14.042 ;
      RECT 4.814 15.206 4.866 15.242 ;
      RECT 4.814 16.406 4.866 16.442 ;
      RECT 4.814 17.606 4.866 17.642 ;
      RECT 4.814 18.806 4.866 18.842 ;
      RECT 4.814 20.006 4.866 20.042 ;
      RECT 4.814 21.206 4.866 21.242 ;
      RECT 4.814 22.406 4.866 22.442 ;
      RECT 4.814 23.606 4.866 23.642 ;
      RECT 4.814 24.806 4.866 24.842 ;
      RECT 4.814 26.006 4.866 26.042 ;
      RECT 4.814 27.206 4.866 27.242 ;
      RECT 4.814 28.406 4.866 28.442 ;
      RECT 4.814 29.606 4.866 29.642 ;
      RECT 4.814 30.806 4.866 30.842 ;
      RECT 4.814 32.622 4.866 32.658 ;
      RECT 4.814 32.862 4.866 32.898 ;
      RECT 4.814 38.622 4.866 38.658 ;
      RECT 4.814 38.862 4.866 38.898 ;
      RECT 4.814 39.926 4.866 39.962 ;
      RECT 4.814 41.126 4.866 41.162 ;
      RECT 4.814 42.326 4.866 42.362 ;
      RECT 4.814 43.526 4.866 43.562 ;
      RECT 4.814 44.726 4.866 44.762 ;
      RECT 4.814 45.926 4.866 45.962 ;
      RECT 4.814 47.126 4.866 47.162 ;
      RECT 4.814 48.326 4.866 48.362 ;
      RECT 4.814 49.526 4.866 49.562 ;
      RECT 4.814 50.726 4.866 50.762 ;
      RECT 4.814 51.926 4.866 51.962 ;
      RECT 4.814 53.126 4.866 53.162 ;
      RECT 4.814 54.326 4.866 54.362 ;
      RECT 4.814 55.526 4.866 55.562 ;
      RECT 4.814 56.726 4.866 56.762 ;
      RECT 4.814 57.926 4.866 57.962 ;
      RECT 4.814 59.126 4.866 59.162 ;
      RECT 4.814 60.326 4.866 60.362 ;
      RECT 4.814 61.526 4.866 61.562 ;
      RECT 4.814 62.726 4.866 62.762 ;
      RECT 4.814 63.926 4.866 63.962 ;
      RECT 4.814 65.126 4.866 65.162 ;
      RECT 4.814 66.326 4.866 66.362 ;
      RECT 4.814 67.526 4.866 67.562 ;
      RECT 4.814 68.726 4.866 68.762 ;
      RECT 4.814 69.926 4.866 69.962 ;
      RECT 4.814 71.126 4.866 71.162 ;
      RECT 4.894 1.558 4.946 1.594 ;
      RECT 4.894 2.758 4.946 2.794 ;
      RECT 4.894 3.958 4.946 3.994 ;
      RECT 4.894 5.158 4.946 5.194 ;
      RECT 4.894 6.358 4.946 6.394 ;
      RECT 4.894 7.558 4.946 7.594 ;
      RECT 4.894 8.758 4.946 8.794 ;
      RECT 4.894 9.958 4.946 9.994 ;
      RECT 4.894 11.158 4.946 11.194 ;
      RECT 4.894 12.358 4.946 12.394 ;
      RECT 4.894 13.558 4.946 13.594 ;
      RECT 4.894 14.758 4.946 14.794 ;
      RECT 4.894 15.958 4.946 15.994 ;
      RECT 4.894 17.158 4.946 17.194 ;
      RECT 4.894 18.358 4.946 18.394 ;
      RECT 4.894 19.558 4.946 19.594 ;
      RECT 4.894 20.758 4.946 20.794 ;
      RECT 4.894 21.958 4.946 21.994 ;
      RECT 4.894 23.158 4.946 23.194 ;
      RECT 4.894 24.358 4.946 24.394 ;
      RECT 4.894 25.558 4.946 25.594 ;
      RECT 4.894 26.758 4.946 26.794 ;
      RECT 4.894 27.958 4.946 27.994 ;
      RECT 4.894 29.158 4.946 29.194 ;
      RECT 4.894 30.358 4.946 30.394 ;
      RECT 4.894 31.558 4.946 31.594 ;
      RECT 4.894 33.342 4.946 33.378 ;
      RECT 4.894 33.582 4.946 33.618 ;
      RECT 4.894 37.902 4.946 37.938 ;
      RECT 4.894 38.142 4.946 38.178 ;
      RECT 4.894 40.678 4.946 40.714 ;
      RECT 4.894 41.878 4.946 41.914 ;
      RECT 4.894 43.078 4.946 43.114 ;
      RECT 4.894 44.278 4.946 44.314 ;
      RECT 4.894 45.478 4.946 45.514 ;
      RECT 4.894 46.678 4.946 46.714 ;
      RECT 4.894 47.878 4.946 47.914 ;
      RECT 4.894 49.078 4.946 49.114 ;
      RECT 4.894 50.278 4.946 50.314 ;
      RECT 4.894 51.478 4.946 51.514 ;
      RECT 4.894 52.678 4.946 52.714 ;
      RECT 4.894 53.878 4.946 53.914 ;
      RECT 4.894 55.078 4.946 55.114 ;
      RECT 4.894 56.278 4.946 56.314 ;
      RECT 4.894 57.478 4.946 57.514 ;
      RECT 4.894 58.678 4.946 58.714 ;
      RECT 4.894 59.878 4.946 59.914 ;
      RECT 4.894 61.078 4.946 61.114 ;
      RECT 4.894 62.278 4.946 62.314 ;
      RECT 4.894 63.478 4.946 63.514 ;
      RECT 4.894 64.678 4.946 64.714 ;
      RECT 4.894 65.878 4.946 65.914 ;
      RECT 4.894 67.078 4.946 67.114 ;
      RECT 4.894 68.278 4.946 68.314 ;
      RECT 4.894 69.478 4.946 69.514 ;
      RECT 4.894 70.678 4.946 70.714 ;
      RECT 4.894 71.878 4.946 71.914 ;
      RECT 4.974 0.281 5.026 0.317 ;
      RECT 4.974 72.403 5.026 72.439 ;
      RECT 5.054 0.806 5.106 0.842 ;
      RECT 5.054 2.006 5.106 2.042 ;
      RECT 5.054 3.206 5.106 3.242 ;
      RECT 5.054 4.406 5.106 4.442 ;
      RECT 5.054 5.606 5.106 5.642 ;
      RECT 5.054 6.806 5.106 6.842 ;
      RECT 5.054 8.006 5.106 8.042 ;
      RECT 5.054 9.206 5.106 9.242 ;
      RECT 5.054 10.406 5.106 10.442 ;
      RECT 5.054 11.606 5.106 11.642 ;
      RECT 5.054 12.806 5.106 12.842 ;
      RECT 5.054 14.006 5.106 14.042 ;
      RECT 5.054 15.206 5.106 15.242 ;
      RECT 5.054 16.406 5.106 16.442 ;
      RECT 5.054 17.606 5.106 17.642 ;
      RECT 5.054 18.806 5.106 18.842 ;
      RECT 5.054 20.006 5.106 20.042 ;
      RECT 5.054 21.206 5.106 21.242 ;
      RECT 5.054 22.406 5.106 22.442 ;
      RECT 5.054 23.606 5.106 23.642 ;
      RECT 5.054 24.806 5.106 24.842 ;
      RECT 5.054 26.006 5.106 26.042 ;
      RECT 5.054 27.206 5.106 27.242 ;
      RECT 5.054 28.406 5.106 28.442 ;
      RECT 5.054 29.606 5.106 29.642 ;
      RECT 5.054 30.806 5.106 30.842 ;
      RECT 5.054 32.622 5.106 32.658 ;
      RECT 5.054 32.862 5.106 32.898 ;
      RECT 5.054 34.302 5.106 34.338 ;
      RECT 5.054 34.782 5.106 34.818 ;
      RECT 5.054 36.702 5.106 36.738 ;
      RECT 5.054 37.182 5.106 37.218 ;
      RECT 5.054 38.622 5.106 38.658 ;
      RECT 5.054 38.862 5.106 38.898 ;
      RECT 5.054 39.926 5.106 39.962 ;
      RECT 5.054 41.126 5.106 41.162 ;
      RECT 5.054 42.326 5.106 42.362 ;
      RECT 5.054 43.526 5.106 43.562 ;
      RECT 5.054 44.726 5.106 44.762 ;
      RECT 5.054 45.926 5.106 45.962 ;
      RECT 5.054 47.126 5.106 47.162 ;
      RECT 5.054 48.326 5.106 48.362 ;
      RECT 5.054 49.526 5.106 49.562 ;
      RECT 5.054 50.726 5.106 50.762 ;
      RECT 5.054 51.926 5.106 51.962 ;
      RECT 5.054 53.126 5.106 53.162 ;
      RECT 5.054 54.326 5.106 54.362 ;
      RECT 5.054 55.526 5.106 55.562 ;
      RECT 5.054 56.726 5.106 56.762 ;
      RECT 5.054 57.926 5.106 57.962 ;
      RECT 5.054 59.126 5.106 59.162 ;
      RECT 5.054 60.326 5.106 60.362 ;
      RECT 5.054 61.526 5.106 61.562 ;
      RECT 5.054 62.726 5.106 62.762 ;
      RECT 5.054 63.926 5.106 63.962 ;
      RECT 5.054 65.126 5.106 65.162 ;
      RECT 5.054 66.326 5.106 66.362 ;
      RECT 5.054 67.526 5.106 67.562 ;
      RECT 5.054 68.726 5.106 68.762 ;
      RECT 5.054 69.926 5.106 69.962 ;
      RECT 5.054 71.126 5.106 71.162 ;
      RECT 5.134 1.558 5.186 1.594 ;
      RECT 5.134 2.758 5.186 2.794 ;
      RECT 5.134 3.958 5.186 3.994 ;
      RECT 5.134 5.158 5.186 5.194 ;
      RECT 5.134 6.358 5.186 6.394 ;
      RECT 5.134 7.558 5.186 7.594 ;
      RECT 5.134 8.758 5.186 8.794 ;
      RECT 5.134 9.958 5.186 9.994 ;
      RECT 5.134 11.158 5.186 11.194 ;
      RECT 5.134 12.358 5.186 12.394 ;
      RECT 5.134 13.558 5.186 13.594 ;
      RECT 5.134 14.758 5.186 14.794 ;
      RECT 5.134 15.958 5.186 15.994 ;
      RECT 5.134 17.158 5.186 17.194 ;
      RECT 5.134 18.358 5.186 18.394 ;
      RECT 5.134 19.558 5.186 19.594 ;
      RECT 5.134 20.758 5.186 20.794 ;
      RECT 5.134 21.958 5.186 21.994 ;
      RECT 5.134 23.158 5.186 23.194 ;
      RECT 5.134 24.358 5.186 24.394 ;
      RECT 5.134 25.558 5.186 25.594 ;
      RECT 5.134 26.758 5.186 26.794 ;
      RECT 5.134 27.958 5.186 27.994 ;
      RECT 5.134 29.158 5.186 29.194 ;
      RECT 5.134 30.358 5.186 30.394 ;
      RECT 5.134 31.558 5.186 31.594 ;
      RECT 5.134 33.342 5.186 33.378 ;
      RECT 5.134 33.582 5.186 33.618 ;
      RECT 5.134 37.902 5.186 37.938 ;
      RECT 5.134 38.142 5.186 38.178 ;
      RECT 5.134 40.678 5.186 40.714 ;
      RECT 5.134 41.878 5.186 41.914 ;
      RECT 5.134 43.078 5.186 43.114 ;
      RECT 5.134 44.278 5.186 44.314 ;
      RECT 5.134 45.478 5.186 45.514 ;
      RECT 5.134 46.678 5.186 46.714 ;
      RECT 5.134 47.878 5.186 47.914 ;
      RECT 5.134 49.078 5.186 49.114 ;
      RECT 5.134 50.278 5.186 50.314 ;
      RECT 5.134 51.478 5.186 51.514 ;
      RECT 5.134 52.678 5.186 52.714 ;
      RECT 5.134 53.878 5.186 53.914 ;
      RECT 5.134 55.078 5.186 55.114 ;
      RECT 5.134 56.278 5.186 56.314 ;
      RECT 5.134 57.478 5.186 57.514 ;
      RECT 5.134 58.678 5.186 58.714 ;
      RECT 5.134 59.878 5.186 59.914 ;
      RECT 5.134 61.078 5.186 61.114 ;
      RECT 5.134 62.278 5.186 62.314 ;
      RECT 5.134 63.478 5.186 63.514 ;
      RECT 5.134 64.678 5.186 64.714 ;
      RECT 5.134 65.878 5.186 65.914 ;
      RECT 5.134 67.078 5.186 67.114 ;
      RECT 5.134 68.278 5.186 68.314 ;
      RECT 5.134 69.478 5.186 69.514 ;
      RECT 5.134 70.678 5.186 70.714 ;
      RECT 5.134 71.878 5.186 71.914 ;
      RECT 5.214 0.806 5.266 0.842 ;
      RECT 5.214 2.006 5.266 2.042 ;
      RECT 5.214 3.206 5.266 3.242 ;
      RECT 5.214 4.406 5.266 4.442 ;
      RECT 5.214 5.606 5.266 5.642 ;
      RECT 5.214 6.806 5.266 6.842 ;
      RECT 5.214 8.006 5.266 8.042 ;
      RECT 5.214 9.206 5.266 9.242 ;
      RECT 5.214 10.406 5.266 10.442 ;
      RECT 5.214 11.606 5.266 11.642 ;
      RECT 5.214 12.806 5.266 12.842 ;
      RECT 5.214 14.006 5.266 14.042 ;
      RECT 5.214 15.206 5.266 15.242 ;
      RECT 5.214 16.406 5.266 16.442 ;
      RECT 5.214 17.606 5.266 17.642 ;
      RECT 5.214 18.806 5.266 18.842 ;
      RECT 5.214 20.006 5.266 20.042 ;
      RECT 5.214 21.206 5.266 21.242 ;
      RECT 5.214 22.406 5.266 22.442 ;
      RECT 5.214 23.606 5.266 23.642 ;
      RECT 5.214 24.806 5.266 24.842 ;
      RECT 5.214 26.006 5.266 26.042 ;
      RECT 5.214 27.206 5.266 27.242 ;
      RECT 5.214 28.406 5.266 28.442 ;
      RECT 5.214 29.606 5.266 29.642 ;
      RECT 5.214 30.806 5.266 30.842 ;
      RECT 5.214 32.622 5.266 32.658 ;
      RECT 5.214 32.862 5.266 32.898 ;
      RECT 5.214 38.622 5.266 38.658 ;
      RECT 5.214 38.862 5.266 38.898 ;
      RECT 5.214 39.926 5.266 39.962 ;
      RECT 5.214 41.126 5.266 41.162 ;
      RECT 5.214 42.326 5.266 42.362 ;
      RECT 5.214 43.526 5.266 43.562 ;
      RECT 5.214 44.726 5.266 44.762 ;
      RECT 5.214 45.926 5.266 45.962 ;
      RECT 5.214 47.126 5.266 47.162 ;
      RECT 5.214 48.326 5.266 48.362 ;
      RECT 5.214 49.526 5.266 49.562 ;
      RECT 5.214 50.726 5.266 50.762 ;
      RECT 5.214 51.926 5.266 51.962 ;
      RECT 5.214 53.126 5.266 53.162 ;
      RECT 5.214 54.326 5.266 54.362 ;
      RECT 5.214 55.526 5.266 55.562 ;
      RECT 5.214 56.726 5.266 56.762 ;
      RECT 5.214 57.926 5.266 57.962 ;
      RECT 5.214 59.126 5.266 59.162 ;
      RECT 5.214 60.326 5.266 60.362 ;
      RECT 5.214 61.526 5.266 61.562 ;
      RECT 5.214 62.726 5.266 62.762 ;
      RECT 5.214 63.926 5.266 63.962 ;
      RECT 5.214 65.126 5.266 65.162 ;
      RECT 5.214 66.326 5.266 66.362 ;
      RECT 5.214 67.526 5.266 67.562 ;
      RECT 5.214 68.726 5.266 68.762 ;
      RECT 5.214 69.926 5.266 69.962 ;
      RECT 5.214 71.126 5.266 71.162 ;
      RECT 5.294 1.558 5.346 1.594 ;
      RECT 5.294 2.758 5.346 2.794 ;
      RECT 5.294 3.958 5.346 3.994 ;
      RECT 5.294 5.158 5.346 5.194 ;
      RECT 5.294 6.358 5.346 6.394 ;
      RECT 5.294 7.558 5.346 7.594 ;
      RECT 5.294 8.758 5.346 8.794 ;
      RECT 5.294 9.958 5.346 9.994 ;
      RECT 5.294 11.158 5.346 11.194 ;
      RECT 5.294 12.358 5.346 12.394 ;
      RECT 5.294 13.558 5.346 13.594 ;
      RECT 5.294 14.758 5.346 14.794 ;
      RECT 5.294 15.958 5.346 15.994 ;
      RECT 5.294 17.158 5.346 17.194 ;
      RECT 5.294 18.358 5.346 18.394 ;
      RECT 5.294 19.558 5.346 19.594 ;
      RECT 5.294 20.758 5.346 20.794 ;
      RECT 5.294 21.958 5.346 21.994 ;
      RECT 5.294 23.158 5.346 23.194 ;
      RECT 5.294 24.358 5.346 24.394 ;
      RECT 5.294 25.558 5.346 25.594 ;
      RECT 5.294 26.758 5.346 26.794 ;
      RECT 5.294 27.958 5.346 27.994 ;
      RECT 5.294 29.158 5.346 29.194 ;
      RECT 5.294 30.358 5.346 30.394 ;
      RECT 5.294 31.558 5.346 31.594 ;
      RECT 5.294 33.342 5.346 33.378 ;
      RECT 5.294 33.582 5.346 33.618 ;
      RECT 5.294 37.902 5.346 37.938 ;
      RECT 5.294 38.142 5.346 38.178 ;
      RECT 5.294 40.678 5.346 40.714 ;
      RECT 5.294 41.878 5.346 41.914 ;
      RECT 5.294 43.078 5.346 43.114 ;
      RECT 5.294 44.278 5.346 44.314 ;
      RECT 5.294 45.478 5.346 45.514 ;
      RECT 5.294 46.678 5.346 46.714 ;
      RECT 5.294 47.878 5.346 47.914 ;
      RECT 5.294 49.078 5.346 49.114 ;
      RECT 5.294 50.278 5.346 50.314 ;
      RECT 5.294 51.478 5.346 51.514 ;
      RECT 5.294 52.678 5.346 52.714 ;
      RECT 5.294 53.878 5.346 53.914 ;
      RECT 5.294 55.078 5.346 55.114 ;
      RECT 5.294 56.278 5.346 56.314 ;
      RECT 5.294 57.478 5.346 57.514 ;
      RECT 5.294 58.678 5.346 58.714 ;
      RECT 5.294 59.878 5.346 59.914 ;
      RECT 5.294 61.078 5.346 61.114 ;
      RECT 5.294 62.278 5.346 62.314 ;
      RECT 5.294 63.478 5.346 63.514 ;
      RECT 5.294 64.678 5.346 64.714 ;
      RECT 5.294 65.878 5.346 65.914 ;
      RECT 5.294 67.078 5.346 67.114 ;
      RECT 5.294 68.278 5.346 68.314 ;
      RECT 5.294 69.478 5.346 69.514 ;
      RECT 5.294 70.678 5.346 70.714 ;
      RECT 5.294 71.878 5.346 71.914 ;
      RECT 5.374 0.281 5.426 0.317 ;
      RECT 5.374 72.403 5.426 72.439 ;
      RECT 5.454 0.806 5.506 0.842 ;
      RECT 5.454 2.006 5.506 2.042 ;
      RECT 5.454 3.206 5.506 3.242 ;
      RECT 5.454 4.406 5.506 4.442 ;
      RECT 5.454 5.606 5.506 5.642 ;
      RECT 5.454 6.806 5.506 6.842 ;
      RECT 5.454 8.006 5.506 8.042 ;
      RECT 5.454 9.206 5.506 9.242 ;
      RECT 5.454 10.406 5.506 10.442 ;
      RECT 5.454 11.606 5.506 11.642 ;
      RECT 5.454 12.806 5.506 12.842 ;
      RECT 5.454 14.006 5.506 14.042 ;
      RECT 5.454 15.206 5.506 15.242 ;
      RECT 5.454 16.406 5.506 16.442 ;
      RECT 5.454 17.606 5.506 17.642 ;
      RECT 5.454 18.806 5.506 18.842 ;
      RECT 5.454 20.006 5.506 20.042 ;
      RECT 5.454 21.206 5.506 21.242 ;
      RECT 5.454 22.406 5.506 22.442 ;
      RECT 5.454 23.606 5.506 23.642 ;
      RECT 5.454 24.806 5.506 24.842 ;
      RECT 5.454 26.006 5.506 26.042 ;
      RECT 5.454 27.206 5.506 27.242 ;
      RECT 5.454 28.406 5.506 28.442 ;
      RECT 5.454 29.606 5.506 29.642 ;
      RECT 5.454 30.806 5.506 30.842 ;
      RECT 5.454 32.622 5.506 32.658 ;
      RECT 5.454 32.862 5.506 32.898 ;
      RECT 5.454 38.622 5.506 38.658 ;
      RECT 5.454 38.862 5.506 38.898 ;
      RECT 5.454 39.926 5.506 39.962 ;
      RECT 5.454 41.126 5.506 41.162 ;
      RECT 5.454 42.326 5.506 42.362 ;
      RECT 5.454 43.526 5.506 43.562 ;
      RECT 5.454 44.726 5.506 44.762 ;
      RECT 5.454 45.926 5.506 45.962 ;
      RECT 5.454 47.126 5.506 47.162 ;
      RECT 5.454 48.326 5.506 48.362 ;
      RECT 5.454 49.526 5.506 49.562 ;
      RECT 5.454 50.726 5.506 50.762 ;
      RECT 5.454 51.926 5.506 51.962 ;
      RECT 5.454 53.126 5.506 53.162 ;
      RECT 5.454 54.326 5.506 54.362 ;
      RECT 5.454 55.526 5.506 55.562 ;
      RECT 5.454 56.726 5.506 56.762 ;
      RECT 5.454 57.926 5.506 57.962 ;
      RECT 5.454 59.126 5.506 59.162 ;
      RECT 5.454 60.326 5.506 60.362 ;
      RECT 5.454 61.526 5.506 61.562 ;
      RECT 5.454 62.726 5.506 62.762 ;
      RECT 5.454 63.926 5.506 63.962 ;
      RECT 5.454 65.126 5.506 65.162 ;
      RECT 5.454 66.326 5.506 66.362 ;
      RECT 5.454 67.526 5.506 67.562 ;
      RECT 5.454 68.726 5.506 68.762 ;
      RECT 5.454 69.926 5.506 69.962 ;
      RECT 5.454 71.126 5.506 71.162 ;
      RECT 5.534 1.558 5.586 1.594 ;
      RECT 5.534 2.758 5.586 2.794 ;
      RECT 5.534 3.958 5.586 3.994 ;
      RECT 5.534 5.158 5.586 5.194 ;
      RECT 5.534 6.358 5.586 6.394 ;
      RECT 5.534 7.558 5.586 7.594 ;
      RECT 5.534 8.758 5.586 8.794 ;
      RECT 5.534 9.958 5.586 9.994 ;
      RECT 5.534 11.158 5.586 11.194 ;
      RECT 5.534 12.358 5.586 12.394 ;
      RECT 5.534 13.558 5.586 13.594 ;
      RECT 5.534 14.758 5.586 14.794 ;
      RECT 5.534 15.958 5.586 15.994 ;
      RECT 5.534 17.158 5.586 17.194 ;
      RECT 5.534 18.358 5.586 18.394 ;
      RECT 5.534 19.558 5.586 19.594 ;
      RECT 5.534 20.758 5.586 20.794 ;
      RECT 5.534 21.958 5.586 21.994 ;
      RECT 5.534 23.158 5.586 23.194 ;
      RECT 5.534 24.358 5.586 24.394 ;
      RECT 5.534 25.558 5.586 25.594 ;
      RECT 5.534 26.758 5.586 26.794 ;
      RECT 5.534 27.958 5.586 27.994 ;
      RECT 5.534 29.158 5.586 29.194 ;
      RECT 5.534 30.358 5.586 30.394 ;
      RECT 5.534 31.558 5.586 31.594 ;
      RECT 5.534 33.342 5.586 33.378 ;
      RECT 5.534 33.582 5.586 33.618 ;
      RECT 5.534 37.902 5.586 37.938 ;
      RECT 5.534 38.142 5.586 38.178 ;
      RECT 5.534 40.678 5.586 40.714 ;
      RECT 5.534 41.878 5.586 41.914 ;
      RECT 5.534 43.078 5.586 43.114 ;
      RECT 5.534 44.278 5.586 44.314 ;
      RECT 5.534 45.478 5.586 45.514 ;
      RECT 5.534 46.678 5.586 46.714 ;
      RECT 5.534 47.878 5.586 47.914 ;
      RECT 5.534 49.078 5.586 49.114 ;
      RECT 5.534 50.278 5.586 50.314 ;
      RECT 5.534 51.478 5.586 51.514 ;
      RECT 5.534 52.678 5.586 52.714 ;
      RECT 5.534 53.878 5.586 53.914 ;
      RECT 5.534 55.078 5.586 55.114 ;
      RECT 5.534 56.278 5.586 56.314 ;
      RECT 5.534 57.478 5.586 57.514 ;
      RECT 5.534 58.678 5.586 58.714 ;
      RECT 5.534 59.878 5.586 59.914 ;
      RECT 5.534 61.078 5.586 61.114 ;
      RECT 5.534 62.278 5.586 62.314 ;
      RECT 5.534 63.478 5.586 63.514 ;
      RECT 5.534 64.678 5.586 64.714 ;
      RECT 5.534 65.878 5.586 65.914 ;
      RECT 5.534 67.078 5.586 67.114 ;
      RECT 5.534 68.278 5.586 68.314 ;
      RECT 5.534 69.478 5.586 69.514 ;
      RECT 5.534 70.678 5.586 70.714 ;
      RECT 5.534 71.878 5.586 71.914 ;
      RECT 5.614 0.806 5.666 0.842 ;
      RECT 5.614 2.006 5.666 2.042 ;
      RECT 5.614 3.206 5.666 3.242 ;
      RECT 5.614 4.406 5.666 4.442 ;
      RECT 5.614 5.606 5.666 5.642 ;
      RECT 5.614 6.806 5.666 6.842 ;
      RECT 5.614 8.006 5.666 8.042 ;
      RECT 5.614 9.206 5.666 9.242 ;
      RECT 5.614 10.406 5.666 10.442 ;
      RECT 5.614 11.606 5.666 11.642 ;
      RECT 5.614 12.806 5.666 12.842 ;
      RECT 5.614 14.006 5.666 14.042 ;
      RECT 5.614 15.206 5.666 15.242 ;
      RECT 5.614 16.406 5.666 16.442 ;
      RECT 5.614 17.606 5.666 17.642 ;
      RECT 5.614 18.806 5.666 18.842 ;
      RECT 5.614 20.006 5.666 20.042 ;
      RECT 5.614 21.206 5.666 21.242 ;
      RECT 5.614 22.406 5.666 22.442 ;
      RECT 5.614 23.606 5.666 23.642 ;
      RECT 5.614 24.806 5.666 24.842 ;
      RECT 5.614 26.006 5.666 26.042 ;
      RECT 5.614 27.206 5.666 27.242 ;
      RECT 5.614 28.406 5.666 28.442 ;
      RECT 5.614 29.606 5.666 29.642 ;
      RECT 5.614 30.806 5.666 30.842 ;
      RECT 5.614 32.622 5.666 32.658 ;
      RECT 5.614 32.862 5.666 32.898 ;
      RECT 5.614 38.622 5.666 38.658 ;
      RECT 5.614 38.862 5.666 38.898 ;
      RECT 5.614 39.926 5.666 39.962 ;
      RECT 5.614 41.126 5.666 41.162 ;
      RECT 5.614 42.326 5.666 42.362 ;
      RECT 5.614 43.526 5.666 43.562 ;
      RECT 5.614 44.726 5.666 44.762 ;
      RECT 5.614 45.926 5.666 45.962 ;
      RECT 5.614 47.126 5.666 47.162 ;
      RECT 5.614 48.326 5.666 48.362 ;
      RECT 5.614 49.526 5.666 49.562 ;
      RECT 5.614 50.726 5.666 50.762 ;
      RECT 5.614 51.926 5.666 51.962 ;
      RECT 5.614 53.126 5.666 53.162 ;
      RECT 5.614 54.326 5.666 54.362 ;
      RECT 5.614 55.526 5.666 55.562 ;
      RECT 5.614 56.726 5.666 56.762 ;
      RECT 5.614 57.926 5.666 57.962 ;
      RECT 5.614 59.126 5.666 59.162 ;
      RECT 5.614 60.326 5.666 60.362 ;
      RECT 5.614 61.526 5.666 61.562 ;
      RECT 5.614 62.726 5.666 62.762 ;
      RECT 5.614 63.926 5.666 63.962 ;
      RECT 5.614 65.126 5.666 65.162 ;
      RECT 5.614 66.326 5.666 66.362 ;
      RECT 5.614 67.526 5.666 67.562 ;
      RECT 5.614 68.726 5.666 68.762 ;
      RECT 5.614 69.926 5.666 69.962 ;
      RECT 5.614 71.126 5.666 71.162 ;
      RECT 5.694 1.558 5.746 1.594 ;
      RECT 5.694 2.758 5.746 2.794 ;
      RECT 5.694 3.958 5.746 3.994 ;
      RECT 5.694 5.158 5.746 5.194 ;
      RECT 5.694 6.358 5.746 6.394 ;
      RECT 5.694 7.558 5.746 7.594 ;
      RECT 5.694 8.758 5.746 8.794 ;
      RECT 5.694 9.958 5.746 9.994 ;
      RECT 5.694 11.158 5.746 11.194 ;
      RECT 5.694 12.358 5.746 12.394 ;
      RECT 5.694 13.558 5.746 13.594 ;
      RECT 5.694 14.758 5.746 14.794 ;
      RECT 5.694 15.958 5.746 15.994 ;
      RECT 5.694 17.158 5.746 17.194 ;
      RECT 5.694 18.358 5.746 18.394 ;
      RECT 5.694 19.558 5.746 19.594 ;
      RECT 5.694 20.758 5.746 20.794 ;
      RECT 5.694 21.958 5.746 21.994 ;
      RECT 5.694 23.158 5.746 23.194 ;
      RECT 5.694 24.358 5.746 24.394 ;
      RECT 5.694 25.558 5.746 25.594 ;
      RECT 5.694 26.758 5.746 26.794 ;
      RECT 5.694 27.958 5.746 27.994 ;
      RECT 5.694 29.158 5.746 29.194 ;
      RECT 5.694 30.358 5.746 30.394 ;
      RECT 5.694 31.558 5.746 31.594 ;
      RECT 5.694 33.342 5.746 33.378 ;
      RECT 5.694 33.582 5.746 33.618 ;
      RECT 5.694 37.902 5.746 37.938 ;
      RECT 5.694 38.142 5.746 38.178 ;
      RECT 5.694 40.678 5.746 40.714 ;
      RECT 5.694 41.878 5.746 41.914 ;
      RECT 5.694 43.078 5.746 43.114 ;
      RECT 5.694 44.278 5.746 44.314 ;
      RECT 5.694 45.478 5.746 45.514 ;
      RECT 5.694 46.678 5.746 46.714 ;
      RECT 5.694 47.878 5.746 47.914 ;
      RECT 5.694 49.078 5.746 49.114 ;
      RECT 5.694 50.278 5.746 50.314 ;
      RECT 5.694 51.478 5.746 51.514 ;
      RECT 5.694 52.678 5.746 52.714 ;
      RECT 5.694 53.878 5.746 53.914 ;
      RECT 5.694 55.078 5.746 55.114 ;
      RECT 5.694 56.278 5.746 56.314 ;
      RECT 5.694 57.478 5.746 57.514 ;
      RECT 5.694 58.678 5.746 58.714 ;
      RECT 5.694 59.878 5.746 59.914 ;
      RECT 5.694 61.078 5.746 61.114 ;
      RECT 5.694 62.278 5.746 62.314 ;
      RECT 5.694 63.478 5.746 63.514 ;
      RECT 5.694 64.678 5.746 64.714 ;
      RECT 5.694 65.878 5.746 65.914 ;
      RECT 5.694 67.078 5.746 67.114 ;
      RECT 5.694 68.278 5.746 68.314 ;
      RECT 5.694 69.478 5.746 69.514 ;
      RECT 5.694 70.678 5.746 70.714 ;
      RECT 5.694 71.878 5.746 71.914 ;
      RECT 5.774 0.281 5.826 0.317 ;
      RECT 5.774 72.403 5.826 72.439 ;
      RECT 5.854 0.806 5.906 0.842 ;
      RECT 5.854 2.006 5.906 2.042 ;
      RECT 5.854 3.206 5.906 3.242 ;
      RECT 5.854 4.406 5.906 4.442 ;
      RECT 5.854 5.606 5.906 5.642 ;
      RECT 5.854 6.806 5.906 6.842 ;
      RECT 5.854 8.006 5.906 8.042 ;
      RECT 5.854 9.206 5.906 9.242 ;
      RECT 5.854 10.406 5.906 10.442 ;
      RECT 5.854 11.606 5.906 11.642 ;
      RECT 5.854 12.806 5.906 12.842 ;
      RECT 5.854 14.006 5.906 14.042 ;
      RECT 5.854 15.206 5.906 15.242 ;
      RECT 5.854 16.406 5.906 16.442 ;
      RECT 5.854 17.606 5.906 17.642 ;
      RECT 5.854 18.806 5.906 18.842 ;
      RECT 5.854 20.006 5.906 20.042 ;
      RECT 5.854 21.206 5.906 21.242 ;
      RECT 5.854 22.406 5.906 22.442 ;
      RECT 5.854 23.606 5.906 23.642 ;
      RECT 5.854 24.806 5.906 24.842 ;
      RECT 5.854 26.006 5.906 26.042 ;
      RECT 5.854 27.206 5.906 27.242 ;
      RECT 5.854 28.406 5.906 28.442 ;
      RECT 5.854 29.606 5.906 29.642 ;
      RECT 5.854 30.806 5.906 30.842 ;
      RECT 5.854 32.622 5.906 32.658 ;
      RECT 5.854 32.862 5.906 32.898 ;
      RECT 5.854 34.302 5.906 34.338 ;
      RECT 5.854 34.782 5.906 34.818 ;
      RECT 5.854 36.702 5.906 36.738 ;
      RECT 5.854 37.182 5.906 37.218 ;
      RECT 5.854 38.622 5.906 38.658 ;
      RECT 5.854 38.862 5.906 38.898 ;
      RECT 5.854 39.926 5.906 39.962 ;
      RECT 5.854 41.126 5.906 41.162 ;
      RECT 5.854 42.326 5.906 42.362 ;
      RECT 5.854 43.526 5.906 43.562 ;
      RECT 5.854 44.726 5.906 44.762 ;
      RECT 5.854 45.926 5.906 45.962 ;
      RECT 5.854 47.126 5.906 47.162 ;
      RECT 5.854 48.326 5.906 48.362 ;
      RECT 5.854 49.526 5.906 49.562 ;
      RECT 5.854 50.726 5.906 50.762 ;
      RECT 5.854 51.926 5.906 51.962 ;
      RECT 5.854 53.126 5.906 53.162 ;
      RECT 5.854 54.326 5.906 54.362 ;
      RECT 5.854 55.526 5.906 55.562 ;
      RECT 5.854 56.726 5.906 56.762 ;
      RECT 5.854 57.926 5.906 57.962 ;
      RECT 5.854 59.126 5.906 59.162 ;
      RECT 5.854 60.326 5.906 60.362 ;
      RECT 5.854 61.526 5.906 61.562 ;
      RECT 5.854 62.726 5.906 62.762 ;
      RECT 5.854 63.926 5.906 63.962 ;
      RECT 5.854 65.126 5.906 65.162 ;
      RECT 5.854 66.326 5.906 66.362 ;
      RECT 5.854 67.526 5.906 67.562 ;
      RECT 5.854 68.726 5.906 68.762 ;
      RECT 5.854 69.926 5.906 69.962 ;
      RECT 5.854 71.126 5.906 71.162 ;
      RECT 5.934 1.558 5.986 1.594 ;
      RECT 5.934 2.758 5.986 2.794 ;
      RECT 5.934 3.958 5.986 3.994 ;
      RECT 5.934 5.158 5.986 5.194 ;
      RECT 5.934 6.358 5.986 6.394 ;
      RECT 5.934 7.558 5.986 7.594 ;
      RECT 5.934 8.758 5.986 8.794 ;
      RECT 5.934 9.958 5.986 9.994 ;
      RECT 5.934 11.158 5.986 11.194 ;
      RECT 5.934 12.358 5.986 12.394 ;
      RECT 5.934 13.558 5.986 13.594 ;
      RECT 5.934 14.758 5.986 14.794 ;
      RECT 5.934 15.958 5.986 15.994 ;
      RECT 5.934 17.158 5.986 17.194 ;
      RECT 5.934 18.358 5.986 18.394 ;
      RECT 5.934 19.558 5.986 19.594 ;
      RECT 5.934 20.758 5.986 20.794 ;
      RECT 5.934 21.958 5.986 21.994 ;
      RECT 5.934 23.158 5.986 23.194 ;
      RECT 5.934 24.358 5.986 24.394 ;
      RECT 5.934 25.558 5.986 25.594 ;
      RECT 5.934 26.758 5.986 26.794 ;
      RECT 5.934 27.958 5.986 27.994 ;
      RECT 5.934 29.158 5.986 29.194 ;
      RECT 5.934 30.358 5.986 30.394 ;
      RECT 5.934 31.558 5.986 31.594 ;
      RECT 5.934 33.342 5.986 33.378 ;
      RECT 5.934 33.582 5.986 33.618 ;
      RECT 5.934 37.902 5.986 37.938 ;
      RECT 5.934 38.142 5.986 38.178 ;
      RECT 5.934 40.678 5.986 40.714 ;
      RECT 5.934 41.878 5.986 41.914 ;
      RECT 5.934 43.078 5.986 43.114 ;
      RECT 5.934 44.278 5.986 44.314 ;
      RECT 5.934 45.478 5.986 45.514 ;
      RECT 5.934 46.678 5.986 46.714 ;
      RECT 5.934 47.878 5.986 47.914 ;
      RECT 5.934 49.078 5.986 49.114 ;
      RECT 5.934 50.278 5.986 50.314 ;
      RECT 5.934 51.478 5.986 51.514 ;
      RECT 5.934 52.678 5.986 52.714 ;
      RECT 5.934 53.878 5.986 53.914 ;
      RECT 5.934 55.078 5.986 55.114 ;
      RECT 5.934 56.278 5.986 56.314 ;
      RECT 5.934 57.478 5.986 57.514 ;
      RECT 5.934 58.678 5.986 58.714 ;
      RECT 5.934 59.878 5.986 59.914 ;
      RECT 5.934 61.078 5.986 61.114 ;
      RECT 5.934 62.278 5.986 62.314 ;
      RECT 5.934 63.478 5.986 63.514 ;
      RECT 5.934 64.678 5.986 64.714 ;
      RECT 5.934 65.878 5.986 65.914 ;
      RECT 5.934 67.078 5.986 67.114 ;
      RECT 5.934 68.278 5.986 68.314 ;
      RECT 5.934 69.478 5.986 69.514 ;
      RECT 5.934 70.678 5.986 70.714 ;
      RECT 5.934 71.878 5.986 71.914 ;
      RECT 6.014 0.806 6.066 0.842 ;
      RECT 6.014 2.006 6.066 2.042 ;
      RECT 6.014 3.206 6.066 3.242 ;
      RECT 6.014 4.406 6.066 4.442 ;
      RECT 6.014 5.606 6.066 5.642 ;
      RECT 6.014 6.806 6.066 6.842 ;
      RECT 6.014 8.006 6.066 8.042 ;
      RECT 6.014 9.206 6.066 9.242 ;
      RECT 6.014 10.406 6.066 10.442 ;
      RECT 6.014 11.606 6.066 11.642 ;
      RECT 6.014 12.806 6.066 12.842 ;
      RECT 6.014 14.006 6.066 14.042 ;
      RECT 6.014 15.206 6.066 15.242 ;
      RECT 6.014 16.406 6.066 16.442 ;
      RECT 6.014 17.606 6.066 17.642 ;
      RECT 6.014 18.806 6.066 18.842 ;
      RECT 6.014 20.006 6.066 20.042 ;
      RECT 6.014 21.206 6.066 21.242 ;
      RECT 6.014 22.406 6.066 22.442 ;
      RECT 6.014 23.606 6.066 23.642 ;
      RECT 6.014 24.806 6.066 24.842 ;
      RECT 6.014 26.006 6.066 26.042 ;
      RECT 6.014 27.206 6.066 27.242 ;
      RECT 6.014 28.406 6.066 28.442 ;
      RECT 6.014 29.606 6.066 29.642 ;
      RECT 6.014 30.806 6.066 30.842 ;
      RECT 6.014 32.622 6.066 32.658 ;
      RECT 6.014 32.862 6.066 32.898 ;
      RECT 6.014 38.622 6.066 38.658 ;
      RECT 6.014 38.862 6.066 38.898 ;
      RECT 6.014 39.926 6.066 39.962 ;
      RECT 6.014 41.126 6.066 41.162 ;
      RECT 6.014 42.326 6.066 42.362 ;
      RECT 6.014 43.526 6.066 43.562 ;
      RECT 6.014 44.726 6.066 44.762 ;
      RECT 6.014 45.926 6.066 45.962 ;
      RECT 6.014 47.126 6.066 47.162 ;
      RECT 6.014 48.326 6.066 48.362 ;
      RECT 6.014 49.526 6.066 49.562 ;
      RECT 6.014 50.726 6.066 50.762 ;
      RECT 6.014 51.926 6.066 51.962 ;
      RECT 6.014 53.126 6.066 53.162 ;
      RECT 6.014 54.326 6.066 54.362 ;
      RECT 6.014 55.526 6.066 55.562 ;
      RECT 6.014 56.726 6.066 56.762 ;
      RECT 6.014 57.926 6.066 57.962 ;
      RECT 6.014 59.126 6.066 59.162 ;
      RECT 6.014 60.326 6.066 60.362 ;
      RECT 6.014 61.526 6.066 61.562 ;
      RECT 6.014 62.726 6.066 62.762 ;
      RECT 6.014 63.926 6.066 63.962 ;
      RECT 6.014 65.126 6.066 65.162 ;
      RECT 6.014 66.326 6.066 66.362 ;
      RECT 6.014 67.526 6.066 67.562 ;
      RECT 6.014 68.726 6.066 68.762 ;
      RECT 6.014 69.926 6.066 69.962 ;
      RECT 6.014 71.126 6.066 71.162 ;
      RECT 6.094 1.558 6.146 1.594 ;
      RECT 6.094 2.758 6.146 2.794 ;
      RECT 6.094 3.958 6.146 3.994 ;
      RECT 6.094 5.158 6.146 5.194 ;
      RECT 6.094 6.358 6.146 6.394 ;
      RECT 6.094 7.558 6.146 7.594 ;
      RECT 6.094 8.758 6.146 8.794 ;
      RECT 6.094 9.958 6.146 9.994 ;
      RECT 6.094 11.158 6.146 11.194 ;
      RECT 6.094 12.358 6.146 12.394 ;
      RECT 6.094 13.558 6.146 13.594 ;
      RECT 6.094 14.758 6.146 14.794 ;
      RECT 6.094 15.958 6.146 15.994 ;
      RECT 6.094 17.158 6.146 17.194 ;
      RECT 6.094 18.358 6.146 18.394 ;
      RECT 6.094 19.558 6.146 19.594 ;
      RECT 6.094 20.758 6.146 20.794 ;
      RECT 6.094 21.958 6.146 21.994 ;
      RECT 6.094 23.158 6.146 23.194 ;
      RECT 6.094 24.358 6.146 24.394 ;
      RECT 6.094 25.558 6.146 25.594 ;
      RECT 6.094 26.758 6.146 26.794 ;
      RECT 6.094 27.958 6.146 27.994 ;
      RECT 6.094 29.158 6.146 29.194 ;
      RECT 6.094 30.358 6.146 30.394 ;
      RECT 6.094 31.558 6.146 31.594 ;
      RECT 6.094 33.342 6.146 33.378 ;
      RECT 6.094 33.582 6.146 33.618 ;
      RECT 6.094 37.902 6.146 37.938 ;
      RECT 6.094 38.142 6.146 38.178 ;
      RECT 6.094 40.678 6.146 40.714 ;
      RECT 6.094 41.878 6.146 41.914 ;
      RECT 6.094 43.078 6.146 43.114 ;
      RECT 6.094 44.278 6.146 44.314 ;
      RECT 6.094 45.478 6.146 45.514 ;
      RECT 6.094 46.678 6.146 46.714 ;
      RECT 6.094 47.878 6.146 47.914 ;
      RECT 6.094 49.078 6.146 49.114 ;
      RECT 6.094 50.278 6.146 50.314 ;
      RECT 6.094 51.478 6.146 51.514 ;
      RECT 6.094 52.678 6.146 52.714 ;
      RECT 6.094 53.878 6.146 53.914 ;
      RECT 6.094 55.078 6.146 55.114 ;
      RECT 6.094 56.278 6.146 56.314 ;
      RECT 6.094 57.478 6.146 57.514 ;
      RECT 6.094 58.678 6.146 58.714 ;
      RECT 6.094 59.878 6.146 59.914 ;
      RECT 6.094 61.078 6.146 61.114 ;
      RECT 6.094 62.278 6.146 62.314 ;
      RECT 6.094 63.478 6.146 63.514 ;
      RECT 6.094 64.678 6.146 64.714 ;
      RECT 6.094 65.878 6.146 65.914 ;
      RECT 6.094 67.078 6.146 67.114 ;
      RECT 6.094 68.278 6.146 68.314 ;
      RECT 6.094 69.478 6.146 69.514 ;
      RECT 6.094 70.678 6.146 70.714 ;
      RECT 6.094 71.878 6.146 71.914 ;
      RECT 6.174 0.281 6.226 0.317 ;
      RECT 6.174 72.403 6.226 72.439 ;
      RECT 6.254 0.806 6.306 0.842 ;
      RECT 6.254 2.006 6.306 2.042 ;
      RECT 6.254 3.206 6.306 3.242 ;
      RECT 6.254 4.406 6.306 4.442 ;
      RECT 6.254 5.606 6.306 5.642 ;
      RECT 6.254 6.806 6.306 6.842 ;
      RECT 6.254 8.006 6.306 8.042 ;
      RECT 6.254 9.206 6.306 9.242 ;
      RECT 6.254 10.406 6.306 10.442 ;
      RECT 6.254 11.606 6.306 11.642 ;
      RECT 6.254 12.806 6.306 12.842 ;
      RECT 6.254 14.006 6.306 14.042 ;
      RECT 6.254 15.206 6.306 15.242 ;
      RECT 6.254 16.406 6.306 16.442 ;
      RECT 6.254 17.606 6.306 17.642 ;
      RECT 6.254 18.806 6.306 18.842 ;
      RECT 6.254 20.006 6.306 20.042 ;
      RECT 6.254 21.206 6.306 21.242 ;
      RECT 6.254 22.406 6.306 22.442 ;
      RECT 6.254 23.606 6.306 23.642 ;
      RECT 6.254 24.806 6.306 24.842 ;
      RECT 6.254 26.006 6.306 26.042 ;
      RECT 6.254 27.206 6.306 27.242 ;
      RECT 6.254 28.406 6.306 28.442 ;
      RECT 6.254 29.606 6.306 29.642 ;
      RECT 6.254 30.806 6.306 30.842 ;
      RECT 6.254 32.622 6.306 32.658 ;
      RECT 6.254 32.862 6.306 32.898 ;
      RECT 6.254 38.622 6.306 38.658 ;
      RECT 6.254 38.862 6.306 38.898 ;
      RECT 6.254 39.926 6.306 39.962 ;
      RECT 6.254 41.126 6.306 41.162 ;
      RECT 6.254 42.326 6.306 42.362 ;
      RECT 6.254 43.526 6.306 43.562 ;
      RECT 6.254 44.726 6.306 44.762 ;
      RECT 6.254 45.926 6.306 45.962 ;
      RECT 6.254 47.126 6.306 47.162 ;
      RECT 6.254 48.326 6.306 48.362 ;
      RECT 6.254 49.526 6.306 49.562 ;
      RECT 6.254 50.726 6.306 50.762 ;
      RECT 6.254 51.926 6.306 51.962 ;
      RECT 6.254 53.126 6.306 53.162 ;
      RECT 6.254 54.326 6.306 54.362 ;
      RECT 6.254 55.526 6.306 55.562 ;
      RECT 6.254 56.726 6.306 56.762 ;
      RECT 6.254 57.926 6.306 57.962 ;
      RECT 6.254 59.126 6.306 59.162 ;
      RECT 6.254 60.326 6.306 60.362 ;
      RECT 6.254 61.526 6.306 61.562 ;
      RECT 6.254 62.726 6.306 62.762 ;
      RECT 6.254 63.926 6.306 63.962 ;
      RECT 6.254 65.126 6.306 65.162 ;
      RECT 6.254 66.326 6.306 66.362 ;
      RECT 6.254 67.526 6.306 67.562 ;
      RECT 6.254 68.726 6.306 68.762 ;
      RECT 6.254 69.926 6.306 69.962 ;
      RECT 6.254 71.126 6.306 71.162 ;
      RECT 6.334 1.558 6.386 1.594 ;
      RECT 6.334 2.758 6.386 2.794 ;
      RECT 6.334 3.958 6.386 3.994 ;
      RECT 6.334 5.158 6.386 5.194 ;
      RECT 6.334 6.358 6.386 6.394 ;
      RECT 6.334 7.558 6.386 7.594 ;
      RECT 6.334 8.758 6.386 8.794 ;
      RECT 6.334 9.958 6.386 9.994 ;
      RECT 6.334 11.158 6.386 11.194 ;
      RECT 6.334 12.358 6.386 12.394 ;
      RECT 6.334 13.558 6.386 13.594 ;
      RECT 6.334 14.758 6.386 14.794 ;
      RECT 6.334 15.958 6.386 15.994 ;
      RECT 6.334 17.158 6.386 17.194 ;
      RECT 6.334 18.358 6.386 18.394 ;
      RECT 6.334 19.558 6.386 19.594 ;
      RECT 6.334 20.758 6.386 20.794 ;
      RECT 6.334 21.958 6.386 21.994 ;
      RECT 6.334 23.158 6.386 23.194 ;
      RECT 6.334 24.358 6.386 24.394 ;
      RECT 6.334 25.558 6.386 25.594 ;
      RECT 6.334 26.758 6.386 26.794 ;
      RECT 6.334 27.958 6.386 27.994 ;
      RECT 6.334 29.158 6.386 29.194 ;
      RECT 6.334 30.358 6.386 30.394 ;
      RECT 6.334 31.558 6.386 31.594 ;
      RECT 6.334 33.342 6.386 33.378 ;
      RECT 6.334 33.582 6.386 33.618 ;
      RECT 6.334 37.902 6.386 37.938 ;
      RECT 6.334 38.142 6.386 38.178 ;
      RECT 6.334 40.678 6.386 40.714 ;
      RECT 6.334 41.878 6.386 41.914 ;
      RECT 6.334 43.078 6.386 43.114 ;
      RECT 6.334 44.278 6.386 44.314 ;
      RECT 6.334 45.478 6.386 45.514 ;
      RECT 6.334 46.678 6.386 46.714 ;
      RECT 6.334 47.878 6.386 47.914 ;
      RECT 6.334 49.078 6.386 49.114 ;
      RECT 6.334 50.278 6.386 50.314 ;
      RECT 6.334 51.478 6.386 51.514 ;
      RECT 6.334 52.678 6.386 52.714 ;
      RECT 6.334 53.878 6.386 53.914 ;
      RECT 6.334 55.078 6.386 55.114 ;
      RECT 6.334 56.278 6.386 56.314 ;
      RECT 6.334 57.478 6.386 57.514 ;
      RECT 6.334 58.678 6.386 58.714 ;
      RECT 6.334 59.878 6.386 59.914 ;
      RECT 6.334 61.078 6.386 61.114 ;
      RECT 6.334 62.278 6.386 62.314 ;
      RECT 6.334 63.478 6.386 63.514 ;
      RECT 6.334 64.678 6.386 64.714 ;
      RECT 6.334 65.878 6.386 65.914 ;
      RECT 6.334 67.078 6.386 67.114 ;
      RECT 6.334 68.278 6.386 68.314 ;
      RECT 6.334 69.478 6.386 69.514 ;
      RECT 6.334 70.678 6.386 70.714 ;
      RECT 6.334 71.878 6.386 71.914 ;
      RECT 6.414 0.806 6.466 0.842 ;
      RECT 6.414 2.006 6.466 2.042 ;
      RECT 6.414 3.206 6.466 3.242 ;
      RECT 6.414 4.406 6.466 4.442 ;
      RECT 6.414 5.606 6.466 5.642 ;
      RECT 6.414 6.806 6.466 6.842 ;
      RECT 6.414 8.006 6.466 8.042 ;
      RECT 6.414 9.206 6.466 9.242 ;
      RECT 6.414 10.406 6.466 10.442 ;
      RECT 6.414 11.606 6.466 11.642 ;
      RECT 6.414 12.806 6.466 12.842 ;
      RECT 6.414 14.006 6.466 14.042 ;
      RECT 6.414 15.206 6.466 15.242 ;
      RECT 6.414 16.406 6.466 16.442 ;
      RECT 6.414 17.606 6.466 17.642 ;
      RECT 6.414 18.806 6.466 18.842 ;
      RECT 6.414 20.006 6.466 20.042 ;
      RECT 6.414 21.206 6.466 21.242 ;
      RECT 6.414 22.406 6.466 22.442 ;
      RECT 6.414 23.606 6.466 23.642 ;
      RECT 6.414 24.806 6.466 24.842 ;
      RECT 6.414 26.006 6.466 26.042 ;
      RECT 6.414 27.206 6.466 27.242 ;
      RECT 6.414 28.406 6.466 28.442 ;
      RECT 6.414 29.606 6.466 29.642 ;
      RECT 6.414 30.806 6.466 30.842 ;
      RECT 6.414 32.622 6.466 32.658 ;
      RECT 6.414 32.862 6.466 32.898 ;
      RECT 6.414 38.622 6.466 38.658 ;
      RECT 6.414 38.862 6.466 38.898 ;
      RECT 6.414 39.926 6.466 39.962 ;
      RECT 6.414 41.126 6.466 41.162 ;
      RECT 6.414 42.326 6.466 42.362 ;
      RECT 6.414 43.526 6.466 43.562 ;
      RECT 6.414 44.726 6.466 44.762 ;
      RECT 6.414 45.926 6.466 45.962 ;
      RECT 6.414 47.126 6.466 47.162 ;
      RECT 6.414 48.326 6.466 48.362 ;
      RECT 6.414 49.526 6.466 49.562 ;
      RECT 6.414 50.726 6.466 50.762 ;
      RECT 6.414 51.926 6.466 51.962 ;
      RECT 6.414 53.126 6.466 53.162 ;
      RECT 6.414 54.326 6.466 54.362 ;
      RECT 6.414 55.526 6.466 55.562 ;
      RECT 6.414 56.726 6.466 56.762 ;
      RECT 6.414 57.926 6.466 57.962 ;
      RECT 6.414 59.126 6.466 59.162 ;
      RECT 6.414 60.326 6.466 60.362 ;
      RECT 6.414 61.526 6.466 61.562 ;
      RECT 6.414 62.726 6.466 62.762 ;
      RECT 6.414 63.926 6.466 63.962 ;
      RECT 6.414 65.126 6.466 65.162 ;
      RECT 6.414 66.326 6.466 66.362 ;
      RECT 6.414 67.526 6.466 67.562 ;
      RECT 6.414 68.726 6.466 68.762 ;
      RECT 6.414 69.926 6.466 69.962 ;
      RECT 6.414 71.126 6.466 71.162 ;
      RECT 6.494 1.558 6.546 1.594 ;
      RECT 6.494 2.758 6.546 2.794 ;
      RECT 6.494 3.958 6.546 3.994 ;
      RECT 6.494 5.158 6.546 5.194 ;
      RECT 6.494 6.358 6.546 6.394 ;
      RECT 6.494 7.558 6.546 7.594 ;
      RECT 6.494 8.758 6.546 8.794 ;
      RECT 6.494 9.958 6.546 9.994 ;
      RECT 6.494 11.158 6.546 11.194 ;
      RECT 6.494 12.358 6.546 12.394 ;
      RECT 6.494 13.558 6.546 13.594 ;
      RECT 6.494 14.758 6.546 14.794 ;
      RECT 6.494 15.958 6.546 15.994 ;
      RECT 6.494 17.158 6.546 17.194 ;
      RECT 6.494 18.358 6.546 18.394 ;
      RECT 6.494 19.558 6.546 19.594 ;
      RECT 6.494 20.758 6.546 20.794 ;
      RECT 6.494 21.958 6.546 21.994 ;
      RECT 6.494 23.158 6.546 23.194 ;
      RECT 6.494 24.358 6.546 24.394 ;
      RECT 6.494 25.558 6.546 25.594 ;
      RECT 6.494 26.758 6.546 26.794 ;
      RECT 6.494 27.958 6.546 27.994 ;
      RECT 6.494 29.158 6.546 29.194 ;
      RECT 6.494 30.358 6.546 30.394 ;
      RECT 6.494 31.558 6.546 31.594 ;
      RECT 6.494 33.342 6.546 33.378 ;
      RECT 6.494 33.582 6.546 33.618 ;
      RECT 6.494 37.902 6.546 37.938 ;
      RECT 6.494 38.142 6.546 38.178 ;
      RECT 6.494 40.678 6.546 40.714 ;
      RECT 6.494 41.878 6.546 41.914 ;
      RECT 6.494 43.078 6.546 43.114 ;
      RECT 6.494 44.278 6.546 44.314 ;
      RECT 6.494 45.478 6.546 45.514 ;
      RECT 6.494 46.678 6.546 46.714 ;
      RECT 6.494 47.878 6.546 47.914 ;
      RECT 6.494 49.078 6.546 49.114 ;
      RECT 6.494 50.278 6.546 50.314 ;
      RECT 6.494 51.478 6.546 51.514 ;
      RECT 6.494 52.678 6.546 52.714 ;
      RECT 6.494 53.878 6.546 53.914 ;
      RECT 6.494 55.078 6.546 55.114 ;
      RECT 6.494 56.278 6.546 56.314 ;
      RECT 6.494 57.478 6.546 57.514 ;
      RECT 6.494 58.678 6.546 58.714 ;
      RECT 6.494 59.878 6.546 59.914 ;
      RECT 6.494 61.078 6.546 61.114 ;
      RECT 6.494 62.278 6.546 62.314 ;
      RECT 6.494 63.478 6.546 63.514 ;
      RECT 6.494 64.678 6.546 64.714 ;
      RECT 6.494 65.878 6.546 65.914 ;
      RECT 6.494 67.078 6.546 67.114 ;
      RECT 6.494 68.278 6.546 68.314 ;
      RECT 6.494 69.478 6.546 69.514 ;
      RECT 6.494 70.678 6.546 70.714 ;
      RECT 6.494 71.878 6.546 71.914 ;
      RECT 6.574 0.281 6.626 0.317 ;
      RECT 6.574 72.403 6.626 72.439 ;
      RECT 6.654 0.806 6.706 0.842 ;
      RECT 6.654 2.006 6.706 2.042 ;
      RECT 6.654 3.206 6.706 3.242 ;
      RECT 6.654 4.406 6.706 4.442 ;
      RECT 6.654 5.606 6.706 5.642 ;
      RECT 6.654 6.806 6.706 6.842 ;
      RECT 6.654 8.006 6.706 8.042 ;
      RECT 6.654 9.206 6.706 9.242 ;
      RECT 6.654 10.406 6.706 10.442 ;
      RECT 6.654 11.606 6.706 11.642 ;
      RECT 6.654 12.806 6.706 12.842 ;
      RECT 6.654 14.006 6.706 14.042 ;
      RECT 6.654 15.206 6.706 15.242 ;
      RECT 6.654 16.406 6.706 16.442 ;
      RECT 6.654 17.606 6.706 17.642 ;
      RECT 6.654 18.806 6.706 18.842 ;
      RECT 6.654 20.006 6.706 20.042 ;
      RECT 6.654 21.206 6.706 21.242 ;
      RECT 6.654 22.406 6.706 22.442 ;
      RECT 6.654 23.606 6.706 23.642 ;
      RECT 6.654 24.806 6.706 24.842 ;
      RECT 6.654 26.006 6.706 26.042 ;
      RECT 6.654 27.206 6.706 27.242 ;
      RECT 6.654 28.406 6.706 28.442 ;
      RECT 6.654 29.606 6.706 29.642 ;
      RECT 6.654 30.806 6.706 30.842 ;
      RECT 6.654 32.622 6.706 32.658 ;
      RECT 6.654 32.862 6.706 32.898 ;
      RECT 6.654 34.302 6.706 34.338 ;
      RECT 6.654 34.782 6.706 34.818 ;
      RECT 6.654 36.702 6.706 36.738 ;
      RECT 6.654 37.182 6.706 37.218 ;
      RECT 6.654 38.622 6.706 38.658 ;
      RECT 6.654 38.862 6.706 38.898 ;
      RECT 6.654 39.926 6.706 39.962 ;
      RECT 6.654 41.126 6.706 41.162 ;
      RECT 6.654 42.326 6.706 42.362 ;
      RECT 6.654 43.526 6.706 43.562 ;
      RECT 6.654 44.726 6.706 44.762 ;
      RECT 6.654 45.926 6.706 45.962 ;
      RECT 6.654 47.126 6.706 47.162 ;
      RECT 6.654 48.326 6.706 48.362 ;
      RECT 6.654 49.526 6.706 49.562 ;
      RECT 6.654 50.726 6.706 50.762 ;
      RECT 6.654 51.926 6.706 51.962 ;
      RECT 6.654 53.126 6.706 53.162 ;
      RECT 6.654 54.326 6.706 54.362 ;
      RECT 6.654 55.526 6.706 55.562 ;
      RECT 6.654 56.726 6.706 56.762 ;
      RECT 6.654 57.926 6.706 57.962 ;
      RECT 6.654 59.126 6.706 59.162 ;
      RECT 6.654 60.326 6.706 60.362 ;
      RECT 6.654 61.526 6.706 61.562 ;
      RECT 6.654 62.726 6.706 62.762 ;
      RECT 6.654 63.926 6.706 63.962 ;
      RECT 6.654 65.126 6.706 65.162 ;
      RECT 6.654 66.326 6.706 66.362 ;
      RECT 6.654 67.526 6.706 67.562 ;
      RECT 6.654 68.726 6.706 68.762 ;
      RECT 6.654 69.926 6.706 69.962 ;
      RECT 6.654 71.126 6.706 71.162 ;
      RECT 6.734 1.558 6.786 1.594 ;
      RECT 6.734 2.758 6.786 2.794 ;
      RECT 6.734 3.958 6.786 3.994 ;
      RECT 6.734 5.158 6.786 5.194 ;
      RECT 6.734 6.358 6.786 6.394 ;
      RECT 6.734 7.558 6.786 7.594 ;
      RECT 6.734 8.758 6.786 8.794 ;
      RECT 6.734 9.958 6.786 9.994 ;
      RECT 6.734 11.158 6.786 11.194 ;
      RECT 6.734 12.358 6.786 12.394 ;
      RECT 6.734 13.558 6.786 13.594 ;
      RECT 6.734 14.758 6.786 14.794 ;
      RECT 6.734 15.958 6.786 15.994 ;
      RECT 6.734 17.158 6.786 17.194 ;
      RECT 6.734 18.358 6.786 18.394 ;
      RECT 6.734 19.558 6.786 19.594 ;
      RECT 6.734 20.758 6.786 20.794 ;
      RECT 6.734 21.958 6.786 21.994 ;
      RECT 6.734 23.158 6.786 23.194 ;
      RECT 6.734 24.358 6.786 24.394 ;
      RECT 6.734 25.558 6.786 25.594 ;
      RECT 6.734 26.758 6.786 26.794 ;
      RECT 6.734 27.958 6.786 27.994 ;
      RECT 6.734 29.158 6.786 29.194 ;
      RECT 6.734 30.358 6.786 30.394 ;
      RECT 6.734 31.558 6.786 31.594 ;
      RECT 6.734 33.342 6.786 33.378 ;
      RECT 6.734 33.582 6.786 33.618 ;
      RECT 6.734 37.902 6.786 37.938 ;
      RECT 6.734 38.142 6.786 38.178 ;
      RECT 6.734 40.678 6.786 40.714 ;
      RECT 6.734 41.878 6.786 41.914 ;
      RECT 6.734 43.078 6.786 43.114 ;
      RECT 6.734 44.278 6.786 44.314 ;
      RECT 6.734 45.478 6.786 45.514 ;
      RECT 6.734 46.678 6.786 46.714 ;
      RECT 6.734 47.878 6.786 47.914 ;
      RECT 6.734 49.078 6.786 49.114 ;
      RECT 6.734 50.278 6.786 50.314 ;
      RECT 6.734 51.478 6.786 51.514 ;
      RECT 6.734 52.678 6.786 52.714 ;
      RECT 6.734 53.878 6.786 53.914 ;
      RECT 6.734 55.078 6.786 55.114 ;
      RECT 6.734 56.278 6.786 56.314 ;
      RECT 6.734 57.478 6.786 57.514 ;
      RECT 6.734 58.678 6.786 58.714 ;
      RECT 6.734 59.878 6.786 59.914 ;
      RECT 6.734 61.078 6.786 61.114 ;
      RECT 6.734 62.278 6.786 62.314 ;
      RECT 6.734 63.478 6.786 63.514 ;
      RECT 6.734 64.678 6.786 64.714 ;
      RECT 6.734 65.878 6.786 65.914 ;
      RECT 6.734 67.078 6.786 67.114 ;
      RECT 6.734 68.278 6.786 68.314 ;
      RECT 6.734 69.478 6.786 69.514 ;
      RECT 6.734 70.678 6.786 70.714 ;
      RECT 6.734 71.878 6.786 71.914 ;
      RECT 6.814 0.806 6.866 0.842 ;
      RECT 6.814 2.006 6.866 2.042 ;
      RECT 6.814 3.206 6.866 3.242 ;
      RECT 6.814 4.406 6.866 4.442 ;
      RECT 6.814 5.606 6.866 5.642 ;
      RECT 6.814 6.806 6.866 6.842 ;
      RECT 6.814 8.006 6.866 8.042 ;
      RECT 6.814 9.206 6.866 9.242 ;
      RECT 6.814 10.406 6.866 10.442 ;
      RECT 6.814 11.606 6.866 11.642 ;
      RECT 6.814 12.806 6.866 12.842 ;
      RECT 6.814 14.006 6.866 14.042 ;
      RECT 6.814 15.206 6.866 15.242 ;
      RECT 6.814 16.406 6.866 16.442 ;
      RECT 6.814 17.606 6.866 17.642 ;
      RECT 6.814 18.806 6.866 18.842 ;
      RECT 6.814 20.006 6.866 20.042 ;
      RECT 6.814 21.206 6.866 21.242 ;
      RECT 6.814 22.406 6.866 22.442 ;
      RECT 6.814 23.606 6.866 23.642 ;
      RECT 6.814 24.806 6.866 24.842 ;
      RECT 6.814 26.006 6.866 26.042 ;
      RECT 6.814 27.206 6.866 27.242 ;
      RECT 6.814 28.406 6.866 28.442 ;
      RECT 6.814 29.606 6.866 29.642 ;
      RECT 6.814 30.806 6.866 30.842 ;
      RECT 6.814 32.622 6.866 32.658 ;
      RECT 6.814 32.862 6.866 32.898 ;
      RECT 6.814 38.622 6.866 38.658 ;
      RECT 6.814 38.862 6.866 38.898 ;
      RECT 6.814 39.926 6.866 39.962 ;
      RECT 6.814 41.126 6.866 41.162 ;
      RECT 6.814 42.326 6.866 42.362 ;
      RECT 6.814 43.526 6.866 43.562 ;
      RECT 6.814 44.726 6.866 44.762 ;
      RECT 6.814 45.926 6.866 45.962 ;
      RECT 6.814 47.126 6.866 47.162 ;
      RECT 6.814 48.326 6.866 48.362 ;
      RECT 6.814 49.526 6.866 49.562 ;
      RECT 6.814 50.726 6.866 50.762 ;
      RECT 6.814 51.926 6.866 51.962 ;
      RECT 6.814 53.126 6.866 53.162 ;
      RECT 6.814 54.326 6.866 54.362 ;
      RECT 6.814 55.526 6.866 55.562 ;
      RECT 6.814 56.726 6.866 56.762 ;
      RECT 6.814 57.926 6.866 57.962 ;
      RECT 6.814 59.126 6.866 59.162 ;
      RECT 6.814 60.326 6.866 60.362 ;
      RECT 6.814 61.526 6.866 61.562 ;
      RECT 6.814 62.726 6.866 62.762 ;
      RECT 6.814 63.926 6.866 63.962 ;
      RECT 6.814 65.126 6.866 65.162 ;
      RECT 6.814 66.326 6.866 66.362 ;
      RECT 6.814 67.526 6.866 67.562 ;
      RECT 6.814 68.726 6.866 68.762 ;
      RECT 6.814 69.926 6.866 69.962 ;
      RECT 6.814 71.126 6.866 71.162 ;
      RECT 6.894 1.558 6.946 1.594 ;
      RECT 6.894 2.758 6.946 2.794 ;
      RECT 6.894 3.958 6.946 3.994 ;
      RECT 6.894 5.158 6.946 5.194 ;
      RECT 6.894 6.358 6.946 6.394 ;
      RECT 6.894 7.558 6.946 7.594 ;
      RECT 6.894 8.758 6.946 8.794 ;
      RECT 6.894 9.958 6.946 9.994 ;
      RECT 6.894 11.158 6.946 11.194 ;
      RECT 6.894 12.358 6.946 12.394 ;
      RECT 6.894 13.558 6.946 13.594 ;
      RECT 6.894 14.758 6.946 14.794 ;
      RECT 6.894 15.958 6.946 15.994 ;
      RECT 6.894 17.158 6.946 17.194 ;
      RECT 6.894 18.358 6.946 18.394 ;
      RECT 6.894 19.558 6.946 19.594 ;
      RECT 6.894 20.758 6.946 20.794 ;
      RECT 6.894 21.958 6.946 21.994 ;
      RECT 6.894 23.158 6.946 23.194 ;
      RECT 6.894 24.358 6.946 24.394 ;
      RECT 6.894 25.558 6.946 25.594 ;
      RECT 6.894 26.758 6.946 26.794 ;
      RECT 6.894 27.958 6.946 27.994 ;
      RECT 6.894 29.158 6.946 29.194 ;
      RECT 6.894 30.358 6.946 30.394 ;
      RECT 6.894 31.558 6.946 31.594 ;
      RECT 6.894 33.342 6.946 33.378 ;
      RECT 6.894 33.582 6.946 33.618 ;
      RECT 6.894 37.902 6.946 37.938 ;
      RECT 6.894 38.142 6.946 38.178 ;
      RECT 6.894 40.678 6.946 40.714 ;
      RECT 6.894 41.878 6.946 41.914 ;
      RECT 6.894 43.078 6.946 43.114 ;
      RECT 6.894 44.278 6.946 44.314 ;
      RECT 6.894 45.478 6.946 45.514 ;
      RECT 6.894 46.678 6.946 46.714 ;
      RECT 6.894 47.878 6.946 47.914 ;
      RECT 6.894 49.078 6.946 49.114 ;
      RECT 6.894 50.278 6.946 50.314 ;
      RECT 6.894 51.478 6.946 51.514 ;
      RECT 6.894 52.678 6.946 52.714 ;
      RECT 6.894 53.878 6.946 53.914 ;
      RECT 6.894 55.078 6.946 55.114 ;
      RECT 6.894 56.278 6.946 56.314 ;
      RECT 6.894 57.478 6.946 57.514 ;
      RECT 6.894 58.678 6.946 58.714 ;
      RECT 6.894 59.878 6.946 59.914 ;
      RECT 6.894 61.078 6.946 61.114 ;
      RECT 6.894 62.278 6.946 62.314 ;
      RECT 6.894 63.478 6.946 63.514 ;
      RECT 6.894 64.678 6.946 64.714 ;
      RECT 6.894 65.878 6.946 65.914 ;
      RECT 6.894 67.078 6.946 67.114 ;
      RECT 6.894 68.278 6.946 68.314 ;
      RECT 6.894 69.478 6.946 69.514 ;
      RECT 6.894 70.678 6.946 70.714 ;
      RECT 6.894 71.878 6.946 71.914 ;
      RECT 6.974 0.281 7.026 0.317 ;
      RECT 6.974 72.403 7.026 72.439 ;
      RECT 7.054 0.806 7.106 0.842 ;
      RECT 7.054 2.006 7.106 2.042 ;
      RECT 7.054 3.206 7.106 3.242 ;
      RECT 7.054 4.406 7.106 4.442 ;
      RECT 7.054 5.606 7.106 5.642 ;
      RECT 7.054 6.806 7.106 6.842 ;
      RECT 7.054 8.006 7.106 8.042 ;
      RECT 7.054 9.206 7.106 9.242 ;
      RECT 7.054 10.406 7.106 10.442 ;
      RECT 7.054 11.606 7.106 11.642 ;
      RECT 7.054 12.806 7.106 12.842 ;
      RECT 7.054 14.006 7.106 14.042 ;
      RECT 7.054 15.206 7.106 15.242 ;
      RECT 7.054 16.406 7.106 16.442 ;
      RECT 7.054 17.606 7.106 17.642 ;
      RECT 7.054 18.806 7.106 18.842 ;
      RECT 7.054 20.006 7.106 20.042 ;
      RECT 7.054 21.206 7.106 21.242 ;
      RECT 7.054 22.406 7.106 22.442 ;
      RECT 7.054 23.606 7.106 23.642 ;
      RECT 7.054 24.806 7.106 24.842 ;
      RECT 7.054 26.006 7.106 26.042 ;
      RECT 7.054 27.206 7.106 27.242 ;
      RECT 7.054 28.406 7.106 28.442 ;
      RECT 7.054 29.606 7.106 29.642 ;
      RECT 7.054 30.806 7.106 30.842 ;
      RECT 7.054 32.622 7.106 32.658 ;
      RECT 7.054 32.862 7.106 32.898 ;
      RECT 7.054 38.622 7.106 38.658 ;
      RECT 7.054 38.862 7.106 38.898 ;
      RECT 7.054 39.926 7.106 39.962 ;
      RECT 7.054 41.126 7.106 41.162 ;
      RECT 7.054 42.326 7.106 42.362 ;
      RECT 7.054 43.526 7.106 43.562 ;
      RECT 7.054 44.726 7.106 44.762 ;
      RECT 7.054 45.926 7.106 45.962 ;
      RECT 7.054 47.126 7.106 47.162 ;
      RECT 7.054 48.326 7.106 48.362 ;
      RECT 7.054 49.526 7.106 49.562 ;
      RECT 7.054 50.726 7.106 50.762 ;
      RECT 7.054 51.926 7.106 51.962 ;
      RECT 7.054 53.126 7.106 53.162 ;
      RECT 7.054 54.326 7.106 54.362 ;
      RECT 7.054 55.526 7.106 55.562 ;
      RECT 7.054 56.726 7.106 56.762 ;
      RECT 7.054 57.926 7.106 57.962 ;
      RECT 7.054 59.126 7.106 59.162 ;
      RECT 7.054 60.326 7.106 60.362 ;
      RECT 7.054 61.526 7.106 61.562 ;
      RECT 7.054 62.726 7.106 62.762 ;
      RECT 7.054 63.926 7.106 63.962 ;
      RECT 7.054 65.126 7.106 65.162 ;
      RECT 7.054 66.326 7.106 66.362 ;
      RECT 7.054 67.526 7.106 67.562 ;
      RECT 7.054 68.726 7.106 68.762 ;
      RECT 7.054 69.926 7.106 69.962 ;
      RECT 7.054 71.126 7.106 71.162 ;
      RECT 7.134 1.558 7.186 1.594 ;
      RECT 7.134 2.758 7.186 2.794 ;
      RECT 7.134 3.958 7.186 3.994 ;
      RECT 7.134 5.158 7.186 5.194 ;
      RECT 7.134 6.358 7.186 6.394 ;
      RECT 7.134 7.558 7.186 7.594 ;
      RECT 7.134 8.758 7.186 8.794 ;
      RECT 7.134 9.958 7.186 9.994 ;
      RECT 7.134 11.158 7.186 11.194 ;
      RECT 7.134 12.358 7.186 12.394 ;
      RECT 7.134 13.558 7.186 13.594 ;
      RECT 7.134 14.758 7.186 14.794 ;
      RECT 7.134 15.958 7.186 15.994 ;
      RECT 7.134 17.158 7.186 17.194 ;
      RECT 7.134 18.358 7.186 18.394 ;
      RECT 7.134 19.558 7.186 19.594 ;
      RECT 7.134 20.758 7.186 20.794 ;
      RECT 7.134 21.958 7.186 21.994 ;
      RECT 7.134 23.158 7.186 23.194 ;
      RECT 7.134 24.358 7.186 24.394 ;
      RECT 7.134 25.558 7.186 25.594 ;
      RECT 7.134 26.758 7.186 26.794 ;
      RECT 7.134 27.958 7.186 27.994 ;
      RECT 7.134 29.158 7.186 29.194 ;
      RECT 7.134 30.358 7.186 30.394 ;
      RECT 7.134 31.558 7.186 31.594 ;
      RECT 7.134 33.342 7.186 33.378 ;
      RECT 7.134 33.582 7.186 33.618 ;
      RECT 7.134 37.902 7.186 37.938 ;
      RECT 7.134 38.142 7.186 38.178 ;
      RECT 7.134 40.678 7.186 40.714 ;
      RECT 7.134 41.878 7.186 41.914 ;
      RECT 7.134 43.078 7.186 43.114 ;
      RECT 7.134 44.278 7.186 44.314 ;
      RECT 7.134 45.478 7.186 45.514 ;
      RECT 7.134 46.678 7.186 46.714 ;
      RECT 7.134 47.878 7.186 47.914 ;
      RECT 7.134 49.078 7.186 49.114 ;
      RECT 7.134 50.278 7.186 50.314 ;
      RECT 7.134 51.478 7.186 51.514 ;
      RECT 7.134 52.678 7.186 52.714 ;
      RECT 7.134 53.878 7.186 53.914 ;
      RECT 7.134 55.078 7.186 55.114 ;
      RECT 7.134 56.278 7.186 56.314 ;
      RECT 7.134 57.478 7.186 57.514 ;
      RECT 7.134 58.678 7.186 58.714 ;
      RECT 7.134 59.878 7.186 59.914 ;
      RECT 7.134 61.078 7.186 61.114 ;
      RECT 7.134 62.278 7.186 62.314 ;
      RECT 7.134 63.478 7.186 63.514 ;
      RECT 7.134 64.678 7.186 64.714 ;
      RECT 7.134 65.878 7.186 65.914 ;
      RECT 7.134 67.078 7.186 67.114 ;
      RECT 7.134 68.278 7.186 68.314 ;
      RECT 7.134 69.478 7.186 69.514 ;
      RECT 7.134 70.678 7.186 70.714 ;
      RECT 7.134 71.878 7.186 71.914 ;
      RECT 7.214 0.806 7.266 0.842 ;
      RECT 7.214 2.006 7.266 2.042 ;
      RECT 7.214 3.206 7.266 3.242 ;
      RECT 7.214 4.406 7.266 4.442 ;
      RECT 7.214 5.606 7.266 5.642 ;
      RECT 7.214 6.806 7.266 6.842 ;
      RECT 7.214 8.006 7.266 8.042 ;
      RECT 7.214 9.206 7.266 9.242 ;
      RECT 7.214 10.406 7.266 10.442 ;
      RECT 7.214 11.606 7.266 11.642 ;
      RECT 7.214 12.806 7.266 12.842 ;
      RECT 7.214 14.006 7.266 14.042 ;
      RECT 7.214 15.206 7.266 15.242 ;
      RECT 7.214 16.406 7.266 16.442 ;
      RECT 7.214 17.606 7.266 17.642 ;
      RECT 7.214 18.806 7.266 18.842 ;
      RECT 7.214 20.006 7.266 20.042 ;
      RECT 7.214 21.206 7.266 21.242 ;
      RECT 7.214 22.406 7.266 22.442 ;
      RECT 7.214 23.606 7.266 23.642 ;
      RECT 7.214 24.806 7.266 24.842 ;
      RECT 7.214 26.006 7.266 26.042 ;
      RECT 7.214 27.206 7.266 27.242 ;
      RECT 7.214 28.406 7.266 28.442 ;
      RECT 7.214 29.606 7.266 29.642 ;
      RECT 7.214 30.806 7.266 30.842 ;
      RECT 7.214 32.622 7.266 32.658 ;
      RECT 7.214 32.862 7.266 32.898 ;
      RECT 7.214 38.622 7.266 38.658 ;
      RECT 7.214 38.862 7.266 38.898 ;
      RECT 7.214 39.926 7.266 39.962 ;
      RECT 7.214 41.126 7.266 41.162 ;
      RECT 7.214 42.326 7.266 42.362 ;
      RECT 7.214 43.526 7.266 43.562 ;
      RECT 7.214 44.726 7.266 44.762 ;
      RECT 7.214 45.926 7.266 45.962 ;
      RECT 7.214 47.126 7.266 47.162 ;
      RECT 7.214 48.326 7.266 48.362 ;
      RECT 7.214 49.526 7.266 49.562 ;
      RECT 7.214 50.726 7.266 50.762 ;
      RECT 7.214 51.926 7.266 51.962 ;
      RECT 7.214 53.126 7.266 53.162 ;
      RECT 7.214 54.326 7.266 54.362 ;
      RECT 7.214 55.526 7.266 55.562 ;
      RECT 7.214 56.726 7.266 56.762 ;
      RECT 7.214 57.926 7.266 57.962 ;
      RECT 7.214 59.126 7.266 59.162 ;
      RECT 7.214 60.326 7.266 60.362 ;
      RECT 7.214 61.526 7.266 61.562 ;
      RECT 7.214 62.726 7.266 62.762 ;
      RECT 7.214 63.926 7.266 63.962 ;
      RECT 7.214 65.126 7.266 65.162 ;
      RECT 7.214 66.326 7.266 66.362 ;
      RECT 7.214 67.526 7.266 67.562 ;
      RECT 7.214 68.726 7.266 68.762 ;
      RECT 7.214 69.926 7.266 69.962 ;
      RECT 7.214 71.126 7.266 71.162 ;
      RECT 7.294 1.558 7.346 1.594 ;
      RECT 7.294 2.758 7.346 2.794 ;
      RECT 7.294 3.958 7.346 3.994 ;
      RECT 7.294 5.158 7.346 5.194 ;
      RECT 7.294 6.358 7.346 6.394 ;
      RECT 7.294 7.558 7.346 7.594 ;
      RECT 7.294 8.758 7.346 8.794 ;
      RECT 7.294 9.958 7.346 9.994 ;
      RECT 7.294 11.158 7.346 11.194 ;
      RECT 7.294 12.358 7.346 12.394 ;
      RECT 7.294 13.558 7.346 13.594 ;
      RECT 7.294 14.758 7.346 14.794 ;
      RECT 7.294 15.958 7.346 15.994 ;
      RECT 7.294 17.158 7.346 17.194 ;
      RECT 7.294 18.358 7.346 18.394 ;
      RECT 7.294 19.558 7.346 19.594 ;
      RECT 7.294 20.758 7.346 20.794 ;
      RECT 7.294 21.958 7.346 21.994 ;
      RECT 7.294 23.158 7.346 23.194 ;
      RECT 7.294 24.358 7.346 24.394 ;
      RECT 7.294 25.558 7.346 25.594 ;
      RECT 7.294 26.758 7.346 26.794 ;
      RECT 7.294 27.958 7.346 27.994 ;
      RECT 7.294 29.158 7.346 29.194 ;
      RECT 7.294 30.358 7.346 30.394 ;
      RECT 7.294 31.558 7.346 31.594 ;
      RECT 7.294 33.342 7.346 33.378 ;
      RECT 7.294 33.582 7.346 33.618 ;
      RECT 7.294 37.902 7.346 37.938 ;
      RECT 7.294 38.142 7.346 38.178 ;
      RECT 7.294 40.678 7.346 40.714 ;
      RECT 7.294 41.878 7.346 41.914 ;
      RECT 7.294 43.078 7.346 43.114 ;
      RECT 7.294 44.278 7.346 44.314 ;
      RECT 7.294 45.478 7.346 45.514 ;
      RECT 7.294 46.678 7.346 46.714 ;
      RECT 7.294 47.878 7.346 47.914 ;
      RECT 7.294 49.078 7.346 49.114 ;
      RECT 7.294 50.278 7.346 50.314 ;
      RECT 7.294 51.478 7.346 51.514 ;
      RECT 7.294 52.678 7.346 52.714 ;
      RECT 7.294 53.878 7.346 53.914 ;
      RECT 7.294 55.078 7.346 55.114 ;
      RECT 7.294 56.278 7.346 56.314 ;
      RECT 7.294 57.478 7.346 57.514 ;
      RECT 7.294 58.678 7.346 58.714 ;
      RECT 7.294 59.878 7.346 59.914 ;
      RECT 7.294 61.078 7.346 61.114 ;
      RECT 7.294 62.278 7.346 62.314 ;
      RECT 7.294 63.478 7.346 63.514 ;
      RECT 7.294 64.678 7.346 64.714 ;
      RECT 7.294 65.878 7.346 65.914 ;
      RECT 7.294 67.078 7.346 67.114 ;
      RECT 7.294 68.278 7.346 68.314 ;
      RECT 7.294 69.478 7.346 69.514 ;
      RECT 7.294 70.678 7.346 70.714 ;
      RECT 7.294 71.878 7.346 71.914 ;
      RECT 7.374 0.281 7.426 0.317 ;
      RECT 7.374 72.403 7.426 72.439 ;
      RECT 7.454 0.806 7.506 0.842 ;
      RECT 7.454 2.006 7.506 2.042 ;
      RECT 7.454 3.206 7.506 3.242 ;
      RECT 7.454 4.406 7.506 4.442 ;
      RECT 7.454 5.606 7.506 5.642 ;
      RECT 7.454 6.806 7.506 6.842 ;
      RECT 7.454 8.006 7.506 8.042 ;
      RECT 7.454 9.206 7.506 9.242 ;
      RECT 7.454 10.406 7.506 10.442 ;
      RECT 7.454 11.606 7.506 11.642 ;
      RECT 7.454 12.806 7.506 12.842 ;
      RECT 7.454 14.006 7.506 14.042 ;
      RECT 7.454 15.206 7.506 15.242 ;
      RECT 7.454 16.406 7.506 16.442 ;
      RECT 7.454 17.606 7.506 17.642 ;
      RECT 7.454 18.806 7.506 18.842 ;
      RECT 7.454 20.006 7.506 20.042 ;
      RECT 7.454 21.206 7.506 21.242 ;
      RECT 7.454 22.406 7.506 22.442 ;
      RECT 7.454 23.606 7.506 23.642 ;
      RECT 7.454 24.806 7.506 24.842 ;
      RECT 7.454 26.006 7.506 26.042 ;
      RECT 7.454 27.206 7.506 27.242 ;
      RECT 7.454 28.406 7.506 28.442 ;
      RECT 7.454 29.606 7.506 29.642 ;
      RECT 7.454 30.806 7.506 30.842 ;
      RECT 7.454 32.622 7.506 32.658 ;
      RECT 7.454 32.862 7.506 32.898 ;
      RECT 7.454 34.302 7.506 34.338 ;
      RECT 7.454 34.782 7.506 34.818 ;
      RECT 7.454 36.702 7.506 36.738 ;
      RECT 7.454 37.182 7.506 37.218 ;
      RECT 7.454 38.622 7.506 38.658 ;
      RECT 7.454 38.862 7.506 38.898 ;
      RECT 7.454 39.926 7.506 39.962 ;
      RECT 7.454 41.126 7.506 41.162 ;
      RECT 7.454 42.326 7.506 42.362 ;
      RECT 7.454 43.526 7.506 43.562 ;
      RECT 7.454 44.726 7.506 44.762 ;
      RECT 7.454 45.926 7.506 45.962 ;
      RECT 7.454 47.126 7.506 47.162 ;
      RECT 7.454 48.326 7.506 48.362 ;
      RECT 7.454 49.526 7.506 49.562 ;
      RECT 7.454 50.726 7.506 50.762 ;
      RECT 7.454 51.926 7.506 51.962 ;
      RECT 7.454 53.126 7.506 53.162 ;
      RECT 7.454 54.326 7.506 54.362 ;
      RECT 7.454 55.526 7.506 55.562 ;
      RECT 7.454 56.726 7.506 56.762 ;
      RECT 7.454 57.926 7.506 57.962 ;
      RECT 7.454 59.126 7.506 59.162 ;
      RECT 7.454 60.326 7.506 60.362 ;
      RECT 7.454 61.526 7.506 61.562 ;
      RECT 7.454 62.726 7.506 62.762 ;
      RECT 7.454 63.926 7.506 63.962 ;
      RECT 7.454 65.126 7.506 65.162 ;
      RECT 7.454 66.326 7.506 66.362 ;
      RECT 7.454 67.526 7.506 67.562 ;
      RECT 7.454 68.726 7.506 68.762 ;
      RECT 7.454 69.926 7.506 69.962 ;
      RECT 7.454 71.126 7.506 71.162 ;
      RECT 7.534 1.558 7.586 1.594 ;
      RECT 7.534 2.758 7.586 2.794 ;
      RECT 7.534 3.958 7.586 3.994 ;
      RECT 7.534 5.158 7.586 5.194 ;
      RECT 7.534 6.358 7.586 6.394 ;
      RECT 7.534 7.558 7.586 7.594 ;
      RECT 7.534 8.758 7.586 8.794 ;
      RECT 7.534 9.958 7.586 9.994 ;
      RECT 7.534 11.158 7.586 11.194 ;
      RECT 7.534 12.358 7.586 12.394 ;
      RECT 7.534 13.558 7.586 13.594 ;
      RECT 7.534 14.758 7.586 14.794 ;
      RECT 7.534 15.958 7.586 15.994 ;
      RECT 7.534 17.158 7.586 17.194 ;
      RECT 7.534 18.358 7.586 18.394 ;
      RECT 7.534 19.558 7.586 19.594 ;
      RECT 7.534 20.758 7.586 20.794 ;
      RECT 7.534 21.958 7.586 21.994 ;
      RECT 7.534 23.158 7.586 23.194 ;
      RECT 7.534 24.358 7.586 24.394 ;
      RECT 7.534 25.558 7.586 25.594 ;
      RECT 7.534 26.758 7.586 26.794 ;
      RECT 7.534 27.958 7.586 27.994 ;
      RECT 7.534 29.158 7.586 29.194 ;
      RECT 7.534 30.358 7.586 30.394 ;
      RECT 7.534 31.558 7.586 31.594 ;
      RECT 7.534 33.342 7.586 33.378 ;
      RECT 7.534 33.582 7.586 33.618 ;
      RECT 7.534 37.902 7.586 37.938 ;
      RECT 7.534 38.142 7.586 38.178 ;
      RECT 7.534 40.678 7.586 40.714 ;
      RECT 7.534 41.878 7.586 41.914 ;
      RECT 7.534 43.078 7.586 43.114 ;
      RECT 7.534 44.278 7.586 44.314 ;
      RECT 7.534 45.478 7.586 45.514 ;
      RECT 7.534 46.678 7.586 46.714 ;
      RECT 7.534 47.878 7.586 47.914 ;
      RECT 7.534 49.078 7.586 49.114 ;
      RECT 7.534 50.278 7.586 50.314 ;
      RECT 7.534 51.478 7.586 51.514 ;
      RECT 7.534 52.678 7.586 52.714 ;
      RECT 7.534 53.878 7.586 53.914 ;
      RECT 7.534 55.078 7.586 55.114 ;
      RECT 7.534 56.278 7.586 56.314 ;
      RECT 7.534 57.478 7.586 57.514 ;
      RECT 7.534 58.678 7.586 58.714 ;
      RECT 7.534 59.878 7.586 59.914 ;
      RECT 7.534 61.078 7.586 61.114 ;
      RECT 7.534 62.278 7.586 62.314 ;
      RECT 7.534 63.478 7.586 63.514 ;
      RECT 7.534 64.678 7.586 64.714 ;
      RECT 7.534 65.878 7.586 65.914 ;
      RECT 7.534 67.078 7.586 67.114 ;
      RECT 7.534 68.278 7.586 68.314 ;
      RECT 7.534 69.478 7.586 69.514 ;
      RECT 7.534 70.678 7.586 70.714 ;
      RECT 7.534 71.878 7.586 71.914 ;
      RECT 7.614 0.806 7.666 0.842 ;
      RECT 7.614 2.006 7.666 2.042 ;
      RECT 7.614 3.206 7.666 3.242 ;
      RECT 7.614 4.406 7.666 4.442 ;
      RECT 7.614 5.606 7.666 5.642 ;
      RECT 7.614 6.806 7.666 6.842 ;
      RECT 7.614 8.006 7.666 8.042 ;
      RECT 7.614 9.206 7.666 9.242 ;
      RECT 7.614 10.406 7.666 10.442 ;
      RECT 7.614 11.606 7.666 11.642 ;
      RECT 7.614 12.806 7.666 12.842 ;
      RECT 7.614 14.006 7.666 14.042 ;
      RECT 7.614 15.206 7.666 15.242 ;
      RECT 7.614 16.406 7.666 16.442 ;
      RECT 7.614 17.606 7.666 17.642 ;
      RECT 7.614 18.806 7.666 18.842 ;
      RECT 7.614 20.006 7.666 20.042 ;
      RECT 7.614 21.206 7.666 21.242 ;
      RECT 7.614 22.406 7.666 22.442 ;
      RECT 7.614 23.606 7.666 23.642 ;
      RECT 7.614 24.806 7.666 24.842 ;
      RECT 7.614 26.006 7.666 26.042 ;
      RECT 7.614 27.206 7.666 27.242 ;
      RECT 7.614 28.406 7.666 28.442 ;
      RECT 7.614 29.606 7.666 29.642 ;
      RECT 7.614 30.806 7.666 30.842 ;
      RECT 7.614 32.622 7.666 32.658 ;
      RECT 7.614 32.862 7.666 32.898 ;
      RECT 7.614 38.622 7.666 38.658 ;
      RECT 7.614 38.862 7.666 38.898 ;
      RECT 7.614 39.926 7.666 39.962 ;
      RECT 7.614 41.126 7.666 41.162 ;
      RECT 7.614 42.326 7.666 42.362 ;
      RECT 7.614 43.526 7.666 43.562 ;
      RECT 7.614 44.726 7.666 44.762 ;
      RECT 7.614 45.926 7.666 45.962 ;
      RECT 7.614 47.126 7.666 47.162 ;
      RECT 7.614 48.326 7.666 48.362 ;
      RECT 7.614 49.526 7.666 49.562 ;
      RECT 7.614 50.726 7.666 50.762 ;
      RECT 7.614 51.926 7.666 51.962 ;
      RECT 7.614 53.126 7.666 53.162 ;
      RECT 7.614 54.326 7.666 54.362 ;
      RECT 7.614 55.526 7.666 55.562 ;
      RECT 7.614 56.726 7.666 56.762 ;
      RECT 7.614 57.926 7.666 57.962 ;
      RECT 7.614 59.126 7.666 59.162 ;
      RECT 7.614 60.326 7.666 60.362 ;
      RECT 7.614 61.526 7.666 61.562 ;
      RECT 7.614 62.726 7.666 62.762 ;
      RECT 7.614 63.926 7.666 63.962 ;
      RECT 7.614 65.126 7.666 65.162 ;
      RECT 7.614 66.326 7.666 66.362 ;
      RECT 7.614 67.526 7.666 67.562 ;
      RECT 7.614 68.726 7.666 68.762 ;
      RECT 7.614 69.926 7.666 69.962 ;
      RECT 7.614 71.126 7.666 71.162 ;
      RECT 7.694 1.558 7.746 1.594 ;
      RECT 7.694 2.758 7.746 2.794 ;
      RECT 7.694 3.958 7.746 3.994 ;
      RECT 7.694 5.158 7.746 5.194 ;
      RECT 7.694 6.358 7.746 6.394 ;
      RECT 7.694 7.558 7.746 7.594 ;
      RECT 7.694 8.758 7.746 8.794 ;
      RECT 7.694 9.958 7.746 9.994 ;
      RECT 7.694 11.158 7.746 11.194 ;
      RECT 7.694 12.358 7.746 12.394 ;
      RECT 7.694 13.558 7.746 13.594 ;
      RECT 7.694 14.758 7.746 14.794 ;
      RECT 7.694 15.958 7.746 15.994 ;
      RECT 7.694 17.158 7.746 17.194 ;
      RECT 7.694 18.358 7.746 18.394 ;
      RECT 7.694 19.558 7.746 19.594 ;
      RECT 7.694 20.758 7.746 20.794 ;
      RECT 7.694 21.958 7.746 21.994 ;
      RECT 7.694 23.158 7.746 23.194 ;
      RECT 7.694 24.358 7.746 24.394 ;
      RECT 7.694 25.558 7.746 25.594 ;
      RECT 7.694 26.758 7.746 26.794 ;
      RECT 7.694 27.958 7.746 27.994 ;
      RECT 7.694 29.158 7.746 29.194 ;
      RECT 7.694 30.358 7.746 30.394 ;
      RECT 7.694 31.558 7.746 31.594 ;
      RECT 7.694 33.342 7.746 33.378 ;
      RECT 7.694 33.582 7.746 33.618 ;
      RECT 7.694 37.902 7.746 37.938 ;
      RECT 7.694 38.142 7.746 38.178 ;
      RECT 7.694 40.678 7.746 40.714 ;
      RECT 7.694 41.878 7.746 41.914 ;
      RECT 7.694 43.078 7.746 43.114 ;
      RECT 7.694 44.278 7.746 44.314 ;
      RECT 7.694 45.478 7.746 45.514 ;
      RECT 7.694 46.678 7.746 46.714 ;
      RECT 7.694 47.878 7.746 47.914 ;
      RECT 7.694 49.078 7.746 49.114 ;
      RECT 7.694 50.278 7.746 50.314 ;
      RECT 7.694 51.478 7.746 51.514 ;
      RECT 7.694 52.678 7.746 52.714 ;
      RECT 7.694 53.878 7.746 53.914 ;
      RECT 7.694 55.078 7.746 55.114 ;
      RECT 7.694 56.278 7.746 56.314 ;
      RECT 7.694 57.478 7.746 57.514 ;
      RECT 7.694 58.678 7.746 58.714 ;
      RECT 7.694 59.878 7.746 59.914 ;
      RECT 7.694 61.078 7.746 61.114 ;
      RECT 7.694 62.278 7.746 62.314 ;
      RECT 7.694 63.478 7.746 63.514 ;
      RECT 7.694 64.678 7.746 64.714 ;
      RECT 7.694 65.878 7.746 65.914 ;
      RECT 7.694 67.078 7.746 67.114 ;
      RECT 7.694 68.278 7.746 68.314 ;
      RECT 7.694 69.478 7.746 69.514 ;
      RECT 7.694 70.678 7.746 70.714 ;
      RECT 7.694 71.878 7.746 71.914 ;
      RECT 7.774 0.281 7.826 0.317 ;
      RECT 7.774 72.403 7.826 72.439 ;
      RECT 7.854 0.806 7.906 0.842 ;
      RECT 7.854 2.006 7.906 2.042 ;
      RECT 7.854 3.206 7.906 3.242 ;
      RECT 7.854 4.406 7.906 4.442 ;
      RECT 7.854 5.606 7.906 5.642 ;
      RECT 7.854 6.806 7.906 6.842 ;
      RECT 7.854 8.006 7.906 8.042 ;
      RECT 7.854 9.206 7.906 9.242 ;
      RECT 7.854 10.406 7.906 10.442 ;
      RECT 7.854 11.606 7.906 11.642 ;
      RECT 7.854 12.806 7.906 12.842 ;
      RECT 7.854 14.006 7.906 14.042 ;
      RECT 7.854 15.206 7.906 15.242 ;
      RECT 7.854 16.406 7.906 16.442 ;
      RECT 7.854 17.606 7.906 17.642 ;
      RECT 7.854 18.806 7.906 18.842 ;
      RECT 7.854 20.006 7.906 20.042 ;
      RECT 7.854 21.206 7.906 21.242 ;
      RECT 7.854 22.406 7.906 22.442 ;
      RECT 7.854 23.606 7.906 23.642 ;
      RECT 7.854 24.806 7.906 24.842 ;
      RECT 7.854 26.006 7.906 26.042 ;
      RECT 7.854 27.206 7.906 27.242 ;
      RECT 7.854 28.406 7.906 28.442 ;
      RECT 7.854 29.606 7.906 29.642 ;
      RECT 7.854 30.806 7.906 30.842 ;
      RECT 7.854 32.622 7.906 32.658 ;
      RECT 7.854 32.862 7.906 32.898 ;
      RECT 7.854 38.622 7.906 38.658 ;
      RECT 7.854 38.862 7.906 38.898 ;
      RECT 7.854 39.926 7.906 39.962 ;
      RECT 7.854 41.126 7.906 41.162 ;
      RECT 7.854 42.326 7.906 42.362 ;
      RECT 7.854 43.526 7.906 43.562 ;
      RECT 7.854 44.726 7.906 44.762 ;
      RECT 7.854 45.926 7.906 45.962 ;
      RECT 7.854 47.126 7.906 47.162 ;
      RECT 7.854 48.326 7.906 48.362 ;
      RECT 7.854 49.526 7.906 49.562 ;
      RECT 7.854 50.726 7.906 50.762 ;
      RECT 7.854 51.926 7.906 51.962 ;
      RECT 7.854 53.126 7.906 53.162 ;
      RECT 7.854 54.326 7.906 54.362 ;
      RECT 7.854 55.526 7.906 55.562 ;
      RECT 7.854 56.726 7.906 56.762 ;
      RECT 7.854 57.926 7.906 57.962 ;
      RECT 7.854 59.126 7.906 59.162 ;
      RECT 7.854 60.326 7.906 60.362 ;
      RECT 7.854 61.526 7.906 61.562 ;
      RECT 7.854 62.726 7.906 62.762 ;
      RECT 7.854 63.926 7.906 63.962 ;
      RECT 7.854 65.126 7.906 65.162 ;
      RECT 7.854 66.326 7.906 66.362 ;
      RECT 7.854 67.526 7.906 67.562 ;
      RECT 7.854 68.726 7.906 68.762 ;
      RECT 7.854 69.926 7.906 69.962 ;
      RECT 7.854 71.126 7.906 71.162 ;
      RECT 7.934 1.558 7.986 1.594 ;
      RECT 7.934 2.758 7.986 2.794 ;
      RECT 7.934 3.958 7.986 3.994 ;
      RECT 7.934 5.158 7.986 5.194 ;
      RECT 7.934 6.358 7.986 6.394 ;
      RECT 7.934 7.558 7.986 7.594 ;
      RECT 7.934 8.758 7.986 8.794 ;
      RECT 7.934 9.958 7.986 9.994 ;
      RECT 7.934 11.158 7.986 11.194 ;
      RECT 7.934 12.358 7.986 12.394 ;
      RECT 7.934 13.558 7.986 13.594 ;
      RECT 7.934 14.758 7.986 14.794 ;
      RECT 7.934 15.958 7.986 15.994 ;
      RECT 7.934 17.158 7.986 17.194 ;
      RECT 7.934 18.358 7.986 18.394 ;
      RECT 7.934 19.558 7.986 19.594 ;
      RECT 7.934 20.758 7.986 20.794 ;
      RECT 7.934 21.958 7.986 21.994 ;
      RECT 7.934 23.158 7.986 23.194 ;
      RECT 7.934 24.358 7.986 24.394 ;
      RECT 7.934 25.558 7.986 25.594 ;
      RECT 7.934 26.758 7.986 26.794 ;
      RECT 7.934 27.958 7.986 27.994 ;
      RECT 7.934 29.158 7.986 29.194 ;
      RECT 7.934 30.358 7.986 30.394 ;
      RECT 7.934 31.558 7.986 31.594 ;
      RECT 7.934 33.342 7.986 33.378 ;
      RECT 7.934 33.582 7.986 33.618 ;
      RECT 7.934 37.902 7.986 37.938 ;
      RECT 7.934 38.142 7.986 38.178 ;
      RECT 7.934 40.678 7.986 40.714 ;
      RECT 7.934 41.878 7.986 41.914 ;
      RECT 7.934 43.078 7.986 43.114 ;
      RECT 7.934 44.278 7.986 44.314 ;
      RECT 7.934 45.478 7.986 45.514 ;
      RECT 7.934 46.678 7.986 46.714 ;
      RECT 7.934 47.878 7.986 47.914 ;
      RECT 7.934 49.078 7.986 49.114 ;
      RECT 7.934 50.278 7.986 50.314 ;
      RECT 7.934 51.478 7.986 51.514 ;
      RECT 7.934 52.678 7.986 52.714 ;
      RECT 7.934 53.878 7.986 53.914 ;
      RECT 7.934 55.078 7.986 55.114 ;
      RECT 7.934 56.278 7.986 56.314 ;
      RECT 7.934 57.478 7.986 57.514 ;
      RECT 7.934 58.678 7.986 58.714 ;
      RECT 7.934 59.878 7.986 59.914 ;
      RECT 7.934 61.078 7.986 61.114 ;
      RECT 7.934 62.278 7.986 62.314 ;
      RECT 7.934 63.478 7.986 63.514 ;
      RECT 7.934 64.678 7.986 64.714 ;
      RECT 7.934 65.878 7.986 65.914 ;
      RECT 7.934 67.078 7.986 67.114 ;
      RECT 7.934 68.278 7.986 68.314 ;
      RECT 7.934 69.478 7.986 69.514 ;
      RECT 7.934 70.678 7.986 70.714 ;
      RECT 7.934 71.878 7.986 71.914 ;
      RECT 8.014 0.806 8.066 0.842 ;
      RECT 8.014 2.006 8.066 2.042 ;
      RECT 8.014 3.206 8.066 3.242 ;
      RECT 8.014 4.406 8.066 4.442 ;
      RECT 8.014 5.606 8.066 5.642 ;
      RECT 8.014 6.806 8.066 6.842 ;
      RECT 8.014 8.006 8.066 8.042 ;
      RECT 8.014 9.206 8.066 9.242 ;
      RECT 8.014 10.406 8.066 10.442 ;
      RECT 8.014 11.606 8.066 11.642 ;
      RECT 8.014 12.806 8.066 12.842 ;
      RECT 8.014 14.006 8.066 14.042 ;
      RECT 8.014 15.206 8.066 15.242 ;
      RECT 8.014 16.406 8.066 16.442 ;
      RECT 8.014 17.606 8.066 17.642 ;
      RECT 8.014 18.806 8.066 18.842 ;
      RECT 8.014 20.006 8.066 20.042 ;
      RECT 8.014 21.206 8.066 21.242 ;
      RECT 8.014 22.406 8.066 22.442 ;
      RECT 8.014 23.606 8.066 23.642 ;
      RECT 8.014 24.806 8.066 24.842 ;
      RECT 8.014 26.006 8.066 26.042 ;
      RECT 8.014 27.206 8.066 27.242 ;
      RECT 8.014 28.406 8.066 28.442 ;
      RECT 8.014 29.606 8.066 29.642 ;
      RECT 8.014 30.806 8.066 30.842 ;
      RECT 8.014 32.622 8.066 32.658 ;
      RECT 8.014 32.862 8.066 32.898 ;
      RECT 8.014 38.622 8.066 38.658 ;
      RECT 8.014 38.862 8.066 38.898 ;
      RECT 8.014 39.926 8.066 39.962 ;
      RECT 8.014 41.126 8.066 41.162 ;
      RECT 8.014 42.326 8.066 42.362 ;
      RECT 8.014 43.526 8.066 43.562 ;
      RECT 8.014 44.726 8.066 44.762 ;
      RECT 8.014 45.926 8.066 45.962 ;
      RECT 8.014 47.126 8.066 47.162 ;
      RECT 8.014 48.326 8.066 48.362 ;
      RECT 8.014 49.526 8.066 49.562 ;
      RECT 8.014 50.726 8.066 50.762 ;
      RECT 8.014 51.926 8.066 51.962 ;
      RECT 8.014 53.126 8.066 53.162 ;
      RECT 8.014 54.326 8.066 54.362 ;
      RECT 8.014 55.526 8.066 55.562 ;
      RECT 8.014 56.726 8.066 56.762 ;
      RECT 8.014 57.926 8.066 57.962 ;
      RECT 8.014 59.126 8.066 59.162 ;
      RECT 8.014 60.326 8.066 60.362 ;
      RECT 8.014 61.526 8.066 61.562 ;
      RECT 8.014 62.726 8.066 62.762 ;
      RECT 8.014 63.926 8.066 63.962 ;
      RECT 8.014 65.126 8.066 65.162 ;
      RECT 8.014 66.326 8.066 66.362 ;
      RECT 8.014 67.526 8.066 67.562 ;
      RECT 8.014 68.726 8.066 68.762 ;
      RECT 8.014 69.926 8.066 69.962 ;
      RECT 8.014 71.126 8.066 71.162 ;
      RECT 8.094 1.558 8.146 1.594 ;
      RECT 8.094 2.758 8.146 2.794 ;
      RECT 8.094 3.958 8.146 3.994 ;
      RECT 8.094 5.158 8.146 5.194 ;
      RECT 8.094 6.358 8.146 6.394 ;
      RECT 8.094 7.558 8.146 7.594 ;
      RECT 8.094 8.758 8.146 8.794 ;
      RECT 8.094 9.958 8.146 9.994 ;
      RECT 8.094 11.158 8.146 11.194 ;
      RECT 8.094 12.358 8.146 12.394 ;
      RECT 8.094 13.558 8.146 13.594 ;
      RECT 8.094 14.758 8.146 14.794 ;
      RECT 8.094 15.958 8.146 15.994 ;
      RECT 8.094 17.158 8.146 17.194 ;
      RECT 8.094 18.358 8.146 18.394 ;
      RECT 8.094 19.558 8.146 19.594 ;
      RECT 8.094 20.758 8.146 20.794 ;
      RECT 8.094 21.958 8.146 21.994 ;
      RECT 8.094 23.158 8.146 23.194 ;
      RECT 8.094 24.358 8.146 24.394 ;
      RECT 8.094 25.558 8.146 25.594 ;
      RECT 8.094 26.758 8.146 26.794 ;
      RECT 8.094 27.958 8.146 27.994 ;
      RECT 8.094 29.158 8.146 29.194 ;
      RECT 8.094 30.358 8.146 30.394 ;
      RECT 8.094 31.558 8.146 31.594 ;
      RECT 8.094 33.342 8.146 33.378 ;
      RECT 8.094 33.582 8.146 33.618 ;
      RECT 8.094 37.902 8.146 37.938 ;
      RECT 8.094 38.142 8.146 38.178 ;
      RECT 8.094 40.678 8.146 40.714 ;
      RECT 8.094 41.878 8.146 41.914 ;
      RECT 8.094 43.078 8.146 43.114 ;
      RECT 8.094 44.278 8.146 44.314 ;
      RECT 8.094 45.478 8.146 45.514 ;
      RECT 8.094 46.678 8.146 46.714 ;
      RECT 8.094 47.878 8.146 47.914 ;
      RECT 8.094 49.078 8.146 49.114 ;
      RECT 8.094 50.278 8.146 50.314 ;
      RECT 8.094 51.478 8.146 51.514 ;
      RECT 8.094 52.678 8.146 52.714 ;
      RECT 8.094 53.878 8.146 53.914 ;
      RECT 8.094 55.078 8.146 55.114 ;
      RECT 8.094 56.278 8.146 56.314 ;
      RECT 8.094 57.478 8.146 57.514 ;
      RECT 8.094 58.678 8.146 58.714 ;
      RECT 8.094 59.878 8.146 59.914 ;
      RECT 8.094 61.078 8.146 61.114 ;
      RECT 8.094 62.278 8.146 62.314 ;
      RECT 8.094 63.478 8.146 63.514 ;
      RECT 8.094 64.678 8.146 64.714 ;
      RECT 8.094 65.878 8.146 65.914 ;
      RECT 8.094 67.078 8.146 67.114 ;
      RECT 8.094 68.278 8.146 68.314 ;
      RECT 8.094 69.478 8.146 69.514 ;
      RECT 8.094 70.678 8.146 70.714 ;
      RECT 8.094 71.878 8.146 71.914 ;
      RECT 8.174 0.281 8.226 0.317 ;
      RECT 8.174 72.403 8.226 72.439 ;
      RECT 8.254 0.806 8.306 0.842 ;
      RECT 8.254 2.006 8.306 2.042 ;
      RECT 8.254 3.206 8.306 3.242 ;
      RECT 8.254 4.406 8.306 4.442 ;
      RECT 8.254 5.606 8.306 5.642 ;
      RECT 8.254 6.806 8.306 6.842 ;
      RECT 8.254 8.006 8.306 8.042 ;
      RECT 8.254 9.206 8.306 9.242 ;
      RECT 8.254 10.406 8.306 10.442 ;
      RECT 8.254 11.606 8.306 11.642 ;
      RECT 8.254 12.806 8.306 12.842 ;
      RECT 8.254 14.006 8.306 14.042 ;
      RECT 8.254 15.206 8.306 15.242 ;
      RECT 8.254 16.406 8.306 16.442 ;
      RECT 8.254 17.606 8.306 17.642 ;
      RECT 8.254 18.806 8.306 18.842 ;
      RECT 8.254 20.006 8.306 20.042 ;
      RECT 8.254 21.206 8.306 21.242 ;
      RECT 8.254 22.406 8.306 22.442 ;
      RECT 8.254 23.606 8.306 23.642 ;
      RECT 8.254 24.806 8.306 24.842 ;
      RECT 8.254 26.006 8.306 26.042 ;
      RECT 8.254 27.206 8.306 27.242 ;
      RECT 8.254 28.406 8.306 28.442 ;
      RECT 8.254 29.606 8.306 29.642 ;
      RECT 8.254 30.806 8.306 30.842 ;
      RECT 8.254 32.622 8.306 32.658 ;
      RECT 8.254 32.862 8.306 32.898 ;
      RECT 8.254 34.302 8.306 34.338 ;
      RECT 8.254 34.782 8.306 34.818 ;
      RECT 8.254 36.702 8.306 36.738 ;
      RECT 8.254 37.182 8.306 37.218 ;
      RECT 8.254 38.622 8.306 38.658 ;
      RECT 8.254 38.862 8.306 38.898 ;
      RECT 8.254 39.926 8.306 39.962 ;
      RECT 8.254 41.126 8.306 41.162 ;
      RECT 8.254 42.326 8.306 42.362 ;
      RECT 8.254 43.526 8.306 43.562 ;
      RECT 8.254 44.726 8.306 44.762 ;
      RECT 8.254 45.926 8.306 45.962 ;
      RECT 8.254 47.126 8.306 47.162 ;
      RECT 8.254 48.326 8.306 48.362 ;
      RECT 8.254 49.526 8.306 49.562 ;
      RECT 8.254 50.726 8.306 50.762 ;
      RECT 8.254 51.926 8.306 51.962 ;
      RECT 8.254 53.126 8.306 53.162 ;
      RECT 8.254 54.326 8.306 54.362 ;
      RECT 8.254 55.526 8.306 55.562 ;
      RECT 8.254 56.726 8.306 56.762 ;
      RECT 8.254 57.926 8.306 57.962 ;
      RECT 8.254 59.126 8.306 59.162 ;
      RECT 8.254 60.326 8.306 60.362 ;
      RECT 8.254 61.526 8.306 61.562 ;
      RECT 8.254 62.726 8.306 62.762 ;
      RECT 8.254 63.926 8.306 63.962 ;
      RECT 8.254 65.126 8.306 65.162 ;
      RECT 8.254 66.326 8.306 66.362 ;
      RECT 8.254 67.526 8.306 67.562 ;
      RECT 8.254 68.726 8.306 68.762 ;
      RECT 8.254 69.926 8.306 69.962 ;
      RECT 8.254 71.126 8.306 71.162 ;
      RECT 8.334 1.558 8.386 1.594 ;
      RECT 8.334 2.758 8.386 2.794 ;
      RECT 8.334 3.958 8.386 3.994 ;
      RECT 8.334 5.158 8.386 5.194 ;
      RECT 8.334 6.358 8.386 6.394 ;
      RECT 8.334 7.558 8.386 7.594 ;
      RECT 8.334 8.758 8.386 8.794 ;
      RECT 8.334 9.958 8.386 9.994 ;
      RECT 8.334 11.158 8.386 11.194 ;
      RECT 8.334 12.358 8.386 12.394 ;
      RECT 8.334 13.558 8.386 13.594 ;
      RECT 8.334 14.758 8.386 14.794 ;
      RECT 8.334 15.958 8.386 15.994 ;
      RECT 8.334 17.158 8.386 17.194 ;
      RECT 8.334 18.358 8.386 18.394 ;
      RECT 8.334 19.558 8.386 19.594 ;
      RECT 8.334 20.758 8.386 20.794 ;
      RECT 8.334 21.958 8.386 21.994 ;
      RECT 8.334 23.158 8.386 23.194 ;
      RECT 8.334 24.358 8.386 24.394 ;
      RECT 8.334 25.558 8.386 25.594 ;
      RECT 8.334 26.758 8.386 26.794 ;
      RECT 8.334 27.958 8.386 27.994 ;
      RECT 8.334 29.158 8.386 29.194 ;
      RECT 8.334 30.358 8.386 30.394 ;
      RECT 8.334 31.558 8.386 31.594 ;
      RECT 8.334 33.342 8.386 33.378 ;
      RECT 8.334 33.582 8.386 33.618 ;
      RECT 8.334 37.902 8.386 37.938 ;
      RECT 8.334 38.142 8.386 38.178 ;
      RECT 8.334 40.678 8.386 40.714 ;
      RECT 8.334 41.878 8.386 41.914 ;
      RECT 8.334 43.078 8.386 43.114 ;
      RECT 8.334 44.278 8.386 44.314 ;
      RECT 8.334 45.478 8.386 45.514 ;
      RECT 8.334 46.678 8.386 46.714 ;
      RECT 8.334 47.878 8.386 47.914 ;
      RECT 8.334 49.078 8.386 49.114 ;
      RECT 8.334 50.278 8.386 50.314 ;
      RECT 8.334 51.478 8.386 51.514 ;
      RECT 8.334 52.678 8.386 52.714 ;
      RECT 8.334 53.878 8.386 53.914 ;
      RECT 8.334 55.078 8.386 55.114 ;
      RECT 8.334 56.278 8.386 56.314 ;
      RECT 8.334 57.478 8.386 57.514 ;
      RECT 8.334 58.678 8.386 58.714 ;
      RECT 8.334 59.878 8.386 59.914 ;
      RECT 8.334 61.078 8.386 61.114 ;
      RECT 8.334 62.278 8.386 62.314 ;
      RECT 8.334 63.478 8.386 63.514 ;
      RECT 8.334 64.678 8.386 64.714 ;
      RECT 8.334 65.878 8.386 65.914 ;
      RECT 8.334 67.078 8.386 67.114 ;
      RECT 8.334 68.278 8.386 68.314 ;
      RECT 8.334 69.478 8.386 69.514 ;
      RECT 8.334 70.678 8.386 70.714 ;
      RECT 8.334 71.878 8.386 71.914 ;
      RECT 8.414 0.806 8.466 0.842 ;
      RECT 8.414 2.006 8.466 2.042 ;
      RECT 8.414 3.206 8.466 3.242 ;
      RECT 8.414 4.406 8.466 4.442 ;
      RECT 8.414 5.606 8.466 5.642 ;
      RECT 8.414 6.806 8.466 6.842 ;
      RECT 8.414 8.006 8.466 8.042 ;
      RECT 8.414 9.206 8.466 9.242 ;
      RECT 8.414 10.406 8.466 10.442 ;
      RECT 8.414 11.606 8.466 11.642 ;
      RECT 8.414 12.806 8.466 12.842 ;
      RECT 8.414 14.006 8.466 14.042 ;
      RECT 8.414 15.206 8.466 15.242 ;
      RECT 8.414 16.406 8.466 16.442 ;
      RECT 8.414 17.606 8.466 17.642 ;
      RECT 8.414 18.806 8.466 18.842 ;
      RECT 8.414 20.006 8.466 20.042 ;
      RECT 8.414 21.206 8.466 21.242 ;
      RECT 8.414 22.406 8.466 22.442 ;
      RECT 8.414 23.606 8.466 23.642 ;
      RECT 8.414 24.806 8.466 24.842 ;
      RECT 8.414 26.006 8.466 26.042 ;
      RECT 8.414 27.206 8.466 27.242 ;
      RECT 8.414 28.406 8.466 28.442 ;
      RECT 8.414 29.606 8.466 29.642 ;
      RECT 8.414 30.806 8.466 30.842 ;
      RECT 8.414 32.622 8.466 32.658 ;
      RECT 8.414 32.862 8.466 32.898 ;
      RECT 8.414 38.622 8.466 38.658 ;
      RECT 8.414 38.862 8.466 38.898 ;
      RECT 8.414 39.926 8.466 39.962 ;
      RECT 8.414 41.126 8.466 41.162 ;
      RECT 8.414 42.326 8.466 42.362 ;
      RECT 8.414 43.526 8.466 43.562 ;
      RECT 8.414 44.726 8.466 44.762 ;
      RECT 8.414 45.926 8.466 45.962 ;
      RECT 8.414 47.126 8.466 47.162 ;
      RECT 8.414 48.326 8.466 48.362 ;
      RECT 8.414 49.526 8.466 49.562 ;
      RECT 8.414 50.726 8.466 50.762 ;
      RECT 8.414 51.926 8.466 51.962 ;
      RECT 8.414 53.126 8.466 53.162 ;
      RECT 8.414 54.326 8.466 54.362 ;
      RECT 8.414 55.526 8.466 55.562 ;
      RECT 8.414 56.726 8.466 56.762 ;
      RECT 8.414 57.926 8.466 57.962 ;
      RECT 8.414 59.126 8.466 59.162 ;
      RECT 8.414 60.326 8.466 60.362 ;
      RECT 8.414 61.526 8.466 61.562 ;
      RECT 8.414 62.726 8.466 62.762 ;
      RECT 8.414 63.926 8.466 63.962 ;
      RECT 8.414 65.126 8.466 65.162 ;
      RECT 8.414 66.326 8.466 66.362 ;
      RECT 8.414 67.526 8.466 67.562 ;
      RECT 8.414 68.726 8.466 68.762 ;
      RECT 8.414 69.926 8.466 69.962 ;
      RECT 8.414 71.126 8.466 71.162 ;
      RECT 8.494 1.558 8.546 1.594 ;
      RECT 8.494 2.758 8.546 2.794 ;
      RECT 8.494 3.958 8.546 3.994 ;
      RECT 8.494 5.158 8.546 5.194 ;
      RECT 8.494 6.358 8.546 6.394 ;
      RECT 8.494 7.558 8.546 7.594 ;
      RECT 8.494 8.758 8.546 8.794 ;
      RECT 8.494 9.958 8.546 9.994 ;
      RECT 8.494 11.158 8.546 11.194 ;
      RECT 8.494 12.358 8.546 12.394 ;
      RECT 8.494 13.558 8.546 13.594 ;
      RECT 8.494 14.758 8.546 14.794 ;
      RECT 8.494 15.958 8.546 15.994 ;
      RECT 8.494 17.158 8.546 17.194 ;
      RECT 8.494 18.358 8.546 18.394 ;
      RECT 8.494 19.558 8.546 19.594 ;
      RECT 8.494 20.758 8.546 20.794 ;
      RECT 8.494 21.958 8.546 21.994 ;
      RECT 8.494 23.158 8.546 23.194 ;
      RECT 8.494 24.358 8.546 24.394 ;
      RECT 8.494 25.558 8.546 25.594 ;
      RECT 8.494 26.758 8.546 26.794 ;
      RECT 8.494 27.958 8.546 27.994 ;
      RECT 8.494 29.158 8.546 29.194 ;
      RECT 8.494 30.358 8.546 30.394 ;
      RECT 8.494 31.558 8.546 31.594 ;
      RECT 8.494 33.342 8.546 33.378 ;
      RECT 8.494 33.582 8.546 33.618 ;
      RECT 8.494 37.902 8.546 37.938 ;
      RECT 8.494 38.142 8.546 38.178 ;
      RECT 8.494 40.678 8.546 40.714 ;
      RECT 8.494 41.878 8.546 41.914 ;
      RECT 8.494 43.078 8.546 43.114 ;
      RECT 8.494 44.278 8.546 44.314 ;
      RECT 8.494 45.478 8.546 45.514 ;
      RECT 8.494 46.678 8.546 46.714 ;
      RECT 8.494 47.878 8.546 47.914 ;
      RECT 8.494 49.078 8.546 49.114 ;
      RECT 8.494 50.278 8.546 50.314 ;
      RECT 8.494 51.478 8.546 51.514 ;
      RECT 8.494 52.678 8.546 52.714 ;
      RECT 8.494 53.878 8.546 53.914 ;
      RECT 8.494 55.078 8.546 55.114 ;
      RECT 8.494 56.278 8.546 56.314 ;
      RECT 8.494 57.478 8.546 57.514 ;
      RECT 8.494 58.678 8.546 58.714 ;
      RECT 8.494 59.878 8.546 59.914 ;
      RECT 8.494 61.078 8.546 61.114 ;
      RECT 8.494 62.278 8.546 62.314 ;
      RECT 8.494 63.478 8.546 63.514 ;
      RECT 8.494 64.678 8.546 64.714 ;
      RECT 8.494 65.878 8.546 65.914 ;
      RECT 8.494 67.078 8.546 67.114 ;
      RECT 8.494 68.278 8.546 68.314 ;
      RECT 8.494 69.478 8.546 69.514 ;
      RECT 8.494 70.678 8.546 70.714 ;
      RECT 8.494 71.878 8.546 71.914 ;
      RECT 8.574 0.281 8.626 0.317 ;
      RECT 8.574 72.403 8.626 72.439 ;
      RECT 8.654 0.806 8.706 0.842 ;
      RECT 8.654 2.006 8.706 2.042 ;
      RECT 8.654 3.206 8.706 3.242 ;
      RECT 8.654 4.406 8.706 4.442 ;
      RECT 8.654 5.606 8.706 5.642 ;
      RECT 8.654 6.806 8.706 6.842 ;
      RECT 8.654 8.006 8.706 8.042 ;
      RECT 8.654 9.206 8.706 9.242 ;
      RECT 8.654 10.406 8.706 10.442 ;
      RECT 8.654 11.606 8.706 11.642 ;
      RECT 8.654 12.806 8.706 12.842 ;
      RECT 8.654 14.006 8.706 14.042 ;
      RECT 8.654 15.206 8.706 15.242 ;
      RECT 8.654 16.406 8.706 16.442 ;
      RECT 8.654 17.606 8.706 17.642 ;
      RECT 8.654 18.806 8.706 18.842 ;
      RECT 8.654 20.006 8.706 20.042 ;
      RECT 8.654 21.206 8.706 21.242 ;
      RECT 8.654 22.406 8.706 22.442 ;
      RECT 8.654 23.606 8.706 23.642 ;
      RECT 8.654 24.806 8.706 24.842 ;
      RECT 8.654 26.006 8.706 26.042 ;
      RECT 8.654 27.206 8.706 27.242 ;
      RECT 8.654 28.406 8.706 28.442 ;
      RECT 8.654 29.606 8.706 29.642 ;
      RECT 8.654 30.806 8.706 30.842 ;
      RECT 8.654 32.622 8.706 32.658 ;
      RECT 8.654 32.862 8.706 32.898 ;
      RECT 8.654 38.622 8.706 38.658 ;
      RECT 8.654 38.862 8.706 38.898 ;
      RECT 8.654 39.926 8.706 39.962 ;
      RECT 8.654 41.126 8.706 41.162 ;
      RECT 8.654 42.326 8.706 42.362 ;
      RECT 8.654 43.526 8.706 43.562 ;
      RECT 8.654 44.726 8.706 44.762 ;
      RECT 8.654 45.926 8.706 45.962 ;
      RECT 8.654 47.126 8.706 47.162 ;
      RECT 8.654 48.326 8.706 48.362 ;
      RECT 8.654 49.526 8.706 49.562 ;
      RECT 8.654 50.726 8.706 50.762 ;
      RECT 8.654 51.926 8.706 51.962 ;
      RECT 8.654 53.126 8.706 53.162 ;
      RECT 8.654 54.326 8.706 54.362 ;
      RECT 8.654 55.526 8.706 55.562 ;
      RECT 8.654 56.726 8.706 56.762 ;
      RECT 8.654 57.926 8.706 57.962 ;
      RECT 8.654 59.126 8.706 59.162 ;
      RECT 8.654 60.326 8.706 60.362 ;
      RECT 8.654 61.526 8.706 61.562 ;
      RECT 8.654 62.726 8.706 62.762 ;
      RECT 8.654 63.926 8.706 63.962 ;
      RECT 8.654 65.126 8.706 65.162 ;
      RECT 8.654 66.326 8.706 66.362 ;
      RECT 8.654 67.526 8.706 67.562 ;
      RECT 8.654 68.726 8.706 68.762 ;
      RECT 8.654 69.926 8.706 69.962 ;
      RECT 8.654 71.126 8.706 71.162 ;
      RECT 8.734 1.558 8.786 1.594 ;
      RECT 8.734 2.758 8.786 2.794 ;
      RECT 8.734 3.958 8.786 3.994 ;
      RECT 8.734 5.158 8.786 5.194 ;
      RECT 8.734 6.358 8.786 6.394 ;
      RECT 8.734 7.558 8.786 7.594 ;
      RECT 8.734 8.758 8.786 8.794 ;
      RECT 8.734 9.958 8.786 9.994 ;
      RECT 8.734 11.158 8.786 11.194 ;
      RECT 8.734 12.358 8.786 12.394 ;
      RECT 8.734 13.558 8.786 13.594 ;
      RECT 8.734 14.758 8.786 14.794 ;
      RECT 8.734 15.958 8.786 15.994 ;
      RECT 8.734 17.158 8.786 17.194 ;
      RECT 8.734 18.358 8.786 18.394 ;
      RECT 8.734 19.558 8.786 19.594 ;
      RECT 8.734 20.758 8.786 20.794 ;
      RECT 8.734 21.958 8.786 21.994 ;
      RECT 8.734 23.158 8.786 23.194 ;
      RECT 8.734 24.358 8.786 24.394 ;
      RECT 8.734 25.558 8.786 25.594 ;
      RECT 8.734 26.758 8.786 26.794 ;
      RECT 8.734 27.958 8.786 27.994 ;
      RECT 8.734 29.158 8.786 29.194 ;
      RECT 8.734 30.358 8.786 30.394 ;
      RECT 8.734 31.558 8.786 31.594 ;
      RECT 8.734 33.342 8.786 33.378 ;
      RECT 8.734 33.582 8.786 33.618 ;
      RECT 8.734 37.902 8.786 37.938 ;
      RECT 8.734 38.142 8.786 38.178 ;
      RECT 8.734 40.678 8.786 40.714 ;
      RECT 8.734 41.878 8.786 41.914 ;
      RECT 8.734 43.078 8.786 43.114 ;
      RECT 8.734 44.278 8.786 44.314 ;
      RECT 8.734 45.478 8.786 45.514 ;
      RECT 8.734 46.678 8.786 46.714 ;
      RECT 8.734 47.878 8.786 47.914 ;
      RECT 8.734 49.078 8.786 49.114 ;
      RECT 8.734 50.278 8.786 50.314 ;
      RECT 8.734 51.478 8.786 51.514 ;
      RECT 8.734 52.678 8.786 52.714 ;
      RECT 8.734 53.878 8.786 53.914 ;
      RECT 8.734 55.078 8.786 55.114 ;
      RECT 8.734 56.278 8.786 56.314 ;
      RECT 8.734 57.478 8.786 57.514 ;
      RECT 8.734 58.678 8.786 58.714 ;
      RECT 8.734 59.878 8.786 59.914 ;
      RECT 8.734 61.078 8.786 61.114 ;
      RECT 8.734 62.278 8.786 62.314 ;
      RECT 8.734 63.478 8.786 63.514 ;
      RECT 8.734 64.678 8.786 64.714 ;
      RECT 8.734 65.878 8.786 65.914 ;
      RECT 8.734 67.078 8.786 67.114 ;
      RECT 8.734 68.278 8.786 68.314 ;
      RECT 8.734 69.478 8.786 69.514 ;
      RECT 8.734 70.678 8.786 70.714 ;
      RECT 8.734 71.878 8.786 71.914 ;
      RECT 8.814 0.806 8.866 0.842 ;
      RECT 8.814 2.006 8.866 2.042 ;
      RECT 8.814 3.206 8.866 3.242 ;
      RECT 8.814 4.406 8.866 4.442 ;
      RECT 8.814 5.606 8.866 5.642 ;
      RECT 8.814 6.806 8.866 6.842 ;
      RECT 8.814 8.006 8.866 8.042 ;
      RECT 8.814 9.206 8.866 9.242 ;
      RECT 8.814 10.406 8.866 10.442 ;
      RECT 8.814 11.606 8.866 11.642 ;
      RECT 8.814 12.806 8.866 12.842 ;
      RECT 8.814 14.006 8.866 14.042 ;
      RECT 8.814 15.206 8.866 15.242 ;
      RECT 8.814 16.406 8.866 16.442 ;
      RECT 8.814 17.606 8.866 17.642 ;
      RECT 8.814 18.806 8.866 18.842 ;
      RECT 8.814 20.006 8.866 20.042 ;
      RECT 8.814 21.206 8.866 21.242 ;
      RECT 8.814 22.406 8.866 22.442 ;
      RECT 8.814 23.606 8.866 23.642 ;
      RECT 8.814 24.806 8.866 24.842 ;
      RECT 8.814 26.006 8.866 26.042 ;
      RECT 8.814 27.206 8.866 27.242 ;
      RECT 8.814 28.406 8.866 28.442 ;
      RECT 8.814 29.606 8.866 29.642 ;
      RECT 8.814 30.806 8.866 30.842 ;
      RECT 8.814 32.622 8.866 32.658 ;
      RECT 8.814 32.862 8.866 32.898 ;
      RECT 8.814 38.622 8.866 38.658 ;
      RECT 8.814 38.862 8.866 38.898 ;
      RECT 8.814 39.926 8.866 39.962 ;
      RECT 8.814 41.126 8.866 41.162 ;
      RECT 8.814 42.326 8.866 42.362 ;
      RECT 8.814 43.526 8.866 43.562 ;
      RECT 8.814 44.726 8.866 44.762 ;
      RECT 8.814 45.926 8.866 45.962 ;
      RECT 8.814 47.126 8.866 47.162 ;
      RECT 8.814 48.326 8.866 48.362 ;
      RECT 8.814 49.526 8.866 49.562 ;
      RECT 8.814 50.726 8.866 50.762 ;
      RECT 8.814 51.926 8.866 51.962 ;
      RECT 8.814 53.126 8.866 53.162 ;
      RECT 8.814 54.326 8.866 54.362 ;
      RECT 8.814 55.526 8.866 55.562 ;
      RECT 8.814 56.726 8.866 56.762 ;
      RECT 8.814 57.926 8.866 57.962 ;
      RECT 8.814 59.126 8.866 59.162 ;
      RECT 8.814 60.326 8.866 60.362 ;
      RECT 8.814 61.526 8.866 61.562 ;
      RECT 8.814 62.726 8.866 62.762 ;
      RECT 8.814 63.926 8.866 63.962 ;
      RECT 8.814 65.126 8.866 65.162 ;
      RECT 8.814 66.326 8.866 66.362 ;
      RECT 8.814 67.526 8.866 67.562 ;
      RECT 8.814 68.726 8.866 68.762 ;
      RECT 8.814 69.926 8.866 69.962 ;
      RECT 8.814 71.126 8.866 71.162 ;
      RECT 8.894 1.558 8.946 1.594 ;
      RECT 8.894 2.758 8.946 2.794 ;
      RECT 8.894 3.958 8.946 3.994 ;
      RECT 8.894 5.158 8.946 5.194 ;
      RECT 8.894 6.358 8.946 6.394 ;
      RECT 8.894 7.558 8.946 7.594 ;
      RECT 8.894 8.758 8.946 8.794 ;
      RECT 8.894 9.958 8.946 9.994 ;
      RECT 8.894 11.158 8.946 11.194 ;
      RECT 8.894 12.358 8.946 12.394 ;
      RECT 8.894 13.558 8.946 13.594 ;
      RECT 8.894 14.758 8.946 14.794 ;
      RECT 8.894 15.958 8.946 15.994 ;
      RECT 8.894 17.158 8.946 17.194 ;
      RECT 8.894 18.358 8.946 18.394 ;
      RECT 8.894 19.558 8.946 19.594 ;
      RECT 8.894 20.758 8.946 20.794 ;
      RECT 8.894 21.958 8.946 21.994 ;
      RECT 8.894 23.158 8.946 23.194 ;
      RECT 8.894 24.358 8.946 24.394 ;
      RECT 8.894 25.558 8.946 25.594 ;
      RECT 8.894 26.758 8.946 26.794 ;
      RECT 8.894 27.958 8.946 27.994 ;
      RECT 8.894 29.158 8.946 29.194 ;
      RECT 8.894 30.358 8.946 30.394 ;
      RECT 8.894 31.558 8.946 31.594 ;
      RECT 8.894 33.342 8.946 33.378 ;
      RECT 8.894 33.582 8.946 33.618 ;
      RECT 8.894 37.902 8.946 37.938 ;
      RECT 8.894 38.142 8.946 38.178 ;
      RECT 8.894 40.678 8.946 40.714 ;
      RECT 8.894 41.878 8.946 41.914 ;
      RECT 8.894 43.078 8.946 43.114 ;
      RECT 8.894 44.278 8.946 44.314 ;
      RECT 8.894 45.478 8.946 45.514 ;
      RECT 8.894 46.678 8.946 46.714 ;
      RECT 8.894 47.878 8.946 47.914 ;
      RECT 8.894 49.078 8.946 49.114 ;
      RECT 8.894 50.278 8.946 50.314 ;
      RECT 8.894 51.478 8.946 51.514 ;
      RECT 8.894 52.678 8.946 52.714 ;
      RECT 8.894 53.878 8.946 53.914 ;
      RECT 8.894 55.078 8.946 55.114 ;
      RECT 8.894 56.278 8.946 56.314 ;
      RECT 8.894 57.478 8.946 57.514 ;
      RECT 8.894 58.678 8.946 58.714 ;
      RECT 8.894 59.878 8.946 59.914 ;
      RECT 8.894 61.078 8.946 61.114 ;
      RECT 8.894 62.278 8.946 62.314 ;
      RECT 8.894 63.478 8.946 63.514 ;
      RECT 8.894 64.678 8.946 64.714 ;
      RECT 8.894 65.878 8.946 65.914 ;
      RECT 8.894 67.078 8.946 67.114 ;
      RECT 8.894 68.278 8.946 68.314 ;
      RECT 8.894 69.478 8.946 69.514 ;
      RECT 8.894 70.678 8.946 70.714 ;
      RECT 8.894 71.878 8.946 71.914 ;
      RECT 8.974 0.281 9.026 0.317 ;
      RECT 8.974 72.403 9.026 72.439 ;
      RECT 9.054 0.806 9.106 0.842 ;
      RECT 9.054 2.006 9.106 2.042 ;
      RECT 9.054 3.206 9.106 3.242 ;
      RECT 9.054 4.406 9.106 4.442 ;
      RECT 9.054 5.606 9.106 5.642 ;
      RECT 9.054 6.806 9.106 6.842 ;
      RECT 9.054 8.006 9.106 8.042 ;
      RECT 9.054 9.206 9.106 9.242 ;
      RECT 9.054 10.406 9.106 10.442 ;
      RECT 9.054 11.606 9.106 11.642 ;
      RECT 9.054 12.806 9.106 12.842 ;
      RECT 9.054 14.006 9.106 14.042 ;
      RECT 9.054 15.206 9.106 15.242 ;
      RECT 9.054 16.406 9.106 16.442 ;
      RECT 9.054 17.606 9.106 17.642 ;
      RECT 9.054 18.806 9.106 18.842 ;
      RECT 9.054 20.006 9.106 20.042 ;
      RECT 9.054 21.206 9.106 21.242 ;
      RECT 9.054 22.406 9.106 22.442 ;
      RECT 9.054 23.606 9.106 23.642 ;
      RECT 9.054 24.806 9.106 24.842 ;
      RECT 9.054 26.006 9.106 26.042 ;
      RECT 9.054 27.206 9.106 27.242 ;
      RECT 9.054 28.406 9.106 28.442 ;
      RECT 9.054 29.606 9.106 29.642 ;
      RECT 9.054 30.806 9.106 30.842 ;
      RECT 9.054 32.622 9.106 32.658 ;
      RECT 9.054 32.862 9.106 32.898 ;
      RECT 9.054 34.302 9.106 34.338 ;
      RECT 9.054 34.782 9.106 34.818 ;
      RECT 9.054 36.702 9.106 36.738 ;
      RECT 9.054 37.182 9.106 37.218 ;
      RECT 9.054 38.622 9.106 38.658 ;
      RECT 9.054 38.862 9.106 38.898 ;
      RECT 9.054 39.926 9.106 39.962 ;
      RECT 9.054 41.126 9.106 41.162 ;
      RECT 9.054 42.326 9.106 42.362 ;
      RECT 9.054 43.526 9.106 43.562 ;
      RECT 9.054 44.726 9.106 44.762 ;
      RECT 9.054 45.926 9.106 45.962 ;
      RECT 9.054 47.126 9.106 47.162 ;
      RECT 9.054 48.326 9.106 48.362 ;
      RECT 9.054 49.526 9.106 49.562 ;
      RECT 9.054 50.726 9.106 50.762 ;
      RECT 9.054 51.926 9.106 51.962 ;
      RECT 9.054 53.126 9.106 53.162 ;
      RECT 9.054 54.326 9.106 54.362 ;
      RECT 9.054 55.526 9.106 55.562 ;
      RECT 9.054 56.726 9.106 56.762 ;
      RECT 9.054 57.926 9.106 57.962 ;
      RECT 9.054 59.126 9.106 59.162 ;
      RECT 9.054 60.326 9.106 60.362 ;
      RECT 9.054 61.526 9.106 61.562 ;
      RECT 9.054 62.726 9.106 62.762 ;
      RECT 9.054 63.926 9.106 63.962 ;
      RECT 9.054 65.126 9.106 65.162 ;
      RECT 9.054 66.326 9.106 66.362 ;
      RECT 9.054 67.526 9.106 67.562 ;
      RECT 9.054 68.726 9.106 68.762 ;
      RECT 9.054 69.926 9.106 69.962 ;
      RECT 9.054 71.126 9.106 71.162 ;
      RECT 9.134 1.558 9.186 1.594 ;
      RECT 9.134 2.758 9.186 2.794 ;
      RECT 9.134 3.958 9.186 3.994 ;
      RECT 9.134 5.158 9.186 5.194 ;
      RECT 9.134 6.358 9.186 6.394 ;
      RECT 9.134 7.558 9.186 7.594 ;
      RECT 9.134 8.758 9.186 8.794 ;
      RECT 9.134 9.958 9.186 9.994 ;
      RECT 9.134 11.158 9.186 11.194 ;
      RECT 9.134 12.358 9.186 12.394 ;
      RECT 9.134 13.558 9.186 13.594 ;
      RECT 9.134 14.758 9.186 14.794 ;
      RECT 9.134 15.958 9.186 15.994 ;
      RECT 9.134 17.158 9.186 17.194 ;
      RECT 9.134 18.358 9.186 18.394 ;
      RECT 9.134 19.558 9.186 19.594 ;
      RECT 9.134 20.758 9.186 20.794 ;
      RECT 9.134 21.958 9.186 21.994 ;
      RECT 9.134 23.158 9.186 23.194 ;
      RECT 9.134 24.358 9.186 24.394 ;
      RECT 9.134 25.558 9.186 25.594 ;
      RECT 9.134 26.758 9.186 26.794 ;
      RECT 9.134 27.958 9.186 27.994 ;
      RECT 9.134 29.158 9.186 29.194 ;
      RECT 9.134 30.358 9.186 30.394 ;
      RECT 9.134 31.558 9.186 31.594 ;
      RECT 9.134 33.342 9.186 33.378 ;
      RECT 9.134 33.582 9.186 33.618 ;
      RECT 9.134 37.902 9.186 37.938 ;
      RECT 9.134 38.142 9.186 38.178 ;
      RECT 9.134 40.678 9.186 40.714 ;
      RECT 9.134 41.878 9.186 41.914 ;
      RECT 9.134 43.078 9.186 43.114 ;
      RECT 9.134 44.278 9.186 44.314 ;
      RECT 9.134 45.478 9.186 45.514 ;
      RECT 9.134 46.678 9.186 46.714 ;
      RECT 9.134 47.878 9.186 47.914 ;
      RECT 9.134 49.078 9.186 49.114 ;
      RECT 9.134 50.278 9.186 50.314 ;
      RECT 9.134 51.478 9.186 51.514 ;
      RECT 9.134 52.678 9.186 52.714 ;
      RECT 9.134 53.878 9.186 53.914 ;
      RECT 9.134 55.078 9.186 55.114 ;
      RECT 9.134 56.278 9.186 56.314 ;
      RECT 9.134 57.478 9.186 57.514 ;
      RECT 9.134 58.678 9.186 58.714 ;
      RECT 9.134 59.878 9.186 59.914 ;
      RECT 9.134 61.078 9.186 61.114 ;
      RECT 9.134 62.278 9.186 62.314 ;
      RECT 9.134 63.478 9.186 63.514 ;
      RECT 9.134 64.678 9.186 64.714 ;
      RECT 9.134 65.878 9.186 65.914 ;
      RECT 9.134 67.078 9.186 67.114 ;
      RECT 9.134 68.278 9.186 68.314 ;
      RECT 9.134 69.478 9.186 69.514 ;
      RECT 9.134 70.678 9.186 70.714 ;
      RECT 9.134 71.878 9.186 71.914 ;
      RECT 9.214 0.806 9.266 0.842 ;
      RECT 9.214 2.006 9.266 2.042 ;
      RECT 9.214 3.206 9.266 3.242 ;
      RECT 9.214 4.406 9.266 4.442 ;
      RECT 9.214 5.606 9.266 5.642 ;
      RECT 9.214 6.806 9.266 6.842 ;
      RECT 9.214 8.006 9.266 8.042 ;
      RECT 9.214 9.206 9.266 9.242 ;
      RECT 9.214 10.406 9.266 10.442 ;
      RECT 9.214 11.606 9.266 11.642 ;
      RECT 9.214 12.806 9.266 12.842 ;
      RECT 9.214 14.006 9.266 14.042 ;
      RECT 9.214 15.206 9.266 15.242 ;
      RECT 9.214 16.406 9.266 16.442 ;
      RECT 9.214 17.606 9.266 17.642 ;
      RECT 9.214 18.806 9.266 18.842 ;
      RECT 9.214 20.006 9.266 20.042 ;
      RECT 9.214 21.206 9.266 21.242 ;
      RECT 9.214 22.406 9.266 22.442 ;
      RECT 9.214 23.606 9.266 23.642 ;
      RECT 9.214 24.806 9.266 24.842 ;
      RECT 9.214 26.006 9.266 26.042 ;
      RECT 9.214 27.206 9.266 27.242 ;
      RECT 9.214 28.406 9.266 28.442 ;
      RECT 9.214 29.606 9.266 29.642 ;
      RECT 9.214 30.806 9.266 30.842 ;
      RECT 9.214 32.622 9.266 32.658 ;
      RECT 9.214 32.862 9.266 32.898 ;
      RECT 9.214 38.622 9.266 38.658 ;
      RECT 9.214 38.862 9.266 38.898 ;
      RECT 9.214 39.926 9.266 39.962 ;
      RECT 9.214 41.126 9.266 41.162 ;
      RECT 9.214 42.326 9.266 42.362 ;
      RECT 9.214 43.526 9.266 43.562 ;
      RECT 9.214 44.726 9.266 44.762 ;
      RECT 9.214 45.926 9.266 45.962 ;
      RECT 9.214 47.126 9.266 47.162 ;
      RECT 9.214 48.326 9.266 48.362 ;
      RECT 9.214 49.526 9.266 49.562 ;
      RECT 9.214 50.726 9.266 50.762 ;
      RECT 9.214 51.926 9.266 51.962 ;
      RECT 9.214 53.126 9.266 53.162 ;
      RECT 9.214 54.326 9.266 54.362 ;
      RECT 9.214 55.526 9.266 55.562 ;
      RECT 9.214 56.726 9.266 56.762 ;
      RECT 9.214 57.926 9.266 57.962 ;
      RECT 9.214 59.126 9.266 59.162 ;
      RECT 9.214 60.326 9.266 60.362 ;
      RECT 9.214 61.526 9.266 61.562 ;
      RECT 9.214 62.726 9.266 62.762 ;
      RECT 9.214 63.926 9.266 63.962 ;
      RECT 9.214 65.126 9.266 65.162 ;
      RECT 9.214 66.326 9.266 66.362 ;
      RECT 9.214 67.526 9.266 67.562 ;
      RECT 9.214 68.726 9.266 68.762 ;
      RECT 9.214 69.926 9.266 69.962 ;
      RECT 9.214 71.126 9.266 71.162 ;
      RECT 9.294 1.558 9.346 1.594 ;
      RECT 9.294 2.758 9.346 2.794 ;
      RECT 9.294 3.958 9.346 3.994 ;
      RECT 9.294 5.158 9.346 5.194 ;
      RECT 9.294 6.358 9.346 6.394 ;
      RECT 9.294 7.558 9.346 7.594 ;
      RECT 9.294 8.758 9.346 8.794 ;
      RECT 9.294 9.958 9.346 9.994 ;
      RECT 9.294 11.158 9.346 11.194 ;
      RECT 9.294 12.358 9.346 12.394 ;
      RECT 9.294 13.558 9.346 13.594 ;
      RECT 9.294 14.758 9.346 14.794 ;
      RECT 9.294 15.958 9.346 15.994 ;
      RECT 9.294 17.158 9.346 17.194 ;
      RECT 9.294 18.358 9.346 18.394 ;
      RECT 9.294 19.558 9.346 19.594 ;
      RECT 9.294 20.758 9.346 20.794 ;
      RECT 9.294 21.958 9.346 21.994 ;
      RECT 9.294 23.158 9.346 23.194 ;
      RECT 9.294 24.358 9.346 24.394 ;
      RECT 9.294 25.558 9.346 25.594 ;
      RECT 9.294 26.758 9.346 26.794 ;
      RECT 9.294 27.958 9.346 27.994 ;
      RECT 9.294 29.158 9.346 29.194 ;
      RECT 9.294 30.358 9.346 30.394 ;
      RECT 9.294 31.558 9.346 31.594 ;
      RECT 9.294 33.342 9.346 33.378 ;
      RECT 9.294 33.582 9.346 33.618 ;
      RECT 9.294 37.902 9.346 37.938 ;
      RECT 9.294 38.142 9.346 38.178 ;
      RECT 9.294 40.678 9.346 40.714 ;
      RECT 9.294 41.878 9.346 41.914 ;
      RECT 9.294 43.078 9.346 43.114 ;
      RECT 9.294 44.278 9.346 44.314 ;
      RECT 9.294 45.478 9.346 45.514 ;
      RECT 9.294 46.678 9.346 46.714 ;
      RECT 9.294 47.878 9.346 47.914 ;
      RECT 9.294 49.078 9.346 49.114 ;
      RECT 9.294 50.278 9.346 50.314 ;
      RECT 9.294 51.478 9.346 51.514 ;
      RECT 9.294 52.678 9.346 52.714 ;
      RECT 9.294 53.878 9.346 53.914 ;
      RECT 9.294 55.078 9.346 55.114 ;
      RECT 9.294 56.278 9.346 56.314 ;
      RECT 9.294 57.478 9.346 57.514 ;
      RECT 9.294 58.678 9.346 58.714 ;
      RECT 9.294 59.878 9.346 59.914 ;
      RECT 9.294 61.078 9.346 61.114 ;
      RECT 9.294 62.278 9.346 62.314 ;
      RECT 9.294 63.478 9.346 63.514 ;
      RECT 9.294 64.678 9.346 64.714 ;
      RECT 9.294 65.878 9.346 65.914 ;
      RECT 9.294 67.078 9.346 67.114 ;
      RECT 9.294 68.278 9.346 68.314 ;
      RECT 9.294 69.478 9.346 69.514 ;
      RECT 9.294 70.678 9.346 70.714 ;
      RECT 9.294 71.878 9.346 71.914 ;
      RECT 9.374 0.281 9.426 0.317 ;
      RECT 9.374 72.403 9.426 72.439 ;
      RECT 9.454 0.806 9.506 0.842 ;
      RECT 9.454 2.006 9.506 2.042 ;
      RECT 9.454 3.206 9.506 3.242 ;
      RECT 9.454 4.406 9.506 4.442 ;
      RECT 9.454 5.606 9.506 5.642 ;
      RECT 9.454 6.806 9.506 6.842 ;
      RECT 9.454 8.006 9.506 8.042 ;
      RECT 9.454 9.206 9.506 9.242 ;
      RECT 9.454 10.406 9.506 10.442 ;
      RECT 9.454 11.606 9.506 11.642 ;
      RECT 9.454 12.806 9.506 12.842 ;
      RECT 9.454 14.006 9.506 14.042 ;
      RECT 9.454 15.206 9.506 15.242 ;
      RECT 9.454 16.406 9.506 16.442 ;
      RECT 9.454 17.606 9.506 17.642 ;
      RECT 9.454 18.806 9.506 18.842 ;
      RECT 9.454 20.006 9.506 20.042 ;
      RECT 9.454 21.206 9.506 21.242 ;
      RECT 9.454 22.406 9.506 22.442 ;
      RECT 9.454 23.606 9.506 23.642 ;
      RECT 9.454 24.806 9.506 24.842 ;
      RECT 9.454 26.006 9.506 26.042 ;
      RECT 9.454 27.206 9.506 27.242 ;
      RECT 9.454 28.406 9.506 28.442 ;
      RECT 9.454 29.606 9.506 29.642 ;
      RECT 9.454 30.806 9.506 30.842 ;
      RECT 9.454 32.622 9.506 32.658 ;
      RECT 9.454 32.862 9.506 32.898 ;
      RECT 9.454 38.622 9.506 38.658 ;
      RECT 9.454 38.862 9.506 38.898 ;
      RECT 9.454 39.926 9.506 39.962 ;
      RECT 9.454 41.126 9.506 41.162 ;
      RECT 9.454 42.326 9.506 42.362 ;
      RECT 9.454 43.526 9.506 43.562 ;
      RECT 9.454 44.726 9.506 44.762 ;
      RECT 9.454 45.926 9.506 45.962 ;
      RECT 9.454 47.126 9.506 47.162 ;
      RECT 9.454 48.326 9.506 48.362 ;
      RECT 9.454 49.526 9.506 49.562 ;
      RECT 9.454 50.726 9.506 50.762 ;
      RECT 9.454 51.926 9.506 51.962 ;
      RECT 9.454 53.126 9.506 53.162 ;
      RECT 9.454 54.326 9.506 54.362 ;
      RECT 9.454 55.526 9.506 55.562 ;
      RECT 9.454 56.726 9.506 56.762 ;
      RECT 9.454 57.926 9.506 57.962 ;
      RECT 9.454 59.126 9.506 59.162 ;
      RECT 9.454 60.326 9.506 60.362 ;
      RECT 9.454 61.526 9.506 61.562 ;
      RECT 9.454 62.726 9.506 62.762 ;
      RECT 9.454 63.926 9.506 63.962 ;
      RECT 9.454 65.126 9.506 65.162 ;
      RECT 9.454 66.326 9.506 66.362 ;
      RECT 9.454 67.526 9.506 67.562 ;
      RECT 9.454 68.726 9.506 68.762 ;
      RECT 9.454 69.926 9.506 69.962 ;
      RECT 9.454 71.126 9.506 71.162 ;
      RECT 9.534 1.558 9.586 1.594 ;
      RECT 9.534 2.758 9.586 2.794 ;
      RECT 9.534 3.958 9.586 3.994 ;
      RECT 9.534 5.158 9.586 5.194 ;
      RECT 9.534 6.358 9.586 6.394 ;
      RECT 9.534 7.558 9.586 7.594 ;
      RECT 9.534 8.758 9.586 8.794 ;
      RECT 9.534 9.958 9.586 9.994 ;
      RECT 9.534 11.158 9.586 11.194 ;
      RECT 9.534 12.358 9.586 12.394 ;
      RECT 9.534 13.558 9.586 13.594 ;
      RECT 9.534 14.758 9.586 14.794 ;
      RECT 9.534 15.958 9.586 15.994 ;
      RECT 9.534 17.158 9.586 17.194 ;
      RECT 9.534 18.358 9.586 18.394 ;
      RECT 9.534 19.558 9.586 19.594 ;
      RECT 9.534 20.758 9.586 20.794 ;
      RECT 9.534 21.958 9.586 21.994 ;
      RECT 9.534 23.158 9.586 23.194 ;
      RECT 9.534 24.358 9.586 24.394 ;
      RECT 9.534 25.558 9.586 25.594 ;
      RECT 9.534 26.758 9.586 26.794 ;
      RECT 9.534 27.958 9.586 27.994 ;
      RECT 9.534 29.158 9.586 29.194 ;
      RECT 9.534 30.358 9.586 30.394 ;
      RECT 9.534 31.558 9.586 31.594 ;
      RECT 9.534 33.342 9.586 33.378 ;
      RECT 9.534 33.582 9.586 33.618 ;
      RECT 9.534 37.902 9.586 37.938 ;
      RECT 9.534 38.142 9.586 38.178 ;
      RECT 9.534 40.678 9.586 40.714 ;
      RECT 9.534 41.878 9.586 41.914 ;
      RECT 9.534 43.078 9.586 43.114 ;
      RECT 9.534 44.278 9.586 44.314 ;
      RECT 9.534 45.478 9.586 45.514 ;
      RECT 9.534 46.678 9.586 46.714 ;
      RECT 9.534 47.878 9.586 47.914 ;
      RECT 9.534 49.078 9.586 49.114 ;
      RECT 9.534 50.278 9.586 50.314 ;
      RECT 9.534 51.478 9.586 51.514 ;
      RECT 9.534 52.678 9.586 52.714 ;
      RECT 9.534 53.878 9.586 53.914 ;
      RECT 9.534 55.078 9.586 55.114 ;
      RECT 9.534 56.278 9.586 56.314 ;
      RECT 9.534 57.478 9.586 57.514 ;
      RECT 9.534 58.678 9.586 58.714 ;
      RECT 9.534 59.878 9.586 59.914 ;
      RECT 9.534 61.078 9.586 61.114 ;
      RECT 9.534 62.278 9.586 62.314 ;
      RECT 9.534 63.478 9.586 63.514 ;
      RECT 9.534 64.678 9.586 64.714 ;
      RECT 9.534 65.878 9.586 65.914 ;
      RECT 9.534 67.078 9.586 67.114 ;
      RECT 9.534 68.278 9.586 68.314 ;
      RECT 9.534 69.478 9.586 69.514 ;
      RECT 9.534 70.678 9.586 70.714 ;
      RECT 9.534 71.878 9.586 71.914 ;
      RECT 9.614 0.806 9.666 0.842 ;
      RECT 9.614 2.006 9.666 2.042 ;
      RECT 9.614 3.206 9.666 3.242 ;
      RECT 9.614 4.406 9.666 4.442 ;
      RECT 9.614 5.606 9.666 5.642 ;
      RECT 9.614 6.806 9.666 6.842 ;
      RECT 9.614 8.006 9.666 8.042 ;
      RECT 9.614 9.206 9.666 9.242 ;
      RECT 9.614 10.406 9.666 10.442 ;
      RECT 9.614 11.606 9.666 11.642 ;
      RECT 9.614 12.806 9.666 12.842 ;
      RECT 9.614 14.006 9.666 14.042 ;
      RECT 9.614 15.206 9.666 15.242 ;
      RECT 9.614 16.406 9.666 16.442 ;
      RECT 9.614 17.606 9.666 17.642 ;
      RECT 9.614 18.806 9.666 18.842 ;
      RECT 9.614 20.006 9.666 20.042 ;
      RECT 9.614 21.206 9.666 21.242 ;
      RECT 9.614 22.406 9.666 22.442 ;
      RECT 9.614 23.606 9.666 23.642 ;
      RECT 9.614 24.806 9.666 24.842 ;
      RECT 9.614 26.006 9.666 26.042 ;
      RECT 9.614 27.206 9.666 27.242 ;
      RECT 9.614 28.406 9.666 28.442 ;
      RECT 9.614 29.606 9.666 29.642 ;
      RECT 9.614 30.806 9.666 30.842 ;
      RECT 9.614 32.622 9.666 32.658 ;
      RECT 9.614 32.862 9.666 32.898 ;
      RECT 9.614 38.622 9.666 38.658 ;
      RECT 9.614 38.862 9.666 38.898 ;
      RECT 9.614 39.926 9.666 39.962 ;
      RECT 9.614 41.126 9.666 41.162 ;
      RECT 9.614 42.326 9.666 42.362 ;
      RECT 9.614 43.526 9.666 43.562 ;
      RECT 9.614 44.726 9.666 44.762 ;
      RECT 9.614 45.926 9.666 45.962 ;
      RECT 9.614 47.126 9.666 47.162 ;
      RECT 9.614 48.326 9.666 48.362 ;
      RECT 9.614 49.526 9.666 49.562 ;
      RECT 9.614 50.726 9.666 50.762 ;
      RECT 9.614 51.926 9.666 51.962 ;
      RECT 9.614 53.126 9.666 53.162 ;
      RECT 9.614 54.326 9.666 54.362 ;
      RECT 9.614 55.526 9.666 55.562 ;
      RECT 9.614 56.726 9.666 56.762 ;
      RECT 9.614 57.926 9.666 57.962 ;
      RECT 9.614 59.126 9.666 59.162 ;
      RECT 9.614 60.326 9.666 60.362 ;
      RECT 9.614 61.526 9.666 61.562 ;
      RECT 9.614 62.726 9.666 62.762 ;
      RECT 9.614 63.926 9.666 63.962 ;
      RECT 9.614 65.126 9.666 65.162 ;
      RECT 9.614 66.326 9.666 66.362 ;
      RECT 9.614 67.526 9.666 67.562 ;
      RECT 9.614 68.726 9.666 68.762 ;
      RECT 9.614 69.926 9.666 69.962 ;
      RECT 9.614 71.126 9.666 71.162 ;
      RECT 9.694 1.558 9.746 1.594 ;
      RECT 9.694 2.758 9.746 2.794 ;
      RECT 9.694 3.958 9.746 3.994 ;
      RECT 9.694 5.158 9.746 5.194 ;
      RECT 9.694 6.358 9.746 6.394 ;
      RECT 9.694 7.558 9.746 7.594 ;
      RECT 9.694 8.758 9.746 8.794 ;
      RECT 9.694 9.958 9.746 9.994 ;
      RECT 9.694 11.158 9.746 11.194 ;
      RECT 9.694 12.358 9.746 12.394 ;
      RECT 9.694 13.558 9.746 13.594 ;
      RECT 9.694 14.758 9.746 14.794 ;
      RECT 9.694 15.958 9.746 15.994 ;
      RECT 9.694 17.158 9.746 17.194 ;
      RECT 9.694 18.358 9.746 18.394 ;
      RECT 9.694 19.558 9.746 19.594 ;
      RECT 9.694 20.758 9.746 20.794 ;
      RECT 9.694 21.958 9.746 21.994 ;
      RECT 9.694 23.158 9.746 23.194 ;
      RECT 9.694 24.358 9.746 24.394 ;
      RECT 9.694 25.558 9.746 25.594 ;
      RECT 9.694 26.758 9.746 26.794 ;
      RECT 9.694 27.958 9.746 27.994 ;
      RECT 9.694 29.158 9.746 29.194 ;
      RECT 9.694 30.358 9.746 30.394 ;
      RECT 9.694 31.558 9.746 31.594 ;
      RECT 9.694 33.342 9.746 33.378 ;
      RECT 9.694 33.582 9.746 33.618 ;
      RECT 9.694 37.902 9.746 37.938 ;
      RECT 9.694 38.142 9.746 38.178 ;
      RECT 9.694 40.678 9.746 40.714 ;
      RECT 9.694 41.878 9.746 41.914 ;
      RECT 9.694 43.078 9.746 43.114 ;
      RECT 9.694 44.278 9.746 44.314 ;
      RECT 9.694 45.478 9.746 45.514 ;
      RECT 9.694 46.678 9.746 46.714 ;
      RECT 9.694 47.878 9.746 47.914 ;
      RECT 9.694 49.078 9.746 49.114 ;
      RECT 9.694 50.278 9.746 50.314 ;
      RECT 9.694 51.478 9.746 51.514 ;
      RECT 9.694 52.678 9.746 52.714 ;
      RECT 9.694 53.878 9.746 53.914 ;
      RECT 9.694 55.078 9.746 55.114 ;
      RECT 9.694 56.278 9.746 56.314 ;
      RECT 9.694 57.478 9.746 57.514 ;
      RECT 9.694 58.678 9.746 58.714 ;
      RECT 9.694 59.878 9.746 59.914 ;
      RECT 9.694 61.078 9.746 61.114 ;
      RECT 9.694 62.278 9.746 62.314 ;
      RECT 9.694 63.478 9.746 63.514 ;
      RECT 9.694 64.678 9.746 64.714 ;
      RECT 9.694 65.878 9.746 65.914 ;
      RECT 9.694 67.078 9.746 67.114 ;
      RECT 9.694 68.278 9.746 68.314 ;
      RECT 9.694 69.478 9.746 69.514 ;
      RECT 9.694 70.678 9.746 70.714 ;
      RECT 9.694 71.878 9.746 71.914 ;
      RECT 9.774 0.281 9.826 0.317 ;
      RECT 9.774 72.403 9.826 72.439 ;
      RECT 9.854 0.806 9.906 0.842 ;
      RECT 9.854 2.006 9.906 2.042 ;
      RECT 9.854 3.206 9.906 3.242 ;
      RECT 9.854 4.406 9.906 4.442 ;
      RECT 9.854 5.606 9.906 5.642 ;
      RECT 9.854 6.806 9.906 6.842 ;
      RECT 9.854 8.006 9.906 8.042 ;
      RECT 9.854 9.206 9.906 9.242 ;
      RECT 9.854 10.406 9.906 10.442 ;
      RECT 9.854 11.606 9.906 11.642 ;
      RECT 9.854 12.806 9.906 12.842 ;
      RECT 9.854 14.006 9.906 14.042 ;
      RECT 9.854 15.206 9.906 15.242 ;
      RECT 9.854 16.406 9.906 16.442 ;
      RECT 9.854 17.606 9.906 17.642 ;
      RECT 9.854 18.806 9.906 18.842 ;
      RECT 9.854 20.006 9.906 20.042 ;
      RECT 9.854 21.206 9.906 21.242 ;
      RECT 9.854 22.406 9.906 22.442 ;
      RECT 9.854 23.606 9.906 23.642 ;
      RECT 9.854 24.806 9.906 24.842 ;
      RECT 9.854 26.006 9.906 26.042 ;
      RECT 9.854 27.206 9.906 27.242 ;
      RECT 9.854 28.406 9.906 28.442 ;
      RECT 9.854 29.606 9.906 29.642 ;
      RECT 9.854 30.806 9.906 30.842 ;
      RECT 9.854 32.622 9.906 32.658 ;
      RECT 9.854 32.862 9.906 32.898 ;
      RECT 9.854 34.302 9.906 34.338 ;
      RECT 9.854 34.782 9.906 34.818 ;
      RECT 9.854 36.702 9.906 36.738 ;
      RECT 9.854 37.182 9.906 37.218 ;
      RECT 9.854 38.622 9.906 38.658 ;
      RECT 9.854 38.862 9.906 38.898 ;
      RECT 9.854 39.926 9.906 39.962 ;
      RECT 9.854 41.126 9.906 41.162 ;
      RECT 9.854 42.326 9.906 42.362 ;
      RECT 9.854 43.526 9.906 43.562 ;
      RECT 9.854 44.726 9.906 44.762 ;
      RECT 9.854 45.926 9.906 45.962 ;
      RECT 9.854 47.126 9.906 47.162 ;
      RECT 9.854 48.326 9.906 48.362 ;
      RECT 9.854 49.526 9.906 49.562 ;
      RECT 9.854 50.726 9.906 50.762 ;
      RECT 9.854 51.926 9.906 51.962 ;
      RECT 9.854 53.126 9.906 53.162 ;
      RECT 9.854 54.326 9.906 54.362 ;
      RECT 9.854 55.526 9.906 55.562 ;
      RECT 9.854 56.726 9.906 56.762 ;
      RECT 9.854 57.926 9.906 57.962 ;
      RECT 9.854 59.126 9.906 59.162 ;
      RECT 9.854 60.326 9.906 60.362 ;
      RECT 9.854 61.526 9.906 61.562 ;
      RECT 9.854 62.726 9.906 62.762 ;
      RECT 9.854 63.926 9.906 63.962 ;
      RECT 9.854 65.126 9.906 65.162 ;
      RECT 9.854 66.326 9.906 66.362 ;
      RECT 9.854 67.526 9.906 67.562 ;
      RECT 9.854 68.726 9.906 68.762 ;
      RECT 9.854 69.926 9.906 69.962 ;
      RECT 9.854 71.126 9.906 71.162 ;
      RECT 9.934 1.558 9.986 1.594 ;
      RECT 9.934 2.758 9.986 2.794 ;
      RECT 9.934 3.958 9.986 3.994 ;
      RECT 9.934 5.158 9.986 5.194 ;
      RECT 9.934 6.358 9.986 6.394 ;
      RECT 9.934 7.558 9.986 7.594 ;
      RECT 9.934 8.758 9.986 8.794 ;
      RECT 9.934 9.958 9.986 9.994 ;
      RECT 9.934 11.158 9.986 11.194 ;
      RECT 9.934 12.358 9.986 12.394 ;
      RECT 9.934 13.558 9.986 13.594 ;
      RECT 9.934 14.758 9.986 14.794 ;
      RECT 9.934 15.958 9.986 15.994 ;
      RECT 9.934 17.158 9.986 17.194 ;
      RECT 9.934 18.358 9.986 18.394 ;
      RECT 9.934 19.558 9.986 19.594 ;
      RECT 9.934 20.758 9.986 20.794 ;
      RECT 9.934 21.958 9.986 21.994 ;
      RECT 9.934 23.158 9.986 23.194 ;
      RECT 9.934 24.358 9.986 24.394 ;
      RECT 9.934 25.558 9.986 25.594 ;
      RECT 9.934 26.758 9.986 26.794 ;
      RECT 9.934 27.958 9.986 27.994 ;
      RECT 9.934 29.158 9.986 29.194 ;
      RECT 9.934 30.358 9.986 30.394 ;
      RECT 9.934 31.558 9.986 31.594 ;
      RECT 9.934 33.342 9.986 33.378 ;
      RECT 9.934 33.582 9.986 33.618 ;
      RECT 9.934 37.902 9.986 37.938 ;
      RECT 9.934 38.142 9.986 38.178 ;
      RECT 9.934 40.678 9.986 40.714 ;
      RECT 9.934 41.878 9.986 41.914 ;
      RECT 9.934 43.078 9.986 43.114 ;
      RECT 9.934 44.278 9.986 44.314 ;
      RECT 9.934 45.478 9.986 45.514 ;
      RECT 9.934 46.678 9.986 46.714 ;
      RECT 9.934 47.878 9.986 47.914 ;
      RECT 9.934 49.078 9.986 49.114 ;
      RECT 9.934 50.278 9.986 50.314 ;
      RECT 9.934 51.478 9.986 51.514 ;
      RECT 9.934 52.678 9.986 52.714 ;
      RECT 9.934 53.878 9.986 53.914 ;
      RECT 9.934 55.078 9.986 55.114 ;
      RECT 9.934 56.278 9.986 56.314 ;
      RECT 9.934 57.478 9.986 57.514 ;
      RECT 9.934 58.678 9.986 58.714 ;
      RECT 9.934 59.878 9.986 59.914 ;
      RECT 9.934 61.078 9.986 61.114 ;
      RECT 9.934 62.278 9.986 62.314 ;
      RECT 9.934 63.478 9.986 63.514 ;
      RECT 9.934 64.678 9.986 64.714 ;
      RECT 9.934 65.878 9.986 65.914 ;
      RECT 9.934 67.078 9.986 67.114 ;
      RECT 9.934 68.278 9.986 68.314 ;
      RECT 9.934 69.478 9.986 69.514 ;
      RECT 9.934 70.678 9.986 70.714 ;
      RECT 9.934 71.878 9.986 71.914 ;
      RECT 10.014 0.806 10.066 0.842 ;
      RECT 10.014 2.006 10.066 2.042 ;
      RECT 10.014 3.206 10.066 3.242 ;
      RECT 10.014 4.406 10.066 4.442 ;
      RECT 10.014 5.606 10.066 5.642 ;
      RECT 10.014 6.806 10.066 6.842 ;
      RECT 10.014 8.006 10.066 8.042 ;
      RECT 10.014 9.206 10.066 9.242 ;
      RECT 10.014 10.406 10.066 10.442 ;
      RECT 10.014 11.606 10.066 11.642 ;
      RECT 10.014 12.806 10.066 12.842 ;
      RECT 10.014 14.006 10.066 14.042 ;
      RECT 10.014 15.206 10.066 15.242 ;
      RECT 10.014 16.406 10.066 16.442 ;
      RECT 10.014 17.606 10.066 17.642 ;
      RECT 10.014 18.806 10.066 18.842 ;
      RECT 10.014 20.006 10.066 20.042 ;
      RECT 10.014 21.206 10.066 21.242 ;
      RECT 10.014 22.406 10.066 22.442 ;
      RECT 10.014 23.606 10.066 23.642 ;
      RECT 10.014 24.806 10.066 24.842 ;
      RECT 10.014 26.006 10.066 26.042 ;
      RECT 10.014 27.206 10.066 27.242 ;
      RECT 10.014 28.406 10.066 28.442 ;
      RECT 10.014 29.606 10.066 29.642 ;
      RECT 10.014 30.806 10.066 30.842 ;
      RECT 10.014 32.622 10.066 32.658 ;
      RECT 10.014 32.862 10.066 32.898 ;
      RECT 10.014 38.622 10.066 38.658 ;
      RECT 10.014 38.862 10.066 38.898 ;
      RECT 10.014 39.926 10.066 39.962 ;
      RECT 10.014 41.126 10.066 41.162 ;
      RECT 10.014 42.326 10.066 42.362 ;
      RECT 10.014 43.526 10.066 43.562 ;
      RECT 10.014 44.726 10.066 44.762 ;
      RECT 10.014 45.926 10.066 45.962 ;
      RECT 10.014 47.126 10.066 47.162 ;
      RECT 10.014 48.326 10.066 48.362 ;
      RECT 10.014 49.526 10.066 49.562 ;
      RECT 10.014 50.726 10.066 50.762 ;
      RECT 10.014 51.926 10.066 51.962 ;
      RECT 10.014 53.126 10.066 53.162 ;
      RECT 10.014 54.326 10.066 54.362 ;
      RECT 10.014 55.526 10.066 55.562 ;
      RECT 10.014 56.726 10.066 56.762 ;
      RECT 10.014 57.926 10.066 57.962 ;
      RECT 10.014 59.126 10.066 59.162 ;
      RECT 10.014 60.326 10.066 60.362 ;
      RECT 10.014 61.526 10.066 61.562 ;
      RECT 10.014 62.726 10.066 62.762 ;
      RECT 10.014 63.926 10.066 63.962 ;
      RECT 10.014 65.126 10.066 65.162 ;
      RECT 10.014 66.326 10.066 66.362 ;
      RECT 10.014 67.526 10.066 67.562 ;
      RECT 10.014 68.726 10.066 68.762 ;
      RECT 10.014 69.926 10.066 69.962 ;
      RECT 10.014 71.126 10.066 71.162 ;
      RECT 10.094 1.558 10.146 1.594 ;
      RECT 10.094 2.758 10.146 2.794 ;
      RECT 10.094 3.958 10.146 3.994 ;
      RECT 10.094 5.158 10.146 5.194 ;
      RECT 10.094 6.358 10.146 6.394 ;
      RECT 10.094 7.558 10.146 7.594 ;
      RECT 10.094 8.758 10.146 8.794 ;
      RECT 10.094 9.958 10.146 9.994 ;
      RECT 10.094 11.158 10.146 11.194 ;
      RECT 10.094 12.358 10.146 12.394 ;
      RECT 10.094 13.558 10.146 13.594 ;
      RECT 10.094 14.758 10.146 14.794 ;
      RECT 10.094 15.958 10.146 15.994 ;
      RECT 10.094 17.158 10.146 17.194 ;
      RECT 10.094 18.358 10.146 18.394 ;
      RECT 10.094 19.558 10.146 19.594 ;
      RECT 10.094 20.758 10.146 20.794 ;
      RECT 10.094 21.958 10.146 21.994 ;
      RECT 10.094 23.158 10.146 23.194 ;
      RECT 10.094 24.358 10.146 24.394 ;
      RECT 10.094 25.558 10.146 25.594 ;
      RECT 10.094 26.758 10.146 26.794 ;
      RECT 10.094 27.958 10.146 27.994 ;
      RECT 10.094 29.158 10.146 29.194 ;
      RECT 10.094 30.358 10.146 30.394 ;
      RECT 10.094 31.558 10.146 31.594 ;
      RECT 10.094 33.342 10.146 33.378 ;
      RECT 10.094 33.582 10.146 33.618 ;
      RECT 10.094 37.902 10.146 37.938 ;
      RECT 10.094 38.142 10.146 38.178 ;
      RECT 10.094 40.678 10.146 40.714 ;
      RECT 10.094 41.878 10.146 41.914 ;
      RECT 10.094 43.078 10.146 43.114 ;
      RECT 10.094 44.278 10.146 44.314 ;
      RECT 10.094 45.478 10.146 45.514 ;
      RECT 10.094 46.678 10.146 46.714 ;
      RECT 10.094 47.878 10.146 47.914 ;
      RECT 10.094 49.078 10.146 49.114 ;
      RECT 10.094 50.278 10.146 50.314 ;
      RECT 10.094 51.478 10.146 51.514 ;
      RECT 10.094 52.678 10.146 52.714 ;
      RECT 10.094 53.878 10.146 53.914 ;
      RECT 10.094 55.078 10.146 55.114 ;
      RECT 10.094 56.278 10.146 56.314 ;
      RECT 10.094 57.478 10.146 57.514 ;
      RECT 10.094 58.678 10.146 58.714 ;
      RECT 10.094 59.878 10.146 59.914 ;
      RECT 10.094 61.078 10.146 61.114 ;
      RECT 10.094 62.278 10.146 62.314 ;
      RECT 10.094 63.478 10.146 63.514 ;
      RECT 10.094 64.678 10.146 64.714 ;
      RECT 10.094 65.878 10.146 65.914 ;
      RECT 10.094 67.078 10.146 67.114 ;
      RECT 10.094 68.278 10.146 68.314 ;
      RECT 10.094 69.478 10.146 69.514 ;
      RECT 10.094 70.678 10.146 70.714 ;
      RECT 10.094 71.878 10.146 71.914 ;
      RECT 10.174 0.281 10.226 0.317 ;
      RECT 10.174 72.403 10.226 72.439 ;
      RECT 10.254 0.806 10.306 0.842 ;
      RECT 10.254 2.006 10.306 2.042 ;
      RECT 10.254 3.206 10.306 3.242 ;
      RECT 10.254 4.406 10.306 4.442 ;
      RECT 10.254 5.606 10.306 5.642 ;
      RECT 10.254 6.806 10.306 6.842 ;
      RECT 10.254 8.006 10.306 8.042 ;
      RECT 10.254 9.206 10.306 9.242 ;
      RECT 10.254 10.406 10.306 10.442 ;
      RECT 10.254 11.606 10.306 11.642 ;
      RECT 10.254 12.806 10.306 12.842 ;
      RECT 10.254 14.006 10.306 14.042 ;
      RECT 10.254 15.206 10.306 15.242 ;
      RECT 10.254 16.406 10.306 16.442 ;
      RECT 10.254 17.606 10.306 17.642 ;
      RECT 10.254 18.806 10.306 18.842 ;
      RECT 10.254 20.006 10.306 20.042 ;
      RECT 10.254 21.206 10.306 21.242 ;
      RECT 10.254 22.406 10.306 22.442 ;
      RECT 10.254 23.606 10.306 23.642 ;
      RECT 10.254 24.806 10.306 24.842 ;
      RECT 10.254 26.006 10.306 26.042 ;
      RECT 10.254 27.206 10.306 27.242 ;
      RECT 10.254 28.406 10.306 28.442 ;
      RECT 10.254 29.606 10.306 29.642 ;
      RECT 10.254 30.806 10.306 30.842 ;
      RECT 10.254 32.622 10.306 32.658 ;
      RECT 10.254 32.862 10.306 32.898 ;
      RECT 10.254 38.622 10.306 38.658 ;
      RECT 10.254 38.862 10.306 38.898 ;
      RECT 10.254 39.926 10.306 39.962 ;
      RECT 10.254 41.126 10.306 41.162 ;
      RECT 10.254 42.326 10.306 42.362 ;
      RECT 10.254 43.526 10.306 43.562 ;
      RECT 10.254 44.726 10.306 44.762 ;
      RECT 10.254 45.926 10.306 45.962 ;
      RECT 10.254 47.126 10.306 47.162 ;
      RECT 10.254 48.326 10.306 48.362 ;
      RECT 10.254 49.526 10.306 49.562 ;
      RECT 10.254 50.726 10.306 50.762 ;
      RECT 10.254 51.926 10.306 51.962 ;
      RECT 10.254 53.126 10.306 53.162 ;
      RECT 10.254 54.326 10.306 54.362 ;
      RECT 10.254 55.526 10.306 55.562 ;
      RECT 10.254 56.726 10.306 56.762 ;
      RECT 10.254 57.926 10.306 57.962 ;
      RECT 10.254 59.126 10.306 59.162 ;
      RECT 10.254 60.326 10.306 60.362 ;
      RECT 10.254 61.526 10.306 61.562 ;
      RECT 10.254 62.726 10.306 62.762 ;
      RECT 10.254 63.926 10.306 63.962 ;
      RECT 10.254 65.126 10.306 65.162 ;
      RECT 10.254 66.326 10.306 66.362 ;
      RECT 10.254 67.526 10.306 67.562 ;
      RECT 10.254 68.726 10.306 68.762 ;
      RECT 10.254 69.926 10.306 69.962 ;
      RECT 10.254 71.126 10.306 71.162 ;
      RECT 10.334 1.558 10.386 1.594 ;
      RECT 10.334 2.758 10.386 2.794 ;
      RECT 10.334 3.958 10.386 3.994 ;
      RECT 10.334 5.158 10.386 5.194 ;
      RECT 10.334 6.358 10.386 6.394 ;
      RECT 10.334 7.558 10.386 7.594 ;
      RECT 10.334 8.758 10.386 8.794 ;
      RECT 10.334 9.958 10.386 9.994 ;
      RECT 10.334 11.158 10.386 11.194 ;
      RECT 10.334 12.358 10.386 12.394 ;
      RECT 10.334 13.558 10.386 13.594 ;
      RECT 10.334 14.758 10.386 14.794 ;
      RECT 10.334 15.958 10.386 15.994 ;
      RECT 10.334 17.158 10.386 17.194 ;
      RECT 10.334 18.358 10.386 18.394 ;
      RECT 10.334 19.558 10.386 19.594 ;
      RECT 10.334 20.758 10.386 20.794 ;
      RECT 10.334 21.958 10.386 21.994 ;
      RECT 10.334 23.158 10.386 23.194 ;
      RECT 10.334 24.358 10.386 24.394 ;
      RECT 10.334 25.558 10.386 25.594 ;
      RECT 10.334 26.758 10.386 26.794 ;
      RECT 10.334 27.958 10.386 27.994 ;
      RECT 10.334 29.158 10.386 29.194 ;
      RECT 10.334 30.358 10.386 30.394 ;
      RECT 10.334 31.558 10.386 31.594 ;
      RECT 10.334 33.342 10.386 33.378 ;
      RECT 10.334 33.582 10.386 33.618 ;
      RECT 10.334 37.902 10.386 37.938 ;
      RECT 10.334 38.142 10.386 38.178 ;
      RECT 10.334 40.678 10.386 40.714 ;
      RECT 10.334 41.878 10.386 41.914 ;
      RECT 10.334 43.078 10.386 43.114 ;
      RECT 10.334 44.278 10.386 44.314 ;
      RECT 10.334 45.478 10.386 45.514 ;
      RECT 10.334 46.678 10.386 46.714 ;
      RECT 10.334 47.878 10.386 47.914 ;
      RECT 10.334 49.078 10.386 49.114 ;
      RECT 10.334 50.278 10.386 50.314 ;
      RECT 10.334 51.478 10.386 51.514 ;
      RECT 10.334 52.678 10.386 52.714 ;
      RECT 10.334 53.878 10.386 53.914 ;
      RECT 10.334 55.078 10.386 55.114 ;
      RECT 10.334 56.278 10.386 56.314 ;
      RECT 10.334 57.478 10.386 57.514 ;
      RECT 10.334 58.678 10.386 58.714 ;
      RECT 10.334 59.878 10.386 59.914 ;
      RECT 10.334 61.078 10.386 61.114 ;
      RECT 10.334 62.278 10.386 62.314 ;
      RECT 10.334 63.478 10.386 63.514 ;
      RECT 10.334 64.678 10.386 64.714 ;
      RECT 10.334 65.878 10.386 65.914 ;
      RECT 10.334 67.078 10.386 67.114 ;
      RECT 10.334 68.278 10.386 68.314 ;
      RECT 10.334 69.478 10.386 69.514 ;
      RECT 10.334 70.678 10.386 70.714 ;
      RECT 10.334 71.878 10.386 71.914 ;
      RECT 10.414 0.806 10.466 0.842 ;
      RECT 10.414 2.006 10.466 2.042 ;
      RECT 10.414 3.206 10.466 3.242 ;
      RECT 10.414 4.406 10.466 4.442 ;
      RECT 10.414 5.606 10.466 5.642 ;
      RECT 10.414 6.806 10.466 6.842 ;
      RECT 10.414 8.006 10.466 8.042 ;
      RECT 10.414 9.206 10.466 9.242 ;
      RECT 10.414 10.406 10.466 10.442 ;
      RECT 10.414 11.606 10.466 11.642 ;
      RECT 10.414 12.806 10.466 12.842 ;
      RECT 10.414 14.006 10.466 14.042 ;
      RECT 10.414 15.206 10.466 15.242 ;
      RECT 10.414 16.406 10.466 16.442 ;
      RECT 10.414 17.606 10.466 17.642 ;
      RECT 10.414 18.806 10.466 18.842 ;
      RECT 10.414 20.006 10.466 20.042 ;
      RECT 10.414 21.206 10.466 21.242 ;
      RECT 10.414 22.406 10.466 22.442 ;
      RECT 10.414 23.606 10.466 23.642 ;
      RECT 10.414 24.806 10.466 24.842 ;
      RECT 10.414 26.006 10.466 26.042 ;
      RECT 10.414 27.206 10.466 27.242 ;
      RECT 10.414 28.406 10.466 28.442 ;
      RECT 10.414 29.606 10.466 29.642 ;
      RECT 10.414 30.806 10.466 30.842 ;
      RECT 10.414 32.622 10.466 32.658 ;
      RECT 10.414 32.862 10.466 32.898 ;
      RECT 10.414 38.622 10.466 38.658 ;
      RECT 10.414 38.862 10.466 38.898 ;
      RECT 10.414 39.926 10.466 39.962 ;
      RECT 10.414 41.126 10.466 41.162 ;
      RECT 10.414 42.326 10.466 42.362 ;
      RECT 10.414 43.526 10.466 43.562 ;
      RECT 10.414 44.726 10.466 44.762 ;
      RECT 10.414 45.926 10.466 45.962 ;
      RECT 10.414 47.126 10.466 47.162 ;
      RECT 10.414 48.326 10.466 48.362 ;
      RECT 10.414 49.526 10.466 49.562 ;
      RECT 10.414 50.726 10.466 50.762 ;
      RECT 10.414 51.926 10.466 51.962 ;
      RECT 10.414 53.126 10.466 53.162 ;
      RECT 10.414 54.326 10.466 54.362 ;
      RECT 10.414 55.526 10.466 55.562 ;
      RECT 10.414 56.726 10.466 56.762 ;
      RECT 10.414 57.926 10.466 57.962 ;
      RECT 10.414 59.126 10.466 59.162 ;
      RECT 10.414 60.326 10.466 60.362 ;
      RECT 10.414 61.526 10.466 61.562 ;
      RECT 10.414 62.726 10.466 62.762 ;
      RECT 10.414 63.926 10.466 63.962 ;
      RECT 10.414 65.126 10.466 65.162 ;
      RECT 10.414 66.326 10.466 66.362 ;
      RECT 10.414 67.526 10.466 67.562 ;
      RECT 10.414 68.726 10.466 68.762 ;
      RECT 10.414 69.926 10.466 69.962 ;
      RECT 10.414 71.126 10.466 71.162 ;
      RECT 10.494 1.558 10.546 1.594 ;
      RECT 10.494 2.758 10.546 2.794 ;
      RECT 10.494 3.958 10.546 3.994 ;
      RECT 10.494 5.158 10.546 5.194 ;
      RECT 10.494 6.358 10.546 6.394 ;
      RECT 10.494 7.558 10.546 7.594 ;
      RECT 10.494 8.758 10.546 8.794 ;
      RECT 10.494 9.958 10.546 9.994 ;
      RECT 10.494 11.158 10.546 11.194 ;
      RECT 10.494 12.358 10.546 12.394 ;
      RECT 10.494 13.558 10.546 13.594 ;
      RECT 10.494 14.758 10.546 14.794 ;
      RECT 10.494 15.958 10.546 15.994 ;
      RECT 10.494 17.158 10.546 17.194 ;
      RECT 10.494 18.358 10.546 18.394 ;
      RECT 10.494 19.558 10.546 19.594 ;
      RECT 10.494 20.758 10.546 20.794 ;
      RECT 10.494 21.958 10.546 21.994 ;
      RECT 10.494 23.158 10.546 23.194 ;
      RECT 10.494 24.358 10.546 24.394 ;
      RECT 10.494 25.558 10.546 25.594 ;
      RECT 10.494 26.758 10.546 26.794 ;
      RECT 10.494 27.958 10.546 27.994 ;
      RECT 10.494 29.158 10.546 29.194 ;
      RECT 10.494 30.358 10.546 30.394 ;
      RECT 10.494 31.558 10.546 31.594 ;
      RECT 10.494 33.342 10.546 33.378 ;
      RECT 10.494 33.582 10.546 33.618 ;
      RECT 10.494 37.902 10.546 37.938 ;
      RECT 10.494 38.142 10.546 38.178 ;
      RECT 10.494 40.678 10.546 40.714 ;
      RECT 10.494 41.878 10.546 41.914 ;
      RECT 10.494 43.078 10.546 43.114 ;
      RECT 10.494 44.278 10.546 44.314 ;
      RECT 10.494 45.478 10.546 45.514 ;
      RECT 10.494 46.678 10.546 46.714 ;
      RECT 10.494 47.878 10.546 47.914 ;
      RECT 10.494 49.078 10.546 49.114 ;
      RECT 10.494 50.278 10.546 50.314 ;
      RECT 10.494 51.478 10.546 51.514 ;
      RECT 10.494 52.678 10.546 52.714 ;
      RECT 10.494 53.878 10.546 53.914 ;
      RECT 10.494 55.078 10.546 55.114 ;
      RECT 10.494 56.278 10.546 56.314 ;
      RECT 10.494 57.478 10.546 57.514 ;
      RECT 10.494 58.678 10.546 58.714 ;
      RECT 10.494 59.878 10.546 59.914 ;
      RECT 10.494 61.078 10.546 61.114 ;
      RECT 10.494 62.278 10.546 62.314 ;
      RECT 10.494 63.478 10.546 63.514 ;
      RECT 10.494 64.678 10.546 64.714 ;
      RECT 10.494 65.878 10.546 65.914 ;
      RECT 10.494 67.078 10.546 67.114 ;
      RECT 10.494 68.278 10.546 68.314 ;
      RECT 10.494 69.478 10.546 69.514 ;
      RECT 10.494 70.678 10.546 70.714 ;
      RECT 10.494 71.878 10.546 71.914 ;
      RECT 10.574 0.281 10.626 0.317 ;
      RECT 10.574 72.403 10.626 72.439 ;
      RECT 10.654 0.806 10.706 0.842 ;
      RECT 10.654 2.006 10.706 2.042 ;
      RECT 10.654 3.206 10.706 3.242 ;
      RECT 10.654 4.406 10.706 4.442 ;
      RECT 10.654 5.606 10.706 5.642 ;
      RECT 10.654 6.806 10.706 6.842 ;
      RECT 10.654 8.006 10.706 8.042 ;
      RECT 10.654 9.206 10.706 9.242 ;
      RECT 10.654 10.406 10.706 10.442 ;
      RECT 10.654 11.606 10.706 11.642 ;
      RECT 10.654 12.806 10.706 12.842 ;
      RECT 10.654 14.006 10.706 14.042 ;
      RECT 10.654 15.206 10.706 15.242 ;
      RECT 10.654 16.406 10.706 16.442 ;
      RECT 10.654 17.606 10.706 17.642 ;
      RECT 10.654 18.806 10.706 18.842 ;
      RECT 10.654 20.006 10.706 20.042 ;
      RECT 10.654 21.206 10.706 21.242 ;
      RECT 10.654 22.406 10.706 22.442 ;
      RECT 10.654 23.606 10.706 23.642 ;
      RECT 10.654 24.806 10.706 24.842 ;
      RECT 10.654 26.006 10.706 26.042 ;
      RECT 10.654 27.206 10.706 27.242 ;
      RECT 10.654 28.406 10.706 28.442 ;
      RECT 10.654 29.606 10.706 29.642 ;
      RECT 10.654 30.806 10.706 30.842 ;
      RECT 10.654 32.622 10.706 32.658 ;
      RECT 10.654 32.862 10.706 32.898 ;
      RECT 10.654 34.302 10.706 34.338 ;
      RECT 10.654 34.782 10.706 34.818 ;
      RECT 10.654 36.702 10.706 36.738 ;
      RECT 10.654 37.182 10.706 37.218 ;
      RECT 10.654 38.622 10.706 38.658 ;
      RECT 10.654 38.862 10.706 38.898 ;
      RECT 10.654 39.926 10.706 39.962 ;
      RECT 10.654 41.126 10.706 41.162 ;
      RECT 10.654 42.326 10.706 42.362 ;
      RECT 10.654 43.526 10.706 43.562 ;
      RECT 10.654 44.726 10.706 44.762 ;
      RECT 10.654 45.926 10.706 45.962 ;
      RECT 10.654 47.126 10.706 47.162 ;
      RECT 10.654 48.326 10.706 48.362 ;
      RECT 10.654 49.526 10.706 49.562 ;
      RECT 10.654 50.726 10.706 50.762 ;
      RECT 10.654 51.926 10.706 51.962 ;
      RECT 10.654 53.126 10.706 53.162 ;
      RECT 10.654 54.326 10.706 54.362 ;
      RECT 10.654 55.526 10.706 55.562 ;
      RECT 10.654 56.726 10.706 56.762 ;
      RECT 10.654 57.926 10.706 57.962 ;
      RECT 10.654 59.126 10.706 59.162 ;
      RECT 10.654 60.326 10.706 60.362 ;
      RECT 10.654 61.526 10.706 61.562 ;
      RECT 10.654 62.726 10.706 62.762 ;
      RECT 10.654 63.926 10.706 63.962 ;
      RECT 10.654 65.126 10.706 65.162 ;
      RECT 10.654 66.326 10.706 66.362 ;
      RECT 10.654 67.526 10.706 67.562 ;
      RECT 10.654 68.726 10.706 68.762 ;
      RECT 10.654 69.926 10.706 69.962 ;
      RECT 10.654 71.126 10.706 71.162 ;
      RECT 10.734 1.558 10.786 1.594 ;
      RECT 10.734 2.758 10.786 2.794 ;
      RECT 10.734 3.958 10.786 3.994 ;
      RECT 10.734 5.158 10.786 5.194 ;
      RECT 10.734 6.358 10.786 6.394 ;
      RECT 10.734 7.558 10.786 7.594 ;
      RECT 10.734 8.758 10.786 8.794 ;
      RECT 10.734 9.958 10.786 9.994 ;
      RECT 10.734 11.158 10.786 11.194 ;
      RECT 10.734 12.358 10.786 12.394 ;
      RECT 10.734 13.558 10.786 13.594 ;
      RECT 10.734 14.758 10.786 14.794 ;
      RECT 10.734 15.958 10.786 15.994 ;
      RECT 10.734 17.158 10.786 17.194 ;
      RECT 10.734 18.358 10.786 18.394 ;
      RECT 10.734 19.558 10.786 19.594 ;
      RECT 10.734 20.758 10.786 20.794 ;
      RECT 10.734 21.958 10.786 21.994 ;
      RECT 10.734 23.158 10.786 23.194 ;
      RECT 10.734 24.358 10.786 24.394 ;
      RECT 10.734 25.558 10.786 25.594 ;
      RECT 10.734 26.758 10.786 26.794 ;
      RECT 10.734 27.958 10.786 27.994 ;
      RECT 10.734 29.158 10.786 29.194 ;
      RECT 10.734 30.358 10.786 30.394 ;
      RECT 10.734 31.558 10.786 31.594 ;
      RECT 10.734 33.342 10.786 33.378 ;
      RECT 10.734 33.582 10.786 33.618 ;
      RECT 10.734 37.902 10.786 37.938 ;
      RECT 10.734 38.142 10.786 38.178 ;
      RECT 10.734 40.678 10.786 40.714 ;
      RECT 10.734 41.878 10.786 41.914 ;
      RECT 10.734 43.078 10.786 43.114 ;
      RECT 10.734 44.278 10.786 44.314 ;
      RECT 10.734 45.478 10.786 45.514 ;
      RECT 10.734 46.678 10.786 46.714 ;
      RECT 10.734 47.878 10.786 47.914 ;
      RECT 10.734 49.078 10.786 49.114 ;
      RECT 10.734 50.278 10.786 50.314 ;
      RECT 10.734 51.478 10.786 51.514 ;
      RECT 10.734 52.678 10.786 52.714 ;
      RECT 10.734 53.878 10.786 53.914 ;
      RECT 10.734 55.078 10.786 55.114 ;
      RECT 10.734 56.278 10.786 56.314 ;
      RECT 10.734 57.478 10.786 57.514 ;
      RECT 10.734 58.678 10.786 58.714 ;
      RECT 10.734 59.878 10.786 59.914 ;
      RECT 10.734 61.078 10.786 61.114 ;
      RECT 10.734 62.278 10.786 62.314 ;
      RECT 10.734 63.478 10.786 63.514 ;
      RECT 10.734 64.678 10.786 64.714 ;
      RECT 10.734 65.878 10.786 65.914 ;
      RECT 10.734 67.078 10.786 67.114 ;
      RECT 10.734 68.278 10.786 68.314 ;
      RECT 10.734 69.478 10.786 69.514 ;
      RECT 10.734 70.678 10.786 70.714 ;
      RECT 10.734 71.878 10.786 71.914 ;
      RECT 10.814 0.806 10.866 0.842 ;
      RECT 10.814 2.006 10.866 2.042 ;
      RECT 10.814 3.206 10.866 3.242 ;
      RECT 10.814 4.406 10.866 4.442 ;
      RECT 10.814 5.606 10.866 5.642 ;
      RECT 10.814 6.806 10.866 6.842 ;
      RECT 10.814 8.006 10.866 8.042 ;
      RECT 10.814 9.206 10.866 9.242 ;
      RECT 10.814 10.406 10.866 10.442 ;
      RECT 10.814 11.606 10.866 11.642 ;
      RECT 10.814 12.806 10.866 12.842 ;
      RECT 10.814 14.006 10.866 14.042 ;
      RECT 10.814 15.206 10.866 15.242 ;
      RECT 10.814 16.406 10.866 16.442 ;
      RECT 10.814 17.606 10.866 17.642 ;
      RECT 10.814 18.806 10.866 18.842 ;
      RECT 10.814 20.006 10.866 20.042 ;
      RECT 10.814 21.206 10.866 21.242 ;
      RECT 10.814 22.406 10.866 22.442 ;
      RECT 10.814 23.606 10.866 23.642 ;
      RECT 10.814 24.806 10.866 24.842 ;
      RECT 10.814 26.006 10.866 26.042 ;
      RECT 10.814 27.206 10.866 27.242 ;
      RECT 10.814 28.406 10.866 28.442 ;
      RECT 10.814 29.606 10.866 29.642 ;
      RECT 10.814 30.806 10.866 30.842 ;
      RECT 10.814 32.622 10.866 32.658 ;
      RECT 10.814 32.862 10.866 32.898 ;
      RECT 10.814 38.622 10.866 38.658 ;
      RECT 10.814 38.862 10.866 38.898 ;
      RECT 10.814 39.926 10.866 39.962 ;
      RECT 10.814 41.126 10.866 41.162 ;
      RECT 10.814 42.326 10.866 42.362 ;
      RECT 10.814 43.526 10.866 43.562 ;
      RECT 10.814 44.726 10.866 44.762 ;
      RECT 10.814 45.926 10.866 45.962 ;
      RECT 10.814 47.126 10.866 47.162 ;
      RECT 10.814 48.326 10.866 48.362 ;
      RECT 10.814 49.526 10.866 49.562 ;
      RECT 10.814 50.726 10.866 50.762 ;
      RECT 10.814 51.926 10.866 51.962 ;
      RECT 10.814 53.126 10.866 53.162 ;
      RECT 10.814 54.326 10.866 54.362 ;
      RECT 10.814 55.526 10.866 55.562 ;
      RECT 10.814 56.726 10.866 56.762 ;
      RECT 10.814 57.926 10.866 57.962 ;
      RECT 10.814 59.126 10.866 59.162 ;
      RECT 10.814 60.326 10.866 60.362 ;
      RECT 10.814 61.526 10.866 61.562 ;
      RECT 10.814 62.726 10.866 62.762 ;
      RECT 10.814 63.926 10.866 63.962 ;
      RECT 10.814 65.126 10.866 65.162 ;
      RECT 10.814 66.326 10.866 66.362 ;
      RECT 10.814 67.526 10.866 67.562 ;
      RECT 10.814 68.726 10.866 68.762 ;
      RECT 10.814 69.926 10.866 69.962 ;
      RECT 10.814 71.126 10.866 71.162 ;
      RECT 10.894 1.558 10.946 1.594 ;
      RECT 10.894 2.758 10.946 2.794 ;
      RECT 10.894 3.958 10.946 3.994 ;
      RECT 10.894 5.158 10.946 5.194 ;
      RECT 10.894 6.358 10.946 6.394 ;
      RECT 10.894 7.558 10.946 7.594 ;
      RECT 10.894 8.758 10.946 8.794 ;
      RECT 10.894 9.958 10.946 9.994 ;
      RECT 10.894 11.158 10.946 11.194 ;
      RECT 10.894 12.358 10.946 12.394 ;
      RECT 10.894 13.558 10.946 13.594 ;
      RECT 10.894 14.758 10.946 14.794 ;
      RECT 10.894 15.958 10.946 15.994 ;
      RECT 10.894 17.158 10.946 17.194 ;
      RECT 10.894 18.358 10.946 18.394 ;
      RECT 10.894 19.558 10.946 19.594 ;
      RECT 10.894 20.758 10.946 20.794 ;
      RECT 10.894 21.958 10.946 21.994 ;
      RECT 10.894 23.158 10.946 23.194 ;
      RECT 10.894 24.358 10.946 24.394 ;
      RECT 10.894 25.558 10.946 25.594 ;
      RECT 10.894 26.758 10.946 26.794 ;
      RECT 10.894 27.958 10.946 27.994 ;
      RECT 10.894 29.158 10.946 29.194 ;
      RECT 10.894 30.358 10.946 30.394 ;
      RECT 10.894 31.558 10.946 31.594 ;
      RECT 10.894 33.342 10.946 33.378 ;
      RECT 10.894 33.582 10.946 33.618 ;
      RECT 10.894 37.902 10.946 37.938 ;
      RECT 10.894 38.142 10.946 38.178 ;
      RECT 10.894 40.678 10.946 40.714 ;
      RECT 10.894 41.878 10.946 41.914 ;
      RECT 10.894 43.078 10.946 43.114 ;
      RECT 10.894 44.278 10.946 44.314 ;
      RECT 10.894 45.478 10.946 45.514 ;
      RECT 10.894 46.678 10.946 46.714 ;
      RECT 10.894 47.878 10.946 47.914 ;
      RECT 10.894 49.078 10.946 49.114 ;
      RECT 10.894 50.278 10.946 50.314 ;
      RECT 10.894 51.478 10.946 51.514 ;
      RECT 10.894 52.678 10.946 52.714 ;
      RECT 10.894 53.878 10.946 53.914 ;
      RECT 10.894 55.078 10.946 55.114 ;
      RECT 10.894 56.278 10.946 56.314 ;
      RECT 10.894 57.478 10.946 57.514 ;
      RECT 10.894 58.678 10.946 58.714 ;
      RECT 10.894 59.878 10.946 59.914 ;
      RECT 10.894 61.078 10.946 61.114 ;
      RECT 10.894 62.278 10.946 62.314 ;
      RECT 10.894 63.478 10.946 63.514 ;
      RECT 10.894 64.678 10.946 64.714 ;
      RECT 10.894 65.878 10.946 65.914 ;
      RECT 10.894 67.078 10.946 67.114 ;
      RECT 10.894 68.278 10.946 68.314 ;
      RECT 10.894 69.478 10.946 69.514 ;
      RECT 10.894 70.678 10.946 70.714 ;
      RECT 10.894 71.878 10.946 71.914 ;
      RECT 10.974 0.281 11.026 0.317 ;
      RECT 10.974 72.403 11.026 72.439 ;
      RECT 11.054 0.806 11.106 0.842 ;
      RECT 11.054 2.006 11.106 2.042 ;
      RECT 11.054 3.206 11.106 3.242 ;
      RECT 11.054 4.406 11.106 4.442 ;
      RECT 11.054 5.606 11.106 5.642 ;
      RECT 11.054 6.806 11.106 6.842 ;
      RECT 11.054 8.006 11.106 8.042 ;
      RECT 11.054 9.206 11.106 9.242 ;
      RECT 11.054 10.406 11.106 10.442 ;
      RECT 11.054 11.606 11.106 11.642 ;
      RECT 11.054 12.806 11.106 12.842 ;
      RECT 11.054 14.006 11.106 14.042 ;
      RECT 11.054 15.206 11.106 15.242 ;
      RECT 11.054 16.406 11.106 16.442 ;
      RECT 11.054 17.606 11.106 17.642 ;
      RECT 11.054 18.806 11.106 18.842 ;
      RECT 11.054 20.006 11.106 20.042 ;
      RECT 11.054 21.206 11.106 21.242 ;
      RECT 11.054 22.406 11.106 22.442 ;
      RECT 11.054 23.606 11.106 23.642 ;
      RECT 11.054 24.806 11.106 24.842 ;
      RECT 11.054 26.006 11.106 26.042 ;
      RECT 11.054 27.206 11.106 27.242 ;
      RECT 11.054 28.406 11.106 28.442 ;
      RECT 11.054 29.606 11.106 29.642 ;
      RECT 11.054 30.806 11.106 30.842 ;
      RECT 11.054 32.622 11.106 32.658 ;
      RECT 11.054 32.862 11.106 32.898 ;
      RECT 11.054 38.622 11.106 38.658 ;
      RECT 11.054 38.862 11.106 38.898 ;
      RECT 11.054 39.926 11.106 39.962 ;
      RECT 11.054 41.126 11.106 41.162 ;
      RECT 11.054 42.326 11.106 42.362 ;
      RECT 11.054 43.526 11.106 43.562 ;
      RECT 11.054 44.726 11.106 44.762 ;
      RECT 11.054 45.926 11.106 45.962 ;
      RECT 11.054 47.126 11.106 47.162 ;
      RECT 11.054 48.326 11.106 48.362 ;
      RECT 11.054 49.526 11.106 49.562 ;
      RECT 11.054 50.726 11.106 50.762 ;
      RECT 11.054 51.926 11.106 51.962 ;
      RECT 11.054 53.126 11.106 53.162 ;
      RECT 11.054 54.326 11.106 54.362 ;
      RECT 11.054 55.526 11.106 55.562 ;
      RECT 11.054 56.726 11.106 56.762 ;
      RECT 11.054 57.926 11.106 57.962 ;
      RECT 11.054 59.126 11.106 59.162 ;
      RECT 11.054 60.326 11.106 60.362 ;
      RECT 11.054 61.526 11.106 61.562 ;
      RECT 11.054 62.726 11.106 62.762 ;
      RECT 11.054 63.926 11.106 63.962 ;
      RECT 11.054 65.126 11.106 65.162 ;
      RECT 11.054 66.326 11.106 66.362 ;
      RECT 11.054 67.526 11.106 67.562 ;
      RECT 11.054 68.726 11.106 68.762 ;
      RECT 11.054 69.926 11.106 69.962 ;
      RECT 11.054 71.126 11.106 71.162 ;
      RECT 11.134 1.558 11.186 1.594 ;
      RECT 11.134 2.758 11.186 2.794 ;
      RECT 11.134 3.958 11.186 3.994 ;
      RECT 11.134 5.158 11.186 5.194 ;
      RECT 11.134 6.358 11.186 6.394 ;
      RECT 11.134 7.558 11.186 7.594 ;
      RECT 11.134 8.758 11.186 8.794 ;
      RECT 11.134 9.958 11.186 9.994 ;
      RECT 11.134 11.158 11.186 11.194 ;
      RECT 11.134 12.358 11.186 12.394 ;
      RECT 11.134 13.558 11.186 13.594 ;
      RECT 11.134 14.758 11.186 14.794 ;
      RECT 11.134 15.958 11.186 15.994 ;
      RECT 11.134 17.158 11.186 17.194 ;
      RECT 11.134 18.358 11.186 18.394 ;
      RECT 11.134 19.558 11.186 19.594 ;
      RECT 11.134 20.758 11.186 20.794 ;
      RECT 11.134 21.958 11.186 21.994 ;
      RECT 11.134 23.158 11.186 23.194 ;
      RECT 11.134 24.358 11.186 24.394 ;
      RECT 11.134 25.558 11.186 25.594 ;
      RECT 11.134 26.758 11.186 26.794 ;
      RECT 11.134 27.958 11.186 27.994 ;
      RECT 11.134 29.158 11.186 29.194 ;
      RECT 11.134 30.358 11.186 30.394 ;
      RECT 11.134 31.558 11.186 31.594 ;
      RECT 11.134 33.342 11.186 33.378 ;
      RECT 11.134 33.582 11.186 33.618 ;
      RECT 11.134 37.902 11.186 37.938 ;
      RECT 11.134 38.142 11.186 38.178 ;
      RECT 11.134 40.678 11.186 40.714 ;
      RECT 11.134 41.878 11.186 41.914 ;
      RECT 11.134 43.078 11.186 43.114 ;
      RECT 11.134 44.278 11.186 44.314 ;
      RECT 11.134 45.478 11.186 45.514 ;
      RECT 11.134 46.678 11.186 46.714 ;
      RECT 11.134 47.878 11.186 47.914 ;
      RECT 11.134 49.078 11.186 49.114 ;
      RECT 11.134 50.278 11.186 50.314 ;
      RECT 11.134 51.478 11.186 51.514 ;
      RECT 11.134 52.678 11.186 52.714 ;
      RECT 11.134 53.878 11.186 53.914 ;
      RECT 11.134 55.078 11.186 55.114 ;
      RECT 11.134 56.278 11.186 56.314 ;
      RECT 11.134 57.478 11.186 57.514 ;
      RECT 11.134 58.678 11.186 58.714 ;
      RECT 11.134 59.878 11.186 59.914 ;
      RECT 11.134 61.078 11.186 61.114 ;
      RECT 11.134 62.278 11.186 62.314 ;
      RECT 11.134 63.478 11.186 63.514 ;
      RECT 11.134 64.678 11.186 64.714 ;
      RECT 11.134 65.878 11.186 65.914 ;
      RECT 11.134 67.078 11.186 67.114 ;
      RECT 11.134 68.278 11.186 68.314 ;
      RECT 11.134 69.478 11.186 69.514 ;
      RECT 11.134 70.678 11.186 70.714 ;
      RECT 11.134 71.878 11.186 71.914 ;
      RECT 11.214 0.806 11.266 0.842 ;
      RECT 11.214 2.006 11.266 2.042 ;
      RECT 11.214 3.206 11.266 3.242 ;
      RECT 11.214 4.406 11.266 4.442 ;
      RECT 11.214 5.606 11.266 5.642 ;
      RECT 11.214 6.806 11.266 6.842 ;
      RECT 11.214 8.006 11.266 8.042 ;
      RECT 11.214 9.206 11.266 9.242 ;
      RECT 11.214 10.406 11.266 10.442 ;
      RECT 11.214 11.606 11.266 11.642 ;
      RECT 11.214 12.806 11.266 12.842 ;
      RECT 11.214 14.006 11.266 14.042 ;
      RECT 11.214 15.206 11.266 15.242 ;
      RECT 11.214 16.406 11.266 16.442 ;
      RECT 11.214 17.606 11.266 17.642 ;
      RECT 11.214 18.806 11.266 18.842 ;
      RECT 11.214 20.006 11.266 20.042 ;
      RECT 11.214 21.206 11.266 21.242 ;
      RECT 11.214 22.406 11.266 22.442 ;
      RECT 11.214 23.606 11.266 23.642 ;
      RECT 11.214 24.806 11.266 24.842 ;
      RECT 11.214 26.006 11.266 26.042 ;
      RECT 11.214 27.206 11.266 27.242 ;
      RECT 11.214 28.406 11.266 28.442 ;
      RECT 11.214 29.606 11.266 29.642 ;
      RECT 11.214 30.806 11.266 30.842 ;
      RECT 11.214 32.622 11.266 32.658 ;
      RECT 11.214 32.862 11.266 32.898 ;
      RECT 11.214 38.622 11.266 38.658 ;
      RECT 11.214 38.862 11.266 38.898 ;
      RECT 11.214 39.926 11.266 39.962 ;
      RECT 11.214 41.126 11.266 41.162 ;
      RECT 11.214 42.326 11.266 42.362 ;
      RECT 11.214 43.526 11.266 43.562 ;
      RECT 11.214 44.726 11.266 44.762 ;
      RECT 11.214 45.926 11.266 45.962 ;
      RECT 11.214 47.126 11.266 47.162 ;
      RECT 11.214 48.326 11.266 48.362 ;
      RECT 11.214 49.526 11.266 49.562 ;
      RECT 11.214 50.726 11.266 50.762 ;
      RECT 11.214 51.926 11.266 51.962 ;
      RECT 11.214 53.126 11.266 53.162 ;
      RECT 11.214 54.326 11.266 54.362 ;
      RECT 11.214 55.526 11.266 55.562 ;
      RECT 11.214 56.726 11.266 56.762 ;
      RECT 11.214 57.926 11.266 57.962 ;
      RECT 11.214 59.126 11.266 59.162 ;
      RECT 11.214 60.326 11.266 60.362 ;
      RECT 11.214 61.526 11.266 61.562 ;
      RECT 11.214 62.726 11.266 62.762 ;
      RECT 11.214 63.926 11.266 63.962 ;
      RECT 11.214 65.126 11.266 65.162 ;
      RECT 11.214 66.326 11.266 66.362 ;
      RECT 11.214 67.526 11.266 67.562 ;
      RECT 11.214 68.726 11.266 68.762 ;
      RECT 11.214 69.926 11.266 69.962 ;
      RECT 11.214 71.126 11.266 71.162 ;
      RECT 11.294 1.558 11.346 1.594 ;
      RECT 11.294 2.758 11.346 2.794 ;
      RECT 11.294 3.958 11.346 3.994 ;
      RECT 11.294 5.158 11.346 5.194 ;
      RECT 11.294 6.358 11.346 6.394 ;
      RECT 11.294 7.558 11.346 7.594 ;
      RECT 11.294 8.758 11.346 8.794 ;
      RECT 11.294 9.958 11.346 9.994 ;
      RECT 11.294 11.158 11.346 11.194 ;
      RECT 11.294 12.358 11.346 12.394 ;
      RECT 11.294 13.558 11.346 13.594 ;
      RECT 11.294 14.758 11.346 14.794 ;
      RECT 11.294 15.958 11.346 15.994 ;
      RECT 11.294 17.158 11.346 17.194 ;
      RECT 11.294 18.358 11.346 18.394 ;
      RECT 11.294 19.558 11.346 19.594 ;
      RECT 11.294 20.758 11.346 20.794 ;
      RECT 11.294 21.958 11.346 21.994 ;
      RECT 11.294 23.158 11.346 23.194 ;
      RECT 11.294 24.358 11.346 24.394 ;
      RECT 11.294 25.558 11.346 25.594 ;
      RECT 11.294 26.758 11.346 26.794 ;
      RECT 11.294 27.958 11.346 27.994 ;
      RECT 11.294 29.158 11.346 29.194 ;
      RECT 11.294 30.358 11.346 30.394 ;
      RECT 11.294 31.558 11.346 31.594 ;
      RECT 11.294 33.342 11.346 33.378 ;
      RECT 11.294 33.582 11.346 33.618 ;
      RECT 11.294 37.902 11.346 37.938 ;
      RECT 11.294 38.142 11.346 38.178 ;
      RECT 11.294 40.678 11.346 40.714 ;
      RECT 11.294 41.878 11.346 41.914 ;
      RECT 11.294 43.078 11.346 43.114 ;
      RECT 11.294 44.278 11.346 44.314 ;
      RECT 11.294 45.478 11.346 45.514 ;
      RECT 11.294 46.678 11.346 46.714 ;
      RECT 11.294 47.878 11.346 47.914 ;
      RECT 11.294 49.078 11.346 49.114 ;
      RECT 11.294 50.278 11.346 50.314 ;
      RECT 11.294 51.478 11.346 51.514 ;
      RECT 11.294 52.678 11.346 52.714 ;
      RECT 11.294 53.878 11.346 53.914 ;
      RECT 11.294 55.078 11.346 55.114 ;
      RECT 11.294 56.278 11.346 56.314 ;
      RECT 11.294 57.478 11.346 57.514 ;
      RECT 11.294 58.678 11.346 58.714 ;
      RECT 11.294 59.878 11.346 59.914 ;
      RECT 11.294 61.078 11.346 61.114 ;
      RECT 11.294 62.278 11.346 62.314 ;
      RECT 11.294 63.478 11.346 63.514 ;
      RECT 11.294 64.678 11.346 64.714 ;
      RECT 11.294 65.878 11.346 65.914 ;
      RECT 11.294 67.078 11.346 67.114 ;
      RECT 11.294 68.278 11.346 68.314 ;
      RECT 11.294 69.478 11.346 69.514 ;
      RECT 11.294 70.678 11.346 70.714 ;
      RECT 11.294 71.878 11.346 71.914 ;
      RECT 11.374 0.281 11.426 0.317 ;
      RECT 11.374 72.403 11.426 72.439 ;
      RECT 11.454 0.806 11.506 0.842 ;
      RECT 11.454 2.006 11.506 2.042 ;
      RECT 11.454 3.206 11.506 3.242 ;
      RECT 11.454 4.406 11.506 4.442 ;
      RECT 11.454 5.606 11.506 5.642 ;
      RECT 11.454 6.806 11.506 6.842 ;
      RECT 11.454 8.006 11.506 8.042 ;
      RECT 11.454 9.206 11.506 9.242 ;
      RECT 11.454 10.406 11.506 10.442 ;
      RECT 11.454 11.606 11.506 11.642 ;
      RECT 11.454 12.806 11.506 12.842 ;
      RECT 11.454 14.006 11.506 14.042 ;
      RECT 11.454 15.206 11.506 15.242 ;
      RECT 11.454 16.406 11.506 16.442 ;
      RECT 11.454 17.606 11.506 17.642 ;
      RECT 11.454 18.806 11.506 18.842 ;
      RECT 11.454 20.006 11.506 20.042 ;
      RECT 11.454 21.206 11.506 21.242 ;
      RECT 11.454 22.406 11.506 22.442 ;
      RECT 11.454 23.606 11.506 23.642 ;
      RECT 11.454 24.806 11.506 24.842 ;
      RECT 11.454 26.006 11.506 26.042 ;
      RECT 11.454 27.206 11.506 27.242 ;
      RECT 11.454 28.406 11.506 28.442 ;
      RECT 11.454 29.606 11.506 29.642 ;
      RECT 11.454 30.806 11.506 30.842 ;
      RECT 11.454 32.622 11.506 32.658 ;
      RECT 11.454 32.862 11.506 32.898 ;
      RECT 11.454 34.302 11.506 34.338 ;
      RECT 11.454 34.782 11.506 34.818 ;
      RECT 11.454 36.702 11.506 36.738 ;
      RECT 11.454 37.182 11.506 37.218 ;
      RECT 11.454 38.622 11.506 38.658 ;
      RECT 11.454 38.862 11.506 38.898 ;
      RECT 11.454 39.926 11.506 39.962 ;
      RECT 11.454 41.126 11.506 41.162 ;
      RECT 11.454 42.326 11.506 42.362 ;
      RECT 11.454 43.526 11.506 43.562 ;
      RECT 11.454 44.726 11.506 44.762 ;
      RECT 11.454 45.926 11.506 45.962 ;
      RECT 11.454 47.126 11.506 47.162 ;
      RECT 11.454 48.326 11.506 48.362 ;
      RECT 11.454 49.526 11.506 49.562 ;
      RECT 11.454 50.726 11.506 50.762 ;
      RECT 11.454 51.926 11.506 51.962 ;
      RECT 11.454 53.126 11.506 53.162 ;
      RECT 11.454 54.326 11.506 54.362 ;
      RECT 11.454 55.526 11.506 55.562 ;
      RECT 11.454 56.726 11.506 56.762 ;
      RECT 11.454 57.926 11.506 57.962 ;
      RECT 11.454 59.126 11.506 59.162 ;
      RECT 11.454 60.326 11.506 60.362 ;
      RECT 11.454 61.526 11.506 61.562 ;
      RECT 11.454 62.726 11.506 62.762 ;
      RECT 11.454 63.926 11.506 63.962 ;
      RECT 11.454 65.126 11.506 65.162 ;
      RECT 11.454 66.326 11.506 66.362 ;
      RECT 11.454 67.526 11.506 67.562 ;
      RECT 11.454 68.726 11.506 68.762 ;
      RECT 11.454 69.926 11.506 69.962 ;
      RECT 11.454 71.126 11.506 71.162 ;
      RECT 11.534 1.558 11.586 1.594 ;
      RECT 11.534 2.758 11.586 2.794 ;
      RECT 11.534 3.958 11.586 3.994 ;
      RECT 11.534 5.158 11.586 5.194 ;
      RECT 11.534 6.358 11.586 6.394 ;
      RECT 11.534 7.558 11.586 7.594 ;
      RECT 11.534 8.758 11.586 8.794 ;
      RECT 11.534 9.958 11.586 9.994 ;
      RECT 11.534 11.158 11.586 11.194 ;
      RECT 11.534 12.358 11.586 12.394 ;
      RECT 11.534 13.558 11.586 13.594 ;
      RECT 11.534 14.758 11.586 14.794 ;
      RECT 11.534 15.958 11.586 15.994 ;
      RECT 11.534 17.158 11.586 17.194 ;
      RECT 11.534 18.358 11.586 18.394 ;
      RECT 11.534 19.558 11.586 19.594 ;
      RECT 11.534 20.758 11.586 20.794 ;
      RECT 11.534 21.958 11.586 21.994 ;
      RECT 11.534 23.158 11.586 23.194 ;
      RECT 11.534 24.358 11.586 24.394 ;
      RECT 11.534 25.558 11.586 25.594 ;
      RECT 11.534 26.758 11.586 26.794 ;
      RECT 11.534 27.958 11.586 27.994 ;
      RECT 11.534 29.158 11.586 29.194 ;
      RECT 11.534 30.358 11.586 30.394 ;
      RECT 11.534 31.558 11.586 31.594 ;
      RECT 11.534 33.342 11.586 33.378 ;
      RECT 11.534 33.582 11.586 33.618 ;
      RECT 11.534 37.902 11.586 37.938 ;
      RECT 11.534 38.142 11.586 38.178 ;
      RECT 11.534 40.678 11.586 40.714 ;
      RECT 11.534 41.878 11.586 41.914 ;
      RECT 11.534 43.078 11.586 43.114 ;
      RECT 11.534 44.278 11.586 44.314 ;
      RECT 11.534 45.478 11.586 45.514 ;
      RECT 11.534 46.678 11.586 46.714 ;
      RECT 11.534 47.878 11.586 47.914 ;
      RECT 11.534 49.078 11.586 49.114 ;
      RECT 11.534 50.278 11.586 50.314 ;
      RECT 11.534 51.478 11.586 51.514 ;
      RECT 11.534 52.678 11.586 52.714 ;
      RECT 11.534 53.878 11.586 53.914 ;
      RECT 11.534 55.078 11.586 55.114 ;
      RECT 11.534 56.278 11.586 56.314 ;
      RECT 11.534 57.478 11.586 57.514 ;
      RECT 11.534 58.678 11.586 58.714 ;
      RECT 11.534 59.878 11.586 59.914 ;
      RECT 11.534 61.078 11.586 61.114 ;
      RECT 11.534 62.278 11.586 62.314 ;
      RECT 11.534 63.478 11.586 63.514 ;
      RECT 11.534 64.678 11.586 64.714 ;
      RECT 11.534 65.878 11.586 65.914 ;
      RECT 11.534 67.078 11.586 67.114 ;
      RECT 11.534 68.278 11.586 68.314 ;
      RECT 11.534 69.478 11.586 69.514 ;
      RECT 11.534 70.678 11.586 70.714 ;
      RECT 11.534 71.878 11.586 71.914 ;
      RECT 11.614 0.806 11.666 0.842 ;
      RECT 11.614 2.006 11.666 2.042 ;
      RECT 11.614 3.206 11.666 3.242 ;
      RECT 11.614 4.406 11.666 4.442 ;
      RECT 11.614 5.606 11.666 5.642 ;
      RECT 11.614 6.806 11.666 6.842 ;
      RECT 11.614 8.006 11.666 8.042 ;
      RECT 11.614 9.206 11.666 9.242 ;
      RECT 11.614 10.406 11.666 10.442 ;
      RECT 11.614 11.606 11.666 11.642 ;
      RECT 11.614 12.806 11.666 12.842 ;
      RECT 11.614 14.006 11.666 14.042 ;
      RECT 11.614 15.206 11.666 15.242 ;
      RECT 11.614 16.406 11.666 16.442 ;
      RECT 11.614 17.606 11.666 17.642 ;
      RECT 11.614 18.806 11.666 18.842 ;
      RECT 11.614 20.006 11.666 20.042 ;
      RECT 11.614 21.206 11.666 21.242 ;
      RECT 11.614 22.406 11.666 22.442 ;
      RECT 11.614 23.606 11.666 23.642 ;
      RECT 11.614 24.806 11.666 24.842 ;
      RECT 11.614 26.006 11.666 26.042 ;
      RECT 11.614 27.206 11.666 27.242 ;
      RECT 11.614 28.406 11.666 28.442 ;
      RECT 11.614 29.606 11.666 29.642 ;
      RECT 11.614 30.806 11.666 30.842 ;
      RECT 11.614 32.622 11.666 32.658 ;
      RECT 11.614 32.862 11.666 32.898 ;
      RECT 11.614 38.622 11.666 38.658 ;
      RECT 11.614 38.862 11.666 38.898 ;
      RECT 11.614 39.926 11.666 39.962 ;
      RECT 11.614 41.126 11.666 41.162 ;
      RECT 11.614 42.326 11.666 42.362 ;
      RECT 11.614 43.526 11.666 43.562 ;
      RECT 11.614 44.726 11.666 44.762 ;
      RECT 11.614 45.926 11.666 45.962 ;
      RECT 11.614 47.126 11.666 47.162 ;
      RECT 11.614 48.326 11.666 48.362 ;
      RECT 11.614 49.526 11.666 49.562 ;
      RECT 11.614 50.726 11.666 50.762 ;
      RECT 11.614 51.926 11.666 51.962 ;
      RECT 11.614 53.126 11.666 53.162 ;
      RECT 11.614 54.326 11.666 54.362 ;
      RECT 11.614 55.526 11.666 55.562 ;
      RECT 11.614 56.726 11.666 56.762 ;
      RECT 11.614 57.926 11.666 57.962 ;
      RECT 11.614 59.126 11.666 59.162 ;
      RECT 11.614 60.326 11.666 60.362 ;
      RECT 11.614 61.526 11.666 61.562 ;
      RECT 11.614 62.726 11.666 62.762 ;
      RECT 11.614 63.926 11.666 63.962 ;
      RECT 11.614 65.126 11.666 65.162 ;
      RECT 11.614 66.326 11.666 66.362 ;
      RECT 11.614 67.526 11.666 67.562 ;
      RECT 11.614 68.726 11.666 68.762 ;
      RECT 11.614 69.926 11.666 69.962 ;
      RECT 11.614 71.126 11.666 71.162 ;
      RECT 11.694 1.558 11.746 1.594 ;
      RECT 11.694 2.758 11.746 2.794 ;
      RECT 11.694 3.958 11.746 3.994 ;
      RECT 11.694 5.158 11.746 5.194 ;
      RECT 11.694 6.358 11.746 6.394 ;
      RECT 11.694 7.558 11.746 7.594 ;
      RECT 11.694 8.758 11.746 8.794 ;
      RECT 11.694 9.958 11.746 9.994 ;
      RECT 11.694 11.158 11.746 11.194 ;
      RECT 11.694 12.358 11.746 12.394 ;
      RECT 11.694 13.558 11.746 13.594 ;
      RECT 11.694 14.758 11.746 14.794 ;
      RECT 11.694 15.958 11.746 15.994 ;
      RECT 11.694 17.158 11.746 17.194 ;
      RECT 11.694 18.358 11.746 18.394 ;
      RECT 11.694 19.558 11.746 19.594 ;
      RECT 11.694 20.758 11.746 20.794 ;
      RECT 11.694 21.958 11.746 21.994 ;
      RECT 11.694 23.158 11.746 23.194 ;
      RECT 11.694 24.358 11.746 24.394 ;
      RECT 11.694 25.558 11.746 25.594 ;
      RECT 11.694 26.758 11.746 26.794 ;
      RECT 11.694 27.958 11.746 27.994 ;
      RECT 11.694 29.158 11.746 29.194 ;
      RECT 11.694 30.358 11.746 30.394 ;
      RECT 11.694 31.558 11.746 31.594 ;
      RECT 11.694 33.342 11.746 33.378 ;
      RECT 11.694 33.582 11.746 33.618 ;
      RECT 11.694 37.902 11.746 37.938 ;
      RECT 11.694 38.142 11.746 38.178 ;
      RECT 11.694 40.678 11.746 40.714 ;
      RECT 11.694 41.878 11.746 41.914 ;
      RECT 11.694 43.078 11.746 43.114 ;
      RECT 11.694 44.278 11.746 44.314 ;
      RECT 11.694 45.478 11.746 45.514 ;
      RECT 11.694 46.678 11.746 46.714 ;
      RECT 11.694 47.878 11.746 47.914 ;
      RECT 11.694 49.078 11.746 49.114 ;
      RECT 11.694 50.278 11.746 50.314 ;
      RECT 11.694 51.478 11.746 51.514 ;
      RECT 11.694 52.678 11.746 52.714 ;
      RECT 11.694 53.878 11.746 53.914 ;
      RECT 11.694 55.078 11.746 55.114 ;
      RECT 11.694 56.278 11.746 56.314 ;
      RECT 11.694 57.478 11.746 57.514 ;
      RECT 11.694 58.678 11.746 58.714 ;
      RECT 11.694 59.878 11.746 59.914 ;
      RECT 11.694 61.078 11.746 61.114 ;
      RECT 11.694 62.278 11.746 62.314 ;
      RECT 11.694 63.478 11.746 63.514 ;
      RECT 11.694 64.678 11.746 64.714 ;
      RECT 11.694 65.878 11.746 65.914 ;
      RECT 11.694 67.078 11.746 67.114 ;
      RECT 11.694 68.278 11.746 68.314 ;
      RECT 11.694 69.478 11.746 69.514 ;
      RECT 11.694 70.678 11.746 70.714 ;
      RECT 11.694 71.878 11.746 71.914 ;
      RECT 11.774 0.281 11.826 0.317 ;
      RECT 11.774 72.403 11.826 72.439 ;
      RECT 11.854 0.806 11.906 0.842 ;
      RECT 11.854 2.006 11.906 2.042 ;
      RECT 11.854 3.206 11.906 3.242 ;
      RECT 11.854 4.406 11.906 4.442 ;
      RECT 11.854 5.606 11.906 5.642 ;
      RECT 11.854 6.806 11.906 6.842 ;
      RECT 11.854 8.006 11.906 8.042 ;
      RECT 11.854 9.206 11.906 9.242 ;
      RECT 11.854 10.406 11.906 10.442 ;
      RECT 11.854 11.606 11.906 11.642 ;
      RECT 11.854 12.806 11.906 12.842 ;
      RECT 11.854 14.006 11.906 14.042 ;
      RECT 11.854 15.206 11.906 15.242 ;
      RECT 11.854 16.406 11.906 16.442 ;
      RECT 11.854 17.606 11.906 17.642 ;
      RECT 11.854 18.806 11.906 18.842 ;
      RECT 11.854 20.006 11.906 20.042 ;
      RECT 11.854 21.206 11.906 21.242 ;
      RECT 11.854 22.406 11.906 22.442 ;
      RECT 11.854 23.606 11.906 23.642 ;
      RECT 11.854 24.806 11.906 24.842 ;
      RECT 11.854 26.006 11.906 26.042 ;
      RECT 11.854 27.206 11.906 27.242 ;
      RECT 11.854 28.406 11.906 28.442 ;
      RECT 11.854 29.606 11.906 29.642 ;
      RECT 11.854 30.806 11.906 30.842 ;
      RECT 11.854 32.622 11.906 32.658 ;
      RECT 11.854 32.862 11.906 32.898 ;
      RECT 11.854 38.622 11.906 38.658 ;
      RECT 11.854 38.862 11.906 38.898 ;
      RECT 11.854 39.926 11.906 39.962 ;
      RECT 11.854 41.126 11.906 41.162 ;
      RECT 11.854 42.326 11.906 42.362 ;
      RECT 11.854 43.526 11.906 43.562 ;
      RECT 11.854 44.726 11.906 44.762 ;
      RECT 11.854 45.926 11.906 45.962 ;
      RECT 11.854 47.126 11.906 47.162 ;
      RECT 11.854 48.326 11.906 48.362 ;
      RECT 11.854 49.526 11.906 49.562 ;
      RECT 11.854 50.726 11.906 50.762 ;
      RECT 11.854 51.926 11.906 51.962 ;
      RECT 11.854 53.126 11.906 53.162 ;
      RECT 11.854 54.326 11.906 54.362 ;
      RECT 11.854 55.526 11.906 55.562 ;
      RECT 11.854 56.726 11.906 56.762 ;
      RECT 11.854 57.926 11.906 57.962 ;
      RECT 11.854 59.126 11.906 59.162 ;
      RECT 11.854 60.326 11.906 60.362 ;
      RECT 11.854 61.526 11.906 61.562 ;
      RECT 11.854 62.726 11.906 62.762 ;
      RECT 11.854 63.926 11.906 63.962 ;
      RECT 11.854 65.126 11.906 65.162 ;
      RECT 11.854 66.326 11.906 66.362 ;
      RECT 11.854 67.526 11.906 67.562 ;
      RECT 11.854 68.726 11.906 68.762 ;
      RECT 11.854 69.926 11.906 69.962 ;
      RECT 11.854 71.126 11.906 71.162 ;
      RECT 11.934 1.558 11.986 1.594 ;
      RECT 11.934 2.758 11.986 2.794 ;
      RECT 11.934 3.958 11.986 3.994 ;
      RECT 11.934 5.158 11.986 5.194 ;
      RECT 11.934 6.358 11.986 6.394 ;
      RECT 11.934 7.558 11.986 7.594 ;
      RECT 11.934 8.758 11.986 8.794 ;
      RECT 11.934 9.958 11.986 9.994 ;
      RECT 11.934 11.158 11.986 11.194 ;
      RECT 11.934 12.358 11.986 12.394 ;
      RECT 11.934 13.558 11.986 13.594 ;
      RECT 11.934 14.758 11.986 14.794 ;
      RECT 11.934 15.958 11.986 15.994 ;
      RECT 11.934 17.158 11.986 17.194 ;
      RECT 11.934 18.358 11.986 18.394 ;
      RECT 11.934 19.558 11.986 19.594 ;
      RECT 11.934 20.758 11.986 20.794 ;
      RECT 11.934 21.958 11.986 21.994 ;
      RECT 11.934 23.158 11.986 23.194 ;
      RECT 11.934 24.358 11.986 24.394 ;
      RECT 11.934 25.558 11.986 25.594 ;
      RECT 11.934 26.758 11.986 26.794 ;
      RECT 11.934 27.958 11.986 27.994 ;
      RECT 11.934 29.158 11.986 29.194 ;
      RECT 11.934 30.358 11.986 30.394 ;
      RECT 11.934 31.558 11.986 31.594 ;
      RECT 11.934 33.342 11.986 33.378 ;
      RECT 11.934 33.582 11.986 33.618 ;
      RECT 11.934 37.902 11.986 37.938 ;
      RECT 11.934 38.142 11.986 38.178 ;
      RECT 11.934 40.678 11.986 40.714 ;
      RECT 11.934 41.878 11.986 41.914 ;
      RECT 11.934 43.078 11.986 43.114 ;
      RECT 11.934 44.278 11.986 44.314 ;
      RECT 11.934 45.478 11.986 45.514 ;
      RECT 11.934 46.678 11.986 46.714 ;
      RECT 11.934 47.878 11.986 47.914 ;
      RECT 11.934 49.078 11.986 49.114 ;
      RECT 11.934 50.278 11.986 50.314 ;
      RECT 11.934 51.478 11.986 51.514 ;
      RECT 11.934 52.678 11.986 52.714 ;
      RECT 11.934 53.878 11.986 53.914 ;
      RECT 11.934 55.078 11.986 55.114 ;
      RECT 11.934 56.278 11.986 56.314 ;
      RECT 11.934 57.478 11.986 57.514 ;
      RECT 11.934 58.678 11.986 58.714 ;
      RECT 11.934 59.878 11.986 59.914 ;
      RECT 11.934 61.078 11.986 61.114 ;
      RECT 11.934 62.278 11.986 62.314 ;
      RECT 11.934 63.478 11.986 63.514 ;
      RECT 11.934 64.678 11.986 64.714 ;
      RECT 11.934 65.878 11.986 65.914 ;
      RECT 11.934 67.078 11.986 67.114 ;
      RECT 11.934 68.278 11.986 68.314 ;
      RECT 11.934 69.478 11.986 69.514 ;
      RECT 11.934 70.678 11.986 70.714 ;
      RECT 11.934 71.878 11.986 71.914 ;
      RECT 12.014 0.806 12.066 0.842 ;
      RECT 12.014 2.006 12.066 2.042 ;
      RECT 12.014 3.206 12.066 3.242 ;
      RECT 12.014 4.406 12.066 4.442 ;
      RECT 12.014 5.606 12.066 5.642 ;
      RECT 12.014 6.806 12.066 6.842 ;
      RECT 12.014 8.006 12.066 8.042 ;
      RECT 12.014 9.206 12.066 9.242 ;
      RECT 12.014 10.406 12.066 10.442 ;
      RECT 12.014 11.606 12.066 11.642 ;
      RECT 12.014 12.806 12.066 12.842 ;
      RECT 12.014 14.006 12.066 14.042 ;
      RECT 12.014 15.206 12.066 15.242 ;
      RECT 12.014 16.406 12.066 16.442 ;
      RECT 12.014 17.606 12.066 17.642 ;
      RECT 12.014 18.806 12.066 18.842 ;
      RECT 12.014 20.006 12.066 20.042 ;
      RECT 12.014 21.206 12.066 21.242 ;
      RECT 12.014 22.406 12.066 22.442 ;
      RECT 12.014 23.606 12.066 23.642 ;
      RECT 12.014 24.806 12.066 24.842 ;
      RECT 12.014 26.006 12.066 26.042 ;
      RECT 12.014 27.206 12.066 27.242 ;
      RECT 12.014 28.406 12.066 28.442 ;
      RECT 12.014 29.606 12.066 29.642 ;
      RECT 12.014 30.806 12.066 30.842 ;
      RECT 12.014 32.622 12.066 32.658 ;
      RECT 12.014 32.862 12.066 32.898 ;
      RECT 12.014 38.622 12.066 38.658 ;
      RECT 12.014 38.862 12.066 38.898 ;
      RECT 12.014 39.926 12.066 39.962 ;
      RECT 12.014 41.126 12.066 41.162 ;
      RECT 12.014 42.326 12.066 42.362 ;
      RECT 12.014 43.526 12.066 43.562 ;
      RECT 12.014 44.726 12.066 44.762 ;
      RECT 12.014 45.926 12.066 45.962 ;
      RECT 12.014 47.126 12.066 47.162 ;
      RECT 12.014 48.326 12.066 48.362 ;
      RECT 12.014 49.526 12.066 49.562 ;
      RECT 12.014 50.726 12.066 50.762 ;
      RECT 12.014 51.926 12.066 51.962 ;
      RECT 12.014 53.126 12.066 53.162 ;
      RECT 12.014 54.326 12.066 54.362 ;
      RECT 12.014 55.526 12.066 55.562 ;
      RECT 12.014 56.726 12.066 56.762 ;
      RECT 12.014 57.926 12.066 57.962 ;
      RECT 12.014 59.126 12.066 59.162 ;
      RECT 12.014 60.326 12.066 60.362 ;
      RECT 12.014 61.526 12.066 61.562 ;
      RECT 12.014 62.726 12.066 62.762 ;
      RECT 12.014 63.926 12.066 63.962 ;
      RECT 12.014 65.126 12.066 65.162 ;
      RECT 12.014 66.326 12.066 66.362 ;
      RECT 12.014 67.526 12.066 67.562 ;
      RECT 12.014 68.726 12.066 68.762 ;
      RECT 12.014 69.926 12.066 69.962 ;
      RECT 12.014 71.126 12.066 71.162 ;
      RECT 12.094 1.558 12.146 1.594 ;
      RECT 12.094 2.758 12.146 2.794 ;
      RECT 12.094 3.958 12.146 3.994 ;
      RECT 12.094 5.158 12.146 5.194 ;
      RECT 12.094 6.358 12.146 6.394 ;
      RECT 12.094 7.558 12.146 7.594 ;
      RECT 12.094 8.758 12.146 8.794 ;
      RECT 12.094 9.958 12.146 9.994 ;
      RECT 12.094 11.158 12.146 11.194 ;
      RECT 12.094 12.358 12.146 12.394 ;
      RECT 12.094 13.558 12.146 13.594 ;
      RECT 12.094 14.758 12.146 14.794 ;
      RECT 12.094 15.958 12.146 15.994 ;
      RECT 12.094 17.158 12.146 17.194 ;
      RECT 12.094 18.358 12.146 18.394 ;
      RECT 12.094 19.558 12.146 19.594 ;
      RECT 12.094 20.758 12.146 20.794 ;
      RECT 12.094 21.958 12.146 21.994 ;
      RECT 12.094 23.158 12.146 23.194 ;
      RECT 12.094 24.358 12.146 24.394 ;
      RECT 12.094 25.558 12.146 25.594 ;
      RECT 12.094 26.758 12.146 26.794 ;
      RECT 12.094 27.958 12.146 27.994 ;
      RECT 12.094 29.158 12.146 29.194 ;
      RECT 12.094 30.358 12.146 30.394 ;
      RECT 12.094 31.558 12.146 31.594 ;
      RECT 12.094 33.342 12.146 33.378 ;
      RECT 12.094 33.582 12.146 33.618 ;
      RECT 12.094 37.902 12.146 37.938 ;
      RECT 12.094 38.142 12.146 38.178 ;
      RECT 12.094 40.678 12.146 40.714 ;
      RECT 12.094 41.878 12.146 41.914 ;
      RECT 12.094 43.078 12.146 43.114 ;
      RECT 12.094 44.278 12.146 44.314 ;
      RECT 12.094 45.478 12.146 45.514 ;
      RECT 12.094 46.678 12.146 46.714 ;
      RECT 12.094 47.878 12.146 47.914 ;
      RECT 12.094 49.078 12.146 49.114 ;
      RECT 12.094 50.278 12.146 50.314 ;
      RECT 12.094 51.478 12.146 51.514 ;
      RECT 12.094 52.678 12.146 52.714 ;
      RECT 12.094 53.878 12.146 53.914 ;
      RECT 12.094 55.078 12.146 55.114 ;
      RECT 12.094 56.278 12.146 56.314 ;
      RECT 12.094 57.478 12.146 57.514 ;
      RECT 12.094 58.678 12.146 58.714 ;
      RECT 12.094 59.878 12.146 59.914 ;
      RECT 12.094 61.078 12.146 61.114 ;
      RECT 12.094 62.278 12.146 62.314 ;
      RECT 12.094 63.478 12.146 63.514 ;
      RECT 12.094 64.678 12.146 64.714 ;
      RECT 12.094 65.878 12.146 65.914 ;
      RECT 12.094 67.078 12.146 67.114 ;
      RECT 12.094 68.278 12.146 68.314 ;
      RECT 12.094 69.478 12.146 69.514 ;
      RECT 12.094 70.678 12.146 70.714 ;
      RECT 12.094 71.878 12.146 71.914 ;
      RECT 12.174 0.281 12.226 0.317 ;
      RECT 12.174 72.403 12.226 72.439 ;
      RECT 12.254 0.806 12.306 0.842 ;
      RECT 12.254 2.006 12.306 2.042 ;
      RECT 12.254 3.206 12.306 3.242 ;
      RECT 12.254 4.406 12.306 4.442 ;
      RECT 12.254 5.606 12.306 5.642 ;
      RECT 12.254 6.806 12.306 6.842 ;
      RECT 12.254 8.006 12.306 8.042 ;
      RECT 12.254 9.206 12.306 9.242 ;
      RECT 12.254 10.406 12.306 10.442 ;
      RECT 12.254 11.606 12.306 11.642 ;
      RECT 12.254 12.806 12.306 12.842 ;
      RECT 12.254 14.006 12.306 14.042 ;
      RECT 12.254 15.206 12.306 15.242 ;
      RECT 12.254 16.406 12.306 16.442 ;
      RECT 12.254 17.606 12.306 17.642 ;
      RECT 12.254 18.806 12.306 18.842 ;
      RECT 12.254 20.006 12.306 20.042 ;
      RECT 12.254 21.206 12.306 21.242 ;
      RECT 12.254 22.406 12.306 22.442 ;
      RECT 12.254 23.606 12.306 23.642 ;
      RECT 12.254 24.806 12.306 24.842 ;
      RECT 12.254 26.006 12.306 26.042 ;
      RECT 12.254 27.206 12.306 27.242 ;
      RECT 12.254 28.406 12.306 28.442 ;
      RECT 12.254 29.606 12.306 29.642 ;
      RECT 12.254 30.806 12.306 30.842 ;
      RECT 12.254 32.622 12.306 32.658 ;
      RECT 12.254 32.862 12.306 32.898 ;
      RECT 12.254 34.302 12.306 34.338 ;
      RECT 12.254 34.782 12.306 34.818 ;
      RECT 12.254 36.702 12.306 36.738 ;
      RECT 12.254 37.182 12.306 37.218 ;
      RECT 12.254 38.622 12.306 38.658 ;
      RECT 12.254 38.862 12.306 38.898 ;
      RECT 12.254 39.926 12.306 39.962 ;
      RECT 12.254 41.126 12.306 41.162 ;
      RECT 12.254 42.326 12.306 42.362 ;
      RECT 12.254 43.526 12.306 43.562 ;
      RECT 12.254 44.726 12.306 44.762 ;
      RECT 12.254 45.926 12.306 45.962 ;
      RECT 12.254 47.126 12.306 47.162 ;
      RECT 12.254 48.326 12.306 48.362 ;
      RECT 12.254 49.526 12.306 49.562 ;
      RECT 12.254 50.726 12.306 50.762 ;
      RECT 12.254 51.926 12.306 51.962 ;
      RECT 12.254 53.126 12.306 53.162 ;
      RECT 12.254 54.326 12.306 54.362 ;
      RECT 12.254 55.526 12.306 55.562 ;
      RECT 12.254 56.726 12.306 56.762 ;
      RECT 12.254 57.926 12.306 57.962 ;
      RECT 12.254 59.126 12.306 59.162 ;
      RECT 12.254 60.326 12.306 60.362 ;
      RECT 12.254 61.526 12.306 61.562 ;
      RECT 12.254 62.726 12.306 62.762 ;
      RECT 12.254 63.926 12.306 63.962 ;
      RECT 12.254 65.126 12.306 65.162 ;
      RECT 12.254 66.326 12.306 66.362 ;
      RECT 12.254 67.526 12.306 67.562 ;
      RECT 12.254 68.726 12.306 68.762 ;
      RECT 12.254 69.926 12.306 69.962 ;
      RECT 12.254 71.126 12.306 71.162 ;
      RECT 12.334 1.558 12.386 1.594 ;
      RECT 12.334 2.758 12.386 2.794 ;
      RECT 12.334 3.958 12.386 3.994 ;
      RECT 12.334 5.158 12.386 5.194 ;
      RECT 12.334 6.358 12.386 6.394 ;
      RECT 12.334 7.558 12.386 7.594 ;
      RECT 12.334 8.758 12.386 8.794 ;
      RECT 12.334 9.958 12.386 9.994 ;
      RECT 12.334 11.158 12.386 11.194 ;
      RECT 12.334 12.358 12.386 12.394 ;
      RECT 12.334 13.558 12.386 13.594 ;
      RECT 12.334 14.758 12.386 14.794 ;
      RECT 12.334 15.958 12.386 15.994 ;
      RECT 12.334 17.158 12.386 17.194 ;
      RECT 12.334 18.358 12.386 18.394 ;
      RECT 12.334 19.558 12.386 19.594 ;
      RECT 12.334 20.758 12.386 20.794 ;
      RECT 12.334 21.958 12.386 21.994 ;
      RECT 12.334 23.158 12.386 23.194 ;
      RECT 12.334 24.358 12.386 24.394 ;
      RECT 12.334 25.558 12.386 25.594 ;
      RECT 12.334 26.758 12.386 26.794 ;
      RECT 12.334 27.958 12.386 27.994 ;
      RECT 12.334 29.158 12.386 29.194 ;
      RECT 12.334 30.358 12.386 30.394 ;
      RECT 12.334 31.558 12.386 31.594 ;
      RECT 12.334 33.342 12.386 33.378 ;
      RECT 12.334 33.582 12.386 33.618 ;
      RECT 12.334 37.902 12.386 37.938 ;
      RECT 12.334 38.142 12.386 38.178 ;
      RECT 12.334 40.678 12.386 40.714 ;
      RECT 12.334 41.878 12.386 41.914 ;
      RECT 12.334 43.078 12.386 43.114 ;
      RECT 12.334 44.278 12.386 44.314 ;
      RECT 12.334 45.478 12.386 45.514 ;
      RECT 12.334 46.678 12.386 46.714 ;
      RECT 12.334 47.878 12.386 47.914 ;
      RECT 12.334 49.078 12.386 49.114 ;
      RECT 12.334 50.278 12.386 50.314 ;
      RECT 12.334 51.478 12.386 51.514 ;
      RECT 12.334 52.678 12.386 52.714 ;
      RECT 12.334 53.878 12.386 53.914 ;
      RECT 12.334 55.078 12.386 55.114 ;
      RECT 12.334 56.278 12.386 56.314 ;
      RECT 12.334 57.478 12.386 57.514 ;
      RECT 12.334 58.678 12.386 58.714 ;
      RECT 12.334 59.878 12.386 59.914 ;
      RECT 12.334 61.078 12.386 61.114 ;
      RECT 12.334 62.278 12.386 62.314 ;
      RECT 12.334 63.478 12.386 63.514 ;
      RECT 12.334 64.678 12.386 64.714 ;
      RECT 12.334 65.878 12.386 65.914 ;
      RECT 12.334 67.078 12.386 67.114 ;
      RECT 12.334 68.278 12.386 68.314 ;
      RECT 12.334 69.478 12.386 69.514 ;
      RECT 12.334 70.678 12.386 70.714 ;
      RECT 12.334 71.878 12.386 71.914 ;
      RECT 12.414 0.806 12.466 0.842 ;
      RECT 12.414 2.006 12.466 2.042 ;
      RECT 12.414 3.206 12.466 3.242 ;
      RECT 12.414 4.406 12.466 4.442 ;
      RECT 12.414 5.606 12.466 5.642 ;
      RECT 12.414 6.806 12.466 6.842 ;
      RECT 12.414 8.006 12.466 8.042 ;
      RECT 12.414 9.206 12.466 9.242 ;
      RECT 12.414 10.406 12.466 10.442 ;
      RECT 12.414 11.606 12.466 11.642 ;
      RECT 12.414 12.806 12.466 12.842 ;
      RECT 12.414 14.006 12.466 14.042 ;
      RECT 12.414 15.206 12.466 15.242 ;
      RECT 12.414 16.406 12.466 16.442 ;
      RECT 12.414 17.606 12.466 17.642 ;
      RECT 12.414 18.806 12.466 18.842 ;
      RECT 12.414 20.006 12.466 20.042 ;
      RECT 12.414 21.206 12.466 21.242 ;
      RECT 12.414 22.406 12.466 22.442 ;
      RECT 12.414 23.606 12.466 23.642 ;
      RECT 12.414 24.806 12.466 24.842 ;
      RECT 12.414 26.006 12.466 26.042 ;
      RECT 12.414 27.206 12.466 27.242 ;
      RECT 12.414 28.406 12.466 28.442 ;
      RECT 12.414 29.606 12.466 29.642 ;
      RECT 12.414 30.806 12.466 30.842 ;
      RECT 12.414 32.622 12.466 32.658 ;
      RECT 12.414 32.862 12.466 32.898 ;
      RECT 12.414 38.622 12.466 38.658 ;
      RECT 12.414 38.862 12.466 38.898 ;
      RECT 12.414 39.926 12.466 39.962 ;
      RECT 12.414 41.126 12.466 41.162 ;
      RECT 12.414 42.326 12.466 42.362 ;
      RECT 12.414 43.526 12.466 43.562 ;
      RECT 12.414 44.726 12.466 44.762 ;
      RECT 12.414 45.926 12.466 45.962 ;
      RECT 12.414 47.126 12.466 47.162 ;
      RECT 12.414 48.326 12.466 48.362 ;
      RECT 12.414 49.526 12.466 49.562 ;
      RECT 12.414 50.726 12.466 50.762 ;
      RECT 12.414 51.926 12.466 51.962 ;
      RECT 12.414 53.126 12.466 53.162 ;
      RECT 12.414 54.326 12.466 54.362 ;
      RECT 12.414 55.526 12.466 55.562 ;
      RECT 12.414 56.726 12.466 56.762 ;
      RECT 12.414 57.926 12.466 57.962 ;
      RECT 12.414 59.126 12.466 59.162 ;
      RECT 12.414 60.326 12.466 60.362 ;
      RECT 12.414 61.526 12.466 61.562 ;
      RECT 12.414 62.726 12.466 62.762 ;
      RECT 12.414 63.926 12.466 63.962 ;
      RECT 12.414 65.126 12.466 65.162 ;
      RECT 12.414 66.326 12.466 66.362 ;
      RECT 12.414 67.526 12.466 67.562 ;
      RECT 12.414 68.726 12.466 68.762 ;
      RECT 12.414 69.926 12.466 69.962 ;
      RECT 12.414 71.126 12.466 71.162 ;
      RECT 12.494 1.558 12.546 1.594 ;
      RECT 12.494 2.758 12.546 2.794 ;
      RECT 12.494 3.958 12.546 3.994 ;
      RECT 12.494 5.158 12.546 5.194 ;
      RECT 12.494 6.358 12.546 6.394 ;
      RECT 12.494 7.558 12.546 7.594 ;
      RECT 12.494 8.758 12.546 8.794 ;
      RECT 12.494 9.958 12.546 9.994 ;
      RECT 12.494 11.158 12.546 11.194 ;
      RECT 12.494 12.358 12.546 12.394 ;
      RECT 12.494 13.558 12.546 13.594 ;
      RECT 12.494 14.758 12.546 14.794 ;
      RECT 12.494 15.958 12.546 15.994 ;
      RECT 12.494 17.158 12.546 17.194 ;
      RECT 12.494 18.358 12.546 18.394 ;
      RECT 12.494 19.558 12.546 19.594 ;
      RECT 12.494 20.758 12.546 20.794 ;
      RECT 12.494 21.958 12.546 21.994 ;
      RECT 12.494 23.158 12.546 23.194 ;
      RECT 12.494 24.358 12.546 24.394 ;
      RECT 12.494 25.558 12.546 25.594 ;
      RECT 12.494 26.758 12.546 26.794 ;
      RECT 12.494 27.958 12.546 27.994 ;
      RECT 12.494 29.158 12.546 29.194 ;
      RECT 12.494 30.358 12.546 30.394 ;
      RECT 12.494 31.558 12.546 31.594 ;
      RECT 12.494 33.342 12.546 33.378 ;
      RECT 12.494 33.582 12.546 33.618 ;
      RECT 12.494 37.902 12.546 37.938 ;
      RECT 12.494 38.142 12.546 38.178 ;
      RECT 12.494 40.678 12.546 40.714 ;
      RECT 12.494 41.878 12.546 41.914 ;
      RECT 12.494 43.078 12.546 43.114 ;
      RECT 12.494 44.278 12.546 44.314 ;
      RECT 12.494 45.478 12.546 45.514 ;
      RECT 12.494 46.678 12.546 46.714 ;
      RECT 12.494 47.878 12.546 47.914 ;
      RECT 12.494 49.078 12.546 49.114 ;
      RECT 12.494 50.278 12.546 50.314 ;
      RECT 12.494 51.478 12.546 51.514 ;
      RECT 12.494 52.678 12.546 52.714 ;
      RECT 12.494 53.878 12.546 53.914 ;
      RECT 12.494 55.078 12.546 55.114 ;
      RECT 12.494 56.278 12.546 56.314 ;
      RECT 12.494 57.478 12.546 57.514 ;
      RECT 12.494 58.678 12.546 58.714 ;
      RECT 12.494 59.878 12.546 59.914 ;
      RECT 12.494 61.078 12.546 61.114 ;
      RECT 12.494 62.278 12.546 62.314 ;
      RECT 12.494 63.478 12.546 63.514 ;
      RECT 12.494 64.678 12.546 64.714 ;
      RECT 12.494 65.878 12.546 65.914 ;
      RECT 12.494 67.078 12.546 67.114 ;
      RECT 12.494 68.278 12.546 68.314 ;
      RECT 12.494 69.478 12.546 69.514 ;
      RECT 12.494 70.678 12.546 70.714 ;
      RECT 12.494 71.878 12.546 71.914 ;
      RECT 12.574 0.281 12.626 0.317 ;
      RECT 12.574 72.403 12.626 72.439 ;
      RECT 12.654 0.806 12.706 0.842 ;
      RECT 12.654 2.006 12.706 2.042 ;
      RECT 12.654 3.206 12.706 3.242 ;
      RECT 12.654 4.406 12.706 4.442 ;
      RECT 12.654 5.606 12.706 5.642 ;
      RECT 12.654 6.806 12.706 6.842 ;
      RECT 12.654 8.006 12.706 8.042 ;
      RECT 12.654 9.206 12.706 9.242 ;
      RECT 12.654 10.406 12.706 10.442 ;
      RECT 12.654 11.606 12.706 11.642 ;
      RECT 12.654 12.806 12.706 12.842 ;
      RECT 12.654 14.006 12.706 14.042 ;
      RECT 12.654 15.206 12.706 15.242 ;
      RECT 12.654 16.406 12.706 16.442 ;
      RECT 12.654 17.606 12.706 17.642 ;
      RECT 12.654 18.806 12.706 18.842 ;
      RECT 12.654 20.006 12.706 20.042 ;
      RECT 12.654 21.206 12.706 21.242 ;
      RECT 12.654 22.406 12.706 22.442 ;
      RECT 12.654 23.606 12.706 23.642 ;
      RECT 12.654 24.806 12.706 24.842 ;
      RECT 12.654 26.006 12.706 26.042 ;
      RECT 12.654 27.206 12.706 27.242 ;
      RECT 12.654 28.406 12.706 28.442 ;
      RECT 12.654 29.606 12.706 29.642 ;
      RECT 12.654 30.806 12.706 30.842 ;
      RECT 12.654 32.622 12.706 32.658 ;
      RECT 12.654 32.862 12.706 32.898 ;
      RECT 12.654 38.622 12.706 38.658 ;
      RECT 12.654 38.862 12.706 38.898 ;
      RECT 12.654 39.926 12.706 39.962 ;
      RECT 12.654 41.126 12.706 41.162 ;
      RECT 12.654 42.326 12.706 42.362 ;
      RECT 12.654 43.526 12.706 43.562 ;
      RECT 12.654 44.726 12.706 44.762 ;
      RECT 12.654 45.926 12.706 45.962 ;
      RECT 12.654 47.126 12.706 47.162 ;
      RECT 12.654 48.326 12.706 48.362 ;
      RECT 12.654 49.526 12.706 49.562 ;
      RECT 12.654 50.726 12.706 50.762 ;
      RECT 12.654 51.926 12.706 51.962 ;
      RECT 12.654 53.126 12.706 53.162 ;
      RECT 12.654 54.326 12.706 54.362 ;
      RECT 12.654 55.526 12.706 55.562 ;
      RECT 12.654 56.726 12.706 56.762 ;
      RECT 12.654 57.926 12.706 57.962 ;
      RECT 12.654 59.126 12.706 59.162 ;
      RECT 12.654 60.326 12.706 60.362 ;
      RECT 12.654 61.526 12.706 61.562 ;
      RECT 12.654 62.726 12.706 62.762 ;
      RECT 12.654 63.926 12.706 63.962 ;
      RECT 12.654 65.126 12.706 65.162 ;
      RECT 12.654 66.326 12.706 66.362 ;
      RECT 12.654 67.526 12.706 67.562 ;
      RECT 12.654 68.726 12.706 68.762 ;
      RECT 12.654 69.926 12.706 69.962 ;
      RECT 12.654 71.126 12.706 71.162 ;
      RECT 12.734 1.558 12.786 1.594 ;
      RECT 12.734 2.758 12.786 2.794 ;
      RECT 12.734 3.958 12.786 3.994 ;
      RECT 12.734 5.158 12.786 5.194 ;
      RECT 12.734 6.358 12.786 6.394 ;
      RECT 12.734 7.558 12.786 7.594 ;
      RECT 12.734 8.758 12.786 8.794 ;
      RECT 12.734 9.958 12.786 9.994 ;
      RECT 12.734 11.158 12.786 11.194 ;
      RECT 12.734 12.358 12.786 12.394 ;
      RECT 12.734 13.558 12.786 13.594 ;
      RECT 12.734 14.758 12.786 14.794 ;
      RECT 12.734 15.958 12.786 15.994 ;
      RECT 12.734 17.158 12.786 17.194 ;
      RECT 12.734 18.358 12.786 18.394 ;
      RECT 12.734 19.558 12.786 19.594 ;
      RECT 12.734 20.758 12.786 20.794 ;
      RECT 12.734 21.958 12.786 21.994 ;
      RECT 12.734 23.158 12.786 23.194 ;
      RECT 12.734 24.358 12.786 24.394 ;
      RECT 12.734 25.558 12.786 25.594 ;
      RECT 12.734 26.758 12.786 26.794 ;
      RECT 12.734 27.958 12.786 27.994 ;
      RECT 12.734 29.158 12.786 29.194 ;
      RECT 12.734 30.358 12.786 30.394 ;
      RECT 12.734 31.558 12.786 31.594 ;
      RECT 12.734 33.342 12.786 33.378 ;
      RECT 12.734 33.582 12.786 33.618 ;
      RECT 12.734 37.902 12.786 37.938 ;
      RECT 12.734 38.142 12.786 38.178 ;
      RECT 12.734 40.678 12.786 40.714 ;
      RECT 12.734 41.878 12.786 41.914 ;
      RECT 12.734 43.078 12.786 43.114 ;
      RECT 12.734 44.278 12.786 44.314 ;
      RECT 12.734 45.478 12.786 45.514 ;
      RECT 12.734 46.678 12.786 46.714 ;
      RECT 12.734 47.878 12.786 47.914 ;
      RECT 12.734 49.078 12.786 49.114 ;
      RECT 12.734 50.278 12.786 50.314 ;
      RECT 12.734 51.478 12.786 51.514 ;
      RECT 12.734 52.678 12.786 52.714 ;
      RECT 12.734 53.878 12.786 53.914 ;
      RECT 12.734 55.078 12.786 55.114 ;
      RECT 12.734 56.278 12.786 56.314 ;
      RECT 12.734 57.478 12.786 57.514 ;
      RECT 12.734 58.678 12.786 58.714 ;
      RECT 12.734 59.878 12.786 59.914 ;
      RECT 12.734 61.078 12.786 61.114 ;
      RECT 12.734 62.278 12.786 62.314 ;
      RECT 12.734 63.478 12.786 63.514 ;
      RECT 12.734 64.678 12.786 64.714 ;
      RECT 12.734 65.878 12.786 65.914 ;
      RECT 12.734 67.078 12.786 67.114 ;
      RECT 12.734 68.278 12.786 68.314 ;
      RECT 12.734 69.478 12.786 69.514 ;
      RECT 12.734 70.678 12.786 70.714 ;
      RECT 12.734 71.878 12.786 71.914 ;
      RECT 12.814 0.806 12.866 0.842 ;
      RECT 12.814 2.006 12.866 2.042 ;
      RECT 12.814 3.206 12.866 3.242 ;
      RECT 12.814 4.406 12.866 4.442 ;
      RECT 12.814 5.606 12.866 5.642 ;
      RECT 12.814 6.806 12.866 6.842 ;
      RECT 12.814 8.006 12.866 8.042 ;
      RECT 12.814 9.206 12.866 9.242 ;
      RECT 12.814 10.406 12.866 10.442 ;
      RECT 12.814 11.606 12.866 11.642 ;
      RECT 12.814 12.806 12.866 12.842 ;
      RECT 12.814 14.006 12.866 14.042 ;
      RECT 12.814 15.206 12.866 15.242 ;
      RECT 12.814 16.406 12.866 16.442 ;
      RECT 12.814 17.606 12.866 17.642 ;
      RECT 12.814 18.806 12.866 18.842 ;
      RECT 12.814 20.006 12.866 20.042 ;
      RECT 12.814 21.206 12.866 21.242 ;
      RECT 12.814 22.406 12.866 22.442 ;
      RECT 12.814 23.606 12.866 23.642 ;
      RECT 12.814 24.806 12.866 24.842 ;
      RECT 12.814 26.006 12.866 26.042 ;
      RECT 12.814 27.206 12.866 27.242 ;
      RECT 12.814 28.406 12.866 28.442 ;
      RECT 12.814 29.606 12.866 29.642 ;
      RECT 12.814 30.806 12.866 30.842 ;
      RECT 12.814 32.622 12.866 32.658 ;
      RECT 12.814 32.862 12.866 32.898 ;
      RECT 12.814 38.622 12.866 38.658 ;
      RECT 12.814 38.862 12.866 38.898 ;
      RECT 12.814 39.926 12.866 39.962 ;
      RECT 12.814 41.126 12.866 41.162 ;
      RECT 12.814 42.326 12.866 42.362 ;
      RECT 12.814 43.526 12.866 43.562 ;
      RECT 12.814 44.726 12.866 44.762 ;
      RECT 12.814 45.926 12.866 45.962 ;
      RECT 12.814 47.126 12.866 47.162 ;
      RECT 12.814 48.326 12.866 48.362 ;
      RECT 12.814 49.526 12.866 49.562 ;
      RECT 12.814 50.726 12.866 50.762 ;
      RECT 12.814 51.926 12.866 51.962 ;
      RECT 12.814 53.126 12.866 53.162 ;
      RECT 12.814 54.326 12.866 54.362 ;
      RECT 12.814 55.526 12.866 55.562 ;
      RECT 12.814 56.726 12.866 56.762 ;
      RECT 12.814 57.926 12.866 57.962 ;
      RECT 12.814 59.126 12.866 59.162 ;
      RECT 12.814 60.326 12.866 60.362 ;
      RECT 12.814 61.526 12.866 61.562 ;
      RECT 12.814 62.726 12.866 62.762 ;
      RECT 12.814 63.926 12.866 63.962 ;
      RECT 12.814 65.126 12.866 65.162 ;
      RECT 12.814 66.326 12.866 66.362 ;
      RECT 12.814 67.526 12.866 67.562 ;
      RECT 12.814 68.726 12.866 68.762 ;
      RECT 12.814 69.926 12.866 69.962 ;
      RECT 12.814 71.126 12.866 71.162 ;
      RECT 12.894 1.558 12.946 1.594 ;
      RECT 12.894 2.758 12.946 2.794 ;
      RECT 12.894 3.958 12.946 3.994 ;
      RECT 12.894 5.158 12.946 5.194 ;
      RECT 12.894 6.358 12.946 6.394 ;
      RECT 12.894 7.558 12.946 7.594 ;
      RECT 12.894 8.758 12.946 8.794 ;
      RECT 12.894 9.958 12.946 9.994 ;
      RECT 12.894 11.158 12.946 11.194 ;
      RECT 12.894 12.358 12.946 12.394 ;
      RECT 12.894 13.558 12.946 13.594 ;
      RECT 12.894 14.758 12.946 14.794 ;
      RECT 12.894 15.958 12.946 15.994 ;
      RECT 12.894 17.158 12.946 17.194 ;
      RECT 12.894 18.358 12.946 18.394 ;
      RECT 12.894 19.558 12.946 19.594 ;
      RECT 12.894 20.758 12.946 20.794 ;
      RECT 12.894 21.958 12.946 21.994 ;
      RECT 12.894 23.158 12.946 23.194 ;
      RECT 12.894 24.358 12.946 24.394 ;
      RECT 12.894 25.558 12.946 25.594 ;
      RECT 12.894 26.758 12.946 26.794 ;
      RECT 12.894 27.958 12.946 27.994 ;
      RECT 12.894 29.158 12.946 29.194 ;
      RECT 12.894 30.358 12.946 30.394 ;
      RECT 12.894 31.558 12.946 31.594 ;
      RECT 12.894 33.342 12.946 33.378 ;
      RECT 12.894 33.582 12.946 33.618 ;
      RECT 12.894 37.902 12.946 37.938 ;
      RECT 12.894 38.142 12.946 38.178 ;
      RECT 12.894 40.678 12.946 40.714 ;
      RECT 12.894 41.878 12.946 41.914 ;
      RECT 12.894 43.078 12.946 43.114 ;
      RECT 12.894 44.278 12.946 44.314 ;
      RECT 12.894 45.478 12.946 45.514 ;
      RECT 12.894 46.678 12.946 46.714 ;
      RECT 12.894 47.878 12.946 47.914 ;
      RECT 12.894 49.078 12.946 49.114 ;
      RECT 12.894 50.278 12.946 50.314 ;
      RECT 12.894 51.478 12.946 51.514 ;
      RECT 12.894 52.678 12.946 52.714 ;
      RECT 12.894 53.878 12.946 53.914 ;
      RECT 12.894 55.078 12.946 55.114 ;
      RECT 12.894 56.278 12.946 56.314 ;
      RECT 12.894 57.478 12.946 57.514 ;
      RECT 12.894 58.678 12.946 58.714 ;
      RECT 12.894 59.878 12.946 59.914 ;
      RECT 12.894 61.078 12.946 61.114 ;
      RECT 12.894 62.278 12.946 62.314 ;
      RECT 12.894 63.478 12.946 63.514 ;
      RECT 12.894 64.678 12.946 64.714 ;
      RECT 12.894 65.878 12.946 65.914 ;
      RECT 12.894 67.078 12.946 67.114 ;
      RECT 12.894 68.278 12.946 68.314 ;
      RECT 12.894 69.478 12.946 69.514 ;
      RECT 12.894 70.678 12.946 70.714 ;
      RECT 12.894 71.878 12.946 71.914 ;
      RECT 12.974 0.281 13.026 0.317 ;
      RECT 12.974 72.403 13.026 72.439 ;
      RECT 13.054 0.806 13.106 0.842 ;
      RECT 13.054 2.006 13.106 2.042 ;
      RECT 13.054 3.206 13.106 3.242 ;
      RECT 13.054 4.406 13.106 4.442 ;
      RECT 13.054 5.606 13.106 5.642 ;
      RECT 13.054 6.806 13.106 6.842 ;
      RECT 13.054 8.006 13.106 8.042 ;
      RECT 13.054 9.206 13.106 9.242 ;
      RECT 13.054 10.406 13.106 10.442 ;
      RECT 13.054 11.606 13.106 11.642 ;
      RECT 13.054 12.806 13.106 12.842 ;
      RECT 13.054 14.006 13.106 14.042 ;
      RECT 13.054 15.206 13.106 15.242 ;
      RECT 13.054 16.406 13.106 16.442 ;
      RECT 13.054 17.606 13.106 17.642 ;
      RECT 13.054 18.806 13.106 18.842 ;
      RECT 13.054 20.006 13.106 20.042 ;
      RECT 13.054 21.206 13.106 21.242 ;
      RECT 13.054 22.406 13.106 22.442 ;
      RECT 13.054 23.606 13.106 23.642 ;
      RECT 13.054 24.806 13.106 24.842 ;
      RECT 13.054 26.006 13.106 26.042 ;
      RECT 13.054 27.206 13.106 27.242 ;
      RECT 13.054 28.406 13.106 28.442 ;
      RECT 13.054 29.606 13.106 29.642 ;
      RECT 13.054 30.806 13.106 30.842 ;
      RECT 13.054 32.622 13.106 32.658 ;
      RECT 13.054 32.862 13.106 32.898 ;
      RECT 13.054 34.302 13.106 34.338 ;
      RECT 13.054 34.782 13.106 34.818 ;
      RECT 13.054 36.702 13.106 36.738 ;
      RECT 13.054 37.182 13.106 37.218 ;
      RECT 13.054 38.622 13.106 38.658 ;
      RECT 13.054 38.862 13.106 38.898 ;
      RECT 13.054 39.926 13.106 39.962 ;
      RECT 13.054 41.126 13.106 41.162 ;
      RECT 13.054 42.326 13.106 42.362 ;
      RECT 13.054 43.526 13.106 43.562 ;
      RECT 13.054 44.726 13.106 44.762 ;
      RECT 13.054 45.926 13.106 45.962 ;
      RECT 13.054 47.126 13.106 47.162 ;
      RECT 13.054 48.326 13.106 48.362 ;
      RECT 13.054 49.526 13.106 49.562 ;
      RECT 13.054 50.726 13.106 50.762 ;
      RECT 13.054 51.926 13.106 51.962 ;
      RECT 13.054 53.126 13.106 53.162 ;
      RECT 13.054 54.326 13.106 54.362 ;
      RECT 13.054 55.526 13.106 55.562 ;
      RECT 13.054 56.726 13.106 56.762 ;
      RECT 13.054 57.926 13.106 57.962 ;
      RECT 13.054 59.126 13.106 59.162 ;
      RECT 13.054 60.326 13.106 60.362 ;
      RECT 13.054 61.526 13.106 61.562 ;
      RECT 13.054 62.726 13.106 62.762 ;
      RECT 13.054 63.926 13.106 63.962 ;
      RECT 13.054 65.126 13.106 65.162 ;
      RECT 13.054 66.326 13.106 66.362 ;
      RECT 13.054 67.526 13.106 67.562 ;
      RECT 13.054 68.726 13.106 68.762 ;
      RECT 13.054 69.926 13.106 69.962 ;
      RECT 13.054 71.126 13.106 71.162 ;
      RECT 13.134 1.558 13.186 1.594 ;
      RECT 13.134 2.758 13.186 2.794 ;
      RECT 13.134 3.958 13.186 3.994 ;
      RECT 13.134 5.158 13.186 5.194 ;
      RECT 13.134 6.358 13.186 6.394 ;
      RECT 13.134 7.558 13.186 7.594 ;
      RECT 13.134 8.758 13.186 8.794 ;
      RECT 13.134 9.958 13.186 9.994 ;
      RECT 13.134 11.158 13.186 11.194 ;
      RECT 13.134 12.358 13.186 12.394 ;
      RECT 13.134 13.558 13.186 13.594 ;
      RECT 13.134 14.758 13.186 14.794 ;
      RECT 13.134 15.958 13.186 15.994 ;
      RECT 13.134 17.158 13.186 17.194 ;
      RECT 13.134 18.358 13.186 18.394 ;
      RECT 13.134 19.558 13.186 19.594 ;
      RECT 13.134 20.758 13.186 20.794 ;
      RECT 13.134 21.958 13.186 21.994 ;
      RECT 13.134 23.158 13.186 23.194 ;
      RECT 13.134 24.358 13.186 24.394 ;
      RECT 13.134 25.558 13.186 25.594 ;
      RECT 13.134 26.758 13.186 26.794 ;
      RECT 13.134 27.958 13.186 27.994 ;
      RECT 13.134 29.158 13.186 29.194 ;
      RECT 13.134 30.358 13.186 30.394 ;
      RECT 13.134 31.558 13.186 31.594 ;
      RECT 13.134 33.342 13.186 33.378 ;
      RECT 13.134 33.582 13.186 33.618 ;
      RECT 13.134 37.902 13.186 37.938 ;
      RECT 13.134 38.142 13.186 38.178 ;
      RECT 13.134 40.678 13.186 40.714 ;
      RECT 13.134 41.878 13.186 41.914 ;
      RECT 13.134 43.078 13.186 43.114 ;
      RECT 13.134 44.278 13.186 44.314 ;
      RECT 13.134 45.478 13.186 45.514 ;
      RECT 13.134 46.678 13.186 46.714 ;
      RECT 13.134 47.878 13.186 47.914 ;
      RECT 13.134 49.078 13.186 49.114 ;
      RECT 13.134 50.278 13.186 50.314 ;
      RECT 13.134 51.478 13.186 51.514 ;
      RECT 13.134 52.678 13.186 52.714 ;
      RECT 13.134 53.878 13.186 53.914 ;
      RECT 13.134 55.078 13.186 55.114 ;
      RECT 13.134 56.278 13.186 56.314 ;
      RECT 13.134 57.478 13.186 57.514 ;
      RECT 13.134 58.678 13.186 58.714 ;
      RECT 13.134 59.878 13.186 59.914 ;
      RECT 13.134 61.078 13.186 61.114 ;
      RECT 13.134 62.278 13.186 62.314 ;
      RECT 13.134 63.478 13.186 63.514 ;
      RECT 13.134 64.678 13.186 64.714 ;
      RECT 13.134 65.878 13.186 65.914 ;
      RECT 13.134 67.078 13.186 67.114 ;
      RECT 13.134 68.278 13.186 68.314 ;
      RECT 13.134 69.478 13.186 69.514 ;
      RECT 13.134 70.678 13.186 70.714 ;
      RECT 13.134 71.878 13.186 71.914 ;
      RECT 13.214 0.806 13.266 0.842 ;
      RECT 13.214 2.006 13.266 2.042 ;
      RECT 13.214 3.206 13.266 3.242 ;
      RECT 13.214 4.406 13.266 4.442 ;
      RECT 13.214 5.606 13.266 5.642 ;
      RECT 13.214 6.806 13.266 6.842 ;
      RECT 13.214 8.006 13.266 8.042 ;
      RECT 13.214 9.206 13.266 9.242 ;
      RECT 13.214 10.406 13.266 10.442 ;
      RECT 13.214 11.606 13.266 11.642 ;
      RECT 13.214 12.806 13.266 12.842 ;
      RECT 13.214 14.006 13.266 14.042 ;
      RECT 13.214 15.206 13.266 15.242 ;
      RECT 13.214 16.406 13.266 16.442 ;
      RECT 13.214 17.606 13.266 17.642 ;
      RECT 13.214 18.806 13.266 18.842 ;
      RECT 13.214 20.006 13.266 20.042 ;
      RECT 13.214 21.206 13.266 21.242 ;
      RECT 13.214 22.406 13.266 22.442 ;
      RECT 13.214 23.606 13.266 23.642 ;
      RECT 13.214 24.806 13.266 24.842 ;
      RECT 13.214 26.006 13.266 26.042 ;
      RECT 13.214 27.206 13.266 27.242 ;
      RECT 13.214 28.406 13.266 28.442 ;
      RECT 13.214 29.606 13.266 29.642 ;
      RECT 13.214 30.806 13.266 30.842 ;
      RECT 13.214 32.622 13.266 32.658 ;
      RECT 13.214 32.862 13.266 32.898 ;
      RECT 13.214 38.622 13.266 38.658 ;
      RECT 13.214 38.862 13.266 38.898 ;
      RECT 13.214 39.926 13.266 39.962 ;
      RECT 13.214 41.126 13.266 41.162 ;
      RECT 13.214 42.326 13.266 42.362 ;
      RECT 13.214 43.526 13.266 43.562 ;
      RECT 13.214 44.726 13.266 44.762 ;
      RECT 13.214 45.926 13.266 45.962 ;
      RECT 13.214 47.126 13.266 47.162 ;
      RECT 13.214 48.326 13.266 48.362 ;
      RECT 13.214 49.526 13.266 49.562 ;
      RECT 13.214 50.726 13.266 50.762 ;
      RECT 13.214 51.926 13.266 51.962 ;
      RECT 13.214 53.126 13.266 53.162 ;
      RECT 13.214 54.326 13.266 54.362 ;
      RECT 13.214 55.526 13.266 55.562 ;
      RECT 13.214 56.726 13.266 56.762 ;
      RECT 13.214 57.926 13.266 57.962 ;
      RECT 13.214 59.126 13.266 59.162 ;
      RECT 13.214 60.326 13.266 60.362 ;
      RECT 13.214 61.526 13.266 61.562 ;
      RECT 13.214 62.726 13.266 62.762 ;
      RECT 13.214 63.926 13.266 63.962 ;
      RECT 13.214 65.126 13.266 65.162 ;
      RECT 13.214 66.326 13.266 66.362 ;
      RECT 13.214 67.526 13.266 67.562 ;
      RECT 13.214 68.726 13.266 68.762 ;
      RECT 13.214 69.926 13.266 69.962 ;
      RECT 13.214 71.126 13.266 71.162 ;
      RECT 13.294 1.558 13.346 1.594 ;
      RECT 13.294 2.758 13.346 2.794 ;
      RECT 13.294 3.958 13.346 3.994 ;
      RECT 13.294 5.158 13.346 5.194 ;
      RECT 13.294 6.358 13.346 6.394 ;
      RECT 13.294 7.558 13.346 7.594 ;
      RECT 13.294 8.758 13.346 8.794 ;
      RECT 13.294 9.958 13.346 9.994 ;
      RECT 13.294 11.158 13.346 11.194 ;
      RECT 13.294 12.358 13.346 12.394 ;
      RECT 13.294 13.558 13.346 13.594 ;
      RECT 13.294 14.758 13.346 14.794 ;
      RECT 13.294 15.958 13.346 15.994 ;
      RECT 13.294 17.158 13.346 17.194 ;
      RECT 13.294 18.358 13.346 18.394 ;
      RECT 13.294 19.558 13.346 19.594 ;
      RECT 13.294 20.758 13.346 20.794 ;
      RECT 13.294 21.958 13.346 21.994 ;
      RECT 13.294 23.158 13.346 23.194 ;
      RECT 13.294 24.358 13.346 24.394 ;
      RECT 13.294 25.558 13.346 25.594 ;
      RECT 13.294 26.758 13.346 26.794 ;
      RECT 13.294 27.958 13.346 27.994 ;
      RECT 13.294 29.158 13.346 29.194 ;
      RECT 13.294 30.358 13.346 30.394 ;
      RECT 13.294 31.558 13.346 31.594 ;
      RECT 13.294 33.342 13.346 33.378 ;
      RECT 13.294 33.582 13.346 33.618 ;
      RECT 13.294 37.902 13.346 37.938 ;
      RECT 13.294 38.142 13.346 38.178 ;
      RECT 13.294 40.678 13.346 40.714 ;
      RECT 13.294 41.878 13.346 41.914 ;
      RECT 13.294 43.078 13.346 43.114 ;
      RECT 13.294 44.278 13.346 44.314 ;
      RECT 13.294 45.478 13.346 45.514 ;
      RECT 13.294 46.678 13.346 46.714 ;
      RECT 13.294 47.878 13.346 47.914 ;
      RECT 13.294 49.078 13.346 49.114 ;
      RECT 13.294 50.278 13.346 50.314 ;
      RECT 13.294 51.478 13.346 51.514 ;
      RECT 13.294 52.678 13.346 52.714 ;
      RECT 13.294 53.878 13.346 53.914 ;
      RECT 13.294 55.078 13.346 55.114 ;
      RECT 13.294 56.278 13.346 56.314 ;
      RECT 13.294 57.478 13.346 57.514 ;
      RECT 13.294 58.678 13.346 58.714 ;
      RECT 13.294 59.878 13.346 59.914 ;
      RECT 13.294 61.078 13.346 61.114 ;
      RECT 13.294 62.278 13.346 62.314 ;
      RECT 13.294 63.478 13.346 63.514 ;
      RECT 13.294 64.678 13.346 64.714 ;
      RECT 13.294 65.878 13.346 65.914 ;
      RECT 13.294 67.078 13.346 67.114 ;
      RECT 13.294 68.278 13.346 68.314 ;
      RECT 13.294 69.478 13.346 69.514 ;
      RECT 13.294 70.678 13.346 70.714 ;
      RECT 13.294 71.878 13.346 71.914 ;
      RECT 13.374 0.281 13.426 0.317 ;
      RECT 13.374 72.403 13.426 72.439 ;
      RECT 13.778 33.0435 13.814 33.0795 ;
      RECT 13.778 34.182 13.814 34.218 ;
      RECT 13.778 37.302 13.814 37.338 ;
      RECT 13.778 38.4405 13.814 38.4765 ;
      RECT 13.978 0.582 14.022 0.618 ;
      RECT 13.978 1.182 14.022 1.218 ;
      RECT 13.978 1.782 14.022 1.818 ;
      RECT 13.978 2.382 14.022 2.418 ;
      RECT 13.978 2.982 14.022 3.018 ;
      RECT 13.978 3.582 14.022 3.618 ;
      RECT 13.978 4.182 14.022 4.218 ;
      RECT 13.978 4.782 14.022 4.818 ;
      RECT 13.978 5.382 14.022 5.418 ;
      RECT 13.978 5.982 14.022 6.018 ;
      RECT 13.978 6.582 14.022 6.618 ;
      RECT 13.978 7.182 14.022 7.218 ;
      RECT 13.978 7.782 14.022 7.818 ;
      RECT 13.978 8.382 14.022 8.418 ;
      RECT 13.978 8.982 14.022 9.018 ;
      RECT 13.978 9.582 14.022 9.618 ;
      RECT 13.978 10.182 14.022 10.218 ;
      RECT 13.978 10.782 14.022 10.818 ;
      RECT 13.978 11.382 14.022 11.418 ;
      RECT 13.978 11.982 14.022 12.018 ;
      RECT 13.978 12.582 14.022 12.618 ;
      RECT 13.978 13.182 14.022 13.218 ;
      RECT 13.978 13.782 14.022 13.818 ;
      RECT 13.978 14.382 14.022 14.418 ;
      RECT 13.978 14.982 14.022 15.018 ;
      RECT 13.978 15.582 14.022 15.618 ;
      RECT 13.978 16.182 14.022 16.218 ;
      RECT 13.978 16.782 14.022 16.818 ;
      RECT 13.978 17.382 14.022 17.418 ;
      RECT 13.978 17.982 14.022 18.018 ;
      RECT 13.978 18.582 14.022 18.618 ;
      RECT 13.978 19.182 14.022 19.218 ;
      RECT 13.978 19.782 14.022 19.818 ;
      RECT 13.978 20.382 14.022 20.418 ;
      RECT 13.978 20.982 14.022 21.018 ;
      RECT 13.978 21.582 14.022 21.618 ;
      RECT 13.978 22.182 14.022 22.218 ;
      RECT 13.978 22.782 14.022 22.818 ;
      RECT 13.978 23.382 14.022 23.418 ;
      RECT 13.978 23.982 14.022 24.018 ;
      RECT 13.978 24.582 14.022 24.618 ;
      RECT 13.978 25.182 14.022 25.218 ;
      RECT 13.978 25.782 14.022 25.818 ;
      RECT 13.978 26.382 14.022 26.418 ;
      RECT 13.978 26.982 14.022 27.018 ;
      RECT 13.978 27.582 14.022 27.618 ;
      RECT 13.978 28.182 14.022 28.218 ;
      RECT 13.978 28.782 14.022 28.818 ;
      RECT 13.978 29.382 14.022 29.418 ;
      RECT 13.978 29.982 14.022 30.018 ;
      RECT 13.978 30.582 14.022 30.618 ;
      RECT 13.978 31.182 14.022 31.218 ;
      RECT 13.978 31.782 14.022 31.818 ;
      RECT 13.978 32.142 14.022 32.178 ;
      RECT 13.978 32.622 14.022 32.658 ;
      RECT 13.978 33.102 14.022 33.138 ;
      RECT 13.978 33.582 14.022 33.618 ;
      RECT 13.978 34.062 14.022 34.098 ;
      RECT 13.978 34.542 14.022 34.578 ;
      RECT 13.978 35.022 14.022 35.058 ;
      RECT 13.978 35.502 14.022 35.538 ;
      RECT 13.978 35.982 14.022 36.018 ;
      RECT 13.978 36.462 14.022 36.498 ;
      RECT 13.978 36.942 14.022 36.978 ;
      RECT 13.978 37.422 14.022 37.458 ;
      RECT 13.978 37.902 14.022 37.938 ;
      RECT 13.978 38.382 14.022 38.418 ;
      RECT 13.978 38.862 14.022 38.898 ;
      RECT 13.978 39.342 14.022 39.378 ;
      RECT 13.978 39.702 14.022 39.738 ;
      RECT 13.978 40.302 14.022 40.338 ;
      RECT 13.978 40.902 14.022 40.938 ;
      RECT 13.978 41.502 14.022 41.538 ;
      RECT 13.978 42.102 14.022 42.138 ;
      RECT 13.978 42.702 14.022 42.738 ;
      RECT 13.978 43.302 14.022 43.338 ;
      RECT 13.978 43.902 14.022 43.938 ;
      RECT 13.978 44.502 14.022 44.538 ;
      RECT 13.978 45.102 14.022 45.138 ;
      RECT 13.978 45.702 14.022 45.738 ;
      RECT 13.978 46.302 14.022 46.338 ;
      RECT 13.978 46.902 14.022 46.938 ;
      RECT 13.978 47.502 14.022 47.538 ;
      RECT 13.978 48.102 14.022 48.138 ;
      RECT 13.978 48.702 14.022 48.738 ;
      RECT 13.978 49.302 14.022 49.338 ;
      RECT 13.978 49.902 14.022 49.938 ;
      RECT 13.978 50.502 14.022 50.538 ;
      RECT 13.978 51.102 14.022 51.138 ;
      RECT 13.978 51.702 14.022 51.738 ;
      RECT 13.978 52.302 14.022 52.338 ;
      RECT 13.978 52.902 14.022 52.938 ;
      RECT 13.978 53.502 14.022 53.538 ;
      RECT 13.978 54.102 14.022 54.138 ;
      RECT 13.978 54.702 14.022 54.738 ;
      RECT 13.978 55.302 14.022 55.338 ;
      RECT 13.978 55.902 14.022 55.938 ;
      RECT 13.978 56.502 14.022 56.538 ;
      RECT 13.978 57.102 14.022 57.138 ;
      RECT 13.978 57.702 14.022 57.738 ;
      RECT 13.978 58.302 14.022 58.338 ;
      RECT 13.978 58.902 14.022 58.938 ;
      RECT 13.978 59.502 14.022 59.538 ;
      RECT 13.978 60.102 14.022 60.138 ;
      RECT 13.978 60.702 14.022 60.738 ;
      RECT 13.978 61.302 14.022 61.338 ;
      RECT 13.978 61.902 14.022 61.938 ;
      RECT 13.978 62.502 14.022 62.538 ;
      RECT 13.978 63.102 14.022 63.138 ;
      RECT 13.978 63.702 14.022 63.738 ;
      RECT 13.978 64.302 14.022 64.338 ;
      RECT 13.978 64.902 14.022 64.938 ;
      RECT 13.978 65.502 14.022 65.538 ;
      RECT 13.978 66.102 14.022 66.138 ;
      RECT 13.978 66.702 14.022 66.738 ;
      RECT 13.978 67.302 14.022 67.338 ;
      RECT 13.978 67.902 14.022 67.938 ;
      RECT 13.978 68.502 14.022 68.538 ;
      RECT 13.978 69.102 14.022 69.138 ;
      RECT 13.978 69.702 14.022 69.738 ;
      RECT 13.978 70.302 14.022 70.338 ;
      RECT 13.978 70.902 14.022 70.938 ;
      RECT 13.978 71.502 14.022 71.538 ;
      RECT 13.978 72.102 14.022 72.138 ;
      RECT 14.132 1.558 14.186 1.594 ;
      RECT 14.132 2.758 14.186 2.794 ;
      RECT 14.132 3.958 14.186 3.994 ;
      RECT 14.132 5.158 14.186 5.194 ;
      RECT 14.132 6.358 14.186 6.394 ;
      RECT 14.132 7.558 14.186 7.594 ;
      RECT 14.132 8.758 14.186 8.794 ;
      RECT 14.132 9.958 14.186 9.994 ;
      RECT 14.132 11.158 14.186 11.194 ;
      RECT 14.132 12.358 14.186 12.394 ;
      RECT 14.132 13.558 14.186 13.594 ;
      RECT 14.132 14.758 14.186 14.794 ;
      RECT 14.132 15.958 14.186 15.994 ;
      RECT 14.132 17.158 14.186 17.194 ;
      RECT 14.132 18.358 14.186 18.394 ;
      RECT 14.132 19.558 14.186 19.594 ;
      RECT 14.132 20.758 14.186 20.794 ;
      RECT 14.132 21.958 14.186 21.994 ;
      RECT 14.132 23.158 14.186 23.194 ;
      RECT 14.132 24.358 14.186 24.394 ;
      RECT 14.132 25.558 14.186 25.594 ;
      RECT 14.132 26.758 14.186 26.794 ;
      RECT 14.132 27.958 14.186 27.994 ;
      RECT 14.132 29.158 14.186 29.194 ;
      RECT 14.132 30.358 14.186 30.394 ;
      RECT 14.132 31.558 14.186 31.594 ;
      RECT 14.132 34.1205 14.186 34.1565 ;
      RECT 14.132 34.3605 14.186 34.3965 ;
      RECT 14.132 35.9235 14.186 35.9595 ;
      RECT 14.132 37.3635 14.186 37.3995 ;
      RECT 14.132 40.678 14.186 40.714 ;
      RECT 14.132 41.878 14.186 41.914 ;
      RECT 14.132 43.078 14.186 43.114 ;
      RECT 14.132 44.278 14.186 44.314 ;
      RECT 14.132 45.478 14.186 45.514 ;
      RECT 14.132 46.678 14.186 46.714 ;
      RECT 14.132 47.878 14.186 47.914 ;
      RECT 14.132 49.078 14.186 49.114 ;
      RECT 14.132 50.278 14.186 50.314 ;
      RECT 14.132 51.478 14.186 51.514 ;
      RECT 14.132 52.678 14.186 52.714 ;
      RECT 14.132 53.878 14.186 53.914 ;
      RECT 14.132 55.078 14.186 55.114 ;
      RECT 14.132 56.278 14.186 56.314 ;
      RECT 14.132 57.478 14.186 57.514 ;
      RECT 14.132 58.678 14.186 58.714 ;
      RECT 14.132 59.878 14.186 59.914 ;
      RECT 14.132 61.078 14.186 61.114 ;
      RECT 14.132 62.278 14.186 62.314 ;
      RECT 14.132 63.478 14.186 63.514 ;
      RECT 14.132 64.678 14.186 64.714 ;
      RECT 14.132 65.878 14.186 65.914 ;
      RECT 14.132 67.078 14.186 67.114 ;
      RECT 14.132 68.278 14.186 68.314 ;
      RECT 14.132 69.478 14.186 69.514 ;
      RECT 14.132 70.678 14.186 70.714 ;
      RECT 14.132 71.878 14.186 71.914 ;
      RECT 14.214 0.806 14.268 0.842 ;
      RECT 14.214 2.006 14.268 2.042 ;
      RECT 14.214 3.206 14.268 3.242 ;
      RECT 14.214 4.406 14.268 4.442 ;
      RECT 14.214 5.606 14.268 5.642 ;
      RECT 14.214 6.806 14.268 6.842 ;
      RECT 14.214 8.006 14.268 8.042 ;
      RECT 14.214 9.206 14.268 9.242 ;
      RECT 14.214 10.406 14.268 10.442 ;
      RECT 14.214 11.606 14.268 11.642 ;
      RECT 14.214 12.806 14.268 12.842 ;
      RECT 14.214 14.006 14.268 14.042 ;
      RECT 14.214 15.206 14.268 15.242 ;
      RECT 14.214 16.406 14.268 16.442 ;
      RECT 14.214 17.606 14.268 17.642 ;
      RECT 14.214 18.806 14.268 18.842 ;
      RECT 14.214 20.006 14.268 20.042 ;
      RECT 14.214 21.206 14.268 21.242 ;
      RECT 14.214 22.406 14.268 22.442 ;
      RECT 14.214 23.606 14.268 23.642 ;
      RECT 14.214 24.806 14.268 24.842 ;
      RECT 14.214 26.006 14.268 26.042 ;
      RECT 14.214 27.206 14.268 27.242 ;
      RECT 14.214 28.406 14.268 28.442 ;
      RECT 14.214 29.606 14.268 29.642 ;
      RECT 14.214 30.806 14.268 30.842 ;
      RECT 14.214 34.0035 14.268 34.0395 ;
      RECT 14.214 37.0005 14.268 37.0365 ;
      RECT 14.214 39.926 14.268 39.962 ;
      RECT 14.214 41.126 14.268 41.162 ;
      RECT 14.214 42.326 14.268 42.362 ;
      RECT 14.214 43.526 14.268 43.562 ;
      RECT 14.214 44.726 14.268 44.762 ;
      RECT 14.214 45.926 14.268 45.962 ;
      RECT 14.214 47.126 14.268 47.162 ;
      RECT 14.214 48.326 14.268 48.362 ;
      RECT 14.214 49.526 14.268 49.562 ;
      RECT 14.214 50.726 14.268 50.762 ;
      RECT 14.214 51.926 14.268 51.962 ;
      RECT 14.214 53.126 14.268 53.162 ;
      RECT 14.214 54.326 14.268 54.362 ;
      RECT 14.214 55.526 14.268 55.562 ;
      RECT 14.214 56.726 14.268 56.762 ;
      RECT 14.214 57.926 14.268 57.962 ;
      RECT 14.214 59.126 14.268 59.162 ;
      RECT 14.214 60.326 14.268 60.362 ;
      RECT 14.214 61.526 14.268 61.562 ;
      RECT 14.214 62.726 14.268 62.762 ;
      RECT 14.214 63.926 14.268 63.962 ;
      RECT 14.214 65.126 14.268 65.162 ;
      RECT 14.214 66.326 14.268 66.362 ;
      RECT 14.214 67.526 14.268 67.562 ;
      RECT 14.214 68.726 14.268 68.762 ;
      RECT 14.214 69.926 14.268 69.962 ;
      RECT 14.214 71.126 14.268 71.162 ;
      RECT 14.378 34.182 14.422 34.218 ;
      RECT 14.378 34.422 14.422 34.458 ;
      RECT 14.378 36.342 14.422 36.378 ;
      RECT 14.378 37.302 14.422 37.338 ;
      RECT 14.532 1.482 14.586 1.518 ;
      RECT 14.532 2.682 14.586 2.718 ;
      RECT 14.532 3.882 14.586 3.918 ;
      RECT 14.532 5.082 14.586 5.118 ;
      RECT 14.532 6.282 14.586 6.318 ;
      RECT 14.532 7.482 14.586 7.518 ;
      RECT 14.532 8.682 14.586 8.718 ;
      RECT 14.532 9.882 14.586 9.918 ;
      RECT 14.532 11.082 14.586 11.118 ;
      RECT 14.532 12.282 14.586 12.318 ;
      RECT 14.532 13.482 14.586 13.518 ;
      RECT 14.532 14.682 14.586 14.718 ;
      RECT 14.532 15.882 14.586 15.918 ;
      RECT 14.532 17.082 14.586 17.118 ;
      RECT 14.532 18.282 14.586 18.318 ;
      RECT 14.532 19.482 14.586 19.518 ;
      RECT 14.532 20.682 14.586 20.718 ;
      RECT 14.532 21.882 14.586 21.918 ;
      RECT 14.532 23.082 14.586 23.118 ;
      RECT 14.532 24.282 14.586 24.318 ;
      RECT 14.532 25.482 14.586 25.518 ;
      RECT 14.532 26.682 14.586 26.718 ;
      RECT 14.532 27.882 14.586 27.918 ;
      RECT 14.532 29.082 14.586 29.118 ;
      RECT 14.532 30.282 14.586 30.318 ;
      RECT 14.532 31.482 14.586 31.518 ;
      RECT 14.532 32.3235 14.586 32.3595 ;
      RECT 14.532 32.4405 14.586 32.4765 ;
      RECT 14.532 37.6035 14.586 37.6395 ;
      RECT 14.532 38.982 14.586 39.018 ;
      RECT 14.532 39.222 14.586 39.258 ;
      RECT 14.532 40.602 14.586 40.638 ;
      RECT 14.532 41.802 14.586 41.838 ;
      RECT 14.532 43.002 14.586 43.038 ;
      RECT 14.532 44.202 14.586 44.238 ;
      RECT 14.532 45.402 14.586 45.438 ;
      RECT 14.532 46.602 14.586 46.638 ;
      RECT 14.532 47.802 14.586 47.838 ;
      RECT 14.532 49.002 14.586 49.038 ;
      RECT 14.532 50.202 14.586 50.238 ;
      RECT 14.532 51.402 14.586 51.438 ;
      RECT 14.532 52.602 14.586 52.638 ;
      RECT 14.532 53.802 14.586 53.838 ;
      RECT 14.532 55.002 14.586 55.038 ;
      RECT 14.532 56.202 14.586 56.238 ;
      RECT 14.532 57.402 14.586 57.438 ;
      RECT 14.532 58.602 14.586 58.638 ;
      RECT 14.532 59.802 14.586 59.838 ;
      RECT 14.532 61.002 14.586 61.038 ;
      RECT 14.532 62.202 14.586 62.238 ;
      RECT 14.532 63.402 14.586 63.438 ;
      RECT 14.532 64.602 14.586 64.638 ;
      RECT 14.532 65.802 14.586 65.838 ;
      RECT 14.532 67.002 14.586 67.038 ;
      RECT 14.532 68.202 14.586 68.238 ;
      RECT 14.532 69.402 14.586 69.438 ;
      RECT 14.532 70.602 14.586 70.638 ;
      RECT 14.532 71.802 14.586 71.838 ;
      RECT 14.614 0.806 14.668 0.842 ;
      RECT 14.614 2.006 14.668 2.042 ;
      RECT 14.614 3.206 14.668 3.242 ;
      RECT 14.614 4.406 14.668 4.442 ;
      RECT 14.614 5.606 14.668 5.642 ;
      RECT 14.614 6.806 14.668 6.842 ;
      RECT 14.614 8.006 14.668 8.042 ;
      RECT 14.614 9.206 14.668 9.242 ;
      RECT 14.614 10.406 14.668 10.442 ;
      RECT 14.614 11.606 14.668 11.642 ;
      RECT 14.614 12.806 14.668 12.842 ;
      RECT 14.614 14.006 14.668 14.042 ;
      RECT 14.614 15.206 14.668 15.242 ;
      RECT 14.614 16.406 14.668 16.442 ;
      RECT 14.614 17.606 14.668 17.642 ;
      RECT 14.614 18.806 14.668 18.842 ;
      RECT 14.614 20.006 14.668 20.042 ;
      RECT 14.614 21.206 14.668 21.242 ;
      RECT 14.614 22.406 14.668 22.442 ;
      RECT 14.614 23.606 14.668 23.642 ;
      RECT 14.614 24.806 14.668 24.842 ;
      RECT 14.614 26.006 14.668 26.042 ;
      RECT 14.614 27.206 14.668 27.242 ;
      RECT 14.614 28.406 14.668 28.442 ;
      RECT 14.614 29.606 14.668 29.642 ;
      RECT 14.614 30.806 14.668 30.842 ;
      RECT 14.614 32.2005 14.668 32.2365 ;
      RECT 14.614 32.6805 14.668 32.7165 ;
      RECT 14.614 37.8435 14.668 37.8795 ;
      RECT 14.614 38.686 14.668 38.711 ;
      RECT 14.614 38.809 14.668 38.834 ;
      RECT 14.614 39.926 14.668 39.962 ;
      RECT 14.614 41.126 14.668 41.162 ;
      RECT 14.614 42.326 14.668 42.362 ;
      RECT 14.614 43.526 14.668 43.562 ;
      RECT 14.614 44.726 14.668 44.762 ;
      RECT 14.614 45.926 14.668 45.962 ;
      RECT 14.614 47.126 14.668 47.162 ;
      RECT 14.614 48.326 14.668 48.362 ;
      RECT 14.614 49.526 14.668 49.562 ;
      RECT 14.614 50.726 14.668 50.762 ;
      RECT 14.614 51.926 14.668 51.962 ;
      RECT 14.614 53.126 14.668 53.162 ;
      RECT 14.614 54.326 14.668 54.362 ;
      RECT 14.614 55.526 14.668 55.562 ;
      RECT 14.614 56.726 14.668 56.762 ;
      RECT 14.614 57.926 14.668 57.962 ;
      RECT 14.614 59.126 14.668 59.162 ;
      RECT 14.614 60.326 14.668 60.362 ;
      RECT 14.614 61.526 14.668 61.562 ;
      RECT 14.614 62.726 14.668 62.762 ;
      RECT 14.614 63.926 14.668 63.962 ;
      RECT 14.614 65.126 14.668 65.162 ;
      RECT 14.614 66.326 14.668 66.362 ;
      RECT 14.614 67.526 14.668 67.562 ;
      RECT 14.614 68.726 14.668 68.762 ;
      RECT 14.614 69.926 14.668 69.962 ;
      RECT 14.614 71.126 14.668 71.162 ;
      RECT 14.696 1.482 14.75 1.518 ;
      RECT 14.696 2.682 14.75 2.718 ;
      RECT 14.696 3.882 14.75 3.918 ;
      RECT 14.696 5.082 14.75 5.118 ;
      RECT 14.696 6.282 14.75 6.318 ;
      RECT 14.696 7.482 14.75 7.518 ;
      RECT 14.696 8.682 14.75 8.718 ;
      RECT 14.696 9.882 14.75 9.918 ;
      RECT 14.696 11.082 14.75 11.118 ;
      RECT 14.696 12.282 14.75 12.318 ;
      RECT 14.696 13.482 14.75 13.518 ;
      RECT 14.696 14.682 14.75 14.718 ;
      RECT 14.696 15.882 14.75 15.918 ;
      RECT 14.696 17.082 14.75 17.118 ;
      RECT 14.696 18.282 14.75 18.318 ;
      RECT 14.696 19.482 14.75 19.518 ;
      RECT 14.696 20.682 14.75 20.718 ;
      RECT 14.696 21.882 14.75 21.918 ;
      RECT 14.696 23.082 14.75 23.118 ;
      RECT 14.696 24.282 14.75 24.318 ;
      RECT 14.696 25.482 14.75 25.518 ;
      RECT 14.696 26.682 14.75 26.718 ;
      RECT 14.696 27.882 14.75 27.918 ;
      RECT 14.696 29.082 14.75 29.118 ;
      RECT 14.696 30.282 14.75 30.318 ;
      RECT 14.696 31.482 14.75 31.518 ;
      RECT 14.696 32.5635 14.75 32.5995 ;
      RECT 14.696 32.8035 14.75 32.8395 ;
      RECT 14.696 37.6035 14.75 37.6395 ;
      RECT 14.696 38.5635 14.75 38.5995 ;
      RECT 14.696 38.9205 14.75 38.9565 ;
      RECT 14.696 40.602 14.75 40.638 ;
      RECT 14.696 41.802 14.75 41.838 ;
      RECT 14.696 43.002 14.75 43.038 ;
      RECT 14.696 44.202 14.75 44.238 ;
      RECT 14.696 45.402 14.75 45.438 ;
      RECT 14.696 46.602 14.75 46.638 ;
      RECT 14.696 47.802 14.75 47.838 ;
      RECT 14.696 49.002 14.75 49.038 ;
      RECT 14.696 50.202 14.75 50.238 ;
      RECT 14.696 51.402 14.75 51.438 ;
      RECT 14.696 52.602 14.75 52.638 ;
      RECT 14.696 53.802 14.75 53.838 ;
      RECT 14.696 55.002 14.75 55.038 ;
      RECT 14.696 56.202 14.75 56.238 ;
      RECT 14.696 57.402 14.75 57.438 ;
      RECT 14.696 58.602 14.75 58.638 ;
      RECT 14.696 59.802 14.75 59.838 ;
      RECT 14.696 61.002 14.75 61.038 ;
      RECT 14.696 62.202 14.75 62.238 ;
      RECT 14.696 63.402 14.75 63.438 ;
      RECT 14.696 64.602 14.75 64.638 ;
      RECT 14.696 65.802 14.75 65.838 ;
      RECT 14.696 67.002 14.75 67.038 ;
      RECT 14.696 68.202 14.75 68.238 ;
      RECT 14.696 69.402 14.75 69.438 ;
      RECT 14.696 70.602 14.75 70.638 ;
      RECT 14.696 71.802 14.75 71.838 ;
      RECT 14.778 0.806 14.832 0.842 ;
      RECT 14.778 2.006 14.832 2.042 ;
      RECT 14.778 3.206 14.832 3.242 ;
      RECT 14.778 4.406 14.832 4.442 ;
      RECT 14.778 5.606 14.832 5.642 ;
      RECT 14.778 6.806 14.832 6.842 ;
      RECT 14.778 8.006 14.832 8.042 ;
      RECT 14.778 9.206 14.832 9.242 ;
      RECT 14.778 10.406 14.832 10.442 ;
      RECT 14.778 11.606 14.832 11.642 ;
      RECT 14.778 12.806 14.832 12.842 ;
      RECT 14.778 14.006 14.832 14.042 ;
      RECT 14.778 15.206 14.832 15.242 ;
      RECT 14.778 16.406 14.832 16.442 ;
      RECT 14.778 17.606 14.832 17.642 ;
      RECT 14.778 18.806 14.832 18.842 ;
      RECT 14.778 20.006 14.832 20.042 ;
      RECT 14.778 21.206 14.832 21.242 ;
      RECT 14.778 22.406 14.832 22.442 ;
      RECT 14.778 23.606 14.832 23.642 ;
      RECT 14.778 24.806 14.832 24.842 ;
      RECT 14.778 26.006 14.832 26.042 ;
      RECT 14.778 27.206 14.832 27.242 ;
      RECT 14.778 28.406 14.832 28.442 ;
      RECT 14.778 29.606 14.832 29.642 ;
      RECT 14.778 30.806 14.832 30.842 ;
      RECT 14.778 32.9205 14.832 32.9565 ;
      RECT 14.778 33.222 14.832 33.258 ;
      RECT 14.778 37.782 14.832 37.818 ;
      RECT 14.778 38.262 14.832 38.298 ;
      RECT 14.778 38.6805 14.832 38.7165 ;
      RECT 14.778 39.926 14.832 39.962 ;
      RECT 14.778 41.126 14.832 41.162 ;
      RECT 14.778 42.326 14.832 42.362 ;
      RECT 14.778 43.526 14.832 43.562 ;
      RECT 14.778 44.726 14.832 44.762 ;
      RECT 14.778 45.926 14.832 45.962 ;
      RECT 14.778 47.126 14.832 47.162 ;
      RECT 14.778 48.326 14.832 48.362 ;
      RECT 14.778 49.526 14.832 49.562 ;
      RECT 14.778 50.726 14.832 50.762 ;
      RECT 14.778 51.926 14.832 51.962 ;
      RECT 14.778 53.126 14.832 53.162 ;
      RECT 14.778 54.326 14.832 54.362 ;
      RECT 14.778 55.526 14.832 55.562 ;
      RECT 14.778 56.726 14.832 56.762 ;
      RECT 14.778 57.926 14.832 57.962 ;
      RECT 14.778 59.126 14.832 59.162 ;
      RECT 14.778 60.326 14.832 60.362 ;
      RECT 14.778 61.526 14.832 61.562 ;
      RECT 14.778 62.726 14.832 62.762 ;
      RECT 14.778 63.926 14.832 63.962 ;
      RECT 14.778 65.126 14.832 65.162 ;
      RECT 14.778 66.326 14.832 66.362 ;
      RECT 14.778 67.526 14.832 67.562 ;
      RECT 14.778 68.726 14.832 68.762 ;
      RECT 14.778 69.926 14.832 69.962 ;
      RECT 14.778 71.126 14.832 71.162 ;
      RECT 14.86 0.582 14.904 0.618 ;
      RECT 14.86 1.782 14.904 1.818 ;
      RECT 14.86 2.982 14.904 3.018 ;
      RECT 14.86 4.182 14.904 4.218 ;
      RECT 14.86 5.382 14.904 5.418 ;
      RECT 14.86 6.582 14.904 6.618 ;
      RECT 14.86 7.782 14.904 7.818 ;
      RECT 14.86 8.982 14.904 9.018 ;
      RECT 14.86 10.182 14.904 10.218 ;
      RECT 14.86 11.382 14.904 11.418 ;
      RECT 14.86 12.582 14.904 12.618 ;
      RECT 14.86 13.782 14.904 13.818 ;
      RECT 14.86 14.982 14.904 15.018 ;
      RECT 14.86 16.182 14.904 16.218 ;
      RECT 14.86 17.382 14.904 17.418 ;
      RECT 14.86 18.582 14.904 18.618 ;
      RECT 14.86 19.782 14.904 19.818 ;
      RECT 14.86 20.982 14.904 21.018 ;
      RECT 14.86 22.182 14.904 22.218 ;
      RECT 14.86 23.382 14.904 23.418 ;
      RECT 14.86 24.582 14.904 24.618 ;
      RECT 14.86 25.782 14.904 25.818 ;
      RECT 14.86 26.982 14.904 27.018 ;
      RECT 14.86 28.182 14.904 28.218 ;
      RECT 14.86 29.382 14.904 29.418 ;
      RECT 14.86 30.582 14.904 30.618 ;
      RECT 14.86 31.782 14.904 31.818 ;
      RECT 14.86 32.142 14.904 32.178 ;
      RECT 14.86 32.622 14.904 32.658 ;
      RECT 14.86 33.102 14.904 33.138 ;
      RECT 14.86 33.582 14.904 33.618 ;
      RECT 14.86 34.062 14.904 34.098 ;
      RECT 14.86 34.542 14.904 34.578 ;
      RECT 14.86 35.022 14.904 35.058 ;
      RECT 14.86 35.502 14.904 35.538 ;
      RECT 14.86 35.982 14.904 36.018 ;
      RECT 14.86 36.462 14.904 36.498 ;
      RECT 14.86 36.942 14.904 36.978 ;
      RECT 14.86 37.422 14.904 37.458 ;
      RECT 14.86 37.902 14.904 37.938 ;
      RECT 14.86 38.382 14.904 38.418 ;
      RECT 14.86 38.862 14.904 38.898 ;
      RECT 14.86 39.342 14.904 39.378 ;
      RECT 14.86 39.702 14.904 39.738 ;
      RECT 14.86 40.902 14.904 40.938 ;
      RECT 14.86 42.102 14.904 42.138 ;
      RECT 14.86 43.302 14.904 43.338 ;
      RECT 14.86 44.502 14.904 44.538 ;
      RECT 14.86 45.702 14.904 45.738 ;
      RECT 14.86 46.902 14.904 46.938 ;
      RECT 14.86 48.102 14.904 48.138 ;
      RECT 14.86 49.302 14.904 49.338 ;
      RECT 14.86 50.502 14.904 50.538 ;
      RECT 14.86 51.702 14.904 51.738 ;
      RECT 14.86 52.902 14.904 52.938 ;
      RECT 14.86 54.102 14.904 54.138 ;
      RECT 14.86 55.302 14.904 55.338 ;
      RECT 14.86 56.502 14.904 56.538 ;
      RECT 14.86 57.702 14.904 57.738 ;
      RECT 14.86 58.902 14.904 58.938 ;
      RECT 14.86 60.102 14.904 60.138 ;
      RECT 14.86 61.302 14.904 61.338 ;
      RECT 14.86 62.502 14.904 62.538 ;
      RECT 14.86 63.702 14.904 63.738 ;
      RECT 14.86 64.902 14.904 64.938 ;
      RECT 14.86 66.102 14.904 66.138 ;
      RECT 14.86 67.302 14.904 67.338 ;
      RECT 14.86 68.502 14.904 68.538 ;
      RECT 14.86 69.702 14.904 69.738 ;
      RECT 14.86 70.902 14.904 70.938 ;
      RECT 14.86 72.102 14.904 72.138 ;
      RECT 15.014 34.4835 15.068 34.5195 ;
      RECT 15.014 37.3635 15.068 37.3995 ;
      RECT 15.178 0.582 15.222 0.618 ;
      RECT 15.178 1.182 15.222 1.218 ;
      RECT 15.178 1.782 15.222 1.818 ;
      RECT 15.178 2.382 15.222 2.418 ;
      RECT 15.178 2.982 15.222 3.018 ;
      RECT 15.178 3.582 15.222 3.618 ;
      RECT 15.178 4.182 15.222 4.218 ;
      RECT 15.178 4.782 15.222 4.818 ;
      RECT 15.178 5.382 15.222 5.418 ;
      RECT 15.178 5.982 15.222 6.018 ;
      RECT 15.178 6.582 15.222 6.618 ;
      RECT 15.178 7.182 15.222 7.218 ;
      RECT 15.178 7.782 15.222 7.818 ;
      RECT 15.178 8.382 15.222 8.418 ;
      RECT 15.178 8.982 15.222 9.018 ;
      RECT 15.178 9.582 15.222 9.618 ;
      RECT 15.178 10.182 15.222 10.218 ;
      RECT 15.178 10.782 15.222 10.818 ;
      RECT 15.178 11.382 15.222 11.418 ;
      RECT 15.178 11.982 15.222 12.018 ;
      RECT 15.178 12.582 15.222 12.618 ;
      RECT 15.178 13.182 15.222 13.218 ;
      RECT 15.178 13.782 15.222 13.818 ;
      RECT 15.178 14.382 15.222 14.418 ;
      RECT 15.178 14.982 15.222 15.018 ;
      RECT 15.178 15.582 15.222 15.618 ;
      RECT 15.178 16.182 15.222 16.218 ;
      RECT 15.178 16.782 15.222 16.818 ;
      RECT 15.178 17.382 15.222 17.418 ;
      RECT 15.178 17.982 15.222 18.018 ;
      RECT 15.178 18.582 15.222 18.618 ;
      RECT 15.178 19.182 15.222 19.218 ;
      RECT 15.178 19.782 15.222 19.818 ;
      RECT 15.178 20.382 15.222 20.418 ;
      RECT 15.178 20.982 15.222 21.018 ;
      RECT 15.178 21.582 15.222 21.618 ;
      RECT 15.178 22.182 15.222 22.218 ;
      RECT 15.178 22.782 15.222 22.818 ;
      RECT 15.178 23.382 15.222 23.418 ;
      RECT 15.178 23.982 15.222 24.018 ;
      RECT 15.178 24.582 15.222 24.618 ;
      RECT 15.178 25.182 15.222 25.218 ;
      RECT 15.178 25.782 15.222 25.818 ;
      RECT 15.178 26.382 15.222 26.418 ;
      RECT 15.178 26.982 15.222 27.018 ;
      RECT 15.178 27.582 15.222 27.618 ;
      RECT 15.178 28.182 15.222 28.218 ;
      RECT 15.178 28.782 15.222 28.818 ;
      RECT 15.178 29.382 15.222 29.418 ;
      RECT 15.178 29.982 15.222 30.018 ;
      RECT 15.178 30.582 15.222 30.618 ;
      RECT 15.178 31.182 15.222 31.218 ;
      RECT 15.178 31.782 15.222 31.818 ;
      RECT 15.178 32.142 15.222 32.178 ;
      RECT 15.178 32.622 15.222 32.658 ;
      RECT 15.178 33.102 15.222 33.138 ;
      RECT 15.178 33.2835 15.222 33.3195 ;
      RECT 15.178 33.582 15.222 33.618 ;
      RECT 15.178 34.062 15.222 34.098 ;
      RECT 15.178 34.542 15.222 34.578 ;
      RECT 15.178 35.022 15.222 35.058 ;
      RECT 15.178 35.502 15.222 35.538 ;
      RECT 15.178 35.982 15.222 36.018 ;
      RECT 15.178 36.462 15.222 36.498 ;
      RECT 15.178 36.942 15.222 36.978 ;
      RECT 15.178 37.4275 15.222 37.4525 ;
      RECT 15.178 37.9075 15.222 37.9325 ;
      RECT 15.178 38.382 15.222 38.418 ;
      RECT 15.178 38.8675 15.222 38.8925 ;
      RECT 15.178 39.342 15.222 39.378 ;
      RECT 15.178 39.702 15.222 39.738 ;
      RECT 15.178 40.302 15.222 40.338 ;
      RECT 15.178 40.902 15.222 40.938 ;
      RECT 15.178 41.502 15.222 41.538 ;
      RECT 15.178 42.102 15.222 42.138 ;
      RECT 15.178 42.702 15.222 42.738 ;
      RECT 15.178 43.302 15.222 43.338 ;
      RECT 15.178 43.902 15.222 43.938 ;
      RECT 15.178 44.502 15.222 44.538 ;
      RECT 15.178 45.102 15.222 45.138 ;
      RECT 15.178 45.702 15.222 45.738 ;
      RECT 15.178 46.302 15.222 46.338 ;
      RECT 15.178 46.902 15.222 46.938 ;
      RECT 15.178 47.502 15.222 47.538 ;
      RECT 15.178 48.102 15.222 48.138 ;
      RECT 15.178 48.702 15.222 48.738 ;
      RECT 15.178 49.302 15.222 49.338 ;
      RECT 15.178 49.902 15.222 49.938 ;
      RECT 15.178 50.502 15.222 50.538 ;
      RECT 15.178 51.102 15.222 51.138 ;
      RECT 15.178 51.702 15.222 51.738 ;
      RECT 15.178 52.302 15.222 52.338 ;
      RECT 15.178 52.902 15.222 52.938 ;
      RECT 15.178 53.502 15.222 53.538 ;
      RECT 15.178 54.102 15.222 54.138 ;
      RECT 15.178 54.702 15.222 54.738 ;
      RECT 15.178 55.302 15.222 55.338 ;
      RECT 15.178 55.902 15.222 55.938 ;
      RECT 15.178 56.502 15.222 56.538 ;
      RECT 15.178 57.102 15.222 57.138 ;
      RECT 15.178 57.702 15.222 57.738 ;
      RECT 15.178 58.302 15.222 58.338 ;
      RECT 15.178 58.902 15.222 58.938 ;
      RECT 15.178 59.502 15.222 59.538 ;
      RECT 15.178 60.102 15.222 60.138 ;
      RECT 15.178 60.702 15.222 60.738 ;
      RECT 15.178 61.302 15.222 61.338 ;
      RECT 15.178 61.902 15.222 61.938 ;
      RECT 15.178 62.502 15.222 62.538 ;
      RECT 15.178 63.102 15.222 63.138 ;
      RECT 15.178 63.702 15.222 63.738 ;
      RECT 15.178 64.302 15.222 64.338 ;
      RECT 15.178 64.902 15.222 64.938 ;
      RECT 15.178 65.502 15.222 65.538 ;
      RECT 15.178 66.102 15.222 66.138 ;
      RECT 15.178 66.702 15.222 66.738 ;
      RECT 15.178 67.302 15.222 67.338 ;
      RECT 15.178 67.902 15.222 67.938 ;
      RECT 15.178 68.502 15.222 68.538 ;
      RECT 15.178 69.102 15.222 69.138 ;
      RECT 15.178 69.702 15.222 69.738 ;
      RECT 15.178 70.302 15.222 70.338 ;
      RECT 15.178 70.902 15.222 70.938 ;
      RECT 15.178 71.502 15.222 71.538 ;
      RECT 15.178 72.102 15.222 72.138 ;
      RECT 15.398 34.6005 15.45 34.6365 ;
      RECT 15.398 36.102 15.45 36.138 ;
      RECT 15.478 33.702 15.53 33.738 ;
      RECT 15.478 38.0835 15.53 38.1195 ;
      RECT 15.558 1.3345 15.63 1.3595 ;
      RECT 15.558 2.5345 15.63 2.5595 ;
      RECT 15.558 3.7345 15.63 3.7595 ;
      RECT 15.558 4.9345 15.63 4.9595 ;
      RECT 15.558 6.1345 15.63 6.1595 ;
      RECT 15.558 7.3345 15.63 7.3595 ;
      RECT 15.558 8.5345 15.63 8.5595 ;
      RECT 15.558 9.7345 15.63 9.7595 ;
      RECT 15.558 10.9345 15.63 10.9595 ;
      RECT 15.558 12.1345 15.63 12.1595 ;
      RECT 15.558 13.3345 15.63 13.3595 ;
      RECT 15.558 14.5345 15.63 14.5595 ;
      RECT 15.558 15.7345 15.63 15.7595 ;
      RECT 15.558 16.9345 15.63 16.9595 ;
      RECT 15.558 18.1345 15.63 18.1595 ;
      RECT 15.558 19.3345 15.63 19.3595 ;
      RECT 15.558 20.5345 15.63 20.5595 ;
      RECT 15.558 21.7345 15.63 21.7595 ;
      RECT 15.558 22.9345 15.63 22.9595 ;
      RECT 15.558 24.1345 15.63 24.1595 ;
      RECT 15.558 25.3345 15.63 25.3595 ;
      RECT 15.558 26.5345 15.63 26.5595 ;
      RECT 15.558 27.7345 15.63 27.7595 ;
      RECT 15.558 28.9345 15.63 28.9595 ;
      RECT 15.558 30.1345 15.63 30.1595 ;
      RECT 15.558 31.3345 15.63 31.3595 ;
      RECT 15.558 32.2675 15.63 32.2925 ;
      RECT 15.558 33.4675 15.63 33.4925 ;
      RECT 15.558 37.7875 15.63 37.8125 ;
      RECT 15.558 39.2275 15.63 39.2525 ;
      RECT 15.558 40.4545 15.63 40.4795 ;
      RECT 15.558 41.6545 15.63 41.6795 ;
      RECT 15.558 42.8545 15.63 42.8795 ;
      RECT 15.558 44.0545 15.63 44.0795 ;
      RECT 15.558 45.2545 15.63 45.2795 ;
      RECT 15.558 46.4545 15.63 46.4795 ;
      RECT 15.558 47.6545 15.63 47.6795 ;
      RECT 15.558 48.8545 15.63 48.8795 ;
      RECT 15.558 50.0545 15.63 50.0795 ;
      RECT 15.558 51.2545 15.63 51.2795 ;
      RECT 15.558 52.4545 15.63 52.4795 ;
      RECT 15.558 53.6545 15.63 53.6795 ;
      RECT 15.558 54.8545 15.63 54.8795 ;
      RECT 15.558 56.0545 15.63 56.0795 ;
      RECT 15.558 57.2545 15.63 57.2795 ;
      RECT 15.558 58.4545 15.63 58.4795 ;
      RECT 15.558 59.6545 15.63 59.6795 ;
      RECT 15.558 60.8545 15.63 60.8795 ;
      RECT 15.558 62.0545 15.63 62.0795 ;
      RECT 15.558 63.2545 15.63 63.2795 ;
      RECT 15.558 64.4545 15.63 64.4795 ;
      RECT 15.558 65.6545 15.63 65.6795 ;
      RECT 15.558 66.8545 15.63 66.8795 ;
      RECT 15.558 68.0545 15.63 68.0795 ;
      RECT 15.558 69.2545 15.63 69.2795 ;
      RECT 15.558 70.4545 15.63 70.4795 ;
      RECT 15.558 71.6545 15.63 71.6795 ;
      RECT 15.738 33.222 15.778 33.258 ;
      RECT 15.738 35.6835 15.778 35.7195 ;
      RECT 15.738 38.262 15.778 38.298 ;
      RECT 15.806 32.982 15.846 33.018 ;
      RECT 15.806 37.302 15.846 37.338 ;
      RECT 16.114 1.558 16.162 1.594 ;
      RECT 16.114 2.758 16.162 2.794 ;
      RECT 16.114 3.958 16.162 3.994 ;
      RECT 16.114 5.158 16.162 5.194 ;
      RECT 16.114 6.358 16.162 6.394 ;
      RECT 16.114 7.558 16.162 7.594 ;
      RECT 16.114 8.758 16.162 8.794 ;
      RECT 16.114 9.958 16.162 9.994 ;
      RECT 16.114 11.158 16.162 11.194 ;
      RECT 16.114 12.358 16.162 12.394 ;
      RECT 16.114 13.558 16.162 13.594 ;
      RECT 16.114 14.758 16.162 14.794 ;
      RECT 16.114 15.958 16.162 15.994 ;
      RECT 16.114 17.158 16.162 17.194 ;
      RECT 16.114 18.358 16.162 18.394 ;
      RECT 16.114 19.558 16.162 19.594 ;
      RECT 16.114 20.758 16.162 20.794 ;
      RECT 16.114 21.958 16.162 21.994 ;
      RECT 16.114 23.158 16.162 23.194 ;
      RECT 16.114 24.358 16.162 24.394 ;
      RECT 16.114 25.558 16.162 25.594 ;
      RECT 16.114 26.758 16.162 26.794 ;
      RECT 16.114 27.958 16.162 27.994 ;
      RECT 16.114 29.158 16.162 29.194 ;
      RECT 16.114 30.358 16.162 30.394 ;
      RECT 16.114 31.558 16.162 31.594 ;
      RECT 16.114 32.742 16.162 32.778 ;
      RECT 16.114 38.9205 16.162 38.9565 ;
      RECT 16.114 40.678 16.162 40.714 ;
      RECT 16.114 41.878 16.162 41.914 ;
      RECT 16.114 43.078 16.162 43.114 ;
      RECT 16.114 44.278 16.162 44.314 ;
      RECT 16.114 45.478 16.162 45.514 ;
      RECT 16.114 46.678 16.162 46.714 ;
      RECT 16.114 47.878 16.162 47.914 ;
      RECT 16.114 49.078 16.162 49.114 ;
      RECT 16.114 50.278 16.162 50.314 ;
      RECT 16.114 51.478 16.162 51.514 ;
      RECT 16.114 52.678 16.162 52.714 ;
      RECT 16.114 53.878 16.162 53.914 ;
      RECT 16.114 55.078 16.162 55.114 ;
      RECT 16.114 56.278 16.162 56.314 ;
      RECT 16.114 57.478 16.162 57.514 ;
      RECT 16.114 58.678 16.162 58.714 ;
      RECT 16.114 59.878 16.162 59.914 ;
      RECT 16.114 61.078 16.162 61.114 ;
      RECT 16.114 62.278 16.162 62.314 ;
      RECT 16.114 63.478 16.162 63.514 ;
      RECT 16.114 64.678 16.162 64.714 ;
      RECT 16.114 65.878 16.162 65.914 ;
      RECT 16.114 67.078 16.162 67.114 ;
      RECT 16.114 68.278 16.162 68.314 ;
      RECT 16.114 69.478 16.162 69.514 ;
      RECT 16.114 70.678 16.162 70.714 ;
      RECT 16.114 71.878 16.162 71.914 ;
      RECT 16.19 1.035 16.238 1.071 ;
      RECT 16.19 2.235 16.238 2.271 ;
      RECT 16.19 3.435 16.238 3.471 ;
      RECT 16.19 4.635 16.238 4.671 ;
      RECT 16.19 5.835 16.238 5.871 ;
      RECT 16.19 7.035 16.238 7.071 ;
      RECT 16.19 8.235 16.238 8.271 ;
      RECT 16.19 9.435 16.238 9.471 ;
      RECT 16.19 10.635 16.238 10.671 ;
      RECT 16.19 11.835 16.238 11.871 ;
      RECT 16.19 13.035 16.238 13.071 ;
      RECT 16.19 14.235 16.238 14.271 ;
      RECT 16.19 15.435 16.238 15.471 ;
      RECT 16.19 16.635 16.238 16.671 ;
      RECT 16.19 17.835 16.238 17.871 ;
      RECT 16.19 19.035 16.238 19.071 ;
      RECT 16.19 20.235 16.238 20.271 ;
      RECT 16.19 21.435 16.238 21.471 ;
      RECT 16.19 22.635 16.238 22.671 ;
      RECT 16.19 23.835 16.238 23.871 ;
      RECT 16.19 25.035 16.238 25.071 ;
      RECT 16.19 26.235 16.238 26.271 ;
      RECT 16.19 27.435 16.238 27.471 ;
      RECT 16.19 28.635 16.238 28.671 ;
      RECT 16.19 29.835 16.238 29.871 ;
      RECT 16.19 31.035 16.238 31.071 ;
      RECT 16.19 32.502 16.238 32.538 ;
      RECT 16.19 33.222 16.238 33.258 ;
      RECT 16.19 37.2405 16.238 37.2765 ;
      RECT 16.19 38.4405 16.238 38.4765 ;
      RECT 16.19 38.742 16.238 38.778 ;
      RECT 16.19 40.155 16.238 40.191 ;
      RECT 16.19 41.355 16.238 41.391 ;
      RECT 16.19 42.555 16.238 42.591 ;
      RECT 16.19 43.755 16.238 43.791 ;
      RECT 16.19 44.955 16.238 44.991 ;
      RECT 16.19 46.155 16.238 46.191 ;
      RECT 16.19 47.355 16.238 47.391 ;
      RECT 16.19 48.555 16.238 48.591 ;
      RECT 16.19 49.755 16.238 49.791 ;
      RECT 16.19 50.955 16.238 50.991 ;
      RECT 16.19 52.155 16.238 52.191 ;
      RECT 16.19 53.355 16.238 53.391 ;
      RECT 16.19 54.555 16.238 54.591 ;
      RECT 16.19 55.755 16.238 55.791 ;
      RECT 16.19 56.955 16.238 56.991 ;
      RECT 16.19 58.155 16.238 58.191 ;
      RECT 16.19 59.355 16.238 59.391 ;
      RECT 16.19 60.555 16.238 60.591 ;
      RECT 16.19 61.755 16.238 61.791 ;
      RECT 16.19 62.955 16.238 62.991 ;
      RECT 16.19 64.155 16.238 64.191 ;
      RECT 16.19 65.355 16.238 65.391 ;
      RECT 16.19 66.555 16.238 66.591 ;
      RECT 16.19 67.755 16.238 67.791 ;
      RECT 16.19 68.955 16.238 68.991 ;
      RECT 16.19 70.155 16.238 70.191 ;
      RECT 16.19 71.355 16.238 71.391 ;
      RECT 16.346 1.329 16.394 1.365 ;
      RECT 16.346 2.529 16.394 2.565 ;
      RECT 16.346 3.729 16.394 3.765 ;
      RECT 16.346 4.929 16.394 4.965 ;
      RECT 16.346 6.129 16.394 6.165 ;
      RECT 16.346 7.329 16.394 7.365 ;
      RECT 16.346 8.529 16.394 8.565 ;
      RECT 16.346 9.729 16.394 9.765 ;
      RECT 16.346 10.929 16.394 10.965 ;
      RECT 16.346 12.129 16.394 12.165 ;
      RECT 16.346 13.329 16.394 13.365 ;
      RECT 16.346 14.529 16.394 14.565 ;
      RECT 16.346 15.729 16.394 15.765 ;
      RECT 16.346 16.929 16.394 16.965 ;
      RECT 16.346 18.129 16.394 18.165 ;
      RECT 16.346 19.329 16.394 19.365 ;
      RECT 16.346 20.529 16.394 20.565 ;
      RECT 16.346 21.729 16.394 21.765 ;
      RECT 16.346 22.929 16.394 22.965 ;
      RECT 16.346 24.129 16.394 24.165 ;
      RECT 16.346 25.329 16.394 25.365 ;
      RECT 16.346 26.529 16.394 26.565 ;
      RECT 16.346 27.729 16.394 27.765 ;
      RECT 16.346 28.929 16.394 28.965 ;
      RECT 16.346 30.129 16.394 30.165 ;
      RECT 16.346 31.329 16.394 31.365 ;
      RECT 16.346 32.6805 16.394 32.7165 ;
      RECT 16.346 33.222 16.394 33.258 ;
      RECT 16.346 35.622 16.394 35.658 ;
      RECT 16.346 38.262 16.394 38.298 ;
      RECT 16.346 38.982 16.394 39.018 ;
      RECT 16.346 40.449 16.394 40.485 ;
      RECT 16.346 41.649 16.394 41.685 ;
      RECT 16.346 42.849 16.394 42.885 ;
      RECT 16.346 44.049 16.394 44.085 ;
      RECT 16.346 45.249 16.394 45.285 ;
      RECT 16.346 46.449 16.394 46.485 ;
      RECT 16.346 47.649 16.394 47.685 ;
      RECT 16.346 48.849 16.394 48.885 ;
      RECT 16.346 50.049 16.394 50.085 ;
      RECT 16.346 51.249 16.394 51.285 ;
      RECT 16.346 52.449 16.394 52.485 ;
      RECT 16.346 53.649 16.394 53.685 ;
      RECT 16.346 54.849 16.394 54.885 ;
      RECT 16.346 56.049 16.394 56.085 ;
      RECT 16.346 57.249 16.394 57.285 ;
      RECT 16.346 58.449 16.394 58.485 ;
      RECT 16.346 59.649 16.394 59.685 ;
      RECT 16.346 60.849 16.394 60.885 ;
      RECT 16.346 62.049 16.394 62.085 ;
      RECT 16.346 63.249 16.394 63.285 ;
      RECT 16.346 64.449 16.394 64.485 ;
      RECT 16.346 65.649 16.394 65.685 ;
      RECT 16.346 66.849 16.394 66.885 ;
      RECT 16.346 68.049 16.394 68.085 ;
      RECT 16.346 69.249 16.394 69.285 ;
      RECT 16.346 70.449 16.394 70.485 ;
      RECT 16.346 71.649 16.394 71.685 ;
      RECT 16.422 1.558 16.47 1.594 ;
      RECT 16.422 2.758 16.47 2.794 ;
      RECT 16.422 3.958 16.47 3.994 ;
      RECT 16.422 5.158 16.47 5.194 ;
      RECT 16.422 6.358 16.47 6.394 ;
      RECT 16.422 7.558 16.47 7.594 ;
      RECT 16.422 8.758 16.47 8.794 ;
      RECT 16.422 9.958 16.47 9.994 ;
      RECT 16.422 11.158 16.47 11.194 ;
      RECT 16.422 12.358 16.47 12.394 ;
      RECT 16.422 13.558 16.47 13.594 ;
      RECT 16.422 14.758 16.47 14.794 ;
      RECT 16.422 15.958 16.47 15.994 ;
      RECT 16.422 17.158 16.47 17.194 ;
      RECT 16.422 18.358 16.47 18.394 ;
      RECT 16.422 19.558 16.47 19.594 ;
      RECT 16.422 20.758 16.47 20.794 ;
      RECT 16.422 21.958 16.47 21.994 ;
      RECT 16.422 23.158 16.47 23.194 ;
      RECT 16.422 24.358 16.47 24.394 ;
      RECT 16.422 25.558 16.47 25.594 ;
      RECT 16.422 26.758 16.47 26.794 ;
      RECT 16.422 27.958 16.47 27.994 ;
      RECT 16.422 29.158 16.47 29.194 ;
      RECT 16.422 30.358 16.47 30.394 ;
      RECT 16.422 31.558 16.47 31.594 ;
      RECT 16.422 32.4405 16.47 32.4765 ;
      RECT 16.422 34.902 16.47 34.938 ;
      RECT 16.422 37.1235 16.47 37.1595 ;
      RECT 16.422 38.6805 16.47 38.7165 ;
      RECT 16.422 40.678 16.47 40.714 ;
      RECT 16.422 41.878 16.47 41.914 ;
      RECT 16.422 43.078 16.47 43.114 ;
      RECT 16.422 44.278 16.47 44.314 ;
      RECT 16.422 45.478 16.47 45.514 ;
      RECT 16.422 46.678 16.47 46.714 ;
      RECT 16.422 47.878 16.47 47.914 ;
      RECT 16.422 49.078 16.47 49.114 ;
      RECT 16.422 50.278 16.47 50.314 ;
      RECT 16.422 51.478 16.47 51.514 ;
      RECT 16.422 52.678 16.47 52.714 ;
      RECT 16.422 53.878 16.47 53.914 ;
      RECT 16.422 55.078 16.47 55.114 ;
      RECT 16.422 56.278 16.47 56.314 ;
      RECT 16.422 57.478 16.47 57.514 ;
      RECT 16.422 58.678 16.47 58.714 ;
      RECT 16.422 59.878 16.47 59.914 ;
      RECT 16.422 61.078 16.47 61.114 ;
      RECT 16.422 62.278 16.47 62.314 ;
      RECT 16.422 63.478 16.47 63.514 ;
      RECT 16.422 64.678 16.47 64.714 ;
      RECT 16.422 65.878 16.47 65.914 ;
      RECT 16.422 67.078 16.47 67.114 ;
      RECT 16.422 68.278 16.47 68.314 ;
      RECT 16.422 69.478 16.47 69.514 ;
      RECT 16.422 70.678 16.47 70.714 ;
      RECT 16.422 71.878 16.47 71.914 ;
      RECT 16.65 32.9205 16.69 32.9565 ;
      RECT 16.718 1.329 16.772 1.365 ;
      RECT 16.718 2.529 16.772 2.565 ;
      RECT 16.718 3.729 16.772 3.765 ;
      RECT 16.718 4.929 16.772 4.965 ;
      RECT 16.718 6.129 16.772 6.165 ;
      RECT 16.718 7.329 16.772 7.365 ;
      RECT 16.718 8.529 16.772 8.565 ;
      RECT 16.718 9.729 16.772 9.765 ;
      RECT 16.718 10.929 16.772 10.965 ;
      RECT 16.718 12.129 16.772 12.165 ;
      RECT 16.718 13.329 16.772 13.365 ;
      RECT 16.718 14.529 16.772 14.565 ;
      RECT 16.718 15.729 16.772 15.765 ;
      RECT 16.718 16.929 16.772 16.965 ;
      RECT 16.718 18.129 16.772 18.165 ;
      RECT 16.718 19.329 16.772 19.365 ;
      RECT 16.718 20.529 16.772 20.565 ;
      RECT 16.718 21.729 16.772 21.765 ;
      RECT 16.718 22.929 16.772 22.965 ;
      RECT 16.718 24.129 16.772 24.165 ;
      RECT 16.718 25.329 16.772 25.365 ;
      RECT 16.718 26.529 16.772 26.565 ;
      RECT 16.718 27.729 16.772 27.765 ;
      RECT 16.718 28.929 16.772 28.965 ;
      RECT 16.718 30.129 16.772 30.165 ;
      RECT 16.718 31.329 16.772 31.365 ;
      RECT 16.718 32.2005 16.772 32.2365 ;
      RECT 16.718 39.2835 16.772 39.3195 ;
      RECT 16.718 40.449 16.772 40.485 ;
      RECT 16.718 41.649 16.772 41.685 ;
      RECT 16.718 42.849 16.772 42.885 ;
      RECT 16.718 44.049 16.772 44.085 ;
      RECT 16.718 45.249 16.772 45.285 ;
      RECT 16.718 46.449 16.772 46.485 ;
      RECT 16.718 47.649 16.772 47.685 ;
      RECT 16.718 48.849 16.772 48.885 ;
      RECT 16.718 50.049 16.772 50.085 ;
      RECT 16.718 51.249 16.772 51.285 ;
      RECT 16.718 52.449 16.772 52.485 ;
      RECT 16.718 53.649 16.772 53.685 ;
      RECT 16.718 54.849 16.772 54.885 ;
      RECT 16.718 56.049 16.772 56.085 ;
      RECT 16.718 57.249 16.772 57.285 ;
      RECT 16.718 58.449 16.772 58.485 ;
      RECT 16.718 59.649 16.772 59.685 ;
      RECT 16.718 60.849 16.772 60.885 ;
      RECT 16.718 62.049 16.772 62.085 ;
      RECT 16.718 63.249 16.772 63.285 ;
      RECT 16.718 64.449 16.772 64.485 ;
      RECT 16.718 65.649 16.772 65.685 ;
      RECT 16.718 66.849 16.772 66.885 ;
      RECT 16.718 68.049 16.772 68.085 ;
      RECT 16.718 69.249 16.772 69.285 ;
      RECT 16.718 70.449 16.772 70.485 ;
      RECT 16.718 71.649 16.772 71.685 ;
      RECT 16.882 1.558 16.936 1.594 ;
      RECT 16.882 2.758 16.936 2.794 ;
      RECT 16.882 3.958 16.936 3.994 ;
      RECT 16.882 5.158 16.936 5.194 ;
      RECT 16.882 6.358 16.936 6.394 ;
      RECT 16.882 7.558 16.936 7.594 ;
      RECT 16.882 8.758 16.936 8.794 ;
      RECT 16.882 9.958 16.936 9.994 ;
      RECT 16.882 11.158 16.936 11.194 ;
      RECT 16.882 12.358 16.936 12.394 ;
      RECT 16.882 13.558 16.936 13.594 ;
      RECT 16.882 14.758 16.936 14.794 ;
      RECT 16.882 15.958 16.936 15.994 ;
      RECT 16.882 17.158 16.936 17.194 ;
      RECT 16.882 18.358 16.936 18.394 ;
      RECT 16.882 19.558 16.936 19.594 ;
      RECT 16.882 20.758 16.936 20.794 ;
      RECT 16.882 21.958 16.936 21.994 ;
      RECT 16.882 23.158 16.936 23.194 ;
      RECT 16.882 24.358 16.936 24.394 ;
      RECT 16.882 25.558 16.936 25.594 ;
      RECT 16.882 26.758 16.936 26.794 ;
      RECT 16.882 27.958 16.936 27.994 ;
      RECT 16.882 29.158 16.936 29.194 ;
      RECT 16.882 30.358 16.936 30.394 ;
      RECT 16.882 31.558 16.936 31.594 ;
      RECT 16.882 32.2005 16.936 32.2365 ;
      RECT 16.882 39.2835 16.936 39.3195 ;
      RECT 16.882 40.678 16.936 40.714 ;
      RECT 16.882 41.878 16.936 41.914 ;
      RECT 16.882 43.078 16.936 43.114 ;
      RECT 16.882 44.278 16.936 44.314 ;
      RECT 16.882 45.478 16.936 45.514 ;
      RECT 16.882 46.678 16.936 46.714 ;
      RECT 16.882 47.878 16.936 47.914 ;
      RECT 16.882 49.078 16.936 49.114 ;
      RECT 16.882 50.278 16.936 50.314 ;
      RECT 16.882 51.478 16.936 51.514 ;
      RECT 16.882 52.678 16.936 52.714 ;
      RECT 16.882 53.878 16.936 53.914 ;
      RECT 16.882 55.078 16.936 55.114 ;
      RECT 16.882 56.278 16.936 56.314 ;
      RECT 16.882 57.478 16.936 57.514 ;
      RECT 16.882 58.678 16.936 58.714 ;
      RECT 16.882 59.878 16.936 59.914 ;
      RECT 16.882 61.078 16.936 61.114 ;
      RECT 16.882 62.278 16.936 62.314 ;
      RECT 16.882 63.478 16.936 63.514 ;
      RECT 16.882 64.678 16.936 64.714 ;
      RECT 16.882 65.878 16.936 65.914 ;
      RECT 16.882 67.078 16.936 67.114 ;
      RECT 16.882 68.278 16.936 68.314 ;
      RECT 16.882 69.478 16.936 69.514 ;
      RECT 16.882 70.678 16.936 70.714 ;
      RECT 16.882 71.878 16.936 71.914 ;
      RECT 17.136 32.622 17.176 32.658 ;
      RECT 17.136 32.742 17.176 32.778 ;
      RECT 17.548 1.035 17.588 1.071 ;
      RECT 17.548 2.235 17.588 2.271 ;
      RECT 17.548 3.435 17.588 3.471 ;
      RECT 17.548 4.635 17.588 4.671 ;
      RECT 17.548 5.835 17.588 5.871 ;
      RECT 17.548 7.035 17.588 7.071 ;
      RECT 17.548 8.235 17.588 8.271 ;
      RECT 17.548 9.435 17.588 9.471 ;
      RECT 17.548 10.635 17.588 10.671 ;
      RECT 17.548 11.835 17.588 11.871 ;
      RECT 17.548 13.035 17.588 13.071 ;
      RECT 17.548 14.235 17.588 14.271 ;
      RECT 17.548 15.435 17.588 15.471 ;
      RECT 17.548 16.635 17.588 16.671 ;
      RECT 17.548 17.835 17.588 17.871 ;
      RECT 17.548 19.035 17.588 19.071 ;
      RECT 17.548 20.235 17.588 20.271 ;
      RECT 17.548 21.435 17.588 21.471 ;
      RECT 17.548 22.635 17.588 22.671 ;
      RECT 17.548 23.835 17.588 23.871 ;
      RECT 17.548 25.035 17.588 25.071 ;
      RECT 17.548 26.235 17.588 26.271 ;
      RECT 17.548 27.435 17.588 27.471 ;
      RECT 17.548 28.635 17.588 28.671 ;
      RECT 17.548 29.835 17.588 29.871 ;
      RECT 17.548 31.035 17.588 31.071 ;
      RECT 17.548 38.982 17.588 39.018 ;
      RECT 17.548 40.155 17.588 40.191 ;
      RECT 17.548 41.355 17.588 41.391 ;
      RECT 17.548 42.555 17.588 42.591 ;
      RECT 17.548 43.755 17.588 43.791 ;
      RECT 17.548 44.955 17.588 44.991 ;
      RECT 17.548 46.155 17.588 46.191 ;
      RECT 17.548 47.355 17.588 47.391 ;
      RECT 17.548 48.555 17.588 48.591 ;
      RECT 17.548 49.755 17.588 49.791 ;
      RECT 17.548 50.955 17.588 50.991 ;
      RECT 17.548 52.155 17.588 52.191 ;
      RECT 17.548 53.355 17.588 53.391 ;
      RECT 17.548 54.555 17.588 54.591 ;
      RECT 17.548 55.755 17.588 55.791 ;
      RECT 17.548 56.955 17.588 56.991 ;
      RECT 17.548 58.155 17.588 58.191 ;
      RECT 17.548 59.355 17.588 59.391 ;
      RECT 17.548 60.555 17.588 60.591 ;
      RECT 17.548 61.755 17.588 61.791 ;
      RECT 17.548 62.955 17.588 62.991 ;
      RECT 17.548 64.155 17.588 64.191 ;
      RECT 17.548 65.355 17.588 65.391 ;
      RECT 17.548 66.555 17.588 66.591 ;
      RECT 17.548 67.755 17.588 67.791 ;
      RECT 17.548 68.955 17.588 68.991 ;
      RECT 17.548 70.155 17.588 70.191 ;
      RECT 17.548 71.355 17.588 71.391 ;
      RECT 17.616 1.035 17.656 1.071 ;
      RECT 17.616 2.235 17.656 2.271 ;
      RECT 17.616 3.435 17.656 3.471 ;
      RECT 17.616 4.635 17.656 4.671 ;
      RECT 17.616 5.835 17.656 5.871 ;
      RECT 17.616 7.035 17.656 7.071 ;
      RECT 17.616 8.235 17.656 8.271 ;
      RECT 17.616 9.435 17.656 9.471 ;
      RECT 17.616 10.635 17.656 10.671 ;
      RECT 17.616 11.835 17.656 11.871 ;
      RECT 17.616 13.035 17.656 13.071 ;
      RECT 17.616 14.235 17.656 14.271 ;
      RECT 17.616 15.435 17.656 15.471 ;
      RECT 17.616 16.635 17.656 16.671 ;
      RECT 17.616 17.835 17.656 17.871 ;
      RECT 17.616 19.035 17.656 19.071 ;
      RECT 17.616 20.235 17.656 20.271 ;
      RECT 17.616 21.435 17.656 21.471 ;
      RECT 17.616 22.635 17.656 22.671 ;
      RECT 17.616 23.835 17.656 23.871 ;
      RECT 17.616 25.035 17.656 25.071 ;
      RECT 17.616 26.235 17.656 26.271 ;
      RECT 17.616 27.435 17.656 27.471 ;
      RECT 17.616 28.635 17.656 28.671 ;
      RECT 17.616 29.835 17.656 29.871 ;
      RECT 17.616 31.035 17.656 31.071 ;
      RECT 17.616 33.4005 17.656 33.4365 ;
      RECT 17.616 33.582 17.656 33.618 ;
      RECT 17.616 34.062 17.656 34.098 ;
      RECT 17.616 38.982 17.656 39.018 ;
      RECT 17.616 40.155 17.656 40.191 ;
      RECT 17.616 41.355 17.656 41.391 ;
      RECT 17.616 42.555 17.656 42.591 ;
      RECT 17.616 43.755 17.656 43.791 ;
      RECT 17.616 44.955 17.656 44.991 ;
      RECT 17.616 46.155 17.656 46.191 ;
      RECT 17.616 47.355 17.656 47.391 ;
      RECT 17.616 48.555 17.656 48.591 ;
      RECT 17.616 49.755 17.656 49.791 ;
      RECT 17.616 50.955 17.656 50.991 ;
      RECT 17.616 52.155 17.656 52.191 ;
      RECT 17.616 53.355 17.656 53.391 ;
      RECT 17.616 54.555 17.656 54.591 ;
      RECT 17.616 55.755 17.656 55.791 ;
      RECT 17.616 56.955 17.656 56.991 ;
      RECT 17.616 58.155 17.656 58.191 ;
      RECT 17.616 59.355 17.656 59.391 ;
      RECT 17.616 60.555 17.656 60.591 ;
      RECT 17.616 61.755 17.656 61.791 ;
      RECT 17.616 62.955 17.656 62.991 ;
      RECT 17.616 64.155 17.656 64.191 ;
      RECT 17.616 65.355 17.656 65.391 ;
      RECT 17.616 66.555 17.656 66.591 ;
      RECT 17.616 67.755 17.656 67.791 ;
      RECT 17.616 68.955 17.656 68.991 ;
      RECT 17.616 70.155 17.656 70.191 ;
      RECT 17.616 71.355 17.656 71.391 ;
      RECT 17.944 32.502 17.984 32.538 ;
      RECT 17.944 32.622 17.984 32.658 ;
      RECT 17.944 32.9205 17.984 32.9565 ;
      RECT 17.944 34.422 17.984 34.458 ;
      RECT 17.944 34.542 17.984 34.578 ;
      RECT 17.944 35.022 17.984 35.058 ;
      RECT 18.012 1.329 18.052 1.365 ;
      RECT 18.012 2.529 18.052 2.565 ;
      RECT 18.012 3.729 18.052 3.765 ;
      RECT 18.012 4.929 18.052 4.965 ;
      RECT 18.012 6.129 18.052 6.165 ;
      RECT 18.012 7.329 18.052 7.365 ;
      RECT 18.012 8.529 18.052 8.565 ;
      RECT 18.012 9.729 18.052 9.765 ;
      RECT 18.012 10.929 18.052 10.965 ;
      RECT 18.012 12.129 18.052 12.165 ;
      RECT 18.012 13.329 18.052 13.365 ;
      RECT 18.012 14.529 18.052 14.565 ;
      RECT 18.012 15.729 18.052 15.765 ;
      RECT 18.012 16.929 18.052 16.965 ;
      RECT 18.012 18.129 18.052 18.165 ;
      RECT 18.012 19.329 18.052 19.365 ;
      RECT 18.012 20.529 18.052 20.565 ;
      RECT 18.012 21.729 18.052 21.765 ;
      RECT 18.012 22.929 18.052 22.965 ;
      RECT 18.012 24.129 18.052 24.165 ;
      RECT 18.012 25.329 18.052 25.365 ;
      RECT 18.012 26.529 18.052 26.565 ;
      RECT 18.012 27.729 18.052 27.765 ;
      RECT 18.012 28.929 18.052 28.965 ;
      RECT 18.012 30.129 18.052 30.165 ;
      RECT 18.012 31.329 18.052 31.365 ;
      RECT 18.012 38.982 18.052 39.018 ;
      RECT 18.012 40.449 18.052 40.485 ;
      RECT 18.012 41.649 18.052 41.685 ;
      RECT 18.012 42.849 18.052 42.885 ;
      RECT 18.012 44.049 18.052 44.085 ;
      RECT 18.012 45.249 18.052 45.285 ;
      RECT 18.012 46.449 18.052 46.485 ;
      RECT 18.012 47.649 18.052 47.685 ;
      RECT 18.012 48.849 18.052 48.885 ;
      RECT 18.012 50.049 18.052 50.085 ;
      RECT 18.012 51.249 18.052 51.285 ;
      RECT 18.012 52.449 18.052 52.485 ;
      RECT 18.012 53.649 18.052 53.685 ;
      RECT 18.012 54.849 18.052 54.885 ;
      RECT 18.012 56.049 18.052 56.085 ;
      RECT 18.012 57.249 18.052 57.285 ;
      RECT 18.012 58.449 18.052 58.485 ;
      RECT 18.012 59.649 18.052 59.685 ;
      RECT 18.012 60.849 18.052 60.885 ;
      RECT 18.012 62.049 18.052 62.085 ;
      RECT 18.012 63.249 18.052 63.285 ;
      RECT 18.012 64.449 18.052 64.485 ;
      RECT 18.012 65.649 18.052 65.685 ;
      RECT 18.012 66.849 18.052 66.885 ;
      RECT 18.012 68.049 18.052 68.085 ;
      RECT 18.012 69.249 18.052 69.285 ;
      RECT 18.012 70.449 18.052 70.485 ;
      RECT 18.012 71.649 18.052 71.685 ;
      RECT 18.08 1.329 18.12 1.365 ;
      RECT 18.08 2.529 18.12 2.565 ;
      RECT 18.08 3.729 18.12 3.765 ;
      RECT 18.08 4.929 18.12 4.965 ;
      RECT 18.08 6.129 18.12 6.165 ;
      RECT 18.08 7.329 18.12 7.365 ;
      RECT 18.08 8.529 18.12 8.565 ;
      RECT 18.08 9.729 18.12 9.765 ;
      RECT 18.08 10.929 18.12 10.965 ;
      RECT 18.08 12.129 18.12 12.165 ;
      RECT 18.08 13.329 18.12 13.365 ;
      RECT 18.08 14.529 18.12 14.565 ;
      RECT 18.08 15.729 18.12 15.765 ;
      RECT 18.08 16.929 18.12 16.965 ;
      RECT 18.08 18.129 18.12 18.165 ;
      RECT 18.08 19.329 18.12 19.365 ;
      RECT 18.08 20.529 18.12 20.565 ;
      RECT 18.08 21.729 18.12 21.765 ;
      RECT 18.08 22.929 18.12 22.965 ;
      RECT 18.08 24.129 18.12 24.165 ;
      RECT 18.08 25.329 18.12 25.365 ;
      RECT 18.08 26.529 18.12 26.565 ;
      RECT 18.08 27.729 18.12 27.765 ;
      RECT 18.08 28.929 18.12 28.965 ;
      RECT 18.08 30.129 18.12 30.165 ;
      RECT 18.08 31.329 18.12 31.365 ;
      RECT 18.08 38.982 18.12 39.018 ;
      RECT 18.08 40.449 18.12 40.485 ;
      RECT 18.08 41.649 18.12 41.685 ;
      RECT 18.08 42.849 18.12 42.885 ;
      RECT 18.08 44.049 18.12 44.085 ;
      RECT 18.08 45.249 18.12 45.285 ;
      RECT 18.08 46.449 18.12 46.485 ;
      RECT 18.08 47.649 18.12 47.685 ;
      RECT 18.08 48.849 18.12 48.885 ;
      RECT 18.08 50.049 18.12 50.085 ;
      RECT 18.08 51.249 18.12 51.285 ;
      RECT 18.08 52.449 18.12 52.485 ;
      RECT 18.08 53.649 18.12 53.685 ;
      RECT 18.08 54.849 18.12 54.885 ;
      RECT 18.08 56.049 18.12 56.085 ;
      RECT 18.08 57.249 18.12 57.285 ;
      RECT 18.08 58.449 18.12 58.485 ;
      RECT 18.08 59.649 18.12 59.685 ;
      RECT 18.08 60.849 18.12 60.885 ;
      RECT 18.08 62.049 18.12 62.085 ;
      RECT 18.08 63.249 18.12 63.285 ;
      RECT 18.08 64.449 18.12 64.485 ;
      RECT 18.08 65.649 18.12 65.685 ;
      RECT 18.08 66.849 18.12 66.885 ;
      RECT 18.08 68.049 18.12 68.085 ;
      RECT 18.08 69.249 18.12 69.285 ;
      RECT 18.08 70.449 18.12 70.485 ;
      RECT 18.08 71.649 18.12 71.685 ;
      RECT 18.492 32.502 18.536 32.538 ;
      RECT 18.764 1.1875 18.836 1.2125 ;
      RECT 18.764 1.3345 18.836 1.3595 ;
      RECT 18.764 2.3875 18.836 2.4125 ;
      RECT 18.764 2.5345 18.836 2.5595 ;
      RECT 18.764 3.5875 18.836 3.6125 ;
      RECT 18.764 3.7345 18.836 3.7595 ;
      RECT 18.764 4.7875 18.836 4.8125 ;
      RECT 18.764 4.9345 18.836 4.9595 ;
      RECT 18.764 5.9875 18.836 6.0125 ;
      RECT 18.764 6.1345 18.836 6.1595 ;
      RECT 18.764 7.1875 18.836 7.2125 ;
      RECT 18.764 7.3345 18.836 7.3595 ;
      RECT 18.764 8.3875 18.836 8.4125 ;
      RECT 18.764 8.5345 18.836 8.5595 ;
      RECT 18.764 9.5875 18.836 9.6125 ;
      RECT 18.764 9.7345 18.836 9.7595 ;
      RECT 18.764 10.7875 18.836 10.8125 ;
      RECT 18.764 10.9345 18.836 10.9595 ;
      RECT 18.764 11.9875 18.836 12.0125 ;
      RECT 18.764 12.1345 18.836 12.1595 ;
      RECT 18.764 13.1875 18.836 13.2125 ;
      RECT 18.764 13.3345 18.836 13.3595 ;
      RECT 18.764 14.3875 18.836 14.4125 ;
      RECT 18.764 14.5345 18.836 14.5595 ;
      RECT 18.764 15.5875 18.836 15.6125 ;
      RECT 18.764 15.7345 18.836 15.7595 ;
      RECT 18.764 16.7875 18.836 16.8125 ;
      RECT 18.764 16.9345 18.836 16.9595 ;
      RECT 18.764 17.9875 18.836 18.0125 ;
      RECT 18.764 18.1345 18.836 18.1595 ;
      RECT 18.764 19.1875 18.836 19.2125 ;
      RECT 18.764 19.3345 18.836 19.3595 ;
      RECT 18.764 20.3875 18.836 20.4125 ;
      RECT 18.764 20.5345 18.836 20.5595 ;
      RECT 18.764 21.5875 18.836 21.6125 ;
      RECT 18.764 21.7345 18.836 21.7595 ;
      RECT 18.764 22.7875 18.836 22.8125 ;
      RECT 18.764 22.9345 18.836 22.9595 ;
      RECT 18.764 23.9875 18.836 24.0125 ;
      RECT 18.764 24.1345 18.836 24.1595 ;
      RECT 18.764 25.1875 18.836 25.2125 ;
      RECT 18.764 25.3345 18.836 25.3595 ;
      RECT 18.764 26.3875 18.836 26.4125 ;
      RECT 18.764 26.5345 18.836 26.5595 ;
      RECT 18.764 27.5875 18.836 27.6125 ;
      RECT 18.764 27.7345 18.836 27.7595 ;
      RECT 18.764 28.7875 18.836 28.8125 ;
      RECT 18.764 28.9345 18.836 28.9595 ;
      RECT 18.764 29.9875 18.836 30.0125 ;
      RECT 18.764 30.1345 18.836 30.1595 ;
      RECT 18.764 31.1875 18.836 31.2125 ;
      RECT 18.764 31.3345 18.836 31.3595 ;
      RECT 18.764 40.3075 18.836 40.3325 ;
      RECT 18.764 40.4545 18.836 40.4795 ;
      RECT 18.764 41.5075 18.836 41.5325 ;
      RECT 18.764 41.6545 18.836 41.6795 ;
      RECT 18.764 42.7075 18.836 42.7325 ;
      RECT 18.764 42.8545 18.836 42.8795 ;
      RECT 18.764 43.9075 18.836 43.9325 ;
      RECT 18.764 44.0545 18.836 44.0795 ;
      RECT 18.764 45.1075 18.836 45.1325 ;
      RECT 18.764 45.2545 18.836 45.2795 ;
      RECT 18.764 46.3075 18.836 46.3325 ;
      RECT 18.764 46.4545 18.836 46.4795 ;
      RECT 18.764 47.5075 18.836 47.5325 ;
      RECT 18.764 47.6545 18.836 47.6795 ;
      RECT 18.764 48.7075 18.836 48.7325 ;
      RECT 18.764 48.8545 18.836 48.8795 ;
      RECT 18.764 49.9075 18.836 49.9325 ;
      RECT 18.764 50.0545 18.836 50.0795 ;
      RECT 18.764 51.1075 18.836 51.1325 ;
      RECT 18.764 51.2545 18.836 51.2795 ;
      RECT 18.764 52.3075 18.836 52.3325 ;
      RECT 18.764 52.4545 18.836 52.4795 ;
      RECT 18.764 53.5075 18.836 53.5325 ;
      RECT 18.764 53.6545 18.836 53.6795 ;
      RECT 18.764 54.7075 18.836 54.7325 ;
      RECT 18.764 54.8545 18.836 54.8795 ;
      RECT 18.764 55.9075 18.836 55.9325 ;
      RECT 18.764 56.0545 18.836 56.0795 ;
      RECT 18.764 57.1075 18.836 57.1325 ;
      RECT 18.764 57.2545 18.836 57.2795 ;
      RECT 18.764 58.3075 18.836 58.3325 ;
      RECT 18.764 58.4545 18.836 58.4795 ;
      RECT 18.764 59.5075 18.836 59.5325 ;
      RECT 18.764 59.6545 18.836 59.6795 ;
      RECT 18.764 60.7075 18.836 60.7325 ;
      RECT 18.764 60.8545 18.836 60.8795 ;
      RECT 18.764 61.9075 18.836 61.9325 ;
      RECT 18.764 62.0545 18.836 62.0795 ;
      RECT 18.764 63.1075 18.836 63.1325 ;
      RECT 18.764 63.2545 18.836 63.2795 ;
      RECT 18.764 64.3075 18.836 64.3325 ;
      RECT 18.764 64.4545 18.836 64.4795 ;
      RECT 18.764 65.5075 18.836 65.5325 ;
      RECT 18.764 65.6545 18.836 65.6795 ;
      RECT 18.764 66.7075 18.836 66.7325 ;
      RECT 18.764 66.8545 18.836 66.8795 ;
      RECT 18.764 67.9075 18.836 67.9325 ;
      RECT 18.764 68.0545 18.836 68.0795 ;
      RECT 18.764 69.1075 18.836 69.1325 ;
      RECT 18.764 69.2545 18.836 69.2795 ;
      RECT 18.764 70.3075 18.836 70.3325 ;
      RECT 18.764 70.4545 18.836 70.4795 ;
      RECT 18.764 71.5075 18.836 71.5325 ;
      RECT 18.764 71.6545 18.836 71.6795 ;
      RECT 19.53 1.558 19.578 1.594 ;
      RECT 19.53 2.758 19.578 2.794 ;
      RECT 19.53 3.958 19.578 3.994 ;
      RECT 19.53 5.158 19.578 5.194 ;
      RECT 19.53 6.358 19.578 6.394 ;
      RECT 19.53 7.558 19.578 7.594 ;
      RECT 19.53 8.758 19.578 8.794 ;
      RECT 19.53 9.958 19.578 9.994 ;
      RECT 19.53 11.158 19.578 11.194 ;
      RECT 19.53 12.358 19.578 12.394 ;
      RECT 19.53 13.558 19.578 13.594 ;
      RECT 19.53 14.758 19.578 14.794 ;
      RECT 19.53 15.958 19.578 15.994 ;
      RECT 19.53 17.158 19.578 17.194 ;
      RECT 19.53 18.358 19.578 18.394 ;
      RECT 19.53 19.558 19.578 19.594 ;
      RECT 19.53 20.758 19.578 20.794 ;
      RECT 19.53 21.958 19.578 21.994 ;
      RECT 19.53 23.158 19.578 23.194 ;
      RECT 19.53 24.358 19.578 24.394 ;
      RECT 19.53 25.558 19.578 25.594 ;
      RECT 19.53 26.758 19.578 26.794 ;
      RECT 19.53 27.958 19.578 27.994 ;
      RECT 19.53 29.158 19.578 29.194 ;
      RECT 19.53 30.358 19.578 30.394 ;
      RECT 19.53 31.558 19.578 31.594 ;
      RECT 19.53 32.3235 19.578 32.3595 ;
      RECT 19.53 38.6805 19.578 38.7165 ;
      RECT 19.53 40.678 19.578 40.714 ;
      RECT 19.53 41.878 19.578 41.914 ;
      RECT 19.53 43.078 19.578 43.114 ;
      RECT 19.53 44.278 19.578 44.314 ;
      RECT 19.53 45.478 19.578 45.514 ;
      RECT 19.53 46.678 19.578 46.714 ;
      RECT 19.53 47.878 19.578 47.914 ;
      RECT 19.53 49.078 19.578 49.114 ;
      RECT 19.53 50.278 19.578 50.314 ;
      RECT 19.53 51.478 19.578 51.514 ;
      RECT 19.53 52.678 19.578 52.714 ;
      RECT 19.53 53.878 19.578 53.914 ;
      RECT 19.53 55.078 19.578 55.114 ;
      RECT 19.53 56.278 19.578 56.314 ;
      RECT 19.53 57.478 19.578 57.514 ;
      RECT 19.53 58.678 19.578 58.714 ;
      RECT 19.53 59.878 19.578 59.914 ;
      RECT 19.53 61.078 19.578 61.114 ;
      RECT 19.53 62.278 19.578 62.314 ;
      RECT 19.53 63.478 19.578 63.514 ;
      RECT 19.53 64.678 19.578 64.714 ;
      RECT 19.53 65.878 19.578 65.914 ;
      RECT 19.53 67.078 19.578 67.114 ;
      RECT 19.53 68.278 19.578 68.314 ;
      RECT 19.53 69.478 19.578 69.514 ;
      RECT 19.53 70.678 19.578 70.714 ;
      RECT 19.53 71.878 19.578 71.914 ;
      RECT 19.606 1.329 19.654 1.365 ;
      RECT 19.606 2.529 19.654 2.565 ;
      RECT 19.606 3.729 19.654 3.765 ;
      RECT 19.606 4.929 19.654 4.965 ;
      RECT 19.606 6.129 19.654 6.165 ;
      RECT 19.606 7.329 19.654 7.365 ;
      RECT 19.606 8.529 19.654 8.565 ;
      RECT 19.606 9.729 19.654 9.765 ;
      RECT 19.606 10.929 19.654 10.965 ;
      RECT 19.606 12.129 19.654 12.165 ;
      RECT 19.606 13.329 19.654 13.365 ;
      RECT 19.606 14.529 19.654 14.565 ;
      RECT 19.606 15.729 19.654 15.765 ;
      RECT 19.606 16.929 19.654 16.965 ;
      RECT 19.606 18.129 19.654 18.165 ;
      RECT 19.606 19.329 19.654 19.365 ;
      RECT 19.606 20.529 19.654 20.565 ;
      RECT 19.606 21.729 19.654 21.765 ;
      RECT 19.606 22.929 19.654 22.965 ;
      RECT 19.606 24.129 19.654 24.165 ;
      RECT 19.606 25.329 19.654 25.365 ;
      RECT 19.606 26.529 19.654 26.565 ;
      RECT 19.606 27.729 19.654 27.765 ;
      RECT 19.606 28.929 19.654 28.965 ;
      RECT 19.606 30.129 19.654 30.165 ;
      RECT 19.606 31.329 19.654 31.365 ;
      RECT 19.606 32.742 19.654 32.778 ;
      RECT 19.606 33.222 19.654 33.258 ;
      RECT 19.606 35.8005 19.654 35.8365 ;
      RECT 19.606 38.262 19.654 38.298 ;
      RECT 19.606 38.982 19.654 39.018 ;
      RECT 19.606 40.449 19.654 40.485 ;
      RECT 19.606 41.649 19.654 41.685 ;
      RECT 19.606 42.849 19.654 42.885 ;
      RECT 19.606 44.049 19.654 44.085 ;
      RECT 19.606 45.249 19.654 45.285 ;
      RECT 19.606 46.449 19.654 46.485 ;
      RECT 19.606 47.649 19.654 47.685 ;
      RECT 19.606 48.849 19.654 48.885 ;
      RECT 19.606 50.049 19.654 50.085 ;
      RECT 19.606 51.249 19.654 51.285 ;
      RECT 19.606 52.449 19.654 52.485 ;
      RECT 19.606 53.649 19.654 53.685 ;
      RECT 19.606 54.849 19.654 54.885 ;
      RECT 19.606 56.049 19.654 56.085 ;
      RECT 19.606 57.249 19.654 57.285 ;
      RECT 19.606 58.449 19.654 58.485 ;
      RECT 19.606 59.649 19.654 59.685 ;
      RECT 19.606 60.849 19.654 60.885 ;
      RECT 19.606 62.049 19.654 62.085 ;
      RECT 19.606 63.249 19.654 63.285 ;
      RECT 19.606 64.449 19.654 64.485 ;
      RECT 19.606 65.649 19.654 65.685 ;
      RECT 19.606 66.849 19.654 66.885 ;
      RECT 19.606 68.049 19.654 68.085 ;
      RECT 19.606 69.249 19.654 69.285 ;
      RECT 19.606 70.449 19.654 70.485 ;
      RECT 19.606 71.649 19.654 71.685 ;
      RECT 19.762 1.035 19.81 1.071 ;
      RECT 19.762 2.235 19.81 2.271 ;
      RECT 19.762 3.435 19.81 3.471 ;
      RECT 19.762 4.635 19.81 4.671 ;
      RECT 19.762 5.835 19.81 5.871 ;
      RECT 19.762 7.035 19.81 7.071 ;
      RECT 19.762 8.235 19.81 8.271 ;
      RECT 19.762 9.435 19.81 9.471 ;
      RECT 19.762 10.635 19.81 10.671 ;
      RECT 19.762 11.835 19.81 11.871 ;
      RECT 19.762 13.035 19.81 13.071 ;
      RECT 19.762 14.235 19.81 14.271 ;
      RECT 19.762 15.435 19.81 15.471 ;
      RECT 19.762 16.635 19.81 16.671 ;
      RECT 19.762 17.835 19.81 17.871 ;
      RECT 19.762 19.035 19.81 19.071 ;
      RECT 19.762 20.235 19.81 20.271 ;
      RECT 19.762 21.435 19.81 21.471 ;
      RECT 19.762 22.635 19.81 22.671 ;
      RECT 19.762 23.835 19.81 23.871 ;
      RECT 19.762 25.035 19.81 25.071 ;
      RECT 19.762 26.235 19.81 26.271 ;
      RECT 19.762 27.435 19.81 27.471 ;
      RECT 19.762 28.635 19.81 28.671 ;
      RECT 19.762 29.835 19.81 29.871 ;
      RECT 19.762 31.035 19.81 31.071 ;
      RECT 19.762 32.262 19.81 32.298 ;
      RECT 19.762 33.222 19.81 33.258 ;
      RECT 19.762 37.1235 19.81 37.1595 ;
      RECT 19.762 38.4405 19.81 38.4765 ;
      RECT 19.762 38.742 19.81 38.778 ;
      RECT 19.762 40.155 19.81 40.191 ;
      RECT 19.762 41.355 19.81 41.391 ;
      RECT 19.762 42.555 19.81 42.591 ;
      RECT 19.762 43.755 19.81 43.791 ;
      RECT 19.762 44.955 19.81 44.991 ;
      RECT 19.762 46.155 19.81 46.191 ;
      RECT 19.762 47.355 19.81 47.391 ;
      RECT 19.762 48.555 19.81 48.591 ;
      RECT 19.762 49.755 19.81 49.791 ;
      RECT 19.762 50.955 19.81 50.991 ;
      RECT 19.762 52.155 19.81 52.191 ;
      RECT 19.762 53.355 19.81 53.391 ;
      RECT 19.762 54.555 19.81 54.591 ;
      RECT 19.762 55.755 19.81 55.791 ;
      RECT 19.762 56.955 19.81 56.991 ;
      RECT 19.762 58.155 19.81 58.191 ;
      RECT 19.762 59.355 19.81 59.391 ;
      RECT 19.762 60.555 19.81 60.591 ;
      RECT 19.762 61.755 19.81 61.791 ;
      RECT 19.762 62.955 19.81 62.991 ;
      RECT 19.762 64.155 19.81 64.191 ;
      RECT 19.762 65.355 19.81 65.391 ;
      RECT 19.762 66.555 19.81 66.591 ;
      RECT 19.762 67.755 19.81 67.791 ;
      RECT 19.762 68.955 19.81 68.991 ;
      RECT 19.762 70.155 19.81 70.191 ;
      RECT 19.762 71.355 19.81 71.391 ;
      RECT 19.838 1.558 19.886 1.594 ;
      RECT 19.838 2.758 19.886 2.794 ;
      RECT 19.838 3.958 19.886 3.994 ;
      RECT 19.838 5.158 19.886 5.194 ;
      RECT 19.838 6.358 19.886 6.394 ;
      RECT 19.838 7.558 19.886 7.594 ;
      RECT 19.838 8.758 19.886 8.794 ;
      RECT 19.838 9.958 19.886 9.994 ;
      RECT 19.838 11.158 19.886 11.194 ;
      RECT 19.838 12.358 19.886 12.394 ;
      RECT 19.838 13.558 19.886 13.594 ;
      RECT 19.838 14.758 19.886 14.794 ;
      RECT 19.838 15.958 19.886 15.994 ;
      RECT 19.838 17.158 19.886 17.194 ;
      RECT 19.838 18.358 19.886 18.394 ;
      RECT 19.838 19.558 19.886 19.594 ;
      RECT 19.838 20.758 19.886 20.794 ;
      RECT 19.838 21.958 19.886 21.994 ;
      RECT 19.838 23.158 19.886 23.194 ;
      RECT 19.838 24.358 19.886 24.394 ;
      RECT 19.838 25.558 19.886 25.594 ;
      RECT 19.838 26.758 19.886 26.794 ;
      RECT 19.838 27.958 19.886 27.994 ;
      RECT 19.838 29.158 19.886 29.194 ;
      RECT 19.838 30.358 19.886 30.394 ;
      RECT 19.838 31.558 19.886 31.594 ;
      RECT 19.838 32.502 19.886 32.538 ;
      RECT 19.838 34.902 19.886 34.938 ;
      RECT 19.838 35.382 19.886 35.418 ;
      RECT 19.838 37.0005 19.886 37.0365 ;
      RECT 19.838 38.9205 19.886 38.9565 ;
      RECT 19.838 40.678 19.886 40.714 ;
      RECT 19.838 41.878 19.886 41.914 ;
      RECT 19.838 43.078 19.886 43.114 ;
      RECT 19.838 44.278 19.886 44.314 ;
      RECT 19.838 45.478 19.886 45.514 ;
      RECT 19.838 46.678 19.886 46.714 ;
      RECT 19.838 47.878 19.886 47.914 ;
      RECT 19.838 49.078 19.886 49.114 ;
      RECT 19.838 50.278 19.886 50.314 ;
      RECT 19.838 51.478 19.886 51.514 ;
      RECT 19.838 52.678 19.886 52.714 ;
      RECT 19.838 53.878 19.886 53.914 ;
      RECT 19.838 55.078 19.886 55.114 ;
      RECT 19.838 56.278 19.886 56.314 ;
      RECT 19.838 57.478 19.886 57.514 ;
      RECT 19.838 58.678 19.886 58.714 ;
      RECT 19.838 59.878 19.886 59.914 ;
      RECT 19.838 61.078 19.886 61.114 ;
      RECT 19.838 62.278 19.886 62.314 ;
      RECT 19.838 63.478 19.886 63.514 ;
      RECT 19.838 64.678 19.886 64.714 ;
      RECT 19.838 65.878 19.886 65.914 ;
      RECT 19.838 67.078 19.886 67.114 ;
      RECT 19.838 68.278 19.886 68.314 ;
      RECT 19.838 69.478 19.886 69.514 ;
      RECT 19.838 70.678 19.886 70.714 ;
      RECT 19.838 71.878 19.886 71.914 ;
      RECT 20.154 32.982 20.194 33.018 ;
      RECT 20.154 37.302 20.194 37.338 ;
      RECT 20.222 33.222 20.262 33.258 ;
      RECT 20.222 35.6835 20.262 35.7195 ;
      RECT 20.222 38.262 20.262 38.298 ;
      RECT 20.37 1.3345 20.442 1.3595 ;
      RECT 20.37 2.5345 20.442 2.5595 ;
      RECT 20.37 3.7345 20.442 3.7595 ;
      RECT 20.37 4.9345 20.442 4.9595 ;
      RECT 20.37 6.1345 20.442 6.1595 ;
      RECT 20.37 7.3345 20.442 7.3595 ;
      RECT 20.37 8.5345 20.442 8.5595 ;
      RECT 20.37 9.7345 20.442 9.7595 ;
      RECT 20.37 10.9345 20.442 10.9595 ;
      RECT 20.37 12.1345 20.442 12.1595 ;
      RECT 20.37 13.3345 20.442 13.3595 ;
      RECT 20.37 14.5345 20.442 14.5595 ;
      RECT 20.37 15.7345 20.442 15.7595 ;
      RECT 20.37 16.9345 20.442 16.9595 ;
      RECT 20.37 18.1345 20.442 18.1595 ;
      RECT 20.37 19.3345 20.442 19.3595 ;
      RECT 20.37 20.5345 20.442 20.5595 ;
      RECT 20.37 21.7345 20.442 21.7595 ;
      RECT 20.37 22.9345 20.442 22.9595 ;
      RECT 20.37 24.1345 20.442 24.1595 ;
      RECT 20.37 25.3345 20.442 25.3595 ;
      RECT 20.37 26.5345 20.442 26.5595 ;
      RECT 20.37 27.7345 20.442 27.7595 ;
      RECT 20.37 28.9345 20.442 28.9595 ;
      RECT 20.37 30.1345 20.442 30.1595 ;
      RECT 20.37 31.3345 20.442 31.3595 ;
      RECT 20.37 32.2675 20.442 32.2925 ;
      RECT 20.37 33.406 20.442 33.431 ;
      RECT 20.37 37.7875 20.442 37.8125 ;
      RECT 20.37 39.2275 20.442 39.2525 ;
      RECT 20.37 40.4545 20.442 40.4795 ;
      RECT 20.37 41.6545 20.442 41.6795 ;
      RECT 20.37 42.8545 20.442 42.8795 ;
      RECT 20.37 44.0545 20.442 44.0795 ;
      RECT 20.37 45.2545 20.442 45.2795 ;
      RECT 20.37 46.4545 20.442 46.4795 ;
      RECT 20.37 47.6545 20.442 47.6795 ;
      RECT 20.37 48.8545 20.442 48.8795 ;
      RECT 20.37 50.0545 20.442 50.0795 ;
      RECT 20.37 51.2545 20.442 51.2795 ;
      RECT 20.37 52.4545 20.442 52.4795 ;
      RECT 20.37 53.6545 20.442 53.6795 ;
      RECT 20.37 54.8545 20.442 54.8795 ;
      RECT 20.37 56.0545 20.442 56.0795 ;
      RECT 20.37 57.2545 20.442 57.2795 ;
      RECT 20.37 58.4545 20.442 58.4795 ;
      RECT 20.37 59.6545 20.442 59.6795 ;
      RECT 20.37 60.8545 20.442 60.8795 ;
      RECT 20.37 62.0545 20.442 62.0795 ;
      RECT 20.37 63.2545 20.442 63.2795 ;
      RECT 20.37 64.4545 20.442 64.4795 ;
      RECT 20.37 65.6545 20.442 65.6795 ;
      RECT 20.37 66.8545 20.442 66.8795 ;
      RECT 20.37 68.0545 20.442 68.0795 ;
      RECT 20.37 69.2545 20.442 69.2795 ;
      RECT 20.37 70.4545 20.442 70.4795 ;
      RECT 20.37 71.6545 20.442 71.6795 ;
      RECT 20.47 33.702 20.522 33.738 ;
      RECT 20.47 38.0835 20.522 38.1195 ;
      RECT 20.55 34.6005 20.602 34.6365 ;
      RECT 20.55 36.102 20.602 36.138 ;
      RECT 20.778 0.582 20.822 0.618 ;
      RECT 20.778 1.182 20.822 1.218 ;
      RECT 20.778 1.782 20.822 1.818 ;
      RECT 20.778 2.382 20.822 2.418 ;
      RECT 20.778 2.982 20.822 3.018 ;
      RECT 20.778 3.582 20.822 3.618 ;
      RECT 20.778 4.182 20.822 4.218 ;
      RECT 20.778 4.782 20.822 4.818 ;
      RECT 20.778 5.382 20.822 5.418 ;
      RECT 20.778 5.982 20.822 6.018 ;
      RECT 20.778 6.582 20.822 6.618 ;
      RECT 20.778 7.182 20.822 7.218 ;
      RECT 20.778 7.782 20.822 7.818 ;
      RECT 20.778 8.382 20.822 8.418 ;
      RECT 20.778 8.982 20.822 9.018 ;
      RECT 20.778 9.582 20.822 9.618 ;
      RECT 20.778 10.182 20.822 10.218 ;
      RECT 20.778 10.782 20.822 10.818 ;
      RECT 20.778 11.382 20.822 11.418 ;
      RECT 20.778 11.982 20.822 12.018 ;
      RECT 20.778 12.582 20.822 12.618 ;
      RECT 20.778 13.182 20.822 13.218 ;
      RECT 20.778 13.782 20.822 13.818 ;
      RECT 20.778 14.382 20.822 14.418 ;
      RECT 20.778 14.982 20.822 15.018 ;
      RECT 20.778 15.582 20.822 15.618 ;
      RECT 20.778 16.182 20.822 16.218 ;
      RECT 20.778 16.782 20.822 16.818 ;
      RECT 20.778 17.382 20.822 17.418 ;
      RECT 20.778 17.982 20.822 18.018 ;
      RECT 20.778 18.582 20.822 18.618 ;
      RECT 20.778 19.182 20.822 19.218 ;
      RECT 20.778 19.782 20.822 19.818 ;
      RECT 20.778 20.382 20.822 20.418 ;
      RECT 20.778 20.982 20.822 21.018 ;
      RECT 20.778 21.582 20.822 21.618 ;
      RECT 20.778 22.182 20.822 22.218 ;
      RECT 20.778 22.782 20.822 22.818 ;
      RECT 20.778 23.382 20.822 23.418 ;
      RECT 20.778 23.982 20.822 24.018 ;
      RECT 20.778 24.582 20.822 24.618 ;
      RECT 20.778 25.182 20.822 25.218 ;
      RECT 20.778 25.782 20.822 25.818 ;
      RECT 20.778 26.382 20.822 26.418 ;
      RECT 20.778 26.982 20.822 27.018 ;
      RECT 20.778 27.582 20.822 27.618 ;
      RECT 20.778 28.182 20.822 28.218 ;
      RECT 20.778 28.782 20.822 28.818 ;
      RECT 20.778 29.382 20.822 29.418 ;
      RECT 20.778 29.982 20.822 30.018 ;
      RECT 20.778 30.582 20.822 30.618 ;
      RECT 20.778 31.182 20.822 31.218 ;
      RECT 20.778 31.782 20.822 31.818 ;
      RECT 20.778 32.142 20.822 32.178 ;
      RECT 20.778 32.622 20.822 32.658 ;
      RECT 20.778 33.102 20.822 33.138 ;
      RECT 20.778 33.582 20.822 33.618 ;
      RECT 20.778 34.062 20.822 34.098 ;
      RECT 20.778 34.542 20.822 34.578 ;
      RECT 20.778 35.022 20.822 35.058 ;
      RECT 20.778 35.502 20.822 35.538 ;
      RECT 20.778 35.982 20.822 36.018 ;
      RECT 20.778 36.462 20.822 36.498 ;
      RECT 20.778 36.942 20.822 36.978 ;
      RECT 20.778 37.4275 20.822 37.4525 ;
      RECT 20.778 37.9075 20.822 37.9325 ;
      RECT 20.778 38.382 20.822 38.418 ;
      RECT 20.778 38.8675 20.822 38.8925 ;
      RECT 20.778 39.342 20.822 39.378 ;
      RECT 20.778 39.702 20.822 39.738 ;
      RECT 20.778 40.302 20.822 40.338 ;
      RECT 20.778 40.902 20.822 40.938 ;
      RECT 20.778 41.502 20.822 41.538 ;
      RECT 20.778 42.102 20.822 42.138 ;
      RECT 20.778 42.702 20.822 42.738 ;
      RECT 20.778 43.302 20.822 43.338 ;
      RECT 20.778 43.902 20.822 43.938 ;
      RECT 20.778 44.502 20.822 44.538 ;
      RECT 20.778 45.102 20.822 45.138 ;
      RECT 20.778 45.702 20.822 45.738 ;
      RECT 20.778 46.302 20.822 46.338 ;
      RECT 20.778 46.902 20.822 46.938 ;
      RECT 20.778 47.502 20.822 47.538 ;
      RECT 20.778 48.102 20.822 48.138 ;
      RECT 20.778 48.702 20.822 48.738 ;
      RECT 20.778 49.302 20.822 49.338 ;
      RECT 20.778 49.902 20.822 49.938 ;
      RECT 20.778 50.502 20.822 50.538 ;
      RECT 20.778 51.102 20.822 51.138 ;
      RECT 20.778 51.702 20.822 51.738 ;
      RECT 20.778 52.302 20.822 52.338 ;
      RECT 20.778 52.902 20.822 52.938 ;
      RECT 20.778 53.502 20.822 53.538 ;
      RECT 20.778 54.102 20.822 54.138 ;
      RECT 20.778 54.702 20.822 54.738 ;
      RECT 20.778 55.302 20.822 55.338 ;
      RECT 20.778 55.902 20.822 55.938 ;
      RECT 20.778 56.502 20.822 56.538 ;
      RECT 20.778 57.102 20.822 57.138 ;
      RECT 20.778 57.702 20.822 57.738 ;
      RECT 20.778 58.302 20.822 58.338 ;
      RECT 20.778 58.902 20.822 58.938 ;
      RECT 20.778 59.502 20.822 59.538 ;
      RECT 20.778 60.102 20.822 60.138 ;
      RECT 20.778 60.702 20.822 60.738 ;
      RECT 20.778 61.302 20.822 61.338 ;
      RECT 20.778 61.902 20.822 61.938 ;
      RECT 20.778 62.502 20.822 62.538 ;
      RECT 20.778 63.102 20.822 63.138 ;
      RECT 20.778 63.702 20.822 63.738 ;
      RECT 20.778 64.302 20.822 64.338 ;
      RECT 20.778 64.902 20.822 64.938 ;
      RECT 20.778 65.502 20.822 65.538 ;
      RECT 20.778 66.102 20.822 66.138 ;
      RECT 20.778 66.702 20.822 66.738 ;
      RECT 20.778 67.302 20.822 67.338 ;
      RECT 20.778 67.902 20.822 67.938 ;
      RECT 20.778 68.502 20.822 68.538 ;
      RECT 20.778 69.102 20.822 69.138 ;
      RECT 20.778 69.702 20.822 69.738 ;
      RECT 20.778 70.302 20.822 70.338 ;
      RECT 20.778 70.902 20.822 70.938 ;
      RECT 20.778 71.502 20.822 71.538 ;
      RECT 20.778 72.102 20.822 72.138 ;
      RECT 20.932 34.4835 20.986 34.5195 ;
      RECT 20.932 37.3635 20.986 37.3995 ;
      RECT 21.096 0.582 21.14 0.618 ;
      RECT 21.096 1.782 21.14 1.818 ;
      RECT 21.096 2.982 21.14 3.018 ;
      RECT 21.096 4.182 21.14 4.218 ;
      RECT 21.096 5.382 21.14 5.418 ;
      RECT 21.096 6.582 21.14 6.618 ;
      RECT 21.096 7.782 21.14 7.818 ;
      RECT 21.096 8.982 21.14 9.018 ;
      RECT 21.096 10.182 21.14 10.218 ;
      RECT 21.096 11.382 21.14 11.418 ;
      RECT 21.096 12.582 21.14 12.618 ;
      RECT 21.096 13.782 21.14 13.818 ;
      RECT 21.096 14.982 21.14 15.018 ;
      RECT 21.096 16.182 21.14 16.218 ;
      RECT 21.096 17.382 21.14 17.418 ;
      RECT 21.096 18.582 21.14 18.618 ;
      RECT 21.096 19.782 21.14 19.818 ;
      RECT 21.096 20.982 21.14 21.018 ;
      RECT 21.096 22.182 21.14 22.218 ;
      RECT 21.096 23.382 21.14 23.418 ;
      RECT 21.096 24.582 21.14 24.618 ;
      RECT 21.096 25.782 21.14 25.818 ;
      RECT 21.096 26.982 21.14 27.018 ;
      RECT 21.096 28.182 21.14 28.218 ;
      RECT 21.096 29.382 21.14 29.418 ;
      RECT 21.096 30.582 21.14 30.618 ;
      RECT 21.096 31.782 21.14 31.818 ;
      RECT 21.096 32.142 21.14 32.178 ;
      RECT 21.096 32.622 21.14 32.658 ;
      RECT 21.096 33.102 21.14 33.138 ;
      RECT 21.096 33.582 21.14 33.618 ;
      RECT 21.096 34.062 21.14 34.098 ;
      RECT 21.096 34.542 21.14 34.578 ;
      RECT 21.096 35.022 21.14 35.058 ;
      RECT 21.096 35.502 21.14 35.538 ;
      RECT 21.096 35.982 21.14 36.018 ;
      RECT 21.096 36.462 21.14 36.498 ;
      RECT 21.096 36.942 21.14 36.978 ;
      RECT 21.096 37.422 21.14 37.458 ;
      RECT 21.096 37.902 21.14 37.938 ;
      RECT 21.096 38.382 21.14 38.418 ;
      RECT 21.096 38.862 21.14 38.898 ;
      RECT 21.096 39.342 21.14 39.378 ;
      RECT 21.096 39.702 21.14 39.738 ;
      RECT 21.096 40.902 21.14 40.938 ;
      RECT 21.096 42.102 21.14 42.138 ;
      RECT 21.096 43.302 21.14 43.338 ;
      RECT 21.096 44.502 21.14 44.538 ;
      RECT 21.096 45.702 21.14 45.738 ;
      RECT 21.096 46.902 21.14 46.938 ;
      RECT 21.096 48.102 21.14 48.138 ;
      RECT 21.096 49.302 21.14 49.338 ;
      RECT 21.096 50.502 21.14 50.538 ;
      RECT 21.096 51.702 21.14 51.738 ;
      RECT 21.096 52.902 21.14 52.938 ;
      RECT 21.096 54.102 21.14 54.138 ;
      RECT 21.096 55.302 21.14 55.338 ;
      RECT 21.096 56.502 21.14 56.538 ;
      RECT 21.096 57.702 21.14 57.738 ;
      RECT 21.096 58.902 21.14 58.938 ;
      RECT 21.096 60.102 21.14 60.138 ;
      RECT 21.096 61.302 21.14 61.338 ;
      RECT 21.096 62.502 21.14 62.538 ;
      RECT 21.096 63.702 21.14 63.738 ;
      RECT 21.096 64.902 21.14 64.938 ;
      RECT 21.096 66.102 21.14 66.138 ;
      RECT 21.096 67.302 21.14 67.338 ;
      RECT 21.096 68.502 21.14 68.538 ;
      RECT 21.096 69.702 21.14 69.738 ;
      RECT 21.096 70.902 21.14 70.938 ;
      RECT 21.096 72.102 21.14 72.138 ;
      RECT 21.168 0.806 21.222 0.842 ;
      RECT 21.168 2.006 21.222 2.042 ;
      RECT 21.168 3.206 21.222 3.242 ;
      RECT 21.168 4.406 21.222 4.442 ;
      RECT 21.168 5.606 21.222 5.642 ;
      RECT 21.168 6.806 21.222 6.842 ;
      RECT 21.168 8.006 21.222 8.042 ;
      RECT 21.168 9.206 21.222 9.242 ;
      RECT 21.168 10.406 21.222 10.442 ;
      RECT 21.168 11.606 21.222 11.642 ;
      RECT 21.168 12.806 21.222 12.842 ;
      RECT 21.168 14.006 21.222 14.042 ;
      RECT 21.168 15.206 21.222 15.242 ;
      RECT 21.168 16.406 21.222 16.442 ;
      RECT 21.168 17.606 21.222 17.642 ;
      RECT 21.168 18.806 21.222 18.842 ;
      RECT 21.168 20.006 21.222 20.042 ;
      RECT 21.168 21.206 21.222 21.242 ;
      RECT 21.168 22.406 21.222 22.442 ;
      RECT 21.168 23.606 21.222 23.642 ;
      RECT 21.168 24.806 21.222 24.842 ;
      RECT 21.168 26.006 21.222 26.042 ;
      RECT 21.168 27.206 21.222 27.242 ;
      RECT 21.168 28.406 21.222 28.442 ;
      RECT 21.168 29.606 21.222 29.642 ;
      RECT 21.168 30.806 21.222 30.842 ;
      RECT 21.168 32.9205 21.222 32.9565 ;
      RECT 21.168 33.222 21.222 33.258 ;
      RECT 21.168 37.782 21.222 37.818 ;
      RECT 21.168 38.262 21.222 38.298 ;
      RECT 21.168 38.6805 21.222 38.7165 ;
      RECT 21.168 39.926 21.222 39.962 ;
      RECT 21.168 41.126 21.222 41.162 ;
      RECT 21.168 42.326 21.222 42.362 ;
      RECT 21.168 43.526 21.222 43.562 ;
      RECT 21.168 44.726 21.222 44.762 ;
      RECT 21.168 45.926 21.222 45.962 ;
      RECT 21.168 47.126 21.222 47.162 ;
      RECT 21.168 48.326 21.222 48.362 ;
      RECT 21.168 49.526 21.222 49.562 ;
      RECT 21.168 50.726 21.222 50.762 ;
      RECT 21.168 51.926 21.222 51.962 ;
      RECT 21.168 53.126 21.222 53.162 ;
      RECT 21.168 54.326 21.222 54.362 ;
      RECT 21.168 55.526 21.222 55.562 ;
      RECT 21.168 56.726 21.222 56.762 ;
      RECT 21.168 57.926 21.222 57.962 ;
      RECT 21.168 59.126 21.222 59.162 ;
      RECT 21.168 60.326 21.222 60.362 ;
      RECT 21.168 61.526 21.222 61.562 ;
      RECT 21.168 62.726 21.222 62.762 ;
      RECT 21.168 63.926 21.222 63.962 ;
      RECT 21.168 65.126 21.222 65.162 ;
      RECT 21.168 66.326 21.222 66.362 ;
      RECT 21.168 67.526 21.222 67.562 ;
      RECT 21.168 68.726 21.222 68.762 ;
      RECT 21.168 69.926 21.222 69.962 ;
      RECT 21.168 71.126 21.222 71.162 ;
      RECT 21.25 1.482 21.304 1.518 ;
      RECT 21.25 2.682 21.304 2.718 ;
      RECT 21.25 3.882 21.304 3.918 ;
      RECT 21.25 5.082 21.304 5.118 ;
      RECT 21.25 6.282 21.304 6.318 ;
      RECT 21.25 7.482 21.304 7.518 ;
      RECT 21.25 8.682 21.304 8.718 ;
      RECT 21.25 9.882 21.304 9.918 ;
      RECT 21.25 11.082 21.304 11.118 ;
      RECT 21.25 12.282 21.304 12.318 ;
      RECT 21.25 13.482 21.304 13.518 ;
      RECT 21.25 14.682 21.304 14.718 ;
      RECT 21.25 15.882 21.304 15.918 ;
      RECT 21.25 17.082 21.304 17.118 ;
      RECT 21.25 18.282 21.304 18.318 ;
      RECT 21.25 19.482 21.304 19.518 ;
      RECT 21.25 20.682 21.304 20.718 ;
      RECT 21.25 21.882 21.304 21.918 ;
      RECT 21.25 23.082 21.304 23.118 ;
      RECT 21.25 24.282 21.304 24.318 ;
      RECT 21.25 25.482 21.304 25.518 ;
      RECT 21.25 26.682 21.304 26.718 ;
      RECT 21.25 27.882 21.304 27.918 ;
      RECT 21.25 29.082 21.304 29.118 ;
      RECT 21.25 30.282 21.304 30.318 ;
      RECT 21.25 31.482 21.304 31.518 ;
      RECT 21.25 32.5635 21.304 32.5995 ;
      RECT 21.25 32.8035 21.304 32.8395 ;
      RECT 21.25 37.6035 21.304 37.6395 ;
      RECT 21.25 38.5635 21.304 38.5995 ;
      RECT 21.25 38.9205 21.304 38.9565 ;
      RECT 21.25 40.602 21.304 40.638 ;
      RECT 21.25 41.802 21.304 41.838 ;
      RECT 21.25 43.002 21.304 43.038 ;
      RECT 21.25 44.202 21.304 44.238 ;
      RECT 21.25 45.402 21.304 45.438 ;
      RECT 21.25 46.602 21.304 46.638 ;
      RECT 21.25 47.802 21.304 47.838 ;
      RECT 21.25 49.002 21.304 49.038 ;
      RECT 21.25 50.202 21.304 50.238 ;
      RECT 21.25 51.402 21.304 51.438 ;
      RECT 21.25 52.602 21.304 52.638 ;
      RECT 21.25 53.802 21.304 53.838 ;
      RECT 21.25 55.002 21.304 55.038 ;
      RECT 21.25 56.202 21.304 56.238 ;
      RECT 21.25 57.402 21.304 57.438 ;
      RECT 21.25 58.602 21.304 58.638 ;
      RECT 21.25 59.802 21.304 59.838 ;
      RECT 21.25 61.002 21.304 61.038 ;
      RECT 21.25 62.202 21.304 62.238 ;
      RECT 21.25 63.402 21.304 63.438 ;
      RECT 21.25 64.602 21.304 64.638 ;
      RECT 21.25 65.802 21.304 65.838 ;
      RECT 21.25 67.002 21.304 67.038 ;
      RECT 21.25 68.202 21.304 68.238 ;
      RECT 21.25 69.402 21.304 69.438 ;
      RECT 21.25 70.602 21.304 70.638 ;
      RECT 21.25 71.802 21.304 71.838 ;
      RECT 21.332 0.806 21.386 0.842 ;
      RECT 21.332 2.006 21.386 2.042 ;
      RECT 21.332 3.206 21.386 3.242 ;
      RECT 21.332 4.406 21.386 4.442 ;
      RECT 21.332 5.606 21.386 5.642 ;
      RECT 21.332 6.806 21.386 6.842 ;
      RECT 21.332 8.006 21.386 8.042 ;
      RECT 21.332 9.206 21.386 9.242 ;
      RECT 21.332 10.406 21.386 10.442 ;
      RECT 21.332 11.606 21.386 11.642 ;
      RECT 21.332 12.806 21.386 12.842 ;
      RECT 21.332 14.006 21.386 14.042 ;
      RECT 21.332 15.206 21.386 15.242 ;
      RECT 21.332 16.406 21.386 16.442 ;
      RECT 21.332 17.606 21.386 17.642 ;
      RECT 21.332 18.806 21.386 18.842 ;
      RECT 21.332 20.006 21.386 20.042 ;
      RECT 21.332 21.206 21.386 21.242 ;
      RECT 21.332 22.406 21.386 22.442 ;
      RECT 21.332 23.606 21.386 23.642 ;
      RECT 21.332 24.806 21.386 24.842 ;
      RECT 21.332 26.006 21.386 26.042 ;
      RECT 21.332 27.206 21.386 27.242 ;
      RECT 21.332 28.406 21.386 28.442 ;
      RECT 21.332 29.606 21.386 29.642 ;
      RECT 21.332 30.806 21.386 30.842 ;
      RECT 21.332 32.2005 21.386 32.2365 ;
      RECT 21.332 32.6805 21.386 32.7165 ;
      RECT 21.332 37.8435 21.386 37.8795 ;
      RECT 21.332 38.686 21.386 38.711 ;
      RECT 21.332 38.809 21.386 38.834 ;
      RECT 21.332 39.926 21.386 39.962 ;
      RECT 21.332 41.126 21.386 41.162 ;
      RECT 21.332 42.326 21.386 42.362 ;
      RECT 21.332 43.526 21.386 43.562 ;
      RECT 21.332 44.726 21.386 44.762 ;
      RECT 21.332 45.926 21.386 45.962 ;
      RECT 21.332 47.126 21.386 47.162 ;
      RECT 21.332 48.326 21.386 48.362 ;
      RECT 21.332 49.526 21.386 49.562 ;
      RECT 21.332 50.726 21.386 50.762 ;
      RECT 21.332 51.926 21.386 51.962 ;
      RECT 21.332 53.126 21.386 53.162 ;
      RECT 21.332 54.326 21.386 54.362 ;
      RECT 21.332 55.526 21.386 55.562 ;
      RECT 21.332 56.726 21.386 56.762 ;
      RECT 21.332 57.926 21.386 57.962 ;
      RECT 21.332 59.126 21.386 59.162 ;
      RECT 21.332 60.326 21.386 60.362 ;
      RECT 21.332 61.526 21.386 61.562 ;
      RECT 21.332 62.726 21.386 62.762 ;
      RECT 21.332 63.926 21.386 63.962 ;
      RECT 21.332 65.126 21.386 65.162 ;
      RECT 21.332 66.326 21.386 66.362 ;
      RECT 21.332 67.526 21.386 67.562 ;
      RECT 21.332 68.726 21.386 68.762 ;
      RECT 21.332 69.926 21.386 69.962 ;
      RECT 21.332 71.126 21.386 71.162 ;
      RECT 21.414 1.482 21.468 1.518 ;
      RECT 21.414 2.682 21.468 2.718 ;
      RECT 21.414 3.882 21.468 3.918 ;
      RECT 21.414 5.082 21.468 5.118 ;
      RECT 21.414 6.282 21.468 6.318 ;
      RECT 21.414 7.482 21.468 7.518 ;
      RECT 21.414 8.682 21.468 8.718 ;
      RECT 21.414 9.882 21.468 9.918 ;
      RECT 21.414 11.082 21.468 11.118 ;
      RECT 21.414 12.282 21.468 12.318 ;
      RECT 21.414 13.482 21.468 13.518 ;
      RECT 21.414 14.682 21.468 14.718 ;
      RECT 21.414 15.882 21.468 15.918 ;
      RECT 21.414 17.082 21.468 17.118 ;
      RECT 21.414 18.282 21.468 18.318 ;
      RECT 21.414 19.482 21.468 19.518 ;
      RECT 21.414 20.682 21.468 20.718 ;
      RECT 21.414 21.882 21.468 21.918 ;
      RECT 21.414 23.082 21.468 23.118 ;
      RECT 21.414 24.282 21.468 24.318 ;
      RECT 21.414 25.482 21.468 25.518 ;
      RECT 21.414 26.682 21.468 26.718 ;
      RECT 21.414 27.882 21.468 27.918 ;
      RECT 21.414 29.082 21.468 29.118 ;
      RECT 21.414 30.282 21.468 30.318 ;
      RECT 21.414 31.482 21.468 31.518 ;
      RECT 21.414 32.3235 21.468 32.3595 ;
      RECT 21.414 32.4405 21.468 32.4765 ;
      RECT 21.414 37.6035 21.468 37.6395 ;
      RECT 21.414 38.982 21.468 39.018 ;
      RECT 21.414 39.222 21.468 39.258 ;
      RECT 21.414 40.602 21.468 40.638 ;
      RECT 21.414 41.802 21.468 41.838 ;
      RECT 21.414 43.002 21.468 43.038 ;
      RECT 21.414 44.202 21.468 44.238 ;
      RECT 21.414 45.402 21.468 45.438 ;
      RECT 21.414 46.602 21.468 46.638 ;
      RECT 21.414 47.802 21.468 47.838 ;
      RECT 21.414 49.002 21.468 49.038 ;
      RECT 21.414 50.202 21.468 50.238 ;
      RECT 21.414 51.402 21.468 51.438 ;
      RECT 21.414 52.602 21.468 52.638 ;
      RECT 21.414 53.802 21.468 53.838 ;
      RECT 21.414 55.002 21.468 55.038 ;
      RECT 21.414 56.202 21.468 56.238 ;
      RECT 21.414 57.402 21.468 57.438 ;
      RECT 21.414 58.602 21.468 58.638 ;
      RECT 21.414 59.802 21.468 59.838 ;
      RECT 21.414 61.002 21.468 61.038 ;
      RECT 21.414 62.202 21.468 62.238 ;
      RECT 21.414 63.402 21.468 63.438 ;
      RECT 21.414 64.602 21.468 64.638 ;
      RECT 21.414 65.802 21.468 65.838 ;
      RECT 21.414 67.002 21.468 67.038 ;
      RECT 21.414 68.202 21.468 68.238 ;
      RECT 21.414 69.402 21.468 69.438 ;
      RECT 21.414 70.602 21.468 70.638 ;
      RECT 21.414 71.802 21.468 71.838 ;
      RECT 21.578 34.182 21.622 34.218 ;
      RECT 21.578 34.422 21.622 34.458 ;
      RECT 21.578 36.342 21.622 36.378 ;
      RECT 21.578 37.302 21.622 37.338 ;
      RECT 21.732 0.806 21.786 0.842 ;
      RECT 21.732 2.006 21.786 2.042 ;
      RECT 21.732 3.206 21.786 3.242 ;
      RECT 21.732 4.406 21.786 4.442 ;
      RECT 21.732 5.606 21.786 5.642 ;
      RECT 21.732 6.806 21.786 6.842 ;
      RECT 21.732 8.006 21.786 8.042 ;
      RECT 21.732 9.206 21.786 9.242 ;
      RECT 21.732 10.406 21.786 10.442 ;
      RECT 21.732 11.606 21.786 11.642 ;
      RECT 21.732 12.806 21.786 12.842 ;
      RECT 21.732 14.006 21.786 14.042 ;
      RECT 21.732 15.206 21.786 15.242 ;
      RECT 21.732 16.406 21.786 16.442 ;
      RECT 21.732 17.606 21.786 17.642 ;
      RECT 21.732 18.806 21.786 18.842 ;
      RECT 21.732 20.006 21.786 20.042 ;
      RECT 21.732 21.206 21.786 21.242 ;
      RECT 21.732 22.406 21.786 22.442 ;
      RECT 21.732 23.606 21.786 23.642 ;
      RECT 21.732 24.806 21.786 24.842 ;
      RECT 21.732 26.006 21.786 26.042 ;
      RECT 21.732 27.206 21.786 27.242 ;
      RECT 21.732 28.406 21.786 28.442 ;
      RECT 21.732 29.606 21.786 29.642 ;
      RECT 21.732 30.806 21.786 30.842 ;
      RECT 21.732 34.0035 21.786 34.0395 ;
      RECT 21.732 37.0005 21.786 37.0365 ;
      RECT 21.732 39.926 21.786 39.962 ;
      RECT 21.732 41.126 21.786 41.162 ;
      RECT 21.732 42.326 21.786 42.362 ;
      RECT 21.732 43.526 21.786 43.562 ;
      RECT 21.732 44.726 21.786 44.762 ;
      RECT 21.732 45.926 21.786 45.962 ;
      RECT 21.732 47.126 21.786 47.162 ;
      RECT 21.732 48.326 21.786 48.362 ;
      RECT 21.732 49.526 21.786 49.562 ;
      RECT 21.732 50.726 21.786 50.762 ;
      RECT 21.732 51.926 21.786 51.962 ;
      RECT 21.732 53.126 21.786 53.162 ;
      RECT 21.732 54.326 21.786 54.362 ;
      RECT 21.732 55.526 21.786 55.562 ;
      RECT 21.732 56.726 21.786 56.762 ;
      RECT 21.732 57.926 21.786 57.962 ;
      RECT 21.732 59.126 21.786 59.162 ;
      RECT 21.732 60.326 21.786 60.362 ;
      RECT 21.732 61.526 21.786 61.562 ;
      RECT 21.732 62.726 21.786 62.762 ;
      RECT 21.732 63.926 21.786 63.962 ;
      RECT 21.732 65.126 21.786 65.162 ;
      RECT 21.732 66.326 21.786 66.362 ;
      RECT 21.732 67.526 21.786 67.562 ;
      RECT 21.732 68.726 21.786 68.762 ;
      RECT 21.732 69.926 21.786 69.962 ;
      RECT 21.732 71.126 21.786 71.162 ;
      RECT 21.814 1.558 21.868 1.594 ;
      RECT 21.814 2.758 21.868 2.794 ;
      RECT 21.814 3.958 21.868 3.994 ;
      RECT 21.814 5.158 21.868 5.194 ;
      RECT 21.814 6.358 21.868 6.394 ;
      RECT 21.814 7.558 21.868 7.594 ;
      RECT 21.814 8.758 21.868 8.794 ;
      RECT 21.814 9.958 21.868 9.994 ;
      RECT 21.814 11.158 21.868 11.194 ;
      RECT 21.814 12.358 21.868 12.394 ;
      RECT 21.814 13.558 21.868 13.594 ;
      RECT 21.814 14.758 21.868 14.794 ;
      RECT 21.814 15.958 21.868 15.994 ;
      RECT 21.814 17.158 21.868 17.194 ;
      RECT 21.814 18.358 21.868 18.394 ;
      RECT 21.814 19.558 21.868 19.594 ;
      RECT 21.814 20.758 21.868 20.794 ;
      RECT 21.814 21.958 21.868 21.994 ;
      RECT 21.814 23.158 21.868 23.194 ;
      RECT 21.814 24.358 21.868 24.394 ;
      RECT 21.814 25.558 21.868 25.594 ;
      RECT 21.814 26.758 21.868 26.794 ;
      RECT 21.814 27.958 21.868 27.994 ;
      RECT 21.814 29.158 21.868 29.194 ;
      RECT 21.814 30.358 21.868 30.394 ;
      RECT 21.814 31.558 21.868 31.594 ;
      RECT 21.814 34.1205 21.868 34.1565 ;
      RECT 21.814 34.3605 21.868 34.3965 ;
      RECT 21.814 35.9235 21.868 35.9595 ;
      RECT 21.814 37.3635 21.868 37.3995 ;
      RECT 21.814 40.678 21.868 40.714 ;
      RECT 21.814 41.878 21.868 41.914 ;
      RECT 21.814 43.078 21.868 43.114 ;
      RECT 21.814 44.278 21.868 44.314 ;
      RECT 21.814 45.478 21.868 45.514 ;
      RECT 21.814 46.678 21.868 46.714 ;
      RECT 21.814 47.878 21.868 47.914 ;
      RECT 21.814 49.078 21.868 49.114 ;
      RECT 21.814 50.278 21.868 50.314 ;
      RECT 21.814 51.478 21.868 51.514 ;
      RECT 21.814 52.678 21.868 52.714 ;
      RECT 21.814 53.878 21.868 53.914 ;
      RECT 21.814 55.078 21.868 55.114 ;
      RECT 21.814 56.278 21.868 56.314 ;
      RECT 21.814 57.478 21.868 57.514 ;
      RECT 21.814 58.678 21.868 58.714 ;
      RECT 21.814 59.878 21.868 59.914 ;
      RECT 21.814 61.078 21.868 61.114 ;
      RECT 21.814 62.278 21.868 62.314 ;
      RECT 21.814 63.478 21.868 63.514 ;
      RECT 21.814 64.678 21.868 64.714 ;
      RECT 21.814 65.878 21.868 65.914 ;
      RECT 21.814 67.078 21.868 67.114 ;
      RECT 21.814 68.278 21.868 68.314 ;
      RECT 21.814 69.478 21.868 69.514 ;
      RECT 21.814 70.678 21.868 70.714 ;
      RECT 21.814 71.878 21.868 71.914 ;
      RECT 21.978 0.582 22.022 0.618 ;
      RECT 21.978 1.182 22.022 1.218 ;
      RECT 21.978 1.782 22.022 1.818 ;
      RECT 21.978 2.382 22.022 2.418 ;
      RECT 21.978 2.982 22.022 3.018 ;
      RECT 21.978 3.582 22.022 3.618 ;
      RECT 21.978 4.182 22.022 4.218 ;
      RECT 21.978 4.782 22.022 4.818 ;
      RECT 21.978 5.382 22.022 5.418 ;
      RECT 21.978 5.982 22.022 6.018 ;
      RECT 21.978 6.582 22.022 6.618 ;
      RECT 21.978 7.182 22.022 7.218 ;
      RECT 21.978 7.782 22.022 7.818 ;
      RECT 21.978 8.382 22.022 8.418 ;
      RECT 21.978 8.982 22.022 9.018 ;
      RECT 21.978 9.582 22.022 9.618 ;
      RECT 21.978 10.182 22.022 10.218 ;
      RECT 21.978 10.782 22.022 10.818 ;
      RECT 21.978 11.382 22.022 11.418 ;
      RECT 21.978 11.982 22.022 12.018 ;
      RECT 21.978 12.582 22.022 12.618 ;
      RECT 21.978 13.182 22.022 13.218 ;
      RECT 21.978 13.782 22.022 13.818 ;
      RECT 21.978 14.382 22.022 14.418 ;
      RECT 21.978 14.982 22.022 15.018 ;
      RECT 21.978 15.582 22.022 15.618 ;
      RECT 21.978 16.182 22.022 16.218 ;
      RECT 21.978 16.782 22.022 16.818 ;
      RECT 21.978 17.382 22.022 17.418 ;
      RECT 21.978 17.982 22.022 18.018 ;
      RECT 21.978 18.582 22.022 18.618 ;
      RECT 21.978 19.182 22.022 19.218 ;
      RECT 21.978 19.782 22.022 19.818 ;
      RECT 21.978 20.382 22.022 20.418 ;
      RECT 21.978 20.982 22.022 21.018 ;
      RECT 21.978 21.582 22.022 21.618 ;
      RECT 21.978 22.182 22.022 22.218 ;
      RECT 21.978 22.782 22.022 22.818 ;
      RECT 21.978 23.382 22.022 23.418 ;
      RECT 21.978 23.982 22.022 24.018 ;
      RECT 21.978 24.582 22.022 24.618 ;
      RECT 21.978 25.182 22.022 25.218 ;
      RECT 21.978 25.782 22.022 25.818 ;
      RECT 21.978 26.382 22.022 26.418 ;
      RECT 21.978 26.982 22.022 27.018 ;
      RECT 21.978 27.582 22.022 27.618 ;
      RECT 21.978 28.182 22.022 28.218 ;
      RECT 21.978 28.782 22.022 28.818 ;
      RECT 21.978 29.382 22.022 29.418 ;
      RECT 21.978 29.982 22.022 30.018 ;
      RECT 21.978 30.582 22.022 30.618 ;
      RECT 21.978 31.182 22.022 31.218 ;
      RECT 21.978 31.782 22.022 31.818 ;
      RECT 21.978 32.142 22.022 32.178 ;
      RECT 21.978 32.622 22.022 32.658 ;
      RECT 21.978 33.102 22.022 33.138 ;
      RECT 21.978 33.582 22.022 33.618 ;
      RECT 21.978 34.062 22.022 34.098 ;
      RECT 21.978 34.542 22.022 34.578 ;
      RECT 21.978 35.022 22.022 35.058 ;
      RECT 21.978 35.502 22.022 35.538 ;
      RECT 21.978 35.982 22.022 36.018 ;
      RECT 21.978 36.462 22.022 36.498 ;
      RECT 21.978 36.942 22.022 36.978 ;
      RECT 21.978 37.422 22.022 37.458 ;
      RECT 21.978 37.902 22.022 37.938 ;
      RECT 21.978 38.382 22.022 38.418 ;
      RECT 21.978 38.862 22.022 38.898 ;
      RECT 21.978 39.342 22.022 39.378 ;
      RECT 21.978 39.702 22.022 39.738 ;
      RECT 21.978 40.302 22.022 40.338 ;
      RECT 21.978 40.902 22.022 40.938 ;
      RECT 21.978 41.502 22.022 41.538 ;
      RECT 21.978 42.102 22.022 42.138 ;
      RECT 21.978 42.702 22.022 42.738 ;
      RECT 21.978 43.302 22.022 43.338 ;
      RECT 21.978 43.902 22.022 43.938 ;
      RECT 21.978 44.502 22.022 44.538 ;
      RECT 21.978 45.102 22.022 45.138 ;
      RECT 21.978 45.702 22.022 45.738 ;
      RECT 21.978 46.302 22.022 46.338 ;
      RECT 21.978 46.902 22.022 46.938 ;
      RECT 21.978 47.502 22.022 47.538 ;
      RECT 21.978 48.102 22.022 48.138 ;
      RECT 21.978 48.702 22.022 48.738 ;
      RECT 21.978 49.302 22.022 49.338 ;
      RECT 21.978 49.902 22.022 49.938 ;
      RECT 21.978 50.502 22.022 50.538 ;
      RECT 21.978 51.102 22.022 51.138 ;
      RECT 21.978 51.702 22.022 51.738 ;
      RECT 21.978 52.302 22.022 52.338 ;
      RECT 21.978 52.902 22.022 52.938 ;
      RECT 21.978 53.502 22.022 53.538 ;
      RECT 21.978 54.102 22.022 54.138 ;
      RECT 21.978 54.702 22.022 54.738 ;
      RECT 21.978 55.302 22.022 55.338 ;
      RECT 21.978 55.902 22.022 55.938 ;
      RECT 21.978 56.502 22.022 56.538 ;
      RECT 21.978 57.102 22.022 57.138 ;
      RECT 21.978 57.702 22.022 57.738 ;
      RECT 21.978 58.302 22.022 58.338 ;
      RECT 21.978 58.902 22.022 58.938 ;
      RECT 21.978 59.502 22.022 59.538 ;
      RECT 21.978 60.102 22.022 60.138 ;
      RECT 21.978 60.702 22.022 60.738 ;
      RECT 21.978 61.302 22.022 61.338 ;
      RECT 21.978 61.902 22.022 61.938 ;
      RECT 21.978 62.502 22.022 62.538 ;
      RECT 21.978 63.102 22.022 63.138 ;
      RECT 21.978 63.702 22.022 63.738 ;
      RECT 21.978 64.302 22.022 64.338 ;
      RECT 21.978 64.902 22.022 64.938 ;
      RECT 21.978 65.502 22.022 65.538 ;
      RECT 21.978 66.102 22.022 66.138 ;
      RECT 21.978 66.702 22.022 66.738 ;
      RECT 21.978 67.302 22.022 67.338 ;
      RECT 21.978 67.902 22.022 67.938 ;
      RECT 21.978 68.502 22.022 68.538 ;
      RECT 21.978 69.102 22.022 69.138 ;
      RECT 21.978 69.702 22.022 69.738 ;
      RECT 21.978 70.302 22.022 70.338 ;
      RECT 21.978 70.902 22.022 70.938 ;
      RECT 21.978 71.502 22.022 71.538 ;
      RECT 21.978 72.102 22.022 72.138 ;
      RECT 22.186 33.0435 22.222 33.0795 ;
      RECT 22.186 34.182 22.222 34.218 ;
      RECT 22.186 37.302 22.222 37.338 ;
      RECT 22.186 38.4405 22.222 38.4765 ;
      RECT 22.614 1.558 22.666 1.594 ;
      RECT 22.614 2.758 22.666 2.794 ;
      RECT 22.614 3.958 22.666 3.994 ;
      RECT 22.614 5.158 22.666 5.194 ;
      RECT 22.614 6.358 22.666 6.394 ;
      RECT 22.614 7.558 22.666 7.594 ;
      RECT 22.614 8.758 22.666 8.794 ;
      RECT 22.614 9.958 22.666 9.994 ;
      RECT 22.614 11.158 22.666 11.194 ;
      RECT 22.614 12.358 22.666 12.394 ;
      RECT 22.614 13.558 22.666 13.594 ;
      RECT 22.614 14.758 22.666 14.794 ;
      RECT 22.614 15.958 22.666 15.994 ;
      RECT 22.614 17.158 22.666 17.194 ;
      RECT 22.614 18.358 22.666 18.394 ;
      RECT 22.614 19.558 22.666 19.594 ;
      RECT 22.614 20.758 22.666 20.794 ;
      RECT 22.614 21.958 22.666 21.994 ;
      RECT 22.614 23.158 22.666 23.194 ;
      RECT 22.614 24.358 22.666 24.394 ;
      RECT 22.614 25.558 22.666 25.594 ;
      RECT 22.614 26.758 22.666 26.794 ;
      RECT 22.614 27.958 22.666 27.994 ;
      RECT 22.614 29.158 22.666 29.194 ;
      RECT 22.614 30.358 22.666 30.394 ;
      RECT 22.614 31.558 22.666 31.594 ;
      RECT 22.614 32.622 22.666 32.658 ;
      RECT 22.614 32.862 22.666 32.898 ;
      RECT 22.614 38.622 22.666 38.658 ;
      RECT 22.614 38.862 22.666 38.898 ;
      RECT 22.614 40.678 22.666 40.714 ;
      RECT 22.614 41.878 22.666 41.914 ;
      RECT 22.614 43.078 22.666 43.114 ;
      RECT 22.614 44.278 22.666 44.314 ;
      RECT 22.614 45.478 22.666 45.514 ;
      RECT 22.614 46.678 22.666 46.714 ;
      RECT 22.614 47.878 22.666 47.914 ;
      RECT 22.614 49.078 22.666 49.114 ;
      RECT 22.614 50.278 22.666 50.314 ;
      RECT 22.614 51.478 22.666 51.514 ;
      RECT 22.614 52.678 22.666 52.714 ;
      RECT 22.614 53.878 22.666 53.914 ;
      RECT 22.614 55.078 22.666 55.114 ;
      RECT 22.614 56.278 22.666 56.314 ;
      RECT 22.614 57.478 22.666 57.514 ;
      RECT 22.614 58.678 22.666 58.714 ;
      RECT 22.614 59.878 22.666 59.914 ;
      RECT 22.614 61.078 22.666 61.114 ;
      RECT 22.614 62.278 22.666 62.314 ;
      RECT 22.614 63.478 22.666 63.514 ;
      RECT 22.614 64.678 22.666 64.714 ;
      RECT 22.614 65.878 22.666 65.914 ;
      RECT 22.614 67.078 22.666 67.114 ;
      RECT 22.614 68.278 22.666 68.314 ;
      RECT 22.614 69.478 22.666 69.514 ;
      RECT 22.614 70.678 22.666 70.714 ;
      RECT 22.614 71.878 22.666 71.914 ;
      RECT 22.694 0.806 22.746 0.842 ;
      RECT 22.694 2.006 22.746 2.042 ;
      RECT 22.694 3.206 22.746 3.242 ;
      RECT 22.694 4.406 22.746 4.442 ;
      RECT 22.694 5.606 22.746 5.642 ;
      RECT 22.694 6.806 22.746 6.842 ;
      RECT 22.694 8.006 22.746 8.042 ;
      RECT 22.694 9.206 22.746 9.242 ;
      RECT 22.694 10.406 22.746 10.442 ;
      RECT 22.694 11.606 22.746 11.642 ;
      RECT 22.694 12.806 22.746 12.842 ;
      RECT 22.694 14.006 22.746 14.042 ;
      RECT 22.694 15.206 22.746 15.242 ;
      RECT 22.694 16.406 22.746 16.442 ;
      RECT 22.694 17.606 22.746 17.642 ;
      RECT 22.694 18.806 22.746 18.842 ;
      RECT 22.694 20.006 22.746 20.042 ;
      RECT 22.694 21.206 22.746 21.242 ;
      RECT 22.694 22.406 22.746 22.442 ;
      RECT 22.694 23.606 22.746 23.642 ;
      RECT 22.694 24.806 22.746 24.842 ;
      RECT 22.694 26.006 22.746 26.042 ;
      RECT 22.694 27.206 22.746 27.242 ;
      RECT 22.694 28.406 22.746 28.442 ;
      RECT 22.694 29.606 22.746 29.642 ;
      RECT 22.694 30.806 22.746 30.842 ;
      RECT 22.694 33.342 22.746 33.378 ;
      RECT 22.694 33.582 22.746 33.618 ;
      RECT 22.694 37.902 22.746 37.938 ;
      RECT 22.694 38.142 22.746 38.178 ;
      RECT 22.694 39.926 22.746 39.962 ;
      RECT 22.694 41.126 22.746 41.162 ;
      RECT 22.694 42.326 22.746 42.362 ;
      RECT 22.694 43.526 22.746 43.562 ;
      RECT 22.694 44.726 22.746 44.762 ;
      RECT 22.694 45.926 22.746 45.962 ;
      RECT 22.694 47.126 22.746 47.162 ;
      RECT 22.694 48.326 22.746 48.362 ;
      RECT 22.694 49.526 22.746 49.562 ;
      RECT 22.694 50.726 22.746 50.762 ;
      RECT 22.694 51.926 22.746 51.962 ;
      RECT 22.694 53.126 22.746 53.162 ;
      RECT 22.694 54.326 22.746 54.362 ;
      RECT 22.694 55.526 22.746 55.562 ;
      RECT 22.694 56.726 22.746 56.762 ;
      RECT 22.694 57.926 22.746 57.962 ;
      RECT 22.694 59.126 22.746 59.162 ;
      RECT 22.694 60.326 22.746 60.362 ;
      RECT 22.694 61.526 22.746 61.562 ;
      RECT 22.694 62.726 22.746 62.762 ;
      RECT 22.694 63.926 22.746 63.962 ;
      RECT 22.694 65.126 22.746 65.162 ;
      RECT 22.694 66.326 22.746 66.362 ;
      RECT 22.694 67.526 22.746 67.562 ;
      RECT 22.694 68.726 22.746 68.762 ;
      RECT 22.694 69.926 22.746 69.962 ;
      RECT 22.694 71.126 22.746 71.162 ;
      RECT 22.774 0.281 22.826 0.317 ;
      RECT 22.774 72.403 22.826 72.439 ;
      RECT 22.854 0.806 22.906 0.842 ;
      RECT 22.854 2.006 22.906 2.042 ;
      RECT 22.854 3.206 22.906 3.242 ;
      RECT 22.854 4.406 22.906 4.442 ;
      RECT 22.854 5.606 22.906 5.642 ;
      RECT 22.854 6.806 22.906 6.842 ;
      RECT 22.854 8.006 22.906 8.042 ;
      RECT 22.854 9.206 22.906 9.242 ;
      RECT 22.854 10.406 22.906 10.442 ;
      RECT 22.854 11.606 22.906 11.642 ;
      RECT 22.854 12.806 22.906 12.842 ;
      RECT 22.854 14.006 22.906 14.042 ;
      RECT 22.854 15.206 22.906 15.242 ;
      RECT 22.854 16.406 22.906 16.442 ;
      RECT 22.854 17.606 22.906 17.642 ;
      RECT 22.854 18.806 22.906 18.842 ;
      RECT 22.854 20.006 22.906 20.042 ;
      RECT 22.854 21.206 22.906 21.242 ;
      RECT 22.854 22.406 22.906 22.442 ;
      RECT 22.854 23.606 22.906 23.642 ;
      RECT 22.854 24.806 22.906 24.842 ;
      RECT 22.854 26.006 22.906 26.042 ;
      RECT 22.854 27.206 22.906 27.242 ;
      RECT 22.854 28.406 22.906 28.442 ;
      RECT 22.854 29.606 22.906 29.642 ;
      RECT 22.854 30.806 22.906 30.842 ;
      RECT 22.854 32.622 22.906 32.658 ;
      RECT 22.854 32.862 22.906 32.898 ;
      RECT 22.854 38.622 22.906 38.658 ;
      RECT 22.854 38.862 22.906 38.898 ;
      RECT 22.854 39.926 22.906 39.962 ;
      RECT 22.854 41.126 22.906 41.162 ;
      RECT 22.854 42.326 22.906 42.362 ;
      RECT 22.854 43.526 22.906 43.562 ;
      RECT 22.854 44.726 22.906 44.762 ;
      RECT 22.854 45.926 22.906 45.962 ;
      RECT 22.854 47.126 22.906 47.162 ;
      RECT 22.854 48.326 22.906 48.362 ;
      RECT 22.854 49.526 22.906 49.562 ;
      RECT 22.854 50.726 22.906 50.762 ;
      RECT 22.854 51.926 22.906 51.962 ;
      RECT 22.854 53.126 22.906 53.162 ;
      RECT 22.854 54.326 22.906 54.362 ;
      RECT 22.854 55.526 22.906 55.562 ;
      RECT 22.854 56.726 22.906 56.762 ;
      RECT 22.854 57.926 22.906 57.962 ;
      RECT 22.854 59.126 22.906 59.162 ;
      RECT 22.854 60.326 22.906 60.362 ;
      RECT 22.854 61.526 22.906 61.562 ;
      RECT 22.854 62.726 22.906 62.762 ;
      RECT 22.854 63.926 22.906 63.962 ;
      RECT 22.854 65.126 22.906 65.162 ;
      RECT 22.854 66.326 22.906 66.362 ;
      RECT 22.854 67.526 22.906 67.562 ;
      RECT 22.854 68.726 22.906 68.762 ;
      RECT 22.854 69.926 22.906 69.962 ;
      RECT 22.854 71.126 22.906 71.162 ;
      RECT 22.934 1.558 22.986 1.594 ;
      RECT 22.934 2.758 22.986 2.794 ;
      RECT 22.934 3.958 22.986 3.994 ;
      RECT 22.934 5.158 22.986 5.194 ;
      RECT 22.934 6.358 22.986 6.394 ;
      RECT 22.934 7.558 22.986 7.594 ;
      RECT 22.934 8.758 22.986 8.794 ;
      RECT 22.934 9.958 22.986 9.994 ;
      RECT 22.934 11.158 22.986 11.194 ;
      RECT 22.934 12.358 22.986 12.394 ;
      RECT 22.934 13.558 22.986 13.594 ;
      RECT 22.934 14.758 22.986 14.794 ;
      RECT 22.934 15.958 22.986 15.994 ;
      RECT 22.934 17.158 22.986 17.194 ;
      RECT 22.934 18.358 22.986 18.394 ;
      RECT 22.934 19.558 22.986 19.594 ;
      RECT 22.934 20.758 22.986 20.794 ;
      RECT 22.934 21.958 22.986 21.994 ;
      RECT 22.934 23.158 22.986 23.194 ;
      RECT 22.934 24.358 22.986 24.394 ;
      RECT 22.934 25.558 22.986 25.594 ;
      RECT 22.934 26.758 22.986 26.794 ;
      RECT 22.934 27.958 22.986 27.994 ;
      RECT 22.934 29.158 22.986 29.194 ;
      RECT 22.934 30.358 22.986 30.394 ;
      RECT 22.934 31.558 22.986 31.594 ;
      RECT 22.934 33.342 22.986 33.378 ;
      RECT 22.934 33.582 22.986 33.618 ;
      RECT 22.934 37.902 22.986 37.938 ;
      RECT 22.934 38.142 22.986 38.178 ;
      RECT 22.934 40.678 22.986 40.714 ;
      RECT 22.934 41.878 22.986 41.914 ;
      RECT 22.934 43.078 22.986 43.114 ;
      RECT 22.934 44.278 22.986 44.314 ;
      RECT 22.934 45.478 22.986 45.514 ;
      RECT 22.934 46.678 22.986 46.714 ;
      RECT 22.934 47.878 22.986 47.914 ;
      RECT 22.934 49.078 22.986 49.114 ;
      RECT 22.934 50.278 22.986 50.314 ;
      RECT 22.934 51.478 22.986 51.514 ;
      RECT 22.934 52.678 22.986 52.714 ;
      RECT 22.934 53.878 22.986 53.914 ;
      RECT 22.934 55.078 22.986 55.114 ;
      RECT 22.934 56.278 22.986 56.314 ;
      RECT 22.934 57.478 22.986 57.514 ;
      RECT 22.934 58.678 22.986 58.714 ;
      RECT 22.934 59.878 22.986 59.914 ;
      RECT 22.934 61.078 22.986 61.114 ;
      RECT 22.934 62.278 22.986 62.314 ;
      RECT 22.934 63.478 22.986 63.514 ;
      RECT 22.934 64.678 22.986 64.714 ;
      RECT 22.934 65.878 22.986 65.914 ;
      RECT 22.934 67.078 22.986 67.114 ;
      RECT 22.934 68.278 22.986 68.314 ;
      RECT 22.934 69.478 22.986 69.514 ;
      RECT 22.934 70.678 22.986 70.714 ;
      RECT 22.934 71.878 22.986 71.914 ;
      RECT 23.014 0.806 23.066 0.842 ;
      RECT 23.014 2.006 23.066 2.042 ;
      RECT 23.014 3.206 23.066 3.242 ;
      RECT 23.014 4.406 23.066 4.442 ;
      RECT 23.014 5.606 23.066 5.642 ;
      RECT 23.014 6.806 23.066 6.842 ;
      RECT 23.014 8.006 23.066 8.042 ;
      RECT 23.014 9.206 23.066 9.242 ;
      RECT 23.014 10.406 23.066 10.442 ;
      RECT 23.014 11.606 23.066 11.642 ;
      RECT 23.014 12.806 23.066 12.842 ;
      RECT 23.014 14.006 23.066 14.042 ;
      RECT 23.014 15.206 23.066 15.242 ;
      RECT 23.014 16.406 23.066 16.442 ;
      RECT 23.014 17.606 23.066 17.642 ;
      RECT 23.014 18.806 23.066 18.842 ;
      RECT 23.014 20.006 23.066 20.042 ;
      RECT 23.014 21.206 23.066 21.242 ;
      RECT 23.014 22.406 23.066 22.442 ;
      RECT 23.014 23.606 23.066 23.642 ;
      RECT 23.014 24.806 23.066 24.842 ;
      RECT 23.014 26.006 23.066 26.042 ;
      RECT 23.014 27.206 23.066 27.242 ;
      RECT 23.014 28.406 23.066 28.442 ;
      RECT 23.014 29.606 23.066 29.642 ;
      RECT 23.014 30.806 23.066 30.842 ;
      RECT 23.014 32.622 23.066 32.658 ;
      RECT 23.014 32.862 23.066 32.898 ;
      RECT 23.014 38.622 23.066 38.658 ;
      RECT 23.014 38.862 23.066 38.898 ;
      RECT 23.014 39.926 23.066 39.962 ;
      RECT 23.014 41.126 23.066 41.162 ;
      RECT 23.014 42.326 23.066 42.362 ;
      RECT 23.014 43.526 23.066 43.562 ;
      RECT 23.014 44.726 23.066 44.762 ;
      RECT 23.014 45.926 23.066 45.962 ;
      RECT 23.014 47.126 23.066 47.162 ;
      RECT 23.014 48.326 23.066 48.362 ;
      RECT 23.014 49.526 23.066 49.562 ;
      RECT 23.014 50.726 23.066 50.762 ;
      RECT 23.014 51.926 23.066 51.962 ;
      RECT 23.014 53.126 23.066 53.162 ;
      RECT 23.014 54.326 23.066 54.362 ;
      RECT 23.014 55.526 23.066 55.562 ;
      RECT 23.014 56.726 23.066 56.762 ;
      RECT 23.014 57.926 23.066 57.962 ;
      RECT 23.014 59.126 23.066 59.162 ;
      RECT 23.014 60.326 23.066 60.362 ;
      RECT 23.014 61.526 23.066 61.562 ;
      RECT 23.014 62.726 23.066 62.762 ;
      RECT 23.014 63.926 23.066 63.962 ;
      RECT 23.014 65.126 23.066 65.162 ;
      RECT 23.014 66.326 23.066 66.362 ;
      RECT 23.014 67.526 23.066 67.562 ;
      RECT 23.014 68.726 23.066 68.762 ;
      RECT 23.014 69.926 23.066 69.962 ;
      RECT 23.014 71.126 23.066 71.162 ;
      RECT 23.094 1.558 23.146 1.594 ;
      RECT 23.094 2.758 23.146 2.794 ;
      RECT 23.094 3.958 23.146 3.994 ;
      RECT 23.094 5.158 23.146 5.194 ;
      RECT 23.094 6.358 23.146 6.394 ;
      RECT 23.094 7.558 23.146 7.594 ;
      RECT 23.094 8.758 23.146 8.794 ;
      RECT 23.094 9.958 23.146 9.994 ;
      RECT 23.094 11.158 23.146 11.194 ;
      RECT 23.094 12.358 23.146 12.394 ;
      RECT 23.094 13.558 23.146 13.594 ;
      RECT 23.094 14.758 23.146 14.794 ;
      RECT 23.094 15.958 23.146 15.994 ;
      RECT 23.094 17.158 23.146 17.194 ;
      RECT 23.094 18.358 23.146 18.394 ;
      RECT 23.094 19.558 23.146 19.594 ;
      RECT 23.094 20.758 23.146 20.794 ;
      RECT 23.094 21.958 23.146 21.994 ;
      RECT 23.094 23.158 23.146 23.194 ;
      RECT 23.094 24.358 23.146 24.394 ;
      RECT 23.094 25.558 23.146 25.594 ;
      RECT 23.094 26.758 23.146 26.794 ;
      RECT 23.094 27.958 23.146 27.994 ;
      RECT 23.094 29.158 23.146 29.194 ;
      RECT 23.094 30.358 23.146 30.394 ;
      RECT 23.094 31.558 23.146 31.594 ;
      RECT 23.094 33.342 23.146 33.378 ;
      RECT 23.094 33.582 23.146 33.618 ;
      RECT 23.094 37.902 23.146 37.938 ;
      RECT 23.094 38.142 23.146 38.178 ;
      RECT 23.094 40.678 23.146 40.714 ;
      RECT 23.094 41.878 23.146 41.914 ;
      RECT 23.094 43.078 23.146 43.114 ;
      RECT 23.094 44.278 23.146 44.314 ;
      RECT 23.094 45.478 23.146 45.514 ;
      RECT 23.094 46.678 23.146 46.714 ;
      RECT 23.094 47.878 23.146 47.914 ;
      RECT 23.094 49.078 23.146 49.114 ;
      RECT 23.094 50.278 23.146 50.314 ;
      RECT 23.094 51.478 23.146 51.514 ;
      RECT 23.094 52.678 23.146 52.714 ;
      RECT 23.094 53.878 23.146 53.914 ;
      RECT 23.094 55.078 23.146 55.114 ;
      RECT 23.094 56.278 23.146 56.314 ;
      RECT 23.094 57.478 23.146 57.514 ;
      RECT 23.094 58.678 23.146 58.714 ;
      RECT 23.094 59.878 23.146 59.914 ;
      RECT 23.094 61.078 23.146 61.114 ;
      RECT 23.094 62.278 23.146 62.314 ;
      RECT 23.094 63.478 23.146 63.514 ;
      RECT 23.094 64.678 23.146 64.714 ;
      RECT 23.094 65.878 23.146 65.914 ;
      RECT 23.094 67.078 23.146 67.114 ;
      RECT 23.094 68.278 23.146 68.314 ;
      RECT 23.094 69.478 23.146 69.514 ;
      RECT 23.094 70.678 23.146 70.714 ;
      RECT 23.094 71.878 23.146 71.914 ;
      RECT 23.174 0.281 23.226 0.317 ;
      RECT 23.174 72.403 23.226 72.439 ;
      RECT 23.254 0.806 23.306 0.842 ;
      RECT 23.254 2.006 23.306 2.042 ;
      RECT 23.254 3.206 23.306 3.242 ;
      RECT 23.254 4.406 23.306 4.442 ;
      RECT 23.254 5.606 23.306 5.642 ;
      RECT 23.254 6.806 23.306 6.842 ;
      RECT 23.254 8.006 23.306 8.042 ;
      RECT 23.254 9.206 23.306 9.242 ;
      RECT 23.254 10.406 23.306 10.442 ;
      RECT 23.254 11.606 23.306 11.642 ;
      RECT 23.254 12.806 23.306 12.842 ;
      RECT 23.254 14.006 23.306 14.042 ;
      RECT 23.254 15.206 23.306 15.242 ;
      RECT 23.254 16.406 23.306 16.442 ;
      RECT 23.254 17.606 23.306 17.642 ;
      RECT 23.254 18.806 23.306 18.842 ;
      RECT 23.254 20.006 23.306 20.042 ;
      RECT 23.254 21.206 23.306 21.242 ;
      RECT 23.254 22.406 23.306 22.442 ;
      RECT 23.254 23.606 23.306 23.642 ;
      RECT 23.254 24.806 23.306 24.842 ;
      RECT 23.254 26.006 23.306 26.042 ;
      RECT 23.254 27.206 23.306 27.242 ;
      RECT 23.254 28.406 23.306 28.442 ;
      RECT 23.254 29.606 23.306 29.642 ;
      RECT 23.254 30.806 23.306 30.842 ;
      RECT 23.254 32.622 23.306 32.658 ;
      RECT 23.254 32.862 23.306 32.898 ;
      RECT 23.254 34.302 23.306 34.338 ;
      RECT 23.254 34.782 23.306 34.818 ;
      RECT 23.254 36.702 23.306 36.738 ;
      RECT 23.254 37.182 23.306 37.218 ;
      RECT 23.254 38.622 23.306 38.658 ;
      RECT 23.254 38.862 23.306 38.898 ;
      RECT 23.254 39.926 23.306 39.962 ;
      RECT 23.254 41.126 23.306 41.162 ;
      RECT 23.254 42.326 23.306 42.362 ;
      RECT 23.254 43.526 23.306 43.562 ;
      RECT 23.254 44.726 23.306 44.762 ;
      RECT 23.254 45.926 23.306 45.962 ;
      RECT 23.254 47.126 23.306 47.162 ;
      RECT 23.254 48.326 23.306 48.362 ;
      RECT 23.254 49.526 23.306 49.562 ;
      RECT 23.254 50.726 23.306 50.762 ;
      RECT 23.254 51.926 23.306 51.962 ;
      RECT 23.254 53.126 23.306 53.162 ;
      RECT 23.254 54.326 23.306 54.362 ;
      RECT 23.254 55.526 23.306 55.562 ;
      RECT 23.254 56.726 23.306 56.762 ;
      RECT 23.254 57.926 23.306 57.962 ;
      RECT 23.254 59.126 23.306 59.162 ;
      RECT 23.254 60.326 23.306 60.362 ;
      RECT 23.254 61.526 23.306 61.562 ;
      RECT 23.254 62.726 23.306 62.762 ;
      RECT 23.254 63.926 23.306 63.962 ;
      RECT 23.254 65.126 23.306 65.162 ;
      RECT 23.254 66.326 23.306 66.362 ;
      RECT 23.254 67.526 23.306 67.562 ;
      RECT 23.254 68.726 23.306 68.762 ;
      RECT 23.254 69.926 23.306 69.962 ;
      RECT 23.254 71.126 23.306 71.162 ;
      RECT 23.334 1.558 23.386 1.594 ;
      RECT 23.334 2.758 23.386 2.794 ;
      RECT 23.334 3.958 23.386 3.994 ;
      RECT 23.334 5.158 23.386 5.194 ;
      RECT 23.334 6.358 23.386 6.394 ;
      RECT 23.334 7.558 23.386 7.594 ;
      RECT 23.334 8.758 23.386 8.794 ;
      RECT 23.334 9.958 23.386 9.994 ;
      RECT 23.334 11.158 23.386 11.194 ;
      RECT 23.334 12.358 23.386 12.394 ;
      RECT 23.334 13.558 23.386 13.594 ;
      RECT 23.334 14.758 23.386 14.794 ;
      RECT 23.334 15.958 23.386 15.994 ;
      RECT 23.334 17.158 23.386 17.194 ;
      RECT 23.334 18.358 23.386 18.394 ;
      RECT 23.334 19.558 23.386 19.594 ;
      RECT 23.334 20.758 23.386 20.794 ;
      RECT 23.334 21.958 23.386 21.994 ;
      RECT 23.334 23.158 23.386 23.194 ;
      RECT 23.334 24.358 23.386 24.394 ;
      RECT 23.334 25.558 23.386 25.594 ;
      RECT 23.334 26.758 23.386 26.794 ;
      RECT 23.334 27.958 23.386 27.994 ;
      RECT 23.334 29.158 23.386 29.194 ;
      RECT 23.334 30.358 23.386 30.394 ;
      RECT 23.334 31.558 23.386 31.594 ;
      RECT 23.334 33.342 23.386 33.378 ;
      RECT 23.334 33.582 23.386 33.618 ;
      RECT 23.334 37.902 23.386 37.938 ;
      RECT 23.334 38.142 23.386 38.178 ;
      RECT 23.334 40.678 23.386 40.714 ;
      RECT 23.334 41.878 23.386 41.914 ;
      RECT 23.334 43.078 23.386 43.114 ;
      RECT 23.334 44.278 23.386 44.314 ;
      RECT 23.334 45.478 23.386 45.514 ;
      RECT 23.334 46.678 23.386 46.714 ;
      RECT 23.334 47.878 23.386 47.914 ;
      RECT 23.334 49.078 23.386 49.114 ;
      RECT 23.334 50.278 23.386 50.314 ;
      RECT 23.334 51.478 23.386 51.514 ;
      RECT 23.334 52.678 23.386 52.714 ;
      RECT 23.334 53.878 23.386 53.914 ;
      RECT 23.334 55.078 23.386 55.114 ;
      RECT 23.334 56.278 23.386 56.314 ;
      RECT 23.334 57.478 23.386 57.514 ;
      RECT 23.334 58.678 23.386 58.714 ;
      RECT 23.334 59.878 23.386 59.914 ;
      RECT 23.334 61.078 23.386 61.114 ;
      RECT 23.334 62.278 23.386 62.314 ;
      RECT 23.334 63.478 23.386 63.514 ;
      RECT 23.334 64.678 23.386 64.714 ;
      RECT 23.334 65.878 23.386 65.914 ;
      RECT 23.334 67.078 23.386 67.114 ;
      RECT 23.334 68.278 23.386 68.314 ;
      RECT 23.334 69.478 23.386 69.514 ;
      RECT 23.334 70.678 23.386 70.714 ;
      RECT 23.334 71.878 23.386 71.914 ;
      RECT 23.414 0.806 23.466 0.842 ;
      RECT 23.414 2.006 23.466 2.042 ;
      RECT 23.414 3.206 23.466 3.242 ;
      RECT 23.414 4.406 23.466 4.442 ;
      RECT 23.414 5.606 23.466 5.642 ;
      RECT 23.414 6.806 23.466 6.842 ;
      RECT 23.414 8.006 23.466 8.042 ;
      RECT 23.414 9.206 23.466 9.242 ;
      RECT 23.414 10.406 23.466 10.442 ;
      RECT 23.414 11.606 23.466 11.642 ;
      RECT 23.414 12.806 23.466 12.842 ;
      RECT 23.414 14.006 23.466 14.042 ;
      RECT 23.414 15.206 23.466 15.242 ;
      RECT 23.414 16.406 23.466 16.442 ;
      RECT 23.414 17.606 23.466 17.642 ;
      RECT 23.414 18.806 23.466 18.842 ;
      RECT 23.414 20.006 23.466 20.042 ;
      RECT 23.414 21.206 23.466 21.242 ;
      RECT 23.414 22.406 23.466 22.442 ;
      RECT 23.414 23.606 23.466 23.642 ;
      RECT 23.414 24.806 23.466 24.842 ;
      RECT 23.414 26.006 23.466 26.042 ;
      RECT 23.414 27.206 23.466 27.242 ;
      RECT 23.414 28.406 23.466 28.442 ;
      RECT 23.414 29.606 23.466 29.642 ;
      RECT 23.414 30.806 23.466 30.842 ;
      RECT 23.414 32.622 23.466 32.658 ;
      RECT 23.414 32.862 23.466 32.898 ;
      RECT 23.414 38.622 23.466 38.658 ;
      RECT 23.414 38.862 23.466 38.898 ;
      RECT 23.414 39.926 23.466 39.962 ;
      RECT 23.414 41.126 23.466 41.162 ;
      RECT 23.414 42.326 23.466 42.362 ;
      RECT 23.414 43.526 23.466 43.562 ;
      RECT 23.414 44.726 23.466 44.762 ;
      RECT 23.414 45.926 23.466 45.962 ;
      RECT 23.414 47.126 23.466 47.162 ;
      RECT 23.414 48.326 23.466 48.362 ;
      RECT 23.414 49.526 23.466 49.562 ;
      RECT 23.414 50.726 23.466 50.762 ;
      RECT 23.414 51.926 23.466 51.962 ;
      RECT 23.414 53.126 23.466 53.162 ;
      RECT 23.414 54.326 23.466 54.362 ;
      RECT 23.414 55.526 23.466 55.562 ;
      RECT 23.414 56.726 23.466 56.762 ;
      RECT 23.414 57.926 23.466 57.962 ;
      RECT 23.414 59.126 23.466 59.162 ;
      RECT 23.414 60.326 23.466 60.362 ;
      RECT 23.414 61.526 23.466 61.562 ;
      RECT 23.414 62.726 23.466 62.762 ;
      RECT 23.414 63.926 23.466 63.962 ;
      RECT 23.414 65.126 23.466 65.162 ;
      RECT 23.414 66.326 23.466 66.362 ;
      RECT 23.414 67.526 23.466 67.562 ;
      RECT 23.414 68.726 23.466 68.762 ;
      RECT 23.414 69.926 23.466 69.962 ;
      RECT 23.414 71.126 23.466 71.162 ;
      RECT 23.494 1.558 23.546 1.594 ;
      RECT 23.494 2.758 23.546 2.794 ;
      RECT 23.494 3.958 23.546 3.994 ;
      RECT 23.494 5.158 23.546 5.194 ;
      RECT 23.494 6.358 23.546 6.394 ;
      RECT 23.494 7.558 23.546 7.594 ;
      RECT 23.494 8.758 23.546 8.794 ;
      RECT 23.494 9.958 23.546 9.994 ;
      RECT 23.494 11.158 23.546 11.194 ;
      RECT 23.494 12.358 23.546 12.394 ;
      RECT 23.494 13.558 23.546 13.594 ;
      RECT 23.494 14.758 23.546 14.794 ;
      RECT 23.494 15.958 23.546 15.994 ;
      RECT 23.494 17.158 23.546 17.194 ;
      RECT 23.494 18.358 23.546 18.394 ;
      RECT 23.494 19.558 23.546 19.594 ;
      RECT 23.494 20.758 23.546 20.794 ;
      RECT 23.494 21.958 23.546 21.994 ;
      RECT 23.494 23.158 23.546 23.194 ;
      RECT 23.494 24.358 23.546 24.394 ;
      RECT 23.494 25.558 23.546 25.594 ;
      RECT 23.494 26.758 23.546 26.794 ;
      RECT 23.494 27.958 23.546 27.994 ;
      RECT 23.494 29.158 23.546 29.194 ;
      RECT 23.494 30.358 23.546 30.394 ;
      RECT 23.494 31.558 23.546 31.594 ;
      RECT 23.494 33.342 23.546 33.378 ;
      RECT 23.494 33.582 23.546 33.618 ;
      RECT 23.494 37.902 23.546 37.938 ;
      RECT 23.494 38.142 23.546 38.178 ;
      RECT 23.494 40.678 23.546 40.714 ;
      RECT 23.494 41.878 23.546 41.914 ;
      RECT 23.494 43.078 23.546 43.114 ;
      RECT 23.494 44.278 23.546 44.314 ;
      RECT 23.494 45.478 23.546 45.514 ;
      RECT 23.494 46.678 23.546 46.714 ;
      RECT 23.494 47.878 23.546 47.914 ;
      RECT 23.494 49.078 23.546 49.114 ;
      RECT 23.494 50.278 23.546 50.314 ;
      RECT 23.494 51.478 23.546 51.514 ;
      RECT 23.494 52.678 23.546 52.714 ;
      RECT 23.494 53.878 23.546 53.914 ;
      RECT 23.494 55.078 23.546 55.114 ;
      RECT 23.494 56.278 23.546 56.314 ;
      RECT 23.494 57.478 23.546 57.514 ;
      RECT 23.494 58.678 23.546 58.714 ;
      RECT 23.494 59.878 23.546 59.914 ;
      RECT 23.494 61.078 23.546 61.114 ;
      RECT 23.494 62.278 23.546 62.314 ;
      RECT 23.494 63.478 23.546 63.514 ;
      RECT 23.494 64.678 23.546 64.714 ;
      RECT 23.494 65.878 23.546 65.914 ;
      RECT 23.494 67.078 23.546 67.114 ;
      RECT 23.494 68.278 23.546 68.314 ;
      RECT 23.494 69.478 23.546 69.514 ;
      RECT 23.494 70.678 23.546 70.714 ;
      RECT 23.494 71.878 23.546 71.914 ;
      RECT 23.574 0.281 23.626 0.317 ;
      RECT 23.574 72.403 23.626 72.439 ;
      RECT 23.654 0.806 23.706 0.842 ;
      RECT 23.654 2.006 23.706 2.042 ;
      RECT 23.654 3.206 23.706 3.242 ;
      RECT 23.654 4.406 23.706 4.442 ;
      RECT 23.654 5.606 23.706 5.642 ;
      RECT 23.654 6.806 23.706 6.842 ;
      RECT 23.654 8.006 23.706 8.042 ;
      RECT 23.654 9.206 23.706 9.242 ;
      RECT 23.654 10.406 23.706 10.442 ;
      RECT 23.654 11.606 23.706 11.642 ;
      RECT 23.654 12.806 23.706 12.842 ;
      RECT 23.654 14.006 23.706 14.042 ;
      RECT 23.654 15.206 23.706 15.242 ;
      RECT 23.654 16.406 23.706 16.442 ;
      RECT 23.654 17.606 23.706 17.642 ;
      RECT 23.654 18.806 23.706 18.842 ;
      RECT 23.654 20.006 23.706 20.042 ;
      RECT 23.654 21.206 23.706 21.242 ;
      RECT 23.654 22.406 23.706 22.442 ;
      RECT 23.654 23.606 23.706 23.642 ;
      RECT 23.654 24.806 23.706 24.842 ;
      RECT 23.654 26.006 23.706 26.042 ;
      RECT 23.654 27.206 23.706 27.242 ;
      RECT 23.654 28.406 23.706 28.442 ;
      RECT 23.654 29.606 23.706 29.642 ;
      RECT 23.654 30.806 23.706 30.842 ;
      RECT 23.654 32.622 23.706 32.658 ;
      RECT 23.654 32.862 23.706 32.898 ;
      RECT 23.654 38.622 23.706 38.658 ;
      RECT 23.654 38.862 23.706 38.898 ;
      RECT 23.654 39.926 23.706 39.962 ;
      RECT 23.654 41.126 23.706 41.162 ;
      RECT 23.654 42.326 23.706 42.362 ;
      RECT 23.654 43.526 23.706 43.562 ;
      RECT 23.654 44.726 23.706 44.762 ;
      RECT 23.654 45.926 23.706 45.962 ;
      RECT 23.654 47.126 23.706 47.162 ;
      RECT 23.654 48.326 23.706 48.362 ;
      RECT 23.654 49.526 23.706 49.562 ;
      RECT 23.654 50.726 23.706 50.762 ;
      RECT 23.654 51.926 23.706 51.962 ;
      RECT 23.654 53.126 23.706 53.162 ;
      RECT 23.654 54.326 23.706 54.362 ;
      RECT 23.654 55.526 23.706 55.562 ;
      RECT 23.654 56.726 23.706 56.762 ;
      RECT 23.654 57.926 23.706 57.962 ;
      RECT 23.654 59.126 23.706 59.162 ;
      RECT 23.654 60.326 23.706 60.362 ;
      RECT 23.654 61.526 23.706 61.562 ;
      RECT 23.654 62.726 23.706 62.762 ;
      RECT 23.654 63.926 23.706 63.962 ;
      RECT 23.654 65.126 23.706 65.162 ;
      RECT 23.654 66.326 23.706 66.362 ;
      RECT 23.654 67.526 23.706 67.562 ;
      RECT 23.654 68.726 23.706 68.762 ;
      RECT 23.654 69.926 23.706 69.962 ;
      RECT 23.654 71.126 23.706 71.162 ;
      RECT 23.734 1.558 23.786 1.594 ;
      RECT 23.734 2.758 23.786 2.794 ;
      RECT 23.734 3.958 23.786 3.994 ;
      RECT 23.734 5.158 23.786 5.194 ;
      RECT 23.734 6.358 23.786 6.394 ;
      RECT 23.734 7.558 23.786 7.594 ;
      RECT 23.734 8.758 23.786 8.794 ;
      RECT 23.734 9.958 23.786 9.994 ;
      RECT 23.734 11.158 23.786 11.194 ;
      RECT 23.734 12.358 23.786 12.394 ;
      RECT 23.734 13.558 23.786 13.594 ;
      RECT 23.734 14.758 23.786 14.794 ;
      RECT 23.734 15.958 23.786 15.994 ;
      RECT 23.734 17.158 23.786 17.194 ;
      RECT 23.734 18.358 23.786 18.394 ;
      RECT 23.734 19.558 23.786 19.594 ;
      RECT 23.734 20.758 23.786 20.794 ;
      RECT 23.734 21.958 23.786 21.994 ;
      RECT 23.734 23.158 23.786 23.194 ;
      RECT 23.734 24.358 23.786 24.394 ;
      RECT 23.734 25.558 23.786 25.594 ;
      RECT 23.734 26.758 23.786 26.794 ;
      RECT 23.734 27.958 23.786 27.994 ;
      RECT 23.734 29.158 23.786 29.194 ;
      RECT 23.734 30.358 23.786 30.394 ;
      RECT 23.734 31.558 23.786 31.594 ;
      RECT 23.734 33.342 23.786 33.378 ;
      RECT 23.734 33.582 23.786 33.618 ;
      RECT 23.734 37.902 23.786 37.938 ;
      RECT 23.734 38.142 23.786 38.178 ;
      RECT 23.734 40.678 23.786 40.714 ;
      RECT 23.734 41.878 23.786 41.914 ;
      RECT 23.734 43.078 23.786 43.114 ;
      RECT 23.734 44.278 23.786 44.314 ;
      RECT 23.734 45.478 23.786 45.514 ;
      RECT 23.734 46.678 23.786 46.714 ;
      RECT 23.734 47.878 23.786 47.914 ;
      RECT 23.734 49.078 23.786 49.114 ;
      RECT 23.734 50.278 23.786 50.314 ;
      RECT 23.734 51.478 23.786 51.514 ;
      RECT 23.734 52.678 23.786 52.714 ;
      RECT 23.734 53.878 23.786 53.914 ;
      RECT 23.734 55.078 23.786 55.114 ;
      RECT 23.734 56.278 23.786 56.314 ;
      RECT 23.734 57.478 23.786 57.514 ;
      RECT 23.734 58.678 23.786 58.714 ;
      RECT 23.734 59.878 23.786 59.914 ;
      RECT 23.734 61.078 23.786 61.114 ;
      RECT 23.734 62.278 23.786 62.314 ;
      RECT 23.734 63.478 23.786 63.514 ;
      RECT 23.734 64.678 23.786 64.714 ;
      RECT 23.734 65.878 23.786 65.914 ;
      RECT 23.734 67.078 23.786 67.114 ;
      RECT 23.734 68.278 23.786 68.314 ;
      RECT 23.734 69.478 23.786 69.514 ;
      RECT 23.734 70.678 23.786 70.714 ;
      RECT 23.734 71.878 23.786 71.914 ;
      RECT 23.814 0.806 23.866 0.842 ;
      RECT 23.814 2.006 23.866 2.042 ;
      RECT 23.814 3.206 23.866 3.242 ;
      RECT 23.814 4.406 23.866 4.442 ;
      RECT 23.814 5.606 23.866 5.642 ;
      RECT 23.814 6.806 23.866 6.842 ;
      RECT 23.814 8.006 23.866 8.042 ;
      RECT 23.814 9.206 23.866 9.242 ;
      RECT 23.814 10.406 23.866 10.442 ;
      RECT 23.814 11.606 23.866 11.642 ;
      RECT 23.814 12.806 23.866 12.842 ;
      RECT 23.814 14.006 23.866 14.042 ;
      RECT 23.814 15.206 23.866 15.242 ;
      RECT 23.814 16.406 23.866 16.442 ;
      RECT 23.814 17.606 23.866 17.642 ;
      RECT 23.814 18.806 23.866 18.842 ;
      RECT 23.814 20.006 23.866 20.042 ;
      RECT 23.814 21.206 23.866 21.242 ;
      RECT 23.814 22.406 23.866 22.442 ;
      RECT 23.814 23.606 23.866 23.642 ;
      RECT 23.814 24.806 23.866 24.842 ;
      RECT 23.814 26.006 23.866 26.042 ;
      RECT 23.814 27.206 23.866 27.242 ;
      RECT 23.814 28.406 23.866 28.442 ;
      RECT 23.814 29.606 23.866 29.642 ;
      RECT 23.814 30.806 23.866 30.842 ;
      RECT 23.814 32.622 23.866 32.658 ;
      RECT 23.814 32.862 23.866 32.898 ;
      RECT 23.814 38.622 23.866 38.658 ;
      RECT 23.814 38.862 23.866 38.898 ;
      RECT 23.814 39.926 23.866 39.962 ;
      RECT 23.814 41.126 23.866 41.162 ;
      RECT 23.814 42.326 23.866 42.362 ;
      RECT 23.814 43.526 23.866 43.562 ;
      RECT 23.814 44.726 23.866 44.762 ;
      RECT 23.814 45.926 23.866 45.962 ;
      RECT 23.814 47.126 23.866 47.162 ;
      RECT 23.814 48.326 23.866 48.362 ;
      RECT 23.814 49.526 23.866 49.562 ;
      RECT 23.814 50.726 23.866 50.762 ;
      RECT 23.814 51.926 23.866 51.962 ;
      RECT 23.814 53.126 23.866 53.162 ;
      RECT 23.814 54.326 23.866 54.362 ;
      RECT 23.814 55.526 23.866 55.562 ;
      RECT 23.814 56.726 23.866 56.762 ;
      RECT 23.814 57.926 23.866 57.962 ;
      RECT 23.814 59.126 23.866 59.162 ;
      RECT 23.814 60.326 23.866 60.362 ;
      RECT 23.814 61.526 23.866 61.562 ;
      RECT 23.814 62.726 23.866 62.762 ;
      RECT 23.814 63.926 23.866 63.962 ;
      RECT 23.814 65.126 23.866 65.162 ;
      RECT 23.814 66.326 23.866 66.362 ;
      RECT 23.814 67.526 23.866 67.562 ;
      RECT 23.814 68.726 23.866 68.762 ;
      RECT 23.814 69.926 23.866 69.962 ;
      RECT 23.814 71.126 23.866 71.162 ;
      RECT 23.894 1.558 23.946 1.594 ;
      RECT 23.894 2.758 23.946 2.794 ;
      RECT 23.894 3.958 23.946 3.994 ;
      RECT 23.894 5.158 23.946 5.194 ;
      RECT 23.894 6.358 23.946 6.394 ;
      RECT 23.894 7.558 23.946 7.594 ;
      RECT 23.894 8.758 23.946 8.794 ;
      RECT 23.894 9.958 23.946 9.994 ;
      RECT 23.894 11.158 23.946 11.194 ;
      RECT 23.894 12.358 23.946 12.394 ;
      RECT 23.894 13.558 23.946 13.594 ;
      RECT 23.894 14.758 23.946 14.794 ;
      RECT 23.894 15.958 23.946 15.994 ;
      RECT 23.894 17.158 23.946 17.194 ;
      RECT 23.894 18.358 23.946 18.394 ;
      RECT 23.894 19.558 23.946 19.594 ;
      RECT 23.894 20.758 23.946 20.794 ;
      RECT 23.894 21.958 23.946 21.994 ;
      RECT 23.894 23.158 23.946 23.194 ;
      RECT 23.894 24.358 23.946 24.394 ;
      RECT 23.894 25.558 23.946 25.594 ;
      RECT 23.894 26.758 23.946 26.794 ;
      RECT 23.894 27.958 23.946 27.994 ;
      RECT 23.894 29.158 23.946 29.194 ;
      RECT 23.894 30.358 23.946 30.394 ;
      RECT 23.894 31.558 23.946 31.594 ;
      RECT 23.894 33.342 23.946 33.378 ;
      RECT 23.894 33.582 23.946 33.618 ;
      RECT 23.894 37.902 23.946 37.938 ;
      RECT 23.894 38.142 23.946 38.178 ;
      RECT 23.894 40.678 23.946 40.714 ;
      RECT 23.894 41.878 23.946 41.914 ;
      RECT 23.894 43.078 23.946 43.114 ;
      RECT 23.894 44.278 23.946 44.314 ;
      RECT 23.894 45.478 23.946 45.514 ;
      RECT 23.894 46.678 23.946 46.714 ;
      RECT 23.894 47.878 23.946 47.914 ;
      RECT 23.894 49.078 23.946 49.114 ;
      RECT 23.894 50.278 23.946 50.314 ;
      RECT 23.894 51.478 23.946 51.514 ;
      RECT 23.894 52.678 23.946 52.714 ;
      RECT 23.894 53.878 23.946 53.914 ;
      RECT 23.894 55.078 23.946 55.114 ;
      RECT 23.894 56.278 23.946 56.314 ;
      RECT 23.894 57.478 23.946 57.514 ;
      RECT 23.894 58.678 23.946 58.714 ;
      RECT 23.894 59.878 23.946 59.914 ;
      RECT 23.894 61.078 23.946 61.114 ;
      RECT 23.894 62.278 23.946 62.314 ;
      RECT 23.894 63.478 23.946 63.514 ;
      RECT 23.894 64.678 23.946 64.714 ;
      RECT 23.894 65.878 23.946 65.914 ;
      RECT 23.894 67.078 23.946 67.114 ;
      RECT 23.894 68.278 23.946 68.314 ;
      RECT 23.894 69.478 23.946 69.514 ;
      RECT 23.894 70.678 23.946 70.714 ;
      RECT 23.894 71.878 23.946 71.914 ;
      RECT 23.974 0.281 24.026 0.317 ;
      RECT 23.974 72.403 24.026 72.439 ;
      RECT 24.054 0.806 24.106 0.842 ;
      RECT 24.054 2.006 24.106 2.042 ;
      RECT 24.054 3.206 24.106 3.242 ;
      RECT 24.054 4.406 24.106 4.442 ;
      RECT 24.054 5.606 24.106 5.642 ;
      RECT 24.054 6.806 24.106 6.842 ;
      RECT 24.054 8.006 24.106 8.042 ;
      RECT 24.054 9.206 24.106 9.242 ;
      RECT 24.054 10.406 24.106 10.442 ;
      RECT 24.054 11.606 24.106 11.642 ;
      RECT 24.054 12.806 24.106 12.842 ;
      RECT 24.054 14.006 24.106 14.042 ;
      RECT 24.054 15.206 24.106 15.242 ;
      RECT 24.054 16.406 24.106 16.442 ;
      RECT 24.054 17.606 24.106 17.642 ;
      RECT 24.054 18.806 24.106 18.842 ;
      RECT 24.054 20.006 24.106 20.042 ;
      RECT 24.054 21.206 24.106 21.242 ;
      RECT 24.054 22.406 24.106 22.442 ;
      RECT 24.054 23.606 24.106 23.642 ;
      RECT 24.054 24.806 24.106 24.842 ;
      RECT 24.054 26.006 24.106 26.042 ;
      RECT 24.054 27.206 24.106 27.242 ;
      RECT 24.054 28.406 24.106 28.442 ;
      RECT 24.054 29.606 24.106 29.642 ;
      RECT 24.054 30.806 24.106 30.842 ;
      RECT 24.054 32.622 24.106 32.658 ;
      RECT 24.054 32.862 24.106 32.898 ;
      RECT 24.054 34.302 24.106 34.338 ;
      RECT 24.054 34.782 24.106 34.818 ;
      RECT 24.054 36.702 24.106 36.738 ;
      RECT 24.054 37.182 24.106 37.218 ;
      RECT 24.054 38.622 24.106 38.658 ;
      RECT 24.054 38.862 24.106 38.898 ;
      RECT 24.054 39.926 24.106 39.962 ;
      RECT 24.054 41.126 24.106 41.162 ;
      RECT 24.054 42.326 24.106 42.362 ;
      RECT 24.054 43.526 24.106 43.562 ;
      RECT 24.054 44.726 24.106 44.762 ;
      RECT 24.054 45.926 24.106 45.962 ;
      RECT 24.054 47.126 24.106 47.162 ;
      RECT 24.054 48.326 24.106 48.362 ;
      RECT 24.054 49.526 24.106 49.562 ;
      RECT 24.054 50.726 24.106 50.762 ;
      RECT 24.054 51.926 24.106 51.962 ;
      RECT 24.054 53.126 24.106 53.162 ;
      RECT 24.054 54.326 24.106 54.362 ;
      RECT 24.054 55.526 24.106 55.562 ;
      RECT 24.054 56.726 24.106 56.762 ;
      RECT 24.054 57.926 24.106 57.962 ;
      RECT 24.054 59.126 24.106 59.162 ;
      RECT 24.054 60.326 24.106 60.362 ;
      RECT 24.054 61.526 24.106 61.562 ;
      RECT 24.054 62.726 24.106 62.762 ;
      RECT 24.054 63.926 24.106 63.962 ;
      RECT 24.054 65.126 24.106 65.162 ;
      RECT 24.054 66.326 24.106 66.362 ;
      RECT 24.054 67.526 24.106 67.562 ;
      RECT 24.054 68.726 24.106 68.762 ;
      RECT 24.054 69.926 24.106 69.962 ;
      RECT 24.054 71.126 24.106 71.162 ;
      RECT 24.134 1.558 24.186 1.594 ;
      RECT 24.134 2.758 24.186 2.794 ;
      RECT 24.134 3.958 24.186 3.994 ;
      RECT 24.134 5.158 24.186 5.194 ;
      RECT 24.134 6.358 24.186 6.394 ;
      RECT 24.134 7.558 24.186 7.594 ;
      RECT 24.134 8.758 24.186 8.794 ;
      RECT 24.134 9.958 24.186 9.994 ;
      RECT 24.134 11.158 24.186 11.194 ;
      RECT 24.134 12.358 24.186 12.394 ;
      RECT 24.134 13.558 24.186 13.594 ;
      RECT 24.134 14.758 24.186 14.794 ;
      RECT 24.134 15.958 24.186 15.994 ;
      RECT 24.134 17.158 24.186 17.194 ;
      RECT 24.134 18.358 24.186 18.394 ;
      RECT 24.134 19.558 24.186 19.594 ;
      RECT 24.134 20.758 24.186 20.794 ;
      RECT 24.134 21.958 24.186 21.994 ;
      RECT 24.134 23.158 24.186 23.194 ;
      RECT 24.134 24.358 24.186 24.394 ;
      RECT 24.134 25.558 24.186 25.594 ;
      RECT 24.134 26.758 24.186 26.794 ;
      RECT 24.134 27.958 24.186 27.994 ;
      RECT 24.134 29.158 24.186 29.194 ;
      RECT 24.134 30.358 24.186 30.394 ;
      RECT 24.134 31.558 24.186 31.594 ;
      RECT 24.134 33.342 24.186 33.378 ;
      RECT 24.134 33.582 24.186 33.618 ;
      RECT 24.134 37.902 24.186 37.938 ;
      RECT 24.134 38.142 24.186 38.178 ;
      RECT 24.134 40.678 24.186 40.714 ;
      RECT 24.134 41.878 24.186 41.914 ;
      RECT 24.134 43.078 24.186 43.114 ;
      RECT 24.134 44.278 24.186 44.314 ;
      RECT 24.134 45.478 24.186 45.514 ;
      RECT 24.134 46.678 24.186 46.714 ;
      RECT 24.134 47.878 24.186 47.914 ;
      RECT 24.134 49.078 24.186 49.114 ;
      RECT 24.134 50.278 24.186 50.314 ;
      RECT 24.134 51.478 24.186 51.514 ;
      RECT 24.134 52.678 24.186 52.714 ;
      RECT 24.134 53.878 24.186 53.914 ;
      RECT 24.134 55.078 24.186 55.114 ;
      RECT 24.134 56.278 24.186 56.314 ;
      RECT 24.134 57.478 24.186 57.514 ;
      RECT 24.134 58.678 24.186 58.714 ;
      RECT 24.134 59.878 24.186 59.914 ;
      RECT 24.134 61.078 24.186 61.114 ;
      RECT 24.134 62.278 24.186 62.314 ;
      RECT 24.134 63.478 24.186 63.514 ;
      RECT 24.134 64.678 24.186 64.714 ;
      RECT 24.134 65.878 24.186 65.914 ;
      RECT 24.134 67.078 24.186 67.114 ;
      RECT 24.134 68.278 24.186 68.314 ;
      RECT 24.134 69.478 24.186 69.514 ;
      RECT 24.134 70.678 24.186 70.714 ;
      RECT 24.134 71.878 24.186 71.914 ;
      RECT 24.214 0.806 24.266 0.842 ;
      RECT 24.214 2.006 24.266 2.042 ;
      RECT 24.214 3.206 24.266 3.242 ;
      RECT 24.214 4.406 24.266 4.442 ;
      RECT 24.214 5.606 24.266 5.642 ;
      RECT 24.214 6.806 24.266 6.842 ;
      RECT 24.214 8.006 24.266 8.042 ;
      RECT 24.214 9.206 24.266 9.242 ;
      RECT 24.214 10.406 24.266 10.442 ;
      RECT 24.214 11.606 24.266 11.642 ;
      RECT 24.214 12.806 24.266 12.842 ;
      RECT 24.214 14.006 24.266 14.042 ;
      RECT 24.214 15.206 24.266 15.242 ;
      RECT 24.214 16.406 24.266 16.442 ;
      RECT 24.214 17.606 24.266 17.642 ;
      RECT 24.214 18.806 24.266 18.842 ;
      RECT 24.214 20.006 24.266 20.042 ;
      RECT 24.214 21.206 24.266 21.242 ;
      RECT 24.214 22.406 24.266 22.442 ;
      RECT 24.214 23.606 24.266 23.642 ;
      RECT 24.214 24.806 24.266 24.842 ;
      RECT 24.214 26.006 24.266 26.042 ;
      RECT 24.214 27.206 24.266 27.242 ;
      RECT 24.214 28.406 24.266 28.442 ;
      RECT 24.214 29.606 24.266 29.642 ;
      RECT 24.214 30.806 24.266 30.842 ;
      RECT 24.214 32.622 24.266 32.658 ;
      RECT 24.214 32.862 24.266 32.898 ;
      RECT 24.214 38.622 24.266 38.658 ;
      RECT 24.214 38.862 24.266 38.898 ;
      RECT 24.214 39.926 24.266 39.962 ;
      RECT 24.214 41.126 24.266 41.162 ;
      RECT 24.214 42.326 24.266 42.362 ;
      RECT 24.214 43.526 24.266 43.562 ;
      RECT 24.214 44.726 24.266 44.762 ;
      RECT 24.214 45.926 24.266 45.962 ;
      RECT 24.214 47.126 24.266 47.162 ;
      RECT 24.214 48.326 24.266 48.362 ;
      RECT 24.214 49.526 24.266 49.562 ;
      RECT 24.214 50.726 24.266 50.762 ;
      RECT 24.214 51.926 24.266 51.962 ;
      RECT 24.214 53.126 24.266 53.162 ;
      RECT 24.214 54.326 24.266 54.362 ;
      RECT 24.214 55.526 24.266 55.562 ;
      RECT 24.214 56.726 24.266 56.762 ;
      RECT 24.214 57.926 24.266 57.962 ;
      RECT 24.214 59.126 24.266 59.162 ;
      RECT 24.214 60.326 24.266 60.362 ;
      RECT 24.214 61.526 24.266 61.562 ;
      RECT 24.214 62.726 24.266 62.762 ;
      RECT 24.214 63.926 24.266 63.962 ;
      RECT 24.214 65.126 24.266 65.162 ;
      RECT 24.214 66.326 24.266 66.362 ;
      RECT 24.214 67.526 24.266 67.562 ;
      RECT 24.214 68.726 24.266 68.762 ;
      RECT 24.214 69.926 24.266 69.962 ;
      RECT 24.214 71.126 24.266 71.162 ;
      RECT 24.294 1.558 24.346 1.594 ;
      RECT 24.294 2.758 24.346 2.794 ;
      RECT 24.294 3.958 24.346 3.994 ;
      RECT 24.294 5.158 24.346 5.194 ;
      RECT 24.294 6.358 24.346 6.394 ;
      RECT 24.294 7.558 24.346 7.594 ;
      RECT 24.294 8.758 24.346 8.794 ;
      RECT 24.294 9.958 24.346 9.994 ;
      RECT 24.294 11.158 24.346 11.194 ;
      RECT 24.294 12.358 24.346 12.394 ;
      RECT 24.294 13.558 24.346 13.594 ;
      RECT 24.294 14.758 24.346 14.794 ;
      RECT 24.294 15.958 24.346 15.994 ;
      RECT 24.294 17.158 24.346 17.194 ;
      RECT 24.294 18.358 24.346 18.394 ;
      RECT 24.294 19.558 24.346 19.594 ;
      RECT 24.294 20.758 24.346 20.794 ;
      RECT 24.294 21.958 24.346 21.994 ;
      RECT 24.294 23.158 24.346 23.194 ;
      RECT 24.294 24.358 24.346 24.394 ;
      RECT 24.294 25.558 24.346 25.594 ;
      RECT 24.294 26.758 24.346 26.794 ;
      RECT 24.294 27.958 24.346 27.994 ;
      RECT 24.294 29.158 24.346 29.194 ;
      RECT 24.294 30.358 24.346 30.394 ;
      RECT 24.294 31.558 24.346 31.594 ;
      RECT 24.294 33.342 24.346 33.378 ;
      RECT 24.294 33.582 24.346 33.618 ;
      RECT 24.294 37.902 24.346 37.938 ;
      RECT 24.294 38.142 24.346 38.178 ;
      RECT 24.294 40.678 24.346 40.714 ;
      RECT 24.294 41.878 24.346 41.914 ;
      RECT 24.294 43.078 24.346 43.114 ;
      RECT 24.294 44.278 24.346 44.314 ;
      RECT 24.294 45.478 24.346 45.514 ;
      RECT 24.294 46.678 24.346 46.714 ;
      RECT 24.294 47.878 24.346 47.914 ;
      RECT 24.294 49.078 24.346 49.114 ;
      RECT 24.294 50.278 24.346 50.314 ;
      RECT 24.294 51.478 24.346 51.514 ;
      RECT 24.294 52.678 24.346 52.714 ;
      RECT 24.294 53.878 24.346 53.914 ;
      RECT 24.294 55.078 24.346 55.114 ;
      RECT 24.294 56.278 24.346 56.314 ;
      RECT 24.294 57.478 24.346 57.514 ;
      RECT 24.294 58.678 24.346 58.714 ;
      RECT 24.294 59.878 24.346 59.914 ;
      RECT 24.294 61.078 24.346 61.114 ;
      RECT 24.294 62.278 24.346 62.314 ;
      RECT 24.294 63.478 24.346 63.514 ;
      RECT 24.294 64.678 24.346 64.714 ;
      RECT 24.294 65.878 24.346 65.914 ;
      RECT 24.294 67.078 24.346 67.114 ;
      RECT 24.294 68.278 24.346 68.314 ;
      RECT 24.294 69.478 24.346 69.514 ;
      RECT 24.294 70.678 24.346 70.714 ;
      RECT 24.294 71.878 24.346 71.914 ;
      RECT 24.374 0.281 24.426 0.317 ;
      RECT 24.374 72.403 24.426 72.439 ;
      RECT 24.454 0.806 24.506 0.842 ;
      RECT 24.454 2.006 24.506 2.042 ;
      RECT 24.454 3.206 24.506 3.242 ;
      RECT 24.454 4.406 24.506 4.442 ;
      RECT 24.454 5.606 24.506 5.642 ;
      RECT 24.454 6.806 24.506 6.842 ;
      RECT 24.454 8.006 24.506 8.042 ;
      RECT 24.454 9.206 24.506 9.242 ;
      RECT 24.454 10.406 24.506 10.442 ;
      RECT 24.454 11.606 24.506 11.642 ;
      RECT 24.454 12.806 24.506 12.842 ;
      RECT 24.454 14.006 24.506 14.042 ;
      RECT 24.454 15.206 24.506 15.242 ;
      RECT 24.454 16.406 24.506 16.442 ;
      RECT 24.454 17.606 24.506 17.642 ;
      RECT 24.454 18.806 24.506 18.842 ;
      RECT 24.454 20.006 24.506 20.042 ;
      RECT 24.454 21.206 24.506 21.242 ;
      RECT 24.454 22.406 24.506 22.442 ;
      RECT 24.454 23.606 24.506 23.642 ;
      RECT 24.454 24.806 24.506 24.842 ;
      RECT 24.454 26.006 24.506 26.042 ;
      RECT 24.454 27.206 24.506 27.242 ;
      RECT 24.454 28.406 24.506 28.442 ;
      RECT 24.454 29.606 24.506 29.642 ;
      RECT 24.454 30.806 24.506 30.842 ;
      RECT 24.454 32.622 24.506 32.658 ;
      RECT 24.454 32.862 24.506 32.898 ;
      RECT 24.454 38.622 24.506 38.658 ;
      RECT 24.454 38.862 24.506 38.898 ;
      RECT 24.454 39.926 24.506 39.962 ;
      RECT 24.454 41.126 24.506 41.162 ;
      RECT 24.454 42.326 24.506 42.362 ;
      RECT 24.454 43.526 24.506 43.562 ;
      RECT 24.454 44.726 24.506 44.762 ;
      RECT 24.454 45.926 24.506 45.962 ;
      RECT 24.454 47.126 24.506 47.162 ;
      RECT 24.454 48.326 24.506 48.362 ;
      RECT 24.454 49.526 24.506 49.562 ;
      RECT 24.454 50.726 24.506 50.762 ;
      RECT 24.454 51.926 24.506 51.962 ;
      RECT 24.454 53.126 24.506 53.162 ;
      RECT 24.454 54.326 24.506 54.362 ;
      RECT 24.454 55.526 24.506 55.562 ;
      RECT 24.454 56.726 24.506 56.762 ;
      RECT 24.454 57.926 24.506 57.962 ;
      RECT 24.454 59.126 24.506 59.162 ;
      RECT 24.454 60.326 24.506 60.362 ;
      RECT 24.454 61.526 24.506 61.562 ;
      RECT 24.454 62.726 24.506 62.762 ;
      RECT 24.454 63.926 24.506 63.962 ;
      RECT 24.454 65.126 24.506 65.162 ;
      RECT 24.454 66.326 24.506 66.362 ;
      RECT 24.454 67.526 24.506 67.562 ;
      RECT 24.454 68.726 24.506 68.762 ;
      RECT 24.454 69.926 24.506 69.962 ;
      RECT 24.454 71.126 24.506 71.162 ;
      RECT 24.534 1.558 24.586 1.594 ;
      RECT 24.534 2.758 24.586 2.794 ;
      RECT 24.534 3.958 24.586 3.994 ;
      RECT 24.534 5.158 24.586 5.194 ;
      RECT 24.534 6.358 24.586 6.394 ;
      RECT 24.534 7.558 24.586 7.594 ;
      RECT 24.534 8.758 24.586 8.794 ;
      RECT 24.534 9.958 24.586 9.994 ;
      RECT 24.534 11.158 24.586 11.194 ;
      RECT 24.534 12.358 24.586 12.394 ;
      RECT 24.534 13.558 24.586 13.594 ;
      RECT 24.534 14.758 24.586 14.794 ;
      RECT 24.534 15.958 24.586 15.994 ;
      RECT 24.534 17.158 24.586 17.194 ;
      RECT 24.534 18.358 24.586 18.394 ;
      RECT 24.534 19.558 24.586 19.594 ;
      RECT 24.534 20.758 24.586 20.794 ;
      RECT 24.534 21.958 24.586 21.994 ;
      RECT 24.534 23.158 24.586 23.194 ;
      RECT 24.534 24.358 24.586 24.394 ;
      RECT 24.534 25.558 24.586 25.594 ;
      RECT 24.534 26.758 24.586 26.794 ;
      RECT 24.534 27.958 24.586 27.994 ;
      RECT 24.534 29.158 24.586 29.194 ;
      RECT 24.534 30.358 24.586 30.394 ;
      RECT 24.534 31.558 24.586 31.594 ;
      RECT 24.534 33.342 24.586 33.378 ;
      RECT 24.534 33.582 24.586 33.618 ;
      RECT 24.534 37.902 24.586 37.938 ;
      RECT 24.534 38.142 24.586 38.178 ;
      RECT 24.534 40.678 24.586 40.714 ;
      RECT 24.534 41.878 24.586 41.914 ;
      RECT 24.534 43.078 24.586 43.114 ;
      RECT 24.534 44.278 24.586 44.314 ;
      RECT 24.534 45.478 24.586 45.514 ;
      RECT 24.534 46.678 24.586 46.714 ;
      RECT 24.534 47.878 24.586 47.914 ;
      RECT 24.534 49.078 24.586 49.114 ;
      RECT 24.534 50.278 24.586 50.314 ;
      RECT 24.534 51.478 24.586 51.514 ;
      RECT 24.534 52.678 24.586 52.714 ;
      RECT 24.534 53.878 24.586 53.914 ;
      RECT 24.534 55.078 24.586 55.114 ;
      RECT 24.534 56.278 24.586 56.314 ;
      RECT 24.534 57.478 24.586 57.514 ;
      RECT 24.534 58.678 24.586 58.714 ;
      RECT 24.534 59.878 24.586 59.914 ;
      RECT 24.534 61.078 24.586 61.114 ;
      RECT 24.534 62.278 24.586 62.314 ;
      RECT 24.534 63.478 24.586 63.514 ;
      RECT 24.534 64.678 24.586 64.714 ;
      RECT 24.534 65.878 24.586 65.914 ;
      RECT 24.534 67.078 24.586 67.114 ;
      RECT 24.534 68.278 24.586 68.314 ;
      RECT 24.534 69.478 24.586 69.514 ;
      RECT 24.534 70.678 24.586 70.714 ;
      RECT 24.534 71.878 24.586 71.914 ;
      RECT 24.614 0.806 24.666 0.842 ;
      RECT 24.614 2.006 24.666 2.042 ;
      RECT 24.614 3.206 24.666 3.242 ;
      RECT 24.614 4.406 24.666 4.442 ;
      RECT 24.614 5.606 24.666 5.642 ;
      RECT 24.614 6.806 24.666 6.842 ;
      RECT 24.614 8.006 24.666 8.042 ;
      RECT 24.614 9.206 24.666 9.242 ;
      RECT 24.614 10.406 24.666 10.442 ;
      RECT 24.614 11.606 24.666 11.642 ;
      RECT 24.614 12.806 24.666 12.842 ;
      RECT 24.614 14.006 24.666 14.042 ;
      RECT 24.614 15.206 24.666 15.242 ;
      RECT 24.614 16.406 24.666 16.442 ;
      RECT 24.614 17.606 24.666 17.642 ;
      RECT 24.614 18.806 24.666 18.842 ;
      RECT 24.614 20.006 24.666 20.042 ;
      RECT 24.614 21.206 24.666 21.242 ;
      RECT 24.614 22.406 24.666 22.442 ;
      RECT 24.614 23.606 24.666 23.642 ;
      RECT 24.614 24.806 24.666 24.842 ;
      RECT 24.614 26.006 24.666 26.042 ;
      RECT 24.614 27.206 24.666 27.242 ;
      RECT 24.614 28.406 24.666 28.442 ;
      RECT 24.614 29.606 24.666 29.642 ;
      RECT 24.614 30.806 24.666 30.842 ;
      RECT 24.614 32.622 24.666 32.658 ;
      RECT 24.614 32.862 24.666 32.898 ;
      RECT 24.614 38.622 24.666 38.658 ;
      RECT 24.614 38.862 24.666 38.898 ;
      RECT 24.614 39.926 24.666 39.962 ;
      RECT 24.614 41.126 24.666 41.162 ;
      RECT 24.614 42.326 24.666 42.362 ;
      RECT 24.614 43.526 24.666 43.562 ;
      RECT 24.614 44.726 24.666 44.762 ;
      RECT 24.614 45.926 24.666 45.962 ;
      RECT 24.614 47.126 24.666 47.162 ;
      RECT 24.614 48.326 24.666 48.362 ;
      RECT 24.614 49.526 24.666 49.562 ;
      RECT 24.614 50.726 24.666 50.762 ;
      RECT 24.614 51.926 24.666 51.962 ;
      RECT 24.614 53.126 24.666 53.162 ;
      RECT 24.614 54.326 24.666 54.362 ;
      RECT 24.614 55.526 24.666 55.562 ;
      RECT 24.614 56.726 24.666 56.762 ;
      RECT 24.614 57.926 24.666 57.962 ;
      RECT 24.614 59.126 24.666 59.162 ;
      RECT 24.614 60.326 24.666 60.362 ;
      RECT 24.614 61.526 24.666 61.562 ;
      RECT 24.614 62.726 24.666 62.762 ;
      RECT 24.614 63.926 24.666 63.962 ;
      RECT 24.614 65.126 24.666 65.162 ;
      RECT 24.614 66.326 24.666 66.362 ;
      RECT 24.614 67.526 24.666 67.562 ;
      RECT 24.614 68.726 24.666 68.762 ;
      RECT 24.614 69.926 24.666 69.962 ;
      RECT 24.614 71.126 24.666 71.162 ;
      RECT 24.694 1.558 24.746 1.594 ;
      RECT 24.694 2.758 24.746 2.794 ;
      RECT 24.694 3.958 24.746 3.994 ;
      RECT 24.694 5.158 24.746 5.194 ;
      RECT 24.694 6.358 24.746 6.394 ;
      RECT 24.694 7.558 24.746 7.594 ;
      RECT 24.694 8.758 24.746 8.794 ;
      RECT 24.694 9.958 24.746 9.994 ;
      RECT 24.694 11.158 24.746 11.194 ;
      RECT 24.694 12.358 24.746 12.394 ;
      RECT 24.694 13.558 24.746 13.594 ;
      RECT 24.694 14.758 24.746 14.794 ;
      RECT 24.694 15.958 24.746 15.994 ;
      RECT 24.694 17.158 24.746 17.194 ;
      RECT 24.694 18.358 24.746 18.394 ;
      RECT 24.694 19.558 24.746 19.594 ;
      RECT 24.694 20.758 24.746 20.794 ;
      RECT 24.694 21.958 24.746 21.994 ;
      RECT 24.694 23.158 24.746 23.194 ;
      RECT 24.694 24.358 24.746 24.394 ;
      RECT 24.694 25.558 24.746 25.594 ;
      RECT 24.694 26.758 24.746 26.794 ;
      RECT 24.694 27.958 24.746 27.994 ;
      RECT 24.694 29.158 24.746 29.194 ;
      RECT 24.694 30.358 24.746 30.394 ;
      RECT 24.694 31.558 24.746 31.594 ;
      RECT 24.694 33.342 24.746 33.378 ;
      RECT 24.694 33.582 24.746 33.618 ;
      RECT 24.694 37.902 24.746 37.938 ;
      RECT 24.694 38.142 24.746 38.178 ;
      RECT 24.694 40.678 24.746 40.714 ;
      RECT 24.694 41.878 24.746 41.914 ;
      RECT 24.694 43.078 24.746 43.114 ;
      RECT 24.694 44.278 24.746 44.314 ;
      RECT 24.694 45.478 24.746 45.514 ;
      RECT 24.694 46.678 24.746 46.714 ;
      RECT 24.694 47.878 24.746 47.914 ;
      RECT 24.694 49.078 24.746 49.114 ;
      RECT 24.694 50.278 24.746 50.314 ;
      RECT 24.694 51.478 24.746 51.514 ;
      RECT 24.694 52.678 24.746 52.714 ;
      RECT 24.694 53.878 24.746 53.914 ;
      RECT 24.694 55.078 24.746 55.114 ;
      RECT 24.694 56.278 24.746 56.314 ;
      RECT 24.694 57.478 24.746 57.514 ;
      RECT 24.694 58.678 24.746 58.714 ;
      RECT 24.694 59.878 24.746 59.914 ;
      RECT 24.694 61.078 24.746 61.114 ;
      RECT 24.694 62.278 24.746 62.314 ;
      RECT 24.694 63.478 24.746 63.514 ;
      RECT 24.694 64.678 24.746 64.714 ;
      RECT 24.694 65.878 24.746 65.914 ;
      RECT 24.694 67.078 24.746 67.114 ;
      RECT 24.694 68.278 24.746 68.314 ;
      RECT 24.694 69.478 24.746 69.514 ;
      RECT 24.694 70.678 24.746 70.714 ;
      RECT 24.694 71.878 24.746 71.914 ;
      RECT 24.774 0.281 24.826 0.317 ;
      RECT 24.774 72.403 24.826 72.439 ;
      RECT 24.854 0.806 24.906 0.842 ;
      RECT 24.854 2.006 24.906 2.042 ;
      RECT 24.854 3.206 24.906 3.242 ;
      RECT 24.854 4.406 24.906 4.442 ;
      RECT 24.854 5.606 24.906 5.642 ;
      RECT 24.854 6.806 24.906 6.842 ;
      RECT 24.854 8.006 24.906 8.042 ;
      RECT 24.854 9.206 24.906 9.242 ;
      RECT 24.854 10.406 24.906 10.442 ;
      RECT 24.854 11.606 24.906 11.642 ;
      RECT 24.854 12.806 24.906 12.842 ;
      RECT 24.854 14.006 24.906 14.042 ;
      RECT 24.854 15.206 24.906 15.242 ;
      RECT 24.854 16.406 24.906 16.442 ;
      RECT 24.854 17.606 24.906 17.642 ;
      RECT 24.854 18.806 24.906 18.842 ;
      RECT 24.854 20.006 24.906 20.042 ;
      RECT 24.854 21.206 24.906 21.242 ;
      RECT 24.854 22.406 24.906 22.442 ;
      RECT 24.854 23.606 24.906 23.642 ;
      RECT 24.854 24.806 24.906 24.842 ;
      RECT 24.854 26.006 24.906 26.042 ;
      RECT 24.854 27.206 24.906 27.242 ;
      RECT 24.854 28.406 24.906 28.442 ;
      RECT 24.854 29.606 24.906 29.642 ;
      RECT 24.854 30.806 24.906 30.842 ;
      RECT 24.854 32.622 24.906 32.658 ;
      RECT 24.854 32.862 24.906 32.898 ;
      RECT 24.854 34.302 24.906 34.338 ;
      RECT 24.854 34.782 24.906 34.818 ;
      RECT 24.854 36.702 24.906 36.738 ;
      RECT 24.854 37.182 24.906 37.218 ;
      RECT 24.854 38.622 24.906 38.658 ;
      RECT 24.854 38.862 24.906 38.898 ;
      RECT 24.854 39.926 24.906 39.962 ;
      RECT 24.854 41.126 24.906 41.162 ;
      RECT 24.854 42.326 24.906 42.362 ;
      RECT 24.854 43.526 24.906 43.562 ;
      RECT 24.854 44.726 24.906 44.762 ;
      RECT 24.854 45.926 24.906 45.962 ;
      RECT 24.854 47.126 24.906 47.162 ;
      RECT 24.854 48.326 24.906 48.362 ;
      RECT 24.854 49.526 24.906 49.562 ;
      RECT 24.854 50.726 24.906 50.762 ;
      RECT 24.854 51.926 24.906 51.962 ;
      RECT 24.854 53.126 24.906 53.162 ;
      RECT 24.854 54.326 24.906 54.362 ;
      RECT 24.854 55.526 24.906 55.562 ;
      RECT 24.854 56.726 24.906 56.762 ;
      RECT 24.854 57.926 24.906 57.962 ;
      RECT 24.854 59.126 24.906 59.162 ;
      RECT 24.854 60.326 24.906 60.362 ;
      RECT 24.854 61.526 24.906 61.562 ;
      RECT 24.854 62.726 24.906 62.762 ;
      RECT 24.854 63.926 24.906 63.962 ;
      RECT 24.854 65.126 24.906 65.162 ;
      RECT 24.854 66.326 24.906 66.362 ;
      RECT 24.854 67.526 24.906 67.562 ;
      RECT 24.854 68.726 24.906 68.762 ;
      RECT 24.854 69.926 24.906 69.962 ;
      RECT 24.854 71.126 24.906 71.162 ;
      RECT 24.934 1.558 24.986 1.594 ;
      RECT 24.934 2.758 24.986 2.794 ;
      RECT 24.934 3.958 24.986 3.994 ;
      RECT 24.934 5.158 24.986 5.194 ;
      RECT 24.934 6.358 24.986 6.394 ;
      RECT 24.934 7.558 24.986 7.594 ;
      RECT 24.934 8.758 24.986 8.794 ;
      RECT 24.934 9.958 24.986 9.994 ;
      RECT 24.934 11.158 24.986 11.194 ;
      RECT 24.934 12.358 24.986 12.394 ;
      RECT 24.934 13.558 24.986 13.594 ;
      RECT 24.934 14.758 24.986 14.794 ;
      RECT 24.934 15.958 24.986 15.994 ;
      RECT 24.934 17.158 24.986 17.194 ;
      RECT 24.934 18.358 24.986 18.394 ;
      RECT 24.934 19.558 24.986 19.594 ;
      RECT 24.934 20.758 24.986 20.794 ;
      RECT 24.934 21.958 24.986 21.994 ;
      RECT 24.934 23.158 24.986 23.194 ;
      RECT 24.934 24.358 24.986 24.394 ;
      RECT 24.934 25.558 24.986 25.594 ;
      RECT 24.934 26.758 24.986 26.794 ;
      RECT 24.934 27.958 24.986 27.994 ;
      RECT 24.934 29.158 24.986 29.194 ;
      RECT 24.934 30.358 24.986 30.394 ;
      RECT 24.934 31.558 24.986 31.594 ;
      RECT 24.934 33.342 24.986 33.378 ;
      RECT 24.934 33.582 24.986 33.618 ;
      RECT 24.934 37.902 24.986 37.938 ;
      RECT 24.934 38.142 24.986 38.178 ;
      RECT 24.934 40.678 24.986 40.714 ;
      RECT 24.934 41.878 24.986 41.914 ;
      RECT 24.934 43.078 24.986 43.114 ;
      RECT 24.934 44.278 24.986 44.314 ;
      RECT 24.934 45.478 24.986 45.514 ;
      RECT 24.934 46.678 24.986 46.714 ;
      RECT 24.934 47.878 24.986 47.914 ;
      RECT 24.934 49.078 24.986 49.114 ;
      RECT 24.934 50.278 24.986 50.314 ;
      RECT 24.934 51.478 24.986 51.514 ;
      RECT 24.934 52.678 24.986 52.714 ;
      RECT 24.934 53.878 24.986 53.914 ;
      RECT 24.934 55.078 24.986 55.114 ;
      RECT 24.934 56.278 24.986 56.314 ;
      RECT 24.934 57.478 24.986 57.514 ;
      RECT 24.934 58.678 24.986 58.714 ;
      RECT 24.934 59.878 24.986 59.914 ;
      RECT 24.934 61.078 24.986 61.114 ;
      RECT 24.934 62.278 24.986 62.314 ;
      RECT 24.934 63.478 24.986 63.514 ;
      RECT 24.934 64.678 24.986 64.714 ;
      RECT 24.934 65.878 24.986 65.914 ;
      RECT 24.934 67.078 24.986 67.114 ;
      RECT 24.934 68.278 24.986 68.314 ;
      RECT 24.934 69.478 24.986 69.514 ;
      RECT 24.934 70.678 24.986 70.714 ;
      RECT 24.934 71.878 24.986 71.914 ;
      RECT 25.014 0.806 25.066 0.842 ;
      RECT 25.014 2.006 25.066 2.042 ;
      RECT 25.014 3.206 25.066 3.242 ;
      RECT 25.014 4.406 25.066 4.442 ;
      RECT 25.014 5.606 25.066 5.642 ;
      RECT 25.014 6.806 25.066 6.842 ;
      RECT 25.014 8.006 25.066 8.042 ;
      RECT 25.014 9.206 25.066 9.242 ;
      RECT 25.014 10.406 25.066 10.442 ;
      RECT 25.014 11.606 25.066 11.642 ;
      RECT 25.014 12.806 25.066 12.842 ;
      RECT 25.014 14.006 25.066 14.042 ;
      RECT 25.014 15.206 25.066 15.242 ;
      RECT 25.014 16.406 25.066 16.442 ;
      RECT 25.014 17.606 25.066 17.642 ;
      RECT 25.014 18.806 25.066 18.842 ;
      RECT 25.014 20.006 25.066 20.042 ;
      RECT 25.014 21.206 25.066 21.242 ;
      RECT 25.014 22.406 25.066 22.442 ;
      RECT 25.014 23.606 25.066 23.642 ;
      RECT 25.014 24.806 25.066 24.842 ;
      RECT 25.014 26.006 25.066 26.042 ;
      RECT 25.014 27.206 25.066 27.242 ;
      RECT 25.014 28.406 25.066 28.442 ;
      RECT 25.014 29.606 25.066 29.642 ;
      RECT 25.014 30.806 25.066 30.842 ;
      RECT 25.014 32.622 25.066 32.658 ;
      RECT 25.014 32.862 25.066 32.898 ;
      RECT 25.014 38.622 25.066 38.658 ;
      RECT 25.014 38.862 25.066 38.898 ;
      RECT 25.014 39.926 25.066 39.962 ;
      RECT 25.014 41.126 25.066 41.162 ;
      RECT 25.014 42.326 25.066 42.362 ;
      RECT 25.014 43.526 25.066 43.562 ;
      RECT 25.014 44.726 25.066 44.762 ;
      RECT 25.014 45.926 25.066 45.962 ;
      RECT 25.014 47.126 25.066 47.162 ;
      RECT 25.014 48.326 25.066 48.362 ;
      RECT 25.014 49.526 25.066 49.562 ;
      RECT 25.014 50.726 25.066 50.762 ;
      RECT 25.014 51.926 25.066 51.962 ;
      RECT 25.014 53.126 25.066 53.162 ;
      RECT 25.014 54.326 25.066 54.362 ;
      RECT 25.014 55.526 25.066 55.562 ;
      RECT 25.014 56.726 25.066 56.762 ;
      RECT 25.014 57.926 25.066 57.962 ;
      RECT 25.014 59.126 25.066 59.162 ;
      RECT 25.014 60.326 25.066 60.362 ;
      RECT 25.014 61.526 25.066 61.562 ;
      RECT 25.014 62.726 25.066 62.762 ;
      RECT 25.014 63.926 25.066 63.962 ;
      RECT 25.014 65.126 25.066 65.162 ;
      RECT 25.014 66.326 25.066 66.362 ;
      RECT 25.014 67.526 25.066 67.562 ;
      RECT 25.014 68.726 25.066 68.762 ;
      RECT 25.014 69.926 25.066 69.962 ;
      RECT 25.014 71.126 25.066 71.162 ;
      RECT 25.094 1.558 25.146 1.594 ;
      RECT 25.094 2.758 25.146 2.794 ;
      RECT 25.094 3.958 25.146 3.994 ;
      RECT 25.094 5.158 25.146 5.194 ;
      RECT 25.094 6.358 25.146 6.394 ;
      RECT 25.094 7.558 25.146 7.594 ;
      RECT 25.094 8.758 25.146 8.794 ;
      RECT 25.094 9.958 25.146 9.994 ;
      RECT 25.094 11.158 25.146 11.194 ;
      RECT 25.094 12.358 25.146 12.394 ;
      RECT 25.094 13.558 25.146 13.594 ;
      RECT 25.094 14.758 25.146 14.794 ;
      RECT 25.094 15.958 25.146 15.994 ;
      RECT 25.094 17.158 25.146 17.194 ;
      RECT 25.094 18.358 25.146 18.394 ;
      RECT 25.094 19.558 25.146 19.594 ;
      RECT 25.094 20.758 25.146 20.794 ;
      RECT 25.094 21.958 25.146 21.994 ;
      RECT 25.094 23.158 25.146 23.194 ;
      RECT 25.094 24.358 25.146 24.394 ;
      RECT 25.094 25.558 25.146 25.594 ;
      RECT 25.094 26.758 25.146 26.794 ;
      RECT 25.094 27.958 25.146 27.994 ;
      RECT 25.094 29.158 25.146 29.194 ;
      RECT 25.094 30.358 25.146 30.394 ;
      RECT 25.094 31.558 25.146 31.594 ;
      RECT 25.094 33.342 25.146 33.378 ;
      RECT 25.094 33.582 25.146 33.618 ;
      RECT 25.094 37.902 25.146 37.938 ;
      RECT 25.094 38.142 25.146 38.178 ;
      RECT 25.094 40.678 25.146 40.714 ;
      RECT 25.094 41.878 25.146 41.914 ;
      RECT 25.094 43.078 25.146 43.114 ;
      RECT 25.094 44.278 25.146 44.314 ;
      RECT 25.094 45.478 25.146 45.514 ;
      RECT 25.094 46.678 25.146 46.714 ;
      RECT 25.094 47.878 25.146 47.914 ;
      RECT 25.094 49.078 25.146 49.114 ;
      RECT 25.094 50.278 25.146 50.314 ;
      RECT 25.094 51.478 25.146 51.514 ;
      RECT 25.094 52.678 25.146 52.714 ;
      RECT 25.094 53.878 25.146 53.914 ;
      RECT 25.094 55.078 25.146 55.114 ;
      RECT 25.094 56.278 25.146 56.314 ;
      RECT 25.094 57.478 25.146 57.514 ;
      RECT 25.094 58.678 25.146 58.714 ;
      RECT 25.094 59.878 25.146 59.914 ;
      RECT 25.094 61.078 25.146 61.114 ;
      RECT 25.094 62.278 25.146 62.314 ;
      RECT 25.094 63.478 25.146 63.514 ;
      RECT 25.094 64.678 25.146 64.714 ;
      RECT 25.094 65.878 25.146 65.914 ;
      RECT 25.094 67.078 25.146 67.114 ;
      RECT 25.094 68.278 25.146 68.314 ;
      RECT 25.094 69.478 25.146 69.514 ;
      RECT 25.094 70.678 25.146 70.714 ;
      RECT 25.094 71.878 25.146 71.914 ;
      RECT 25.174 0.281 25.226 0.317 ;
      RECT 25.174 72.403 25.226 72.439 ;
      RECT 25.254 0.806 25.306 0.842 ;
      RECT 25.254 2.006 25.306 2.042 ;
      RECT 25.254 3.206 25.306 3.242 ;
      RECT 25.254 4.406 25.306 4.442 ;
      RECT 25.254 5.606 25.306 5.642 ;
      RECT 25.254 6.806 25.306 6.842 ;
      RECT 25.254 8.006 25.306 8.042 ;
      RECT 25.254 9.206 25.306 9.242 ;
      RECT 25.254 10.406 25.306 10.442 ;
      RECT 25.254 11.606 25.306 11.642 ;
      RECT 25.254 12.806 25.306 12.842 ;
      RECT 25.254 14.006 25.306 14.042 ;
      RECT 25.254 15.206 25.306 15.242 ;
      RECT 25.254 16.406 25.306 16.442 ;
      RECT 25.254 17.606 25.306 17.642 ;
      RECT 25.254 18.806 25.306 18.842 ;
      RECT 25.254 20.006 25.306 20.042 ;
      RECT 25.254 21.206 25.306 21.242 ;
      RECT 25.254 22.406 25.306 22.442 ;
      RECT 25.254 23.606 25.306 23.642 ;
      RECT 25.254 24.806 25.306 24.842 ;
      RECT 25.254 26.006 25.306 26.042 ;
      RECT 25.254 27.206 25.306 27.242 ;
      RECT 25.254 28.406 25.306 28.442 ;
      RECT 25.254 29.606 25.306 29.642 ;
      RECT 25.254 30.806 25.306 30.842 ;
      RECT 25.254 32.622 25.306 32.658 ;
      RECT 25.254 32.862 25.306 32.898 ;
      RECT 25.254 38.622 25.306 38.658 ;
      RECT 25.254 38.862 25.306 38.898 ;
      RECT 25.254 39.926 25.306 39.962 ;
      RECT 25.254 41.126 25.306 41.162 ;
      RECT 25.254 42.326 25.306 42.362 ;
      RECT 25.254 43.526 25.306 43.562 ;
      RECT 25.254 44.726 25.306 44.762 ;
      RECT 25.254 45.926 25.306 45.962 ;
      RECT 25.254 47.126 25.306 47.162 ;
      RECT 25.254 48.326 25.306 48.362 ;
      RECT 25.254 49.526 25.306 49.562 ;
      RECT 25.254 50.726 25.306 50.762 ;
      RECT 25.254 51.926 25.306 51.962 ;
      RECT 25.254 53.126 25.306 53.162 ;
      RECT 25.254 54.326 25.306 54.362 ;
      RECT 25.254 55.526 25.306 55.562 ;
      RECT 25.254 56.726 25.306 56.762 ;
      RECT 25.254 57.926 25.306 57.962 ;
      RECT 25.254 59.126 25.306 59.162 ;
      RECT 25.254 60.326 25.306 60.362 ;
      RECT 25.254 61.526 25.306 61.562 ;
      RECT 25.254 62.726 25.306 62.762 ;
      RECT 25.254 63.926 25.306 63.962 ;
      RECT 25.254 65.126 25.306 65.162 ;
      RECT 25.254 66.326 25.306 66.362 ;
      RECT 25.254 67.526 25.306 67.562 ;
      RECT 25.254 68.726 25.306 68.762 ;
      RECT 25.254 69.926 25.306 69.962 ;
      RECT 25.254 71.126 25.306 71.162 ;
      RECT 25.334 1.558 25.386 1.594 ;
      RECT 25.334 2.758 25.386 2.794 ;
      RECT 25.334 3.958 25.386 3.994 ;
      RECT 25.334 5.158 25.386 5.194 ;
      RECT 25.334 6.358 25.386 6.394 ;
      RECT 25.334 7.558 25.386 7.594 ;
      RECT 25.334 8.758 25.386 8.794 ;
      RECT 25.334 9.958 25.386 9.994 ;
      RECT 25.334 11.158 25.386 11.194 ;
      RECT 25.334 12.358 25.386 12.394 ;
      RECT 25.334 13.558 25.386 13.594 ;
      RECT 25.334 14.758 25.386 14.794 ;
      RECT 25.334 15.958 25.386 15.994 ;
      RECT 25.334 17.158 25.386 17.194 ;
      RECT 25.334 18.358 25.386 18.394 ;
      RECT 25.334 19.558 25.386 19.594 ;
      RECT 25.334 20.758 25.386 20.794 ;
      RECT 25.334 21.958 25.386 21.994 ;
      RECT 25.334 23.158 25.386 23.194 ;
      RECT 25.334 24.358 25.386 24.394 ;
      RECT 25.334 25.558 25.386 25.594 ;
      RECT 25.334 26.758 25.386 26.794 ;
      RECT 25.334 27.958 25.386 27.994 ;
      RECT 25.334 29.158 25.386 29.194 ;
      RECT 25.334 30.358 25.386 30.394 ;
      RECT 25.334 31.558 25.386 31.594 ;
      RECT 25.334 33.342 25.386 33.378 ;
      RECT 25.334 33.582 25.386 33.618 ;
      RECT 25.334 37.902 25.386 37.938 ;
      RECT 25.334 38.142 25.386 38.178 ;
      RECT 25.334 40.678 25.386 40.714 ;
      RECT 25.334 41.878 25.386 41.914 ;
      RECT 25.334 43.078 25.386 43.114 ;
      RECT 25.334 44.278 25.386 44.314 ;
      RECT 25.334 45.478 25.386 45.514 ;
      RECT 25.334 46.678 25.386 46.714 ;
      RECT 25.334 47.878 25.386 47.914 ;
      RECT 25.334 49.078 25.386 49.114 ;
      RECT 25.334 50.278 25.386 50.314 ;
      RECT 25.334 51.478 25.386 51.514 ;
      RECT 25.334 52.678 25.386 52.714 ;
      RECT 25.334 53.878 25.386 53.914 ;
      RECT 25.334 55.078 25.386 55.114 ;
      RECT 25.334 56.278 25.386 56.314 ;
      RECT 25.334 57.478 25.386 57.514 ;
      RECT 25.334 58.678 25.386 58.714 ;
      RECT 25.334 59.878 25.386 59.914 ;
      RECT 25.334 61.078 25.386 61.114 ;
      RECT 25.334 62.278 25.386 62.314 ;
      RECT 25.334 63.478 25.386 63.514 ;
      RECT 25.334 64.678 25.386 64.714 ;
      RECT 25.334 65.878 25.386 65.914 ;
      RECT 25.334 67.078 25.386 67.114 ;
      RECT 25.334 68.278 25.386 68.314 ;
      RECT 25.334 69.478 25.386 69.514 ;
      RECT 25.334 70.678 25.386 70.714 ;
      RECT 25.334 71.878 25.386 71.914 ;
      RECT 25.414 0.806 25.466 0.842 ;
      RECT 25.414 2.006 25.466 2.042 ;
      RECT 25.414 3.206 25.466 3.242 ;
      RECT 25.414 4.406 25.466 4.442 ;
      RECT 25.414 5.606 25.466 5.642 ;
      RECT 25.414 6.806 25.466 6.842 ;
      RECT 25.414 8.006 25.466 8.042 ;
      RECT 25.414 9.206 25.466 9.242 ;
      RECT 25.414 10.406 25.466 10.442 ;
      RECT 25.414 11.606 25.466 11.642 ;
      RECT 25.414 12.806 25.466 12.842 ;
      RECT 25.414 14.006 25.466 14.042 ;
      RECT 25.414 15.206 25.466 15.242 ;
      RECT 25.414 16.406 25.466 16.442 ;
      RECT 25.414 17.606 25.466 17.642 ;
      RECT 25.414 18.806 25.466 18.842 ;
      RECT 25.414 20.006 25.466 20.042 ;
      RECT 25.414 21.206 25.466 21.242 ;
      RECT 25.414 22.406 25.466 22.442 ;
      RECT 25.414 23.606 25.466 23.642 ;
      RECT 25.414 24.806 25.466 24.842 ;
      RECT 25.414 26.006 25.466 26.042 ;
      RECT 25.414 27.206 25.466 27.242 ;
      RECT 25.414 28.406 25.466 28.442 ;
      RECT 25.414 29.606 25.466 29.642 ;
      RECT 25.414 30.806 25.466 30.842 ;
      RECT 25.414 32.622 25.466 32.658 ;
      RECT 25.414 32.862 25.466 32.898 ;
      RECT 25.414 38.622 25.466 38.658 ;
      RECT 25.414 38.862 25.466 38.898 ;
      RECT 25.414 39.926 25.466 39.962 ;
      RECT 25.414 41.126 25.466 41.162 ;
      RECT 25.414 42.326 25.466 42.362 ;
      RECT 25.414 43.526 25.466 43.562 ;
      RECT 25.414 44.726 25.466 44.762 ;
      RECT 25.414 45.926 25.466 45.962 ;
      RECT 25.414 47.126 25.466 47.162 ;
      RECT 25.414 48.326 25.466 48.362 ;
      RECT 25.414 49.526 25.466 49.562 ;
      RECT 25.414 50.726 25.466 50.762 ;
      RECT 25.414 51.926 25.466 51.962 ;
      RECT 25.414 53.126 25.466 53.162 ;
      RECT 25.414 54.326 25.466 54.362 ;
      RECT 25.414 55.526 25.466 55.562 ;
      RECT 25.414 56.726 25.466 56.762 ;
      RECT 25.414 57.926 25.466 57.962 ;
      RECT 25.414 59.126 25.466 59.162 ;
      RECT 25.414 60.326 25.466 60.362 ;
      RECT 25.414 61.526 25.466 61.562 ;
      RECT 25.414 62.726 25.466 62.762 ;
      RECT 25.414 63.926 25.466 63.962 ;
      RECT 25.414 65.126 25.466 65.162 ;
      RECT 25.414 66.326 25.466 66.362 ;
      RECT 25.414 67.526 25.466 67.562 ;
      RECT 25.414 68.726 25.466 68.762 ;
      RECT 25.414 69.926 25.466 69.962 ;
      RECT 25.414 71.126 25.466 71.162 ;
      RECT 25.494 1.558 25.546 1.594 ;
      RECT 25.494 2.758 25.546 2.794 ;
      RECT 25.494 3.958 25.546 3.994 ;
      RECT 25.494 5.158 25.546 5.194 ;
      RECT 25.494 6.358 25.546 6.394 ;
      RECT 25.494 7.558 25.546 7.594 ;
      RECT 25.494 8.758 25.546 8.794 ;
      RECT 25.494 9.958 25.546 9.994 ;
      RECT 25.494 11.158 25.546 11.194 ;
      RECT 25.494 12.358 25.546 12.394 ;
      RECT 25.494 13.558 25.546 13.594 ;
      RECT 25.494 14.758 25.546 14.794 ;
      RECT 25.494 15.958 25.546 15.994 ;
      RECT 25.494 17.158 25.546 17.194 ;
      RECT 25.494 18.358 25.546 18.394 ;
      RECT 25.494 19.558 25.546 19.594 ;
      RECT 25.494 20.758 25.546 20.794 ;
      RECT 25.494 21.958 25.546 21.994 ;
      RECT 25.494 23.158 25.546 23.194 ;
      RECT 25.494 24.358 25.546 24.394 ;
      RECT 25.494 25.558 25.546 25.594 ;
      RECT 25.494 26.758 25.546 26.794 ;
      RECT 25.494 27.958 25.546 27.994 ;
      RECT 25.494 29.158 25.546 29.194 ;
      RECT 25.494 30.358 25.546 30.394 ;
      RECT 25.494 31.558 25.546 31.594 ;
      RECT 25.494 33.342 25.546 33.378 ;
      RECT 25.494 33.582 25.546 33.618 ;
      RECT 25.494 37.902 25.546 37.938 ;
      RECT 25.494 38.142 25.546 38.178 ;
      RECT 25.494 40.678 25.546 40.714 ;
      RECT 25.494 41.878 25.546 41.914 ;
      RECT 25.494 43.078 25.546 43.114 ;
      RECT 25.494 44.278 25.546 44.314 ;
      RECT 25.494 45.478 25.546 45.514 ;
      RECT 25.494 46.678 25.546 46.714 ;
      RECT 25.494 47.878 25.546 47.914 ;
      RECT 25.494 49.078 25.546 49.114 ;
      RECT 25.494 50.278 25.546 50.314 ;
      RECT 25.494 51.478 25.546 51.514 ;
      RECT 25.494 52.678 25.546 52.714 ;
      RECT 25.494 53.878 25.546 53.914 ;
      RECT 25.494 55.078 25.546 55.114 ;
      RECT 25.494 56.278 25.546 56.314 ;
      RECT 25.494 57.478 25.546 57.514 ;
      RECT 25.494 58.678 25.546 58.714 ;
      RECT 25.494 59.878 25.546 59.914 ;
      RECT 25.494 61.078 25.546 61.114 ;
      RECT 25.494 62.278 25.546 62.314 ;
      RECT 25.494 63.478 25.546 63.514 ;
      RECT 25.494 64.678 25.546 64.714 ;
      RECT 25.494 65.878 25.546 65.914 ;
      RECT 25.494 67.078 25.546 67.114 ;
      RECT 25.494 68.278 25.546 68.314 ;
      RECT 25.494 69.478 25.546 69.514 ;
      RECT 25.494 70.678 25.546 70.714 ;
      RECT 25.494 71.878 25.546 71.914 ;
      RECT 25.574 0.281 25.626 0.317 ;
      RECT 25.574 72.403 25.626 72.439 ;
      RECT 25.654 0.806 25.706 0.842 ;
      RECT 25.654 2.006 25.706 2.042 ;
      RECT 25.654 3.206 25.706 3.242 ;
      RECT 25.654 4.406 25.706 4.442 ;
      RECT 25.654 5.606 25.706 5.642 ;
      RECT 25.654 6.806 25.706 6.842 ;
      RECT 25.654 8.006 25.706 8.042 ;
      RECT 25.654 9.206 25.706 9.242 ;
      RECT 25.654 10.406 25.706 10.442 ;
      RECT 25.654 11.606 25.706 11.642 ;
      RECT 25.654 12.806 25.706 12.842 ;
      RECT 25.654 14.006 25.706 14.042 ;
      RECT 25.654 15.206 25.706 15.242 ;
      RECT 25.654 16.406 25.706 16.442 ;
      RECT 25.654 17.606 25.706 17.642 ;
      RECT 25.654 18.806 25.706 18.842 ;
      RECT 25.654 20.006 25.706 20.042 ;
      RECT 25.654 21.206 25.706 21.242 ;
      RECT 25.654 22.406 25.706 22.442 ;
      RECT 25.654 23.606 25.706 23.642 ;
      RECT 25.654 24.806 25.706 24.842 ;
      RECT 25.654 26.006 25.706 26.042 ;
      RECT 25.654 27.206 25.706 27.242 ;
      RECT 25.654 28.406 25.706 28.442 ;
      RECT 25.654 29.606 25.706 29.642 ;
      RECT 25.654 30.806 25.706 30.842 ;
      RECT 25.654 32.622 25.706 32.658 ;
      RECT 25.654 32.862 25.706 32.898 ;
      RECT 25.654 34.302 25.706 34.338 ;
      RECT 25.654 34.782 25.706 34.818 ;
      RECT 25.654 36.702 25.706 36.738 ;
      RECT 25.654 37.182 25.706 37.218 ;
      RECT 25.654 38.622 25.706 38.658 ;
      RECT 25.654 38.862 25.706 38.898 ;
      RECT 25.654 39.926 25.706 39.962 ;
      RECT 25.654 41.126 25.706 41.162 ;
      RECT 25.654 42.326 25.706 42.362 ;
      RECT 25.654 43.526 25.706 43.562 ;
      RECT 25.654 44.726 25.706 44.762 ;
      RECT 25.654 45.926 25.706 45.962 ;
      RECT 25.654 47.126 25.706 47.162 ;
      RECT 25.654 48.326 25.706 48.362 ;
      RECT 25.654 49.526 25.706 49.562 ;
      RECT 25.654 50.726 25.706 50.762 ;
      RECT 25.654 51.926 25.706 51.962 ;
      RECT 25.654 53.126 25.706 53.162 ;
      RECT 25.654 54.326 25.706 54.362 ;
      RECT 25.654 55.526 25.706 55.562 ;
      RECT 25.654 56.726 25.706 56.762 ;
      RECT 25.654 57.926 25.706 57.962 ;
      RECT 25.654 59.126 25.706 59.162 ;
      RECT 25.654 60.326 25.706 60.362 ;
      RECT 25.654 61.526 25.706 61.562 ;
      RECT 25.654 62.726 25.706 62.762 ;
      RECT 25.654 63.926 25.706 63.962 ;
      RECT 25.654 65.126 25.706 65.162 ;
      RECT 25.654 66.326 25.706 66.362 ;
      RECT 25.654 67.526 25.706 67.562 ;
      RECT 25.654 68.726 25.706 68.762 ;
      RECT 25.654 69.926 25.706 69.962 ;
      RECT 25.654 71.126 25.706 71.162 ;
      RECT 25.734 1.558 25.786 1.594 ;
      RECT 25.734 2.758 25.786 2.794 ;
      RECT 25.734 3.958 25.786 3.994 ;
      RECT 25.734 5.158 25.786 5.194 ;
      RECT 25.734 6.358 25.786 6.394 ;
      RECT 25.734 7.558 25.786 7.594 ;
      RECT 25.734 8.758 25.786 8.794 ;
      RECT 25.734 9.958 25.786 9.994 ;
      RECT 25.734 11.158 25.786 11.194 ;
      RECT 25.734 12.358 25.786 12.394 ;
      RECT 25.734 13.558 25.786 13.594 ;
      RECT 25.734 14.758 25.786 14.794 ;
      RECT 25.734 15.958 25.786 15.994 ;
      RECT 25.734 17.158 25.786 17.194 ;
      RECT 25.734 18.358 25.786 18.394 ;
      RECT 25.734 19.558 25.786 19.594 ;
      RECT 25.734 20.758 25.786 20.794 ;
      RECT 25.734 21.958 25.786 21.994 ;
      RECT 25.734 23.158 25.786 23.194 ;
      RECT 25.734 24.358 25.786 24.394 ;
      RECT 25.734 25.558 25.786 25.594 ;
      RECT 25.734 26.758 25.786 26.794 ;
      RECT 25.734 27.958 25.786 27.994 ;
      RECT 25.734 29.158 25.786 29.194 ;
      RECT 25.734 30.358 25.786 30.394 ;
      RECT 25.734 31.558 25.786 31.594 ;
      RECT 25.734 33.342 25.786 33.378 ;
      RECT 25.734 33.582 25.786 33.618 ;
      RECT 25.734 37.902 25.786 37.938 ;
      RECT 25.734 38.142 25.786 38.178 ;
      RECT 25.734 40.678 25.786 40.714 ;
      RECT 25.734 41.878 25.786 41.914 ;
      RECT 25.734 43.078 25.786 43.114 ;
      RECT 25.734 44.278 25.786 44.314 ;
      RECT 25.734 45.478 25.786 45.514 ;
      RECT 25.734 46.678 25.786 46.714 ;
      RECT 25.734 47.878 25.786 47.914 ;
      RECT 25.734 49.078 25.786 49.114 ;
      RECT 25.734 50.278 25.786 50.314 ;
      RECT 25.734 51.478 25.786 51.514 ;
      RECT 25.734 52.678 25.786 52.714 ;
      RECT 25.734 53.878 25.786 53.914 ;
      RECT 25.734 55.078 25.786 55.114 ;
      RECT 25.734 56.278 25.786 56.314 ;
      RECT 25.734 57.478 25.786 57.514 ;
      RECT 25.734 58.678 25.786 58.714 ;
      RECT 25.734 59.878 25.786 59.914 ;
      RECT 25.734 61.078 25.786 61.114 ;
      RECT 25.734 62.278 25.786 62.314 ;
      RECT 25.734 63.478 25.786 63.514 ;
      RECT 25.734 64.678 25.786 64.714 ;
      RECT 25.734 65.878 25.786 65.914 ;
      RECT 25.734 67.078 25.786 67.114 ;
      RECT 25.734 68.278 25.786 68.314 ;
      RECT 25.734 69.478 25.786 69.514 ;
      RECT 25.734 70.678 25.786 70.714 ;
      RECT 25.734 71.878 25.786 71.914 ;
      RECT 25.814 0.806 25.866 0.842 ;
      RECT 25.814 2.006 25.866 2.042 ;
      RECT 25.814 3.206 25.866 3.242 ;
      RECT 25.814 4.406 25.866 4.442 ;
      RECT 25.814 5.606 25.866 5.642 ;
      RECT 25.814 6.806 25.866 6.842 ;
      RECT 25.814 8.006 25.866 8.042 ;
      RECT 25.814 9.206 25.866 9.242 ;
      RECT 25.814 10.406 25.866 10.442 ;
      RECT 25.814 11.606 25.866 11.642 ;
      RECT 25.814 12.806 25.866 12.842 ;
      RECT 25.814 14.006 25.866 14.042 ;
      RECT 25.814 15.206 25.866 15.242 ;
      RECT 25.814 16.406 25.866 16.442 ;
      RECT 25.814 17.606 25.866 17.642 ;
      RECT 25.814 18.806 25.866 18.842 ;
      RECT 25.814 20.006 25.866 20.042 ;
      RECT 25.814 21.206 25.866 21.242 ;
      RECT 25.814 22.406 25.866 22.442 ;
      RECT 25.814 23.606 25.866 23.642 ;
      RECT 25.814 24.806 25.866 24.842 ;
      RECT 25.814 26.006 25.866 26.042 ;
      RECT 25.814 27.206 25.866 27.242 ;
      RECT 25.814 28.406 25.866 28.442 ;
      RECT 25.814 29.606 25.866 29.642 ;
      RECT 25.814 30.806 25.866 30.842 ;
      RECT 25.814 32.622 25.866 32.658 ;
      RECT 25.814 32.862 25.866 32.898 ;
      RECT 25.814 38.622 25.866 38.658 ;
      RECT 25.814 38.862 25.866 38.898 ;
      RECT 25.814 39.926 25.866 39.962 ;
      RECT 25.814 41.126 25.866 41.162 ;
      RECT 25.814 42.326 25.866 42.362 ;
      RECT 25.814 43.526 25.866 43.562 ;
      RECT 25.814 44.726 25.866 44.762 ;
      RECT 25.814 45.926 25.866 45.962 ;
      RECT 25.814 47.126 25.866 47.162 ;
      RECT 25.814 48.326 25.866 48.362 ;
      RECT 25.814 49.526 25.866 49.562 ;
      RECT 25.814 50.726 25.866 50.762 ;
      RECT 25.814 51.926 25.866 51.962 ;
      RECT 25.814 53.126 25.866 53.162 ;
      RECT 25.814 54.326 25.866 54.362 ;
      RECT 25.814 55.526 25.866 55.562 ;
      RECT 25.814 56.726 25.866 56.762 ;
      RECT 25.814 57.926 25.866 57.962 ;
      RECT 25.814 59.126 25.866 59.162 ;
      RECT 25.814 60.326 25.866 60.362 ;
      RECT 25.814 61.526 25.866 61.562 ;
      RECT 25.814 62.726 25.866 62.762 ;
      RECT 25.814 63.926 25.866 63.962 ;
      RECT 25.814 65.126 25.866 65.162 ;
      RECT 25.814 66.326 25.866 66.362 ;
      RECT 25.814 67.526 25.866 67.562 ;
      RECT 25.814 68.726 25.866 68.762 ;
      RECT 25.814 69.926 25.866 69.962 ;
      RECT 25.814 71.126 25.866 71.162 ;
      RECT 25.894 1.558 25.946 1.594 ;
      RECT 25.894 2.758 25.946 2.794 ;
      RECT 25.894 3.958 25.946 3.994 ;
      RECT 25.894 5.158 25.946 5.194 ;
      RECT 25.894 6.358 25.946 6.394 ;
      RECT 25.894 7.558 25.946 7.594 ;
      RECT 25.894 8.758 25.946 8.794 ;
      RECT 25.894 9.958 25.946 9.994 ;
      RECT 25.894 11.158 25.946 11.194 ;
      RECT 25.894 12.358 25.946 12.394 ;
      RECT 25.894 13.558 25.946 13.594 ;
      RECT 25.894 14.758 25.946 14.794 ;
      RECT 25.894 15.958 25.946 15.994 ;
      RECT 25.894 17.158 25.946 17.194 ;
      RECT 25.894 18.358 25.946 18.394 ;
      RECT 25.894 19.558 25.946 19.594 ;
      RECT 25.894 20.758 25.946 20.794 ;
      RECT 25.894 21.958 25.946 21.994 ;
      RECT 25.894 23.158 25.946 23.194 ;
      RECT 25.894 24.358 25.946 24.394 ;
      RECT 25.894 25.558 25.946 25.594 ;
      RECT 25.894 26.758 25.946 26.794 ;
      RECT 25.894 27.958 25.946 27.994 ;
      RECT 25.894 29.158 25.946 29.194 ;
      RECT 25.894 30.358 25.946 30.394 ;
      RECT 25.894 31.558 25.946 31.594 ;
      RECT 25.894 33.342 25.946 33.378 ;
      RECT 25.894 33.582 25.946 33.618 ;
      RECT 25.894 37.902 25.946 37.938 ;
      RECT 25.894 38.142 25.946 38.178 ;
      RECT 25.894 40.678 25.946 40.714 ;
      RECT 25.894 41.878 25.946 41.914 ;
      RECT 25.894 43.078 25.946 43.114 ;
      RECT 25.894 44.278 25.946 44.314 ;
      RECT 25.894 45.478 25.946 45.514 ;
      RECT 25.894 46.678 25.946 46.714 ;
      RECT 25.894 47.878 25.946 47.914 ;
      RECT 25.894 49.078 25.946 49.114 ;
      RECT 25.894 50.278 25.946 50.314 ;
      RECT 25.894 51.478 25.946 51.514 ;
      RECT 25.894 52.678 25.946 52.714 ;
      RECT 25.894 53.878 25.946 53.914 ;
      RECT 25.894 55.078 25.946 55.114 ;
      RECT 25.894 56.278 25.946 56.314 ;
      RECT 25.894 57.478 25.946 57.514 ;
      RECT 25.894 58.678 25.946 58.714 ;
      RECT 25.894 59.878 25.946 59.914 ;
      RECT 25.894 61.078 25.946 61.114 ;
      RECT 25.894 62.278 25.946 62.314 ;
      RECT 25.894 63.478 25.946 63.514 ;
      RECT 25.894 64.678 25.946 64.714 ;
      RECT 25.894 65.878 25.946 65.914 ;
      RECT 25.894 67.078 25.946 67.114 ;
      RECT 25.894 68.278 25.946 68.314 ;
      RECT 25.894 69.478 25.946 69.514 ;
      RECT 25.894 70.678 25.946 70.714 ;
      RECT 25.894 71.878 25.946 71.914 ;
      RECT 25.974 0.281 26.026 0.317 ;
      RECT 25.974 72.403 26.026 72.439 ;
      RECT 26.054 0.806 26.106 0.842 ;
      RECT 26.054 2.006 26.106 2.042 ;
      RECT 26.054 3.206 26.106 3.242 ;
      RECT 26.054 4.406 26.106 4.442 ;
      RECT 26.054 5.606 26.106 5.642 ;
      RECT 26.054 6.806 26.106 6.842 ;
      RECT 26.054 8.006 26.106 8.042 ;
      RECT 26.054 9.206 26.106 9.242 ;
      RECT 26.054 10.406 26.106 10.442 ;
      RECT 26.054 11.606 26.106 11.642 ;
      RECT 26.054 12.806 26.106 12.842 ;
      RECT 26.054 14.006 26.106 14.042 ;
      RECT 26.054 15.206 26.106 15.242 ;
      RECT 26.054 16.406 26.106 16.442 ;
      RECT 26.054 17.606 26.106 17.642 ;
      RECT 26.054 18.806 26.106 18.842 ;
      RECT 26.054 20.006 26.106 20.042 ;
      RECT 26.054 21.206 26.106 21.242 ;
      RECT 26.054 22.406 26.106 22.442 ;
      RECT 26.054 23.606 26.106 23.642 ;
      RECT 26.054 24.806 26.106 24.842 ;
      RECT 26.054 26.006 26.106 26.042 ;
      RECT 26.054 27.206 26.106 27.242 ;
      RECT 26.054 28.406 26.106 28.442 ;
      RECT 26.054 29.606 26.106 29.642 ;
      RECT 26.054 30.806 26.106 30.842 ;
      RECT 26.054 32.622 26.106 32.658 ;
      RECT 26.054 32.862 26.106 32.898 ;
      RECT 26.054 38.622 26.106 38.658 ;
      RECT 26.054 38.862 26.106 38.898 ;
      RECT 26.054 39.926 26.106 39.962 ;
      RECT 26.054 41.126 26.106 41.162 ;
      RECT 26.054 42.326 26.106 42.362 ;
      RECT 26.054 43.526 26.106 43.562 ;
      RECT 26.054 44.726 26.106 44.762 ;
      RECT 26.054 45.926 26.106 45.962 ;
      RECT 26.054 47.126 26.106 47.162 ;
      RECT 26.054 48.326 26.106 48.362 ;
      RECT 26.054 49.526 26.106 49.562 ;
      RECT 26.054 50.726 26.106 50.762 ;
      RECT 26.054 51.926 26.106 51.962 ;
      RECT 26.054 53.126 26.106 53.162 ;
      RECT 26.054 54.326 26.106 54.362 ;
      RECT 26.054 55.526 26.106 55.562 ;
      RECT 26.054 56.726 26.106 56.762 ;
      RECT 26.054 57.926 26.106 57.962 ;
      RECT 26.054 59.126 26.106 59.162 ;
      RECT 26.054 60.326 26.106 60.362 ;
      RECT 26.054 61.526 26.106 61.562 ;
      RECT 26.054 62.726 26.106 62.762 ;
      RECT 26.054 63.926 26.106 63.962 ;
      RECT 26.054 65.126 26.106 65.162 ;
      RECT 26.054 66.326 26.106 66.362 ;
      RECT 26.054 67.526 26.106 67.562 ;
      RECT 26.054 68.726 26.106 68.762 ;
      RECT 26.054 69.926 26.106 69.962 ;
      RECT 26.054 71.126 26.106 71.162 ;
      RECT 26.134 1.558 26.186 1.594 ;
      RECT 26.134 2.758 26.186 2.794 ;
      RECT 26.134 3.958 26.186 3.994 ;
      RECT 26.134 5.158 26.186 5.194 ;
      RECT 26.134 6.358 26.186 6.394 ;
      RECT 26.134 7.558 26.186 7.594 ;
      RECT 26.134 8.758 26.186 8.794 ;
      RECT 26.134 9.958 26.186 9.994 ;
      RECT 26.134 11.158 26.186 11.194 ;
      RECT 26.134 12.358 26.186 12.394 ;
      RECT 26.134 13.558 26.186 13.594 ;
      RECT 26.134 14.758 26.186 14.794 ;
      RECT 26.134 15.958 26.186 15.994 ;
      RECT 26.134 17.158 26.186 17.194 ;
      RECT 26.134 18.358 26.186 18.394 ;
      RECT 26.134 19.558 26.186 19.594 ;
      RECT 26.134 20.758 26.186 20.794 ;
      RECT 26.134 21.958 26.186 21.994 ;
      RECT 26.134 23.158 26.186 23.194 ;
      RECT 26.134 24.358 26.186 24.394 ;
      RECT 26.134 25.558 26.186 25.594 ;
      RECT 26.134 26.758 26.186 26.794 ;
      RECT 26.134 27.958 26.186 27.994 ;
      RECT 26.134 29.158 26.186 29.194 ;
      RECT 26.134 30.358 26.186 30.394 ;
      RECT 26.134 31.558 26.186 31.594 ;
      RECT 26.134 33.342 26.186 33.378 ;
      RECT 26.134 33.582 26.186 33.618 ;
      RECT 26.134 37.902 26.186 37.938 ;
      RECT 26.134 38.142 26.186 38.178 ;
      RECT 26.134 40.678 26.186 40.714 ;
      RECT 26.134 41.878 26.186 41.914 ;
      RECT 26.134 43.078 26.186 43.114 ;
      RECT 26.134 44.278 26.186 44.314 ;
      RECT 26.134 45.478 26.186 45.514 ;
      RECT 26.134 46.678 26.186 46.714 ;
      RECT 26.134 47.878 26.186 47.914 ;
      RECT 26.134 49.078 26.186 49.114 ;
      RECT 26.134 50.278 26.186 50.314 ;
      RECT 26.134 51.478 26.186 51.514 ;
      RECT 26.134 52.678 26.186 52.714 ;
      RECT 26.134 53.878 26.186 53.914 ;
      RECT 26.134 55.078 26.186 55.114 ;
      RECT 26.134 56.278 26.186 56.314 ;
      RECT 26.134 57.478 26.186 57.514 ;
      RECT 26.134 58.678 26.186 58.714 ;
      RECT 26.134 59.878 26.186 59.914 ;
      RECT 26.134 61.078 26.186 61.114 ;
      RECT 26.134 62.278 26.186 62.314 ;
      RECT 26.134 63.478 26.186 63.514 ;
      RECT 26.134 64.678 26.186 64.714 ;
      RECT 26.134 65.878 26.186 65.914 ;
      RECT 26.134 67.078 26.186 67.114 ;
      RECT 26.134 68.278 26.186 68.314 ;
      RECT 26.134 69.478 26.186 69.514 ;
      RECT 26.134 70.678 26.186 70.714 ;
      RECT 26.134 71.878 26.186 71.914 ;
      RECT 26.214 0.806 26.266 0.842 ;
      RECT 26.214 2.006 26.266 2.042 ;
      RECT 26.214 3.206 26.266 3.242 ;
      RECT 26.214 4.406 26.266 4.442 ;
      RECT 26.214 5.606 26.266 5.642 ;
      RECT 26.214 6.806 26.266 6.842 ;
      RECT 26.214 8.006 26.266 8.042 ;
      RECT 26.214 9.206 26.266 9.242 ;
      RECT 26.214 10.406 26.266 10.442 ;
      RECT 26.214 11.606 26.266 11.642 ;
      RECT 26.214 12.806 26.266 12.842 ;
      RECT 26.214 14.006 26.266 14.042 ;
      RECT 26.214 15.206 26.266 15.242 ;
      RECT 26.214 16.406 26.266 16.442 ;
      RECT 26.214 17.606 26.266 17.642 ;
      RECT 26.214 18.806 26.266 18.842 ;
      RECT 26.214 20.006 26.266 20.042 ;
      RECT 26.214 21.206 26.266 21.242 ;
      RECT 26.214 22.406 26.266 22.442 ;
      RECT 26.214 23.606 26.266 23.642 ;
      RECT 26.214 24.806 26.266 24.842 ;
      RECT 26.214 26.006 26.266 26.042 ;
      RECT 26.214 27.206 26.266 27.242 ;
      RECT 26.214 28.406 26.266 28.442 ;
      RECT 26.214 29.606 26.266 29.642 ;
      RECT 26.214 30.806 26.266 30.842 ;
      RECT 26.214 32.622 26.266 32.658 ;
      RECT 26.214 32.862 26.266 32.898 ;
      RECT 26.214 38.622 26.266 38.658 ;
      RECT 26.214 38.862 26.266 38.898 ;
      RECT 26.214 39.926 26.266 39.962 ;
      RECT 26.214 41.126 26.266 41.162 ;
      RECT 26.214 42.326 26.266 42.362 ;
      RECT 26.214 43.526 26.266 43.562 ;
      RECT 26.214 44.726 26.266 44.762 ;
      RECT 26.214 45.926 26.266 45.962 ;
      RECT 26.214 47.126 26.266 47.162 ;
      RECT 26.214 48.326 26.266 48.362 ;
      RECT 26.214 49.526 26.266 49.562 ;
      RECT 26.214 50.726 26.266 50.762 ;
      RECT 26.214 51.926 26.266 51.962 ;
      RECT 26.214 53.126 26.266 53.162 ;
      RECT 26.214 54.326 26.266 54.362 ;
      RECT 26.214 55.526 26.266 55.562 ;
      RECT 26.214 56.726 26.266 56.762 ;
      RECT 26.214 57.926 26.266 57.962 ;
      RECT 26.214 59.126 26.266 59.162 ;
      RECT 26.214 60.326 26.266 60.362 ;
      RECT 26.214 61.526 26.266 61.562 ;
      RECT 26.214 62.726 26.266 62.762 ;
      RECT 26.214 63.926 26.266 63.962 ;
      RECT 26.214 65.126 26.266 65.162 ;
      RECT 26.214 66.326 26.266 66.362 ;
      RECT 26.214 67.526 26.266 67.562 ;
      RECT 26.214 68.726 26.266 68.762 ;
      RECT 26.214 69.926 26.266 69.962 ;
      RECT 26.214 71.126 26.266 71.162 ;
      RECT 26.294 1.558 26.346 1.594 ;
      RECT 26.294 2.758 26.346 2.794 ;
      RECT 26.294 3.958 26.346 3.994 ;
      RECT 26.294 5.158 26.346 5.194 ;
      RECT 26.294 6.358 26.346 6.394 ;
      RECT 26.294 7.558 26.346 7.594 ;
      RECT 26.294 8.758 26.346 8.794 ;
      RECT 26.294 9.958 26.346 9.994 ;
      RECT 26.294 11.158 26.346 11.194 ;
      RECT 26.294 12.358 26.346 12.394 ;
      RECT 26.294 13.558 26.346 13.594 ;
      RECT 26.294 14.758 26.346 14.794 ;
      RECT 26.294 15.958 26.346 15.994 ;
      RECT 26.294 17.158 26.346 17.194 ;
      RECT 26.294 18.358 26.346 18.394 ;
      RECT 26.294 19.558 26.346 19.594 ;
      RECT 26.294 20.758 26.346 20.794 ;
      RECT 26.294 21.958 26.346 21.994 ;
      RECT 26.294 23.158 26.346 23.194 ;
      RECT 26.294 24.358 26.346 24.394 ;
      RECT 26.294 25.558 26.346 25.594 ;
      RECT 26.294 26.758 26.346 26.794 ;
      RECT 26.294 27.958 26.346 27.994 ;
      RECT 26.294 29.158 26.346 29.194 ;
      RECT 26.294 30.358 26.346 30.394 ;
      RECT 26.294 31.558 26.346 31.594 ;
      RECT 26.294 33.342 26.346 33.378 ;
      RECT 26.294 33.582 26.346 33.618 ;
      RECT 26.294 37.902 26.346 37.938 ;
      RECT 26.294 38.142 26.346 38.178 ;
      RECT 26.294 40.678 26.346 40.714 ;
      RECT 26.294 41.878 26.346 41.914 ;
      RECT 26.294 43.078 26.346 43.114 ;
      RECT 26.294 44.278 26.346 44.314 ;
      RECT 26.294 45.478 26.346 45.514 ;
      RECT 26.294 46.678 26.346 46.714 ;
      RECT 26.294 47.878 26.346 47.914 ;
      RECT 26.294 49.078 26.346 49.114 ;
      RECT 26.294 50.278 26.346 50.314 ;
      RECT 26.294 51.478 26.346 51.514 ;
      RECT 26.294 52.678 26.346 52.714 ;
      RECT 26.294 53.878 26.346 53.914 ;
      RECT 26.294 55.078 26.346 55.114 ;
      RECT 26.294 56.278 26.346 56.314 ;
      RECT 26.294 57.478 26.346 57.514 ;
      RECT 26.294 58.678 26.346 58.714 ;
      RECT 26.294 59.878 26.346 59.914 ;
      RECT 26.294 61.078 26.346 61.114 ;
      RECT 26.294 62.278 26.346 62.314 ;
      RECT 26.294 63.478 26.346 63.514 ;
      RECT 26.294 64.678 26.346 64.714 ;
      RECT 26.294 65.878 26.346 65.914 ;
      RECT 26.294 67.078 26.346 67.114 ;
      RECT 26.294 68.278 26.346 68.314 ;
      RECT 26.294 69.478 26.346 69.514 ;
      RECT 26.294 70.678 26.346 70.714 ;
      RECT 26.294 71.878 26.346 71.914 ;
      RECT 26.374 0.281 26.426 0.317 ;
      RECT 26.374 72.403 26.426 72.439 ;
      RECT 26.454 0.806 26.506 0.842 ;
      RECT 26.454 2.006 26.506 2.042 ;
      RECT 26.454 3.206 26.506 3.242 ;
      RECT 26.454 4.406 26.506 4.442 ;
      RECT 26.454 5.606 26.506 5.642 ;
      RECT 26.454 6.806 26.506 6.842 ;
      RECT 26.454 8.006 26.506 8.042 ;
      RECT 26.454 9.206 26.506 9.242 ;
      RECT 26.454 10.406 26.506 10.442 ;
      RECT 26.454 11.606 26.506 11.642 ;
      RECT 26.454 12.806 26.506 12.842 ;
      RECT 26.454 14.006 26.506 14.042 ;
      RECT 26.454 15.206 26.506 15.242 ;
      RECT 26.454 16.406 26.506 16.442 ;
      RECT 26.454 17.606 26.506 17.642 ;
      RECT 26.454 18.806 26.506 18.842 ;
      RECT 26.454 20.006 26.506 20.042 ;
      RECT 26.454 21.206 26.506 21.242 ;
      RECT 26.454 22.406 26.506 22.442 ;
      RECT 26.454 23.606 26.506 23.642 ;
      RECT 26.454 24.806 26.506 24.842 ;
      RECT 26.454 26.006 26.506 26.042 ;
      RECT 26.454 27.206 26.506 27.242 ;
      RECT 26.454 28.406 26.506 28.442 ;
      RECT 26.454 29.606 26.506 29.642 ;
      RECT 26.454 30.806 26.506 30.842 ;
      RECT 26.454 32.622 26.506 32.658 ;
      RECT 26.454 32.862 26.506 32.898 ;
      RECT 26.454 34.302 26.506 34.338 ;
      RECT 26.454 34.782 26.506 34.818 ;
      RECT 26.454 36.702 26.506 36.738 ;
      RECT 26.454 37.182 26.506 37.218 ;
      RECT 26.454 38.622 26.506 38.658 ;
      RECT 26.454 38.862 26.506 38.898 ;
      RECT 26.454 39.926 26.506 39.962 ;
      RECT 26.454 41.126 26.506 41.162 ;
      RECT 26.454 42.326 26.506 42.362 ;
      RECT 26.454 43.526 26.506 43.562 ;
      RECT 26.454 44.726 26.506 44.762 ;
      RECT 26.454 45.926 26.506 45.962 ;
      RECT 26.454 47.126 26.506 47.162 ;
      RECT 26.454 48.326 26.506 48.362 ;
      RECT 26.454 49.526 26.506 49.562 ;
      RECT 26.454 50.726 26.506 50.762 ;
      RECT 26.454 51.926 26.506 51.962 ;
      RECT 26.454 53.126 26.506 53.162 ;
      RECT 26.454 54.326 26.506 54.362 ;
      RECT 26.454 55.526 26.506 55.562 ;
      RECT 26.454 56.726 26.506 56.762 ;
      RECT 26.454 57.926 26.506 57.962 ;
      RECT 26.454 59.126 26.506 59.162 ;
      RECT 26.454 60.326 26.506 60.362 ;
      RECT 26.454 61.526 26.506 61.562 ;
      RECT 26.454 62.726 26.506 62.762 ;
      RECT 26.454 63.926 26.506 63.962 ;
      RECT 26.454 65.126 26.506 65.162 ;
      RECT 26.454 66.326 26.506 66.362 ;
      RECT 26.454 67.526 26.506 67.562 ;
      RECT 26.454 68.726 26.506 68.762 ;
      RECT 26.454 69.926 26.506 69.962 ;
      RECT 26.454 71.126 26.506 71.162 ;
      RECT 26.534 1.558 26.586 1.594 ;
      RECT 26.534 2.758 26.586 2.794 ;
      RECT 26.534 3.958 26.586 3.994 ;
      RECT 26.534 5.158 26.586 5.194 ;
      RECT 26.534 6.358 26.586 6.394 ;
      RECT 26.534 7.558 26.586 7.594 ;
      RECT 26.534 8.758 26.586 8.794 ;
      RECT 26.534 9.958 26.586 9.994 ;
      RECT 26.534 11.158 26.586 11.194 ;
      RECT 26.534 12.358 26.586 12.394 ;
      RECT 26.534 13.558 26.586 13.594 ;
      RECT 26.534 14.758 26.586 14.794 ;
      RECT 26.534 15.958 26.586 15.994 ;
      RECT 26.534 17.158 26.586 17.194 ;
      RECT 26.534 18.358 26.586 18.394 ;
      RECT 26.534 19.558 26.586 19.594 ;
      RECT 26.534 20.758 26.586 20.794 ;
      RECT 26.534 21.958 26.586 21.994 ;
      RECT 26.534 23.158 26.586 23.194 ;
      RECT 26.534 24.358 26.586 24.394 ;
      RECT 26.534 25.558 26.586 25.594 ;
      RECT 26.534 26.758 26.586 26.794 ;
      RECT 26.534 27.958 26.586 27.994 ;
      RECT 26.534 29.158 26.586 29.194 ;
      RECT 26.534 30.358 26.586 30.394 ;
      RECT 26.534 31.558 26.586 31.594 ;
      RECT 26.534 33.342 26.586 33.378 ;
      RECT 26.534 33.582 26.586 33.618 ;
      RECT 26.534 37.902 26.586 37.938 ;
      RECT 26.534 38.142 26.586 38.178 ;
      RECT 26.534 40.678 26.586 40.714 ;
      RECT 26.534 41.878 26.586 41.914 ;
      RECT 26.534 43.078 26.586 43.114 ;
      RECT 26.534 44.278 26.586 44.314 ;
      RECT 26.534 45.478 26.586 45.514 ;
      RECT 26.534 46.678 26.586 46.714 ;
      RECT 26.534 47.878 26.586 47.914 ;
      RECT 26.534 49.078 26.586 49.114 ;
      RECT 26.534 50.278 26.586 50.314 ;
      RECT 26.534 51.478 26.586 51.514 ;
      RECT 26.534 52.678 26.586 52.714 ;
      RECT 26.534 53.878 26.586 53.914 ;
      RECT 26.534 55.078 26.586 55.114 ;
      RECT 26.534 56.278 26.586 56.314 ;
      RECT 26.534 57.478 26.586 57.514 ;
      RECT 26.534 58.678 26.586 58.714 ;
      RECT 26.534 59.878 26.586 59.914 ;
      RECT 26.534 61.078 26.586 61.114 ;
      RECT 26.534 62.278 26.586 62.314 ;
      RECT 26.534 63.478 26.586 63.514 ;
      RECT 26.534 64.678 26.586 64.714 ;
      RECT 26.534 65.878 26.586 65.914 ;
      RECT 26.534 67.078 26.586 67.114 ;
      RECT 26.534 68.278 26.586 68.314 ;
      RECT 26.534 69.478 26.586 69.514 ;
      RECT 26.534 70.678 26.586 70.714 ;
      RECT 26.534 71.878 26.586 71.914 ;
      RECT 26.614 0.806 26.666 0.842 ;
      RECT 26.614 2.006 26.666 2.042 ;
      RECT 26.614 3.206 26.666 3.242 ;
      RECT 26.614 4.406 26.666 4.442 ;
      RECT 26.614 5.606 26.666 5.642 ;
      RECT 26.614 6.806 26.666 6.842 ;
      RECT 26.614 8.006 26.666 8.042 ;
      RECT 26.614 9.206 26.666 9.242 ;
      RECT 26.614 10.406 26.666 10.442 ;
      RECT 26.614 11.606 26.666 11.642 ;
      RECT 26.614 12.806 26.666 12.842 ;
      RECT 26.614 14.006 26.666 14.042 ;
      RECT 26.614 15.206 26.666 15.242 ;
      RECT 26.614 16.406 26.666 16.442 ;
      RECT 26.614 17.606 26.666 17.642 ;
      RECT 26.614 18.806 26.666 18.842 ;
      RECT 26.614 20.006 26.666 20.042 ;
      RECT 26.614 21.206 26.666 21.242 ;
      RECT 26.614 22.406 26.666 22.442 ;
      RECT 26.614 23.606 26.666 23.642 ;
      RECT 26.614 24.806 26.666 24.842 ;
      RECT 26.614 26.006 26.666 26.042 ;
      RECT 26.614 27.206 26.666 27.242 ;
      RECT 26.614 28.406 26.666 28.442 ;
      RECT 26.614 29.606 26.666 29.642 ;
      RECT 26.614 30.806 26.666 30.842 ;
      RECT 26.614 32.622 26.666 32.658 ;
      RECT 26.614 32.862 26.666 32.898 ;
      RECT 26.614 38.622 26.666 38.658 ;
      RECT 26.614 38.862 26.666 38.898 ;
      RECT 26.614 39.926 26.666 39.962 ;
      RECT 26.614 41.126 26.666 41.162 ;
      RECT 26.614 42.326 26.666 42.362 ;
      RECT 26.614 43.526 26.666 43.562 ;
      RECT 26.614 44.726 26.666 44.762 ;
      RECT 26.614 45.926 26.666 45.962 ;
      RECT 26.614 47.126 26.666 47.162 ;
      RECT 26.614 48.326 26.666 48.362 ;
      RECT 26.614 49.526 26.666 49.562 ;
      RECT 26.614 50.726 26.666 50.762 ;
      RECT 26.614 51.926 26.666 51.962 ;
      RECT 26.614 53.126 26.666 53.162 ;
      RECT 26.614 54.326 26.666 54.362 ;
      RECT 26.614 55.526 26.666 55.562 ;
      RECT 26.614 56.726 26.666 56.762 ;
      RECT 26.614 57.926 26.666 57.962 ;
      RECT 26.614 59.126 26.666 59.162 ;
      RECT 26.614 60.326 26.666 60.362 ;
      RECT 26.614 61.526 26.666 61.562 ;
      RECT 26.614 62.726 26.666 62.762 ;
      RECT 26.614 63.926 26.666 63.962 ;
      RECT 26.614 65.126 26.666 65.162 ;
      RECT 26.614 66.326 26.666 66.362 ;
      RECT 26.614 67.526 26.666 67.562 ;
      RECT 26.614 68.726 26.666 68.762 ;
      RECT 26.614 69.926 26.666 69.962 ;
      RECT 26.614 71.126 26.666 71.162 ;
      RECT 26.694 1.558 26.746 1.594 ;
      RECT 26.694 2.758 26.746 2.794 ;
      RECT 26.694 3.958 26.746 3.994 ;
      RECT 26.694 5.158 26.746 5.194 ;
      RECT 26.694 6.358 26.746 6.394 ;
      RECT 26.694 7.558 26.746 7.594 ;
      RECT 26.694 8.758 26.746 8.794 ;
      RECT 26.694 9.958 26.746 9.994 ;
      RECT 26.694 11.158 26.746 11.194 ;
      RECT 26.694 12.358 26.746 12.394 ;
      RECT 26.694 13.558 26.746 13.594 ;
      RECT 26.694 14.758 26.746 14.794 ;
      RECT 26.694 15.958 26.746 15.994 ;
      RECT 26.694 17.158 26.746 17.194 ;
      RECT 26.694 18.358 26.746 18.394 ;
      RECT 26.694 19.558 26.746 19.594 ;
      RECT 26.694 20.758 26.746 20.794 ;
      RECT 26.694 21.958 26.746 21.994 ;
      RECT 26.694 23.158 26.746 23.194 ;
      RECT 26.694 24.358 26.746 24.394 ;
      RECT 26.694 25.558 26.746 25.594 ;
      RECT 26.694 26.758 26.746 26.794 ;
      RECT 26.694 27.958 26.746 27.994 ;
      RECT 26.694 29.158 26.746 29.194 ;
      RECT 26.694 30.358 26.746 30.394 ;
      RECT 26.694 31.558 26.746 31.594 ;
      RECT 26.694 33.342 26.746 33.378 ;
      RECT 26.694 33.582 26.746 33.618 ;
      RECT 26.694 37.902 26.746 37.938 ;
      RECT 26.694 38.142 26.746 38.178 ;
      RECT 26.694 40.678 26.746 40.714 ;
      RECT 26.694 41.878 26.746 41.914 ;
      RECT 26.694 43.078 26.746 43.114 ;
      RECT 26.694 44.278 26.746 44.314 ;
      RECT 26.694 45.478 26.746 45.514 ;
      RECT 26.694 46.678 26.746 46.714 ;
      RECT 26.694 47.878 26.746 47.914 ;
      RECT 26.694 49.078 26.746 49.114 ;
      RECT 26.694 50.278 26.746 50.314 ;
      RECT 26.694 51.478 26.746 51.514 ;
      RECT 26.694 52.678 26.746 52.714 ;
      RECT 26.694 53.878 26.746 53.914 ;
      RECT 26.694 55.078 26.746 55.114 ;
      RECT 26.694 56.278 26.746 56.314 ;
      RECT 26.694 57.478 26.746 57.514 ;
      RECT 26.694 58.678 26.746 58.714 ;
      RECT 26.694 59.878 26.746 59.914 ;
      RECT 26.694 61.078 26.746 61.114 ;
      RECT 26.694 62.278 26.746 62.314 ;
      RECT 26.694 63.478 26.746 63.514 ;
      RECT 26.694 64.678 26.746 64.714 ;
      RECT 26.694 65.878 26.746 65.914 ;
      RECT 26.694 67.078 26.746 67.114 ;
      RECT 26.694 68.278 26.746 68.314 ;
      RECT 26.694 69.478 26.746 69.514 ;
      RECT 26.694 70.678 26.746 70.714 ;
      RECT 26.694 71.878 26.746 71.914 ;
      RECT 26.774 0.281 26.826 0.317 ;
      RECT 26.774 72.403 26.826 72.439 ;
      RECT 26.854 0.806 26.906 0.842 ;
      RECT 26.854 2.006 26.906 2.042 ;
      RECT 26.854 3.206 26.906 3.242 ;
      RECT 26.854 4.406 26.906 4.442 ;
      RECT 26.854 5.606 26.906 5.642 ;
      RECT 26.854 6.806 26.906 6.842 ;
      RECT 26.854 8.006 26.906 8.042 ;
      RECT 26.854 9.206 26.906 9.242 ;
      RECT 26.854 10.406 26.906 10.442 ;
      RECT 26.854 11.606 26.906 11.642 ;
      RECT 26.854 12.806 26.906 12.842 ;
      RECT 26.854 14.006 26.906 14.042 ;
      RECT 26.854 15.206 26.906 15.242 ;
      RECT 26.854 16.406 26.906 16.442 ;
      RECT 26.854 17.606 26.906 17.642 ;
      RECT 26.854 18.806 26.906 18.842 ;
      RECT 26.854 20.006 26.906 20.042 ;
      RECT 26.854 21.206 26.906 21.242 ;
      RECT 26.854 22.406 26.906 22.442 ;
      RECT 26.854 23.606 26.906 23.642 ;
      RECT 26.854 24.806 26.906 24.842 ;
      RECT 26.854 26.006 26.906 26.042 ;
      RECT 26.854 27.206 26.906 27.242 ;
      RECT 26.854 28.406 26.906 28.442 ;
      RECT 26.854 29.606 26.906 29.642 ;
      RECT 26.854 30.806 26.906 30.842 ;
      RECT 26.854 32.622 26.906 32.658 ;
      RECT 26.854 32.862 26.906 32.898 ;
      RECT 26.854 38.622 26.906 38.658 ;
      RECT 26.854 38.862 26.906 38.898 ;
      RECT 26.854 39.926 26.906 39.962 ;
      RECT 26.854 41.126 26.906 41.162 ;
      RECT 26.854 42.326 26.906 42.362 ;
      RECT 26.854 43.526 26.906 43.562 ;
      RECT 26.854 44.726 26.906 44.762 ;
      RECT 26.854 45.926 26.906 45.962 ;
      RECT 26.854 47.126 26.906 47.162 ;
      RECT 26.854 48.326 26.906 48.362 ;
      RECT 26.854 49.526 26.906 49.562 ;
      RECT 26.854 50.726 26.906 50.762 ;
      RECT 26.854 51.926 26.906 51.962 ;
      RECT 26.854 53.126 26.906 53.162 ;
      RECT 26.854 54.326 26.906 54.362 ;
      RECT 26.854 55.526 26.906 55.562 ;
      RECT 26.854 56.726 26.906 56.762 ;
      RECT 26.854 57.926 26.906 57.962 ;
      RECT 26.854 59.126 26.906 59.162 ;
      RECT 26.854 60.326 26.906 60.362 ;
      RECT 26.854 61.526 26.906 61.562 ;
      RECT 26.854 62.726 26.906 62.762 ;
      RECT 26.854 63.926 26.906 63.962 ;
      RECT 26.854 65.126 26.906 65.162 ;
      RECT 26.854 66.326 26.906 66.362 ;
      RECT 26.854 67.526 26.906 67.562 ;
      RECT 26.854 68.726 26.906 68.762 ;
      RECT 26.854 69.926 26.906 69.962 ;
      RECT 26.854 71.126 26.906 71.162 ;
      RECT 26.934 1.558 26.986 1.594 ;
      RECT 26.934 2.758 26.986 2.794 ;
      RECT 26.934 3.958 26.986 3.994 ;
      RECT 26.934 5.158 26.986 5.194 ;
      RECT 26.934 6.358 26.986 6.394 ;
      RECT 26.934 7.558 26.986 7.594 ;
      RECT 26.934 8.758 26.986 8.794 ;
      RECT 26.934 9.958 26.986 9.994 ;
      RECT 26.934 11.158 26.986 11.194 ;
      RECT 26.934 12.358 26.986 12.394 ;
      RECT 26.934 13.558 26.986 13.594 ;
      RECT 26.934 14.758 26.986 14.794 ;
      RECT 26.934 15.958 26.986 15.994 ;
      RECT 26.934 17.158 26.986 17.194 ;
      RECT 26.934 18.358 26.986 18.394 ;
      RECT 26.934 19.558 26.986 19.594 ;
      RECT 26.934 20.758 26.986 20.794 ;
      RECT 26.934 21.958 26.986 21.994 ;
      RECT 26.934 23.158 26.986 23.194 ;
      RECT 26.934 24.358 26.986 24.394 ;
      RECT 26.934 25.558 26.986 25.594 ;
      RECT 26.934 26.758 26.986 26.794 ;
      RECT 26.934 27.958 26.986 27.994 ;
      RECT 26.934 29.158 26.986 29.194 ;
      RECT 26.934 30.358 26.986 30.394 ;
      RECT 26.934 31.558 26.986 31.594 ;
      RECT 26.934 33.342 26.986 33.378 ;
      RECT 26.934 33.582 26.986 33.618 ;
      RECT 26.934 37.902 26.986 37.938 ;
      RECT 26.934 38.142 26.986 38.178 ;
      RECT 26.934 40.678 26.986 40.714 ;
      RECT 26.934 41.878 26.986 41.914 ;
      RECT 26.934 43.078 26.986 43.114 ;
      RECT 26.934 44.278 26.986 44.314 ;
      RECT 26.934 45.478 26.986 45.514 ;
      RECT 26.934 46.678 26.986 46.714 ;
      RECT 26.934 47.878 26.986 47.914 ;
      RECT 26.934 49.078 26.986 49.114 ;
      RECT 26.934 50.278 26.986 50.314 ;
      RECT 26.934 51.478 26.986 51.514 ;
      RECT 26.934 52.678 26.986 52.714 ;
      RECT 26.934 53.878 26.986 53.914 ;
      RECT 26.934 55.078 26.986 55.114 ;
      RECT 26.934 56.278 26.986 56.314 ;
      RECT 26.934 57.478 26.986 57.514 ;
      RECT 26.934 58.678 26.986 58.714 ;
      RECT 26.934 59.878 26.986 59.914 ;
      RECT 26.934 61.078 26.986 61.114 ;
      RECT 26.934 62.278 26.986 62.314 ;
      RECT 26.934 63.478 26.986 63.514 ;
      RECT 26.934 64.678 26.986 64.714 ;
      RECT 26.934 65.878 26.986 65.914 ;
      RECT 26.934 67.078 26.986 67.114 ;
      RECT 26.934 68.278 26.986 68.314 ;
      RECT 26.934 69.478 26.986 69.514 ;
      RECT 26.934 70.678 26.986 70.714 ;
      RECT 26.934 71.878 26.986 71.914 ;
      RECT 27.014 0.806 27.066 0.842 ;
      RECT 27.014 2.006 27.066 2.042 ;
      RECT 27.014 3.206 27.066 3.242 ;
      RECT 27.014 4.406 27.066 4.442 ;
      RECT 27.014 5.606 27.066 5.642 ;
      RECT 27.014 6.806 27.066 6.842 ;
      RECT 27.014 8.006 27.066 8.042 ;
      RECT 27.014 9.206 27.066 9.242 ;
      RECT 27.014 10.406 27.066 10.442 ;
      RECT 27.014 11.606 27.066 11.642 ;
      RECT 27.014 12.806 27.066 12.842 ;
      RECT 27.014 14.006 27.066 14.042 ;
      RECT 27.014 15.206 27.066 15.242 ;
      RECT 27.014 16.406 27.066 16.442 ;
      RECT 27.014 17.606 27.066 17.642 ;
      RECT 27.014 18.806 27.066 18.842 ;
      RECT 27.014 20.006 27.066 20.042 ;
      RECT 27.014 21.206 27.066 21.242 ;
      RECT 27.014 22.406 27.066 22.442 ;
      RECT 27.014 23.606 27.066 23.642 ;
      RECT 27.014 24.806 27.066 24.842 ;
      RECT 27.014 26.006 27.066 26.042 ;
      RECT 27.014 27.206 27.066 27.242 ;
      RECT 27.014 28.406 27.066 28.442 ;
      RECT 27.014 29.606 27.066 29.642 ;
      RECT 27.014 30.806 27.066 30.842 ;
      RECT 27.014 32.622 27.066 32.658 ;
      RECT 27.014 32.862 27.066 32.898 ;
      RECT 27.014 38.622 27.066 38.658 ;
      RECT 27.014 38.862 27.066 38.898 ;
      RECT 27.014 39.926 27.066 39.962 ;
      RECT 27.014 41.126 27.066 41.162 ;
      RECT 27.014 42.326 27.066 42.362 ;
      RECT 27.014 43.526 27.066 43.562 ;
      RECT 27.014 44.726 27.066 44.762 ;
      RECT 27.014 45.926 27.066 45.962 ;
      RECT 27.014 47.126 27.066 47.162 ;
      RECT 27.014 48.326 27.066 48.362 ;
      RECT 27.014 49.526 27.066 49.562 ;
      RECT 27.014 50.726 27.066 50.762 ;
      RECT 27.014 51.926 27.066 51.962 ;
      RECT 27.014 53.126 27.066 53.162 ;
      RECT 27.014 54.326 27.066 54.362 ;
      RECT 27.014 55.526 27.066 55.562 ;
      RECT 27.014 56.726 27.066 56.762 ;
      RECT 27.014 57.926 27.066 57.962 ;
      RECT 27.014 59.126 27.066 59.162 ;
      RECT 27.014 60.326 27.066 60.362 ;
      RECT 27.014 61.526 27.066 61.562 ;
      RECT 27.014 62.726 27.066 62.762 ;
      RECT 27.014 63.926 27.066 63.962 ;
      RECT 27.014 65.126 27.066 65.162 ;
      RECT 27.014 66.326 27.066 66.362 ;
      RECT 27.014 67.526 27.066 67.562 ;
      RECT 27.014 68.726 27.066 68.762 ;
      RECT 27.014 69.926 27.066 69.962 ;
      RECT 27.014 71.126 27.066 71.162 ;
      RECT 27.094 1.558 27.146 1.594 ;
      RECT 27.094 2.758 27.146 2.794 ;
      RECT 27.094 3.958 27.146 3.994 ;
      RECT 27.094 5.158 27.146 5.194 ;
      RECT 27.094 6.358 27.146 6.394 ;
      RECT 27.094 7.558 27.146 7.594 ;
      RECT 27.094 8.758 27.146 8.794 ;
      RECT 27.094 9.958 27.146 9.994 ;
      RECT 27.094 11.158 27.146 11.194 ;
      RECT 27.094 12.358 27.146 12.394 ;
      RECT 27.094 13.558 27.146 13.594 ;
      RECT 27.094 14.758 27.146 14.794 ;
      RECT 27.094 15.958 27.146 15.994 ;
      RECT 27.094 17.158 27.146 17.194 ;
      RECT 27.094 18.358 27.146 18.394 ;
      RECT 27.094 19.558 27.146 19.594 ;
      RECT 27.094 20.758 27.146 20.794 ;
      RECT 27.094 21.958 27.146 21.994 ;
      RECT 27.094 23.158 27.146 23.194 ;
      RECT 27.094 24.358 27.146 24.394 ;
      RECT 27.094 25.558 27.146 25.594 ;
      RECT 27.094 26.758 27.146 26.794 ;
      RECT 27.094 27.958 27.146 27.994 ;
      RECT 27.094 29.158 27.146 29.194 ;
      RECT 27.094 30.358 27.146 30.394 ;
      RECT 27.094 31.558 27.146 31.594 ;
      RECT 27.094 33.342 27.146 33.378 ;
      RECT 27.094 33.582 27.146 33.618 ;
      RECT 27.094 37.902 27.146 37.938 ;
      RECT 27.094 38.142 27.146 38.178 ;
      RECT 27.094 40.678 27.146 40.714 ;
      RECT 27.094 41.878 27.146 41.914 ;
      RECT 27.094 43.078 27.146 43.114 ;
      RECT 27.094 44.278 27.146 44.314 ;
      RECT 27.094 45.478 27.146 45.514 ;
      RECT 27.094 46.678 27.146 46.714 ;
      RECT 27.094 47.878 27.146 47.914 ;
      RECT 27.094 49.078 27.146 49.114 ;
      RECT 27.094 50.278 27.146 50.314 ;
      RECT 27.094 51.478 27.146 51.514 ;
      RECT 27.094 52.678 27.146 52.714 ;
      RECT 27.094 53.878 27.146 53.914 ;
      RECT 27.094 55.078 27.146 55.114 ;
      RECT 27.094 56.278 27.146 56.314 ;
      RECT 27.094 57.478 27.146 57.514 ;
      RECT 27.094 58.678 27.146 58.714 ;
      RECT 27.094 59.878 27.146 59.914 ;
      RECT 27.094 61.078 27.146 61.114 ;
      RECT 27.094 62.278 27.146 62.314 ;
      RECT 27.094 63.478 27.146 63.514 ;
      RECT 27.094 64.678 27.146 64.714 ;
      RECT 27.094 65.878 27.146 65.914 ;
      RECT 27.094 67.078 27.146 67.114 ;
      RECT 27.094 68.278 27.146 68.314 ;
      RECT 27.094 69.478 27.146 69.514 ;
      RECT 27.094 70.678 27.146 70.714 ;
      RECT 27.094 71.878 27.146 71.914 ;
      RECT 27.174 0.281 27.226 0.317 ;
      RECT 27.174 72.403 27.226 72.439 ;
      RECT 27.254 0.806 27.306 0.842 ;
      RECT 27.254 2.006 27.306 2.042 ;
      RECT 27.254 3.206 27.306 3.242 ;
      RECT 27.254 4.406 27.306 4.442 ;
      RECT 27.254 5.606 27.306 5.642 ;
      RECT 27.254 6.806 27.306 6.842 ;
      RECT 27.254 8.006 27.306 8.042 ;
      RECT 27.254 9.206 27.306 9.242 ;
      RECT 27.254 10.406 27.306 10.442 ;
      RECT 27.254 11.606 27.306 11.642 ;
      RECT 27.254 12.806 27.306 12.842 ;
      RECT 27.254 14.006 27.306 14.042 ;
      RECT 27.254 15.206 27.306 15.242 ;
      RECT 27.254 16.406 27.306 16.442 ;
      RECT 27.254 17.606 27.306 17.642 ;
      RECT 27.254 18.806 27.306 18.842 ;
      RECT 27.254 20.006 27.306 20.042 ;
      RECT 27.254 21.206 27.306 21.242 ;
      RECT 27.254 22.406 27.306 22.442 ;
      RECT 27.254 23.606 27.306 23.642 ;
      RECT 27.254 24.806 27.306 24.842 ;
      RECT 27.254 26.006 27.306 26.042 ;
      RECT 27.254 27.206 27.306 27.242 ;
      RECT 27.254 28.406 27.306 28.442 ;
      RECT 27.254 29.606 27.306 29.642 ;
      RECT 27.254 30.806 27.306 30.842 ;
      RECT 27.254 32.622 27.306 32.658 ;
      RECT 27.254 32.862 27.306 32.898 ;
      RECT 27.254 34.302 27.306 34.338 ;
      RECT 27.254 34.782 27.306 34.818 ;
      RECT 27.254 36.702 27.306 36.738 ;
      RECT 27.254 37.182 27.306 37.218 ;
      RECT 27.254 38.622 27.306 38.658 ;
      RECT 27.254 38.862 27.306 38.898 ;
      RECT 27.254 39.926 27.306 39.962 ;
      RECT 27.254 41.126 27.306 41.162 ;
      RECT 27.254 42.326 27.306 42.362 ;
      RECT 27.254 43.526 27.306 43.562 ;
      RECT 27.254 44.726 27.306 44.762 ;
      RECT 27.254 45.926 27.306 45.962 ;
      RECT 27.254 47.126 27.306 47.162 ;
      RECT 27.254 48.326 27.306 48.362 ;
      RECT 27.254 49.526 27.306 49.562 ;
      RECT 27.254 50.726 27.306 50.762 ;
      RECT 27.254 51.926 27.306 51.962 ;
      RECT 27.254 53.126 27.306 53.162 ;
      RECT 27.254 54.326 27.306 54.362 ;
      RECT 27.254 55.526 27.306 55.562 ;
      RECT 27.254 56.726 27.306 56.762 ;
      RECT 27.254 57.926 27.306 57.962 ;
      RECT 27.254 59.126 27.306 59.162 ;
      RECT 27.254 60.326 27.306 60.362 ;
      RECT 27.254 61.526 27.306 61.562 ;
      RECT 27.254 62.726 27.306 62.762 ;
      RECT 27.254 63.926 27.306 63.962 ;
      RECT 27.254 65.126 27.306 65.162 ;
      RECT 27.254 66.326 27.306 66.362 ;
      RECT 27.254 67.526 27.306 67.562 ;
      RECT 27.254 68.726 27.306 68.762 ;
      RECT 27.254 69.926 27.306 69.962 ;
      RECT 27.254 71.126 27.306 71.162 ;
      RECT 27.334 1.558 27.386 1.594 ;
      RECT 27.334 2.758 27.386 2.794 ;
      RECT 27.334 3.958 27.386 3.994 ;
      RECT 27.334 5.158 27.386 5.194 ;
      RECT 27.334 6.358 27.386 6.394 ;
      RECT 27.334 7.558 27.386 7.594 ;
      RECT 27.334 8.758 27.386 8.794 ;
      RECT 27.334 9.958 27.386 9.994 ;
      RECT 27.334 11.158 27.386 11.194 ;
      RECT 27.334 12.358 27.386 12.394 ;
      RECT 27.334 13.558 27.386 13.594 ;
      RECT 27.334 14.758 27.386 14.794 ;
      RECT 27.334 15.958 27.386 15.994 ;
      RECT 27.334 17.158 27.386 17.194 ;
      RECT 27.334 18.358 27.386 18.394 ;
      RECT 27.334 19.558 27.386 19.594 ;
      RECT 27.334 20.758 27.386 20.794 ;
      RECT 27.334 21.958 27.386 21.994 ;
      RECT 27.334 23.158 27.386 23.194 ;
      RECT 27.334 24.358 27.386 24.394 ;
      RECT 27.334 25.558 27.386 25.594 ;
      RECT 27.334 26.758 27.386 26.794 ;
      RECT 27.334 27.958 27.386 27.994 ;
      RECT 27.334 29.158 27.386 29.194 ;
      RECT 27.334 30.358 27.386 30.394 ;
      RECT 27.334 31.558 27.386 31.594 ;
      RECT 27.334 33.342 27.386 33.378 ;
      RECT 27.334 33.582 27.386 33.618 ;
      RECT 27.334 37.902 27.386 37.938 ;
      RECT 27.334 38.142 27.386 38.178 ;
      RECT 27.334 40.678 27.386 40.714 ;
      RECT 27.334 41.878 27.386 41.914 ;
      RECT 27.334 43.078 27.386 43.114 ;
      RECT 27.334 44.278 27.386 44.314 ;
      RECT 27.334 45.478 27.386 45.514 ;
      RECT 27.334 46.678 27.386 46.714 ;
      RECT 27.334 47.878 27.386 47.914 ;
      RECT 27.334 49.078 27.386 49.114 ;
      RECT 27.334 50.278 27.386 50.314 ;
      RECT 27.334 51.478 27.386 51.514 ;
      RECT 27.334 52.678 27.386 52.714 ;
      RECT 27.334 53.878 27.386 53.914 ;
      RECT 27.334 55.078 27.386 55.114 ;
      RECT 27.334 56.278 27.386 56.314 ;
      RECT 27.334 57.478 27.386 57.514 ;
      RECT 27.334 58.678 27.386 58.714 ;
      RECT 27.334 59.878 27.386 59.914 ;
      RECT 27.334 61.078 27.386 61.114 ;
      RECT 27.334 62.278 27.386 62.314 ;
      RECT 27.334 63.478 27.386 63.514 ;
      RECT 27.334 64.678 27.386 64.714 ;
      RECT 27.334 65.878 27.386 65.914 ;
      RECT 27.334 67.078 27.386 67.114 ;
      RECT 27.334 68.278 27.386 68.314 ;
      RECT 27.334 69.478 27.386 69.514 ;
      RECT 27.334 70.678 27.386 70.714 ;
      RECT 27.334 71.878 27.386 71.914 ;
      RECT 27.414 0.806 27.466 0.842 ;
      RECT 27.414 2.006 27.466 2.042 ;
      RECT 27.414 3.206 27.466 3.242 ;
      RECT 27.414 4.406 27.466 4.442 ;
      RECT 27.414 5.606 27.466 5.642 ;
      RECT 27.414 6.806 27.466 6.842 ;
      RECT 27.414 8.006 27.466 8.042 ;
      RECT 27.414 9.206 27.466 9.242 ;
      RECT 27.414 10.406 27.466 10.442 ;
      RECT 27.414 11.606 27.466 11.642 ;
      RECT 27.414 12.806 27.466 12.842 ;
      RECT 27.414 14.006 27.466 14.042 ;
      RECT 27.414 15.206 27.466 15.242 ;
      RECT 27.414 16.406 27.466 16.442 ;
      RECT 27.414 17.606 27.466 17.642 ;
      RECT 27.414 18.806 27.466 18.842 ;
      RECT 27.414 20.006 27.466 20.042 ;
      RECT 27.414 21.206 27.466 21.242 ;
      RECT 27.414 22.406 27.466 22.442 ;
      RECT 27.414 23.606 27.466 23.642 ;
      RECT 27.414 24.806 27.466 24.842 ;
      RECT 27.414 26.006 27.466 26.042 ;
      RECT 27.414 27.206 27.466 27.242 ;
      RECT 27.414 28.406 27.466 28.442 ;
      RECT 27.414 29.606 27.466 29.642 ;
      RECT 27.414 30.806 27.466 30.842 ;
      RECT 27.414 32.622 27.466 32.658 ;
      RECT 27.414 32.862 27.466 32.898 ;
      RECT 27.414 38.622 27.466 38.658 ;
      RECT 27.414 38.862 27.466 38.898 ;
      RECT 27.414 39.926 27.466 39.962 ;
      RECT 27.414 41.126 27.466 41.162 ;
      RECT 27.414 42.326 27.466 42.362 ;
      RECT 27.414 43.526 27.466 43.562 ;
      RECT 27.414 44.726 27.466 44.762 ;
      RECT 27.414 45.926 27.466 45.962 ;
      RECT 27.414 47.126 27.466 47.162 ;
      RECT 27.414 48.326 27.466 48.362 ;
      RECT 27.414 49.526 27.466 49.562 ;
      RECT 27.414 50.726 27.466 50.762 ;
      RECT 27.414 51.926 27.466 51.962 ;
      RECT 27.414 53.126 27.466 53.162 ;
      RECT 27.414 54.326 27.466 54.362 ;
      RECT 27.414 55.526 27.466 55.562 ;
      RECT 27.414 56.726 27.466 56.762 ;
      RECT 27.414 57.926 27.466 57.962 ;
      RECT 27.414 59.126 27.466 59.162 ;
      RECT 27.414 60.326 27.466 60.362 ;
      RECT 27.414 61.526 27.466 61.562 ;
      RECT 27.414 62.726 27.466 62.762 ;
      RECT 27.414 63.926 27.466 63.962 ;
      RECT 27.414 65.126 27.466 65.162 ;
      RECT 27.414 66.326 27.466 66.362 ;
      RECT 27.414 67.526 27.466 67.562 ;
      RECT 27.414 68.726 27.466 68.762 ;
      RECT 27.414 69.926 27.466 69.962 ;
      RECT 27.414 71.126 27.466 71.162 ;
      RECT 27.494 1.558 27.546 1.594 ;
      RECT 27.494 2.758 27.546 2.794 ;
      RECT 27.494 3.958 27.546 3.994 ;
      RECT 27.494 5.158 27.546 5.194 ;
      RECT 27.494 6.358 27.546 6.394 ;
      RECT 27.494 7.558 27.546 7.594 ;
      RECT 27.494 8.758 27.546 8.794 ;
      RECT 27.494 9.958 27.546 9.994 ;
      RECT 27.494 11.158 27.546 11.194 ;
      RECT 27.494 12.358 27.546 12.394 ;
      RECT 27.494 13.558 27.546 13.594 ;
      RECT 27.494 14.758 27.546 14.794 ;
      RECT 27.494 15.958 27.546 15.994 ;
      RECT 27.494 17.158 27.546 17.194 ;
      RECT 27.494 18.358 27.546 18.394 ;
      RECT 27.494 19.558 27.546 19.594 ;
      RECT 27.494 20.758 27.546 20.794 ;
      RECT 27.494 21.958 27.546 21.994 ;
      RECT 27.494 23.158 27.546 23.194 ;
      RECT 27.494 24.358 27.546 24.394 ;
      RECT 27.494 25.558 27.546 25.594 ;
      RECT 27.494 26.758 27.546 26.794 ;
      RECT 27.494 27.958 27.546 27.994 ;
      RECT 27.494 29.158 27.546 29.194 ;
      RECT 27.494 30.358 27.546 30.394 ;
      RECT 27.494 31.558 27.546 31.594 ;
      RECT 27.494 33.342 27.546 33.378 ;
      RECT 27.494 33.582 27.546 33.618 ;
      RECT 27.494 37.902 27.546 37.938 ;
      RECT 27.494 38.142 27.546 38.178 ;
      RECT 27.494 40.678 27.546 40.714 ;
      RECT 27.494 41.878 27.546 41.914 ;
      RECT 27.494 43.078 27.546 43.114 ;
      RECT 27.494 44.278 27.546 44.314 ;
      RECT 27.494 45.478 27.546 45.514 ;
      RECT 27.494 46.678 27.546 46.714 ;
      RECT 27.494 47.878 27.546 47.914 ;
      RECT 27.494 49.078 27.546 49.114 ;
      RECT 27.494 50.278 27.546 50.314 ;
      RECT 27.494 51.478 27.546 51.514 ;
      RECT 27.494 52.678 27.546 52.714 ;
      RECT 27.494 53.878 27.546 53.914 ;
      RECT 27.494 55.078 27.546 55.114 ;
      RECT 27.494 56.278 27.546 56.314 ;
      RECT 27.494 57.478 27.546 57.514 ;
      RECT 27.494 58.678 27.546 58.714 ;
      RECT 27.494 59.878 27.546 59.914 ;
      RECT 27.494 61.078 27.546 61.114 ;
      RECT 27.494 62.278 27.546 62.314 ;
      RECT 27.494 63.478 27.546 63.514 ;
      RECT 27.494 64.678 27.546 64.714 ;
      RECT 27.494 65.878 27.546 65.914 ;
      RECT 27.494 67.078 27.546 67.114 ;
      RECT 27.494 68.278 27.546 68.314 ;
      RECT 27.494 69.478 27.546 69.514 ;
      RECT 27.494 70.678 27.546 70.714 ;
      RECT 27.494 71.878 27.546 71.914 ;
      RECT 27.574 0.281 27.626 0.317 ;
      RECT 27.574 72.403 27.626 72.439 ;
      RECT 27.654 0.806 27.706 0.842 ;
      RECT 27.654 2.006 27.706 2.042 ;
      RECT 27.654 3.206 27.706 3.242 ;
      RECT 27.654 4.406 27.706 4.442 ;
      RECT 27.654 5.606 27.706 5.642 ;
      RECT 27.654 6.806 27.706 6.842 ;
      RECT 27.654 8.006 27.706 8.042 ;
      RECT 27.654 9.206 27.706 9.242 ;
      RECT 27.654 10.406 27.706 10.442 ;
      RECT 27.654 11.606 27.706 11.642 ;
      RECT 27.654 12.806 27.706 12.842 ;
      RECT 27.654 14.006 27.706 14.042 ;
      RECT 27.654 15.206 27.706 15.242 ;
      RECT 27.654 16.406 27.706 16.442 ;
      RECT 27.654 17.606 27.706 17.642 ;
      RECT 27.654 18.806 27.706 18.842 ;
      RECT 27.654 20.006 27.706 20.042 ;
      RECT 27.654 21.206 27.706 21.242 ;
      RECT 27.654 22.406 27.706 22.442 ;
      RECT 27.654 23.606 27.706 23.642 ;
      RECT 27.654 24.806 27.706 24.842 ;
      RECT 27.654 26.006 27.706 26.042 ;
      RECT 27.654 27.206 27.706 27.242 ;
      RECT 27.654 28.406 27.706 28.442 ;
      RECT 27.654 29.606 27.706 29.642 ;
      RECT 27.654 30.806 27.706 30.842 ;
      RECT 27.654 32.622 27.706 32.658 ;
      RECT 27.654 32.862 27.706 32.898 ;
      RECT 27.654 38.622 27.706 38.658 ;
      RECT 27.654 38.862 27.706 38.898 ;
      RECT 27.654 39.926 27.706 39.962 ;
      RECT 27.654 41.126 27.706 41.162 ;
      RECT 27.654 42.326 27.706 42.362 ;
      RECT 27.654 43.526 27.706 43.562 ;
      RECT 27.654 44.726 27.706 44.762 ;
      RECT 27.654 45.926 27.706 45.962 ;
      RECT 27.654 47.126 27.706 47.162 ;
      RECT 27.654 48.326 27.706 48.362 ;
      RECT 27.654 49.526 27.706 49.562 ;
      RECT 27.654 50.726 27.706 50.762 ;
      RECT 27.654 51.926 27.706 51.962 ;
      RECT 27.654 53.126 27.706 53.162 ;
      RECT 27.654 54.326 27.706 54.362 ;
      RECT 27.654 55.526 27.706 55.562 ;
      RECT 27.654 56.726 27.706 56.762 ;
      RECT 27.654 57.926 27.706 57.962 ;
      RECT 27.654 59.126 27.706 59.162 ;
      RECT 27.654 60.326 27.706 60.362 ;
      RECT 27.654 61.526 27.706 61.562 ;
      RECT 27.654 62.726 27.706 62.762 ;
      RECT 27.654 63.926 27.706 63.962 ;
      RECT 27.654 65.126 27.706 65.162 ;
      RECT 27.654 66.326 27.706 66.362 ;
      RECT 27.654 67.526 27.706 67.562 ;
      RECT 27.654 68.726 27.706 68.762 ;
      RECT 27.654 69.926 27.706 69.962 ;
      RECT 27.654 71.126 27.706 71.162 ;
      RECT 27.734 1.558 27.786 1.594 ;
      RECT 27.734 2.758 27.786 2.794 ;
      RECT 27.734 3.958 27.786 3.994 ;
      RECT 27.734 5.158 27.786 5.194 ;
      RECT 27.734 6.358 27.786 6.394 ;
      RECT 27.734 7.558 27.786 7.594 ;
      RECT 27.734 8.758 27.786 8.794 ;
      RECT 27.734 9.958 27.786 9.994 ;
      RECT 27.734 11.158 27.786 11.194 ;
      RECT 27.734 12.358 27.786 12.394 ;
      RECT 27.734 13.558 27.786 13.594 ;
      RECT 27.734 14.758 27.786 14.794 ;
      RECT 27.734 15.958 27.786 15.994 ;
      RECT 27.734 17.158 27.786 17.194 ;
      RECT 27.734 18.358 27.786 18.394 ;
      RECT 27.734 19.558 27.786 19.594 ;
      RECT 27.734 20.758 27.786 20.794 ;
      RECT 27.734 21.958 27.786 21.994 ;
      RECT 27.734 23.158 27.786 23.194 ;
      RECT 27.734 24.358 27.786 24.394 ;
      RECT 27.734 25.558 27.786 25.594 ;
      RECT 27.734 26.758 27.786 26.794 ;
      RECT 27.734 27.958 27.786 27.994 ;
      RECT 27.734 29.158 27.786 29.194 ;
      RECT 27.734 30.358 27.786 30.394 ;
      RECT 27.734 31.558 27.786 31.594 ;
      RECT 27.734 33.342 27.786 33.378 ;
      RECT 27.734 33.582 27.786 33.618 ;
      RECT 27.734 37.902 27.786 37.938 ;
      RECT 27.734 38.142 27.786 38.178 ;
      RECT 27.734 40.678 27.786 40.714 ;
      RECT 27.734 41.878 27.786 41.914 ;
      RECT 27.734 43.078 27.786 43.114 ;
      RECT 27.734 44.278 27.786 44.314 ;
      RECT 27.734 45.478 27.786 45.514 ;
      RECT 27.734 46.678 27.786 46.714 ;
      RECT 27.734 47.878 27.786 47.914 ;
      RECT 27.734 49.078 27.786 49.114 ;
      RECT 27.734 50.278 27.786 50.314 ;
      RECT 27.734 51.478 27.786 51.514 ;
      RECT 27.734 52.678 27.786 52.714 ;
      RECT 27.734 53.878 27.786 53.914 ;
      RECT 27.734 55.078 27.786 55.114 ;
      RECT 27.734 56.278 27.786 56.314 ;
      RECT 27.734 57.478 27.786 57.514 ;
      RECT 27.734 58.678 27.786 58.714 ;
      RECT 27.734 59.878 27.786 59.914 ;
      RECT 27.734 61.078 27.786 61.114 ;
      RECT 27.734 62.278 27.786 62.314 ;
      RECT 27.734 63.478 27.786 63.514 ;
      RECT 27.734 64.678 27.786 64.714 ;
      RECT 27.734 65.878 27.786 65.914 ;
      RECT 27.734 67.078 27.786 67.114 ;
      RECT 27.734 68.278 27.786 68.314 ;
      RECT 27.734 69.478 27.786 69.514 ;
      RECT 27.734 70.678 27.786 70.714 ;
      RECT 27.734 71.878 27.786 71.914 ;
      RECT 27.814 0.806 27.866 0.842 ;
      RECT 27.814 2.006 27.866 2.042 ;
      RECT 27.814 3.206 27.866 3.242 ;
      RECT 27.814 4.406 27.866 4.442 ;
      RECT 27.814 5.606 27.866 5.642 ;
      RECT 27.814 6.806 27.866 6.842 ;
      RECT 27.814 8.006 27.866 8.042 ;
      RECT 27.814 9.206 27.866 9.242 ;
      RECT 27.814 10.406 27.866 10.442 ;
      RECT 27.814 11.606 27.866 11.642 ;
      RECT 27.814 12.806 27.866 12.842 ;
      RECT 27.814 14.006 27.866 14.042 ;
      RECT 27.814 15.206 27.866 15.242 ;
      RECT 27.814 16.406 27.866 16.442 ;
      RECT 27.814 17.606 27.866 17.642 ;
      RECT 27.814 18.806 27.866 18.842 ;
      RECT 27.814 20.006 27.866 20.042 ;
      RECT 27.814 21.206 27.866 21.242 ;
      RECT 27.814 22.406 27.866 22.442 ;
      RECT 27.814 23.606 27.866 23.642 ;
      RECT 27.814 24.806 27.866 24.842 ;
      RECT 27.814 26.006 27.866 26.042 ;
      RECT 27.814 27.206 27.866 27.242 ;
      RECT 27.814 28.406 27.866 28.442 ;
      RECT 27.814 29.606 27.866 29.642 ;
      RECT 27.814 30.806 27.866 30.842 ;
      RECT 27.814 32.622 27.866 32.658 ;
      RECT 27.814 32.862 27.866 32.898 ;
      RECT 27.814 38.622 27.866 38.658 ;
      RECT 27.814 38.862 27.866 38.898 ;
      RECT 27.814 39.926 27.866 39.962 ;
      RECT 27.814 41.126 27.866 41.162 ;
      RECT 27.814 42.326 27.866 42.362 ;
      RECT 27.814 43.526 27.866 43.562 ;
      RECT 27.814 44.726 27.866 44.762 ;
      RECT 27.814 45.926 27.866 45.962 ;
      RECT 27.814 47.126 27.866 47.162 ;
      RECT 27.814 48.326 27.866 48.362 ;
      RECT 27.814 49.526 27.866 49.562 ;
      RECT 27.814 50.726 27.866 50.762 ;
      RECT 27.814 51.926 27.866 51.962 ;
      RECT 27.814 53.126 27.866 53.162 ;
      RECT 27.814 54.326 27.866 54.362 ;
      RECT 27.814 55.526 27.866 55.562 ;
      RECT 27.814 56.726 27.866 56.762 ;
      RECT 27.814 57.926 27.866 57.962 ;
      RECT 27.814 59.126 27.866 59.162 ;
      RECT 27.814 60.326 27.866 60.362 ;
      RECT 27.814 61.526 27.866 61.562 ;
      RECT 27.814 62.726 27.866 62.762 ;
      RECT 27.814 63.926 27.866 63.962 ;
      RECT 27.814 65.126 27.866 65.162 ;
      RECT 27.814 66.326 27.866 66.362 ;
      RECT 27.814 67.526 27.866 67.562 ;
      RECT 27.814 68.726 27.866 68.762 ;
      RECT 27.814 69.926 27.866 69.962 ;
      RECT 27.814 71.126 27.866 71.162 ;
      RECT 27.894 1.558 27.946 1.594 ;
      RECT 27.894 2.758 27.946 2.794 ;
      RECT 27.894 3.958 27.946 3.994 ;
      RECT 27.894 5.158 27.946 5.194 ;
      RECT 27.894 6.358 27.946 6.394 ;
      RECT 27.894 7.558 27.946 7.594 ;
      RECT 27.894 8.758 27.946 8.794 ;
      RECT 27.894 9.958 27.946 9.994 ;
      RECT 27.894 11.158 27.946 11.194 ;
      RECT 27.894 12.358 27.946 12.394 ;
      RECT 27.894 13.558 27.946 13.594 ;
      RECT 27.894 14.758 27.946 14.794 ;
      RECT 27.894 15.958 27.946 15.994 ;
      RECT 27.894 17.158 27.946 17.194 ;
      RECT 27.894 18.358 27.946 18.394 ;
      RECT 27.894 19.558 27.946 19.594 ;
      RECT 27.894 20.758 27.946 20.794 ;
      RECT 27.894 21.958 27.946 21.994 ;
      RECT 27.894 23.158 27.946 23.194 ;
      RECT 27.894 24.358 27.946 24.394 ;
      RECT 27.894 25.558 27.946 25.594 ;
      RECT 27.894 26.758 27.946 26.794 ;
      RECT 27.894 27.958 27.946 27.994 ;
      RECT 27.894 29.158 27.946 29.194 ;
      RECT 27.894 30.358 27.946 30.394 ;
      RECT 27.894 31.558 27.946 31.594 ;
      RECT 27.894 33.342 27.946 33.378 ;
      RECT 27.894 33.582 27.946 33.618 ;
      RECT 27.894 37.902 27.946 37.938 ;
      RECT 27.894 38.142 27.946 38.178 ;
      RECT 27.894 40.678 27.946 40.714 ;
      RECT 27.894 41.878 27.946 41.914 ;
      RECT 27.894 43.078 27.946 43.114 ;
      RECT 27.894 44.278 27.946 44.314 ;
      RECT 27.894 45.478 27.946 45.514 ;
      RECT 27.894 46.678 27.946 46.714 ;
      RECT 27.894 47.878 27.946 47.914 ;
      RECT 27.894 49.078 27.946 49.114 ;
      RECT 27.894 50.278 27.946 50.314 ;
      RECT 27.894 51.478 27.946 51.514 ;
      RECT 27.894 52.678 27.946 52.714 ;
      RECT 27.894 53.878 27.946 53.914 ;
      RECT 27.894 55.078 27.946 55.114 ;
      RECT 27.894 56.278 27.946 56.314 ;
      RECT 27.894 57.478 27.946 57.514 ;
      RECT 27.894 58.678 27.946 58.714 ;
      RECT 27.894 59.878 27.946 59.914 ;
      RECT 27.894 61.078 27.946 61.114 ;
      RECT 27.894 62.278 27.946 62.314 ;
      RECT 27.894 63.478 27.946 63.514 ;
      RECT 27.894 64.678 27.946 64.714 ;
      RECT 27.894 65.878 27.946 65.914 ;
      RECT 27.894 67.078 27.946 67.114 ;
      RECT 27.894 68.278 27.946 68.314 ;
      RECT 27.894 69.478 27.946 69.514 ;
      RECT 27.894 70.678 27.946 70.714 ;
      RECT 27.894 71.878 27.946 71.914 ;
      RECT 27.974 0.281 28.026 0.317 ;
      RECT 27.974 72.403 28.026 72.439 ;
      RECT 28.054 0.806 28.106 0.842 ;
      RECT 28.054 2.006 28.106 2.042 ;
      RECT 28.054 3.206 28.106 3.242 ;
      RECT 28.054 4.406 28.106 4.442 ;
      RECT 28.054 5.606 28.106 5.642 ;
      RECT 28.054 6.806 28.106 6.842 ;
      RECT 28.054 8.006 28.106 8.042 ;
      RECT 28.054 9.206 28.106 9.242 ;
      RECT 28.054 10.406 28.106 10.442 ;
      RECT 28.054 11.606 28.106 11.642 ;
      RECT 28.054 12.806 28.106 12.842 ;
      RECT 28.054 14.006 28.106 14.042 ;
      RECT 28.054 15.206 28.106 15.242 ;
      RECT 28.054 16.406 28.106 16.442 ;
      RECT 28.054 17.606 28.106 17.642 ;
      RECT 28.054 18.806 28.106 18.842 ;
      RECT 28.054 20.006 28.106 20.042 ;
      RECT 28.054 21.206 28.106 21.242 ;
      RECT 28.054 22.406 28.106 22.442 ;
      RECT 28.054 23.606 28.106 23.642 ;
      RECT 28.054 24.806 28.106 24.842 ;
      RECT 28.054 26.006 28.106 26.042 ;
      RECT 28.054 27.206 28.106 27.242 ;
      RECT 28.054 28.406 28.106 28.442 ;
      RECT 28.054 29.606 28.106 29.642 ;
      RECT 28.054 30.806 28.106 30.842 ;
      RECT 28.054 32.622 28.106 32.658 ;
      RECT 28.054 32.862 28.106 32.898 ;
      RECT 28.054 34.302 28.106 34.338 ;
      RECT 28.054 34.782 28.106 34.818 ;
      RECT 28.054 36.702 28.106 36.738 ;
      RECT 28.054 37.182 28.106 37.218 ;
      RECT 28.054 38.622 28.106 38.658 ;
      RECT 28.054 38.862 28.106 38.898 ;
      RECT 28.054 39.926 28.106 39.962 ;
      RECT 28.054 41.126 28.106 41.162 ;
      RECT 28.054 42.326 28.106 42.362 ;
      RECT 28.054 43.526 28.106 43.562 ;
      RECT 28.054 44.726 28.106 44.762 ;
      RECT 28.054 45.926 28.106 45.962 ;
      RECT 28.054 47.126 28.106 47.162 ;
      RECT 28.054 48.326 28.106 48.362 ;
      RECT 28.054 49.526 28.106 49.562 ;
      RECT 28.054 50.726 28.106 50.762 ;
      RECT 28.054 51.926 28.106 51.962 ;
      RECT 28.054 53.126 28.106 53.162 ;
      RECT 28.054 54.326 28.106 54.362 ;
      RECT 28.054 55.526 28.106 55.562 ;
      RECT 28.054 56.726 28.106 56.762 ;
      RECT 28.054 57.926 28.106 57.962 ;
      RECT 28.054 59.126 28.106 59.162 ;
      RECT 28.054 60.326 28.106 60.362 ;
      RECT 28.054 61.526 28.106 61.562 ;
      RECT 28.054 62.726 28.106 62.762 ;
      RECT 28.054 63.926 28.106 63.962 ;
      RECT 28.054 65.126 28.106 65.162 ;
      RECT 28.054 66.326 28.106 66.362 ;
      RECT 28.054 67.526 28.106 67.562 ;
      RECT 28.054 68.726 28.106 68.762 ;
      RECT 28.054 69.926 28.106 69.962 ;
      RECT 28.054 71.126 28.106 71.162 ;
      RECT 28.134 1.558 28.186 1.594 ;
      RECT 28.134 2.758 28.186 2.794 ;
      RECT 28.134 3.958 28.186 3.994 ;
      RECT 28.134 5.158 28.186 5.194 ;
      RECT 28.134 6.358 28.186 6.394 ;
      RECT 28.134 7.558 28.186 7.594 ;
      RECT 28.134 8.758 28.186 8.794 ;
      RECT 28.134 9.958 28.186 9.994 ;
      RECT 28.134 11.158 28.186 11.194 ;
      RECT 28.134 12.358 28.186 12.394 ;
      RECT 28.134 13.558 28.186 13.594 ;
      RECT 28.134 14.758 28.186 14.794 ;
      RECT 28.134 15.958 28.186 15.994 ;
      RECT 28.134 17.158 28.186 17.194 ;
      RECT 28.134 18.358 28.186 18.394 ;
      RECT 28.134 19.558 28.186 19.594 ;
      RECT 28.134 20.758 28.186 20.794 ;
      RECT 28.134 21.958 28.186 21.994 ;
      RECT 28.134 23.158 28.186 23.194 ;
      RECT 28.134 24.358 28.186 24.394 ;
      RECT 28.134 25.558 28.186 25.594 ;
      RECT 28.134 26.758 28.186 26.794 ;
      RECT 28.134 27.958 28.186 27.994 ;
      RECT 28.134 29.158 28.186 29.194 ;
      RECT 28.134 30.358 28.186 30.394 ;
      RECT 28.134 31.558 28.186 31.594 ;
      RECT 28.134 33.342 28.186 33.378 ;
      RECT 28.134 33.582 28.186 33.618 ;
      RECT 28.134 37.902 28.186 37.938 ;
      RECT 28.134 38.142 28.186 38.178 ;
      RECT 28.134 40.678 28.186 40.714 ;
      RECT 28.134 41.878 28.186 41.914 ;
      RECT 28.134 43.078 28.186 43.114 ;
      RECT 28.134 44.278 28.186 44.314 ;
      RECT 28.134 45.478 28.186 45.514 ;
      RECT 28.134 46.678 28.186 46.714 ;
      RECT 28.134 47.878 28.186 47.914 ;
      RECT 28.134 49.078 28.186 49.114 ;
      RECT 28.134 50.278 28.186 50.314 ;
      RECT 28.134 51.478 28.186 51.514 ;
      RECT 28.134 52.678 28.186 52.714 ;
      RECT 28.134 53.878 28.186 53.914 ;
      RECT 28.134 55.078 28.186 55.114 ;
      RECT 28.134 56.278 28.186 56.314 ;
      RECT 28.134 57.478 28.186 57.514 ;
      RECT 28.134 58.678 28.186 58.714 ;
      RECT 28.134 59.878 28.186 59.914 ;
      RECT 28.134 61.078 28.186 61.114 ;
      RECT 28.134 62.278 28.186 62.314 ;
      RECT 28.134 63.478 28.186 63.514 ;
      RECT 28.134 64.678 28.186 64.714 ;
      RECT 28.134 65.878 28.186 65.914 ;
      RECT 28.134 67.078 28.186 67.114 ;
      RECT 28.134 68.278 28.186 68.314 ;
      RECT 28.134 69.478 28.186 69.514 ;
      RECT 28.134 70.678 28.186 70.714 ;
      RECT 28.134 71.878 28.186 71.914 ;
      RECT 28.214 0.806 28.266 0.842 ;
      RECT 28.214 2.006 28.266 2.042 ;
      RECT 28.214 3.206 28.266 3.242 ;
      RECT 28.214 4.406 28.266 4.442 ;
      RECT 28.214 5.606 28.266 5.642 ;
      RECT 28.214 6.806 28.266 6.842 ;
      RECT 28.214 8.006 28.266 8.042 ;
      RECT 28.214 9.206 28.266 9.242 ;
      RECT 28.214 10.406 28.266 10.442 ;
      RECT 28.214 11.606 28.266 11.642 ;
      RECT 28.214 12.806 28.266 12.842 ;
      RECT 28.214 14.006 28.266 14.042 ;
      RECT 28.214 15.206 28.266 15.242 ;
      RECT 28.214 16.406 28.266 16.442 ;
      RECT 28.214 17.606 28.266 17.642 ;
      RECT 28.214 18.806 28.266 18.842 ;
      RECT 28.214 20.006 28.266 20.042 ;
      RECT 28.214 21.206 28.266 21.242 ;
      RECT 28.214 22.406 28.266 22.442 ;
      RECT 28.214 23.606 28.266 23.642 ;
      RECT 28.214 24.806 28.266 24.842 ;
      RECT 28.214 26.006 28.266 26.042 ;
      RECT 28.214 27.206 28.266 27.242 ;
      RECT 28.214 28.406 28.266 28.442 ;
      RECT 28.214 29.606 28.266 29.642 ;
      RECT 28.214 30.806 28.266 30.842 ;
      RECT 28.214 32.622 28.266 32.658 ;
      RECT 28.214 32.862 28.266 32.898 ;
      RECT 28.214 38.622 28.266 38.658 ;
      RECT 28.214 38.862 28.266 38.898 ;
      RECT 28.214 39.926 28.266 39.962 ;
      RECT 28.214 41.126 28.266 41.162 ;
      RECT 28.214 42.326 28.266 42.362 ;
      RECT 28.214 43.526 28.266 43.562 ;
      RECT 28.214 44.726 28.266 44.762 ;
      RECT 28.214 45.926 28.266 45.962 ;
      RECT 28.214 47.126 28.266 47.162 ;
      RECT 28.214 48.326 28.266 48.362 ;
      RECT 28.214 49.526 28.266 49.562 ;
      RECT 28.214 50.726 28.266 50.762 ;
      RECT 28.214 51.926 28.266 51.962 ;
      RECT 28.214 53.126 28.266 53.162 ;
      RECT 28.214 54.326 28.266 54.362 ;
      RECT 28.214 55.526 28.266 55.562 ;
      RECT 28.214 56.726 28.266 56.762 ;
      RECT 28.214 57.926 28.266 57.962 ;
      RECT 28.214 59.126 28.266 59.162 ;
      RECT 28.214 60.326 28.266 60.362 ;
      RECT 28.214 61.526 28.266 61.562 ;
      RECT 28.214 62.726 28.266 62.762 ;
      RECT 28.214 63.926 28.266 63.962 ;
      RECT 28.214 65.126 28.266 65.162 ;
      RECT 28.214 66.326 28.266 66.362 ;
      RECT 28.214 67.526 28.266 67.562 ;
      RECT 28.214 68.726 28.266 68.762 ;
      RECT 28.214 69.926 28.266 69.962 ;
      RECT 28.214 71.126 28.266 71.162 ;
      RECT 28.294 1.558 28.346 1.594 ;
      RECT 28.294 2.758 28.346 2.794 ;
      RECT 28.294 3.958 28.346 3.994 ;
      RECT 28.294 5.158 28.346 5.194 ;
      RECT 28.294 6.358 28.346 6.394 ;
      RECT 28.294 7.558 28.346 7.594 ;
      RECT 28.294 8.758 28.346 8.794 ;
      RECT 28.294 9.958 28.346 9.994 ;
      RECT 28.294 11.158 28.346 11.194 ;
      RECT 28.294 12.358 28.346 12.394 ;
      RECT 28.294 13.558 28.346 13.594 ;
      RECT 28.294 14.758 28.346 14.794 ;
      RECT 28.294 15.958 28.346 15.994 ;
      RECT 28.294 17.158 28.346 17.194 ;
      RECT 28.294 18.358 28.346 18.394 ;
      RECT 28.294 19.558 28.346 19.594 ;
      RECT 28.294 20.758 28.346 20.794 ;
      RECT 28.294 21.958 28.346 21.994 ;
      RECT 28.294 23.158 28.346 23.194 ;
      RECT 28.294 24.358 28.346 24.394 ;
      RECT 28.294 25.558 28.346 25.594 ;
      RECT 28.294 26.758 28.346 26.794 ;
      RECT 28.294 27.958 28.346 27.994 ;
      RECT 28.294 29.158 28.346 29.194 ;
      RECT 28.294 30.358 28.346 30.394 ;
      RECT 28.294 31.558 28.346 31.594 ;
      RECT 28.294 33.342 28.346 33.378 ;
      RECT 28.294 33.582 28.346 33.618 ;
      RECT 28.294 37.902 28.346 37.938 ;
      RECT 28.294 38.142 28.346 38.178 ;
      RECT 28.294 40.678 28.346 40.714 ;
      RECT 28.294 41.878 28.346 41.914 ;
      RECT 28.294 43.078 28.346 43.114 ;
      RECT 28.294 44.278 28.346 44.314 ;
      RECT 28.294 45.478 28.346 45.514 ;
      RECT 28.294 46.678 28.346 46.714 ;
      RECT 28.294 47.878 28.346 47.914 ;
      RECT 28.294 49.078 28.346 49.114 ;
      RECT 28.294 50.278 28.346 50.314 ;
      RECT 28.294 51.478 28.346 51.514 ;
      RECT 28.294 52.678 28.346 52.714 ;
      RECT 28.294 53.878 28.346 53.914 ;
      RECT 28.294 55.078 28.346 55.114 ;
      RECT 28.294 56.278 28.346 56.314 ;
      RECT 28.294 57.478 28.346 57.514 ;
      RECT 28.294 58.678 28.346 58.714 ;
      RECT 28.294 59.878 28.346 59.914 ;
      RECT 28.294 61.078 28.346 61.114 ;
      RECT 28.294 62.278 28.346 62.314 ;
      RECT 28.294 63.478 28.346 63.514 ;
      RECT 28.294 64.678 28.346 64.714 ;
      RECT 28.294 65.878 28.346 65.914 ;
      RECT 28.294 67.078 28.346 67.114 ;
      RECT 28.294 68.278 28.346 68.314 ;
      RECT 28.294 69.478 28.346 69.514 ;
      RECT 28.294 70.678 28.346 70.714 ;
      RECT 28.294 71.878 28.346 71.914 ;
      RECT 28.374 0.281 28.426 0.317 ;
      RECT 28.374 72.403 28.426 72.439 ;
      RECT 28.454 0.806 28.506 0.842 ;
      RECT 28.454 2.006 28.506 2.042 ;
      RECT 28.454 3.206 28.506 3.242 ;
      RECT 28.454 4.406 28.506 4.442 ;
      RECT 28.454 5.606 28.506 5.642 ;
      RECT 28.454 6.806 28.506 6.842 ;
      RECT 28.454 8.006 28.506 8.042 ;
      RECT 28.454 9.206 28.506 9.242 ;
      RECT 28.454 10.406 28.506 10.442 ;
      RECT 28.454 11.606 28.506 11.642 ;
      RECT 28.454 12.806 28.506 12.842 ;
      RECT 28.454 14.006 28.506 14.042 ;
      RECT 28.454 15.206 28.506 15.242 ;
      RECT 28.454 16.406 28.506 16.442 ;
      RECT 28.454 17.606 28.506 17.642 ;
      RECT 28.454 18.806 28.506 18.842 ;
      RECT 28.454 20.006 28.506 20.042 ;
      RECT 28.454 21.206 28.506 21.242 ;
      RECT 28.454 22.406 28.506 22.442 ;
      RECT 28.454 23.606 28.506 23.642 ;
      RECT 28.454 24.806 28.506 24.842 ;
      RECT 28.454 26.006 28.506 26.042 ;
      RECT 28.454 27.206 28.506 27.242 ;
      RECT 28.454 28.406 28.506 28.442 ;
      RECT 28.454 29.606 28.506 29.642 ;
      RECT 28.454 30.806 28.506 30.842 ;
      RECT 28.454 32.622 28.506 32.658 ;
      RECT 28.454 32.862 28.506 32.898 ;
      RECT 28.454 38.622 28.506 38.658 ;
      RECT 28.454 38.862 28.506 38.898 ;
      RECT 28.454 39.926 28.506 39.962 ;
      RECT 28.454 41.126 28.506 41.162 ;
      RECT 28.454 42.326 28.506 42.362 ;
      RECT 28.454 43.526 28.506 43.562 ;
      RECT 28.454 44.726 28.506 44.762 ;
      RECT 28.454 45.926 28.506 45.962 ;
      RECT 28.454 47.126 28.506 47.162 ;
      RECT 28.454 48.326 28.506 48.362 ;
      RECT 28.454 49.526 28.506 49.562 ;
      RECT 28.454 50.726 28.506 50.762 ;
      RECT 28.454 51.926 28.506 51.962 ;
      RECT 28.454 53.126 28.506 53.162 ;
      RECT 28.454 54.326 28.506 54.362 ;
      RECT 28.454 55.526 28.506 55.562 ;
      RECT 28.454 56.726 28.506 56.762 ;
      RECT 28.454 57.926 28.506 57.962 ;
      RECT 28.454 59.126 28.506 59.162 ;
      RECT 28.454 60.326 28.506 60.362 ;
      RECT 28.454 61.526 28.506 61.562 ;
      RECT 28.454 62.726 28.506 62.762 ;
      RECT 28.454 63.926 28.506 63.962 ;
      RECT 28.454 65.126 28.506 65.162 ;
      RECT 28.454 66.326 28.506 66.362 ;
      RECT 28.454 67.526 28.506 67.562 ;
      RECT 28.454 68.726 28.506 68.762 ;
      RECT 28.454 69.926 28.506 69.962 ;
      RECT 28.454 71.126 28.506 71.162 ;
      RECT 28.534 1.558 28.586 1.594 ;
      RECT 28.534 2.758 28.586 2.794 ;
      RECT 28.534 3.958 28.586 3.994 ;
      RECT 28.534 5.158 28.586 5.194 ;
      RECT 28.534 6.358 28.586 6.394 ;
      RECT 28.534 7.558 28.586 7.594 ;
      RECT 28.534 8.758 28.586 8.794 ;
      RECT 28.534 9.958 28.586 9.994 ;
      RECT 28.534 11.158 28.586 11.194 ;
      RECT 28.534 12.358 28.586 12.394 ;
      RECT 28.534 13.558 28.586 13.594 ;
      RECT 28.534 14.758 28.586 14.794 ;
      RECT 28.534 15.958 28.586 15.994 ;
      RECT 28.534 17.158 28.586 17.194 ;
      RECT 28.534 18.358 28.586 18.394 ;
      RECT 28.534 19.558 28.586 19.594 ;
      RECT 28.534 20.758 28.586 20.794 ;
      RECT 28.534 21.958 28.586 21.994 ;
      RECT 28.534 23.158 28.586 23.194 ;
      RECT 28.534 24.358 28.586 24.394 ;
      RECT 28.534 25.558 28.586 25.594 ;
      RECT 28.534 26.758 28.586 26.794 ;
      RECT 28.534 27.958 28.586 27.994 ;
      RECT 28.534 29.158 28.586 29.194 ;
      RECT 28.534 30.358 28.586 30.394 ;
      RECT 28.534 31.558 28.586 31.594 ;
      RECT 28.534 33.342 28.586 33.378 ;
      RECT 28.534 33.582 28.586 33.618 ;
      RECT 28.534 37.902 28.586 37.938 ;
      RECT 28.534 38.142 28.586 38.178 ;
      RECT 28.534 40.678 28.586 40.714 ;
      RECT 28.534 41.878 28.586 41.914 ;
      RECT 28.534 43.078 28.586 43.114 ;
      RECT 28.534 44.278 28.586 44.314 ;
      RECT 28.534 45.478 28.586 45.514 ;
      RECT 28.534 46.678 28.586 46.714 ;
      RECT 28.534 47.878 28.586 47.914 ;
      RECT 28.534 49.078 28.586 49.114 ;
      RECT 28.534 50.278 28.586 50.314 ;
      RECT 28.534 51.478 28.586 51.514 ;
      RECT 28.534 52.678 28.586 52.714 ;
      RECT 28.534 53.878 28.586 53.914 ;
      RECT 28.534 55.078 28.586 55.114 ;
      RECT 28.534 56.278 28.586 56.314 ;
      RECT 28.534 57.478 28.586 57.514 ;
      RECT 28.534 58.678 28.586 58.714 ;
      RECT 28.534 59.878 28.586 59.914 ;
      RECT 28.534 61.078 28.586 61.114 ;
      RECT 28.534 62.278 28.586 62.314 ;
      RECT 28.534 63.478 28.586 63.514 ;
      RECT 28.534 64.678 28.586 64.714 ;
      RECT 28.534 65.878 28.586 65.914 ;
      RECT 28.534 67.078 28.586 67.114 ;
      RECT 28.534 68.278 28.586 68.314 ;
      RECT 28.534 69.478 28.586 69.514 ;
      RECT 28.534 70.678 28.586 70.714 ;
      RECT 28.534 71.878 28.586 71.914 ;
      RECT 28.614 0.806 28.666 0.842 ;
      RECT 28.614 2.006 28.666 2.042 ;
      RECT 28.614 3.206 28.666 3.242 ;
      RECT 28.614 4.406 28.666 4.442 ;
      RECT 28.614 5.606 28.666 5.642 ;
      RECT 28.614 6.806 28.666 6.842 ;
      RECT 28.614 8.006 28.666 8.042 ;
      RECT 28.614 9.206 28.666 9.242 ;
      RECT 28.614 10.406 28.666 10.442 ;
      RECT 28.614 11.606 28.666 11.642 ;
      RECT 28.614 12.806 28.666 12.842 ;
      RECT 28.614 14.006 28.666 14.042 ;
      RECT 28.614 15.206 28.666 15.242 ;
      RECT 28.614 16.406 28.666 16.442 ;
      RECT 28.614 17.606 28.666 17.642 ;
      RECT 28.614 18.806 28.666 18.842 ;
      RECT 28.614 20.006 28.666 20.042 ;
      RECT 28.614 21.206 28.666 21.242 ;
      RECT 28.614 22.406 28.666 22.442 ;
      RECT 28.614 23.606 28.666 23.642 ;
      RECT 28.614 24.806 28.666 24.842 ;
      RECT 28.614 26.006 28.666 26.042 ;
      RECT 28.614 27.206 28.666 27.242 ;
      RECT 28.614 28.406 28.666 28.442 ;
      RECT 28.614 29.606 28.666 29.642 ;
      RECT 28.614 30.806 28.666 30.842 ;
      RECT 28.614 32.622 28.666 32.658 ;
      RECT 28.614 32.862 28.666 32.898 ;
      RECT 28.614 38.622 28.666 38.658 ;
      RECT 28.614 38.862 28.666 38.898 ;
      RECT 28.614 39.926 28.666 39.962 ;
      RECT 28.614 41.126 28.666 41.162 ;
      RECT 28.614 42.326 28.666 42.362 ;
      RECT 28.614 43.526 28.666 43.562 ;
      RECT 28.614 44.726 28.666 44.762 ;
      RECT 28.614 45.926 28.666 45.962 ;
      RECT 28.614 47.126 28.666 47.162 ;
      RECT 28.614 48.326 28.666 48.362 ;
      RECT 28.614 49.526 28.666 49.562 ;
      RECT 28.614 50.726 28.666 50.762 ;
      RECT 28.614 51.926 28.666 51.962 ;
      RECT 28.614 53.126 28.666 53.162 ;
      RECT 28.614 54.326 28.666 54.362 ;
      RECT 28.614 55.526 28.666 55.562 ;
      RECT 28.614 56.726 28.666 56.762 ;
      RECT 28.614 57.926 28.666 57.962 ;
      RECT 28.614 59.126 28.666 59.162 ;
      RECT 28.614 60.326 28.666 60.362 ;
      RECT 28.614 61.526 28.666 61.562 ;
      RECT 28.614 62.726 28.666 62.762 ;
      RECT 28.614 63.926 28.666 63.962 ;
      RECT 28.614 65.126 28.666 65.162 ;
      RECT 28.614 66.326 28.666 66.362 ;
      RECT 28.614 67.526 28.666 67.562 ;
      RECT 28.614 68.726 28.666 68.762 ;
      RECT 28.614 69.926 28.666 69.962 ;
      RECT 28.614 71.126 28.666 71.162 ;
      RECT 28.694 1.558 28.746 1.594 ;
      RECT 28.694 2.758 28.746 2.794 ;
      RECT 28.694 3.958 28.746 3.994 ;
      RECT 28.694 5.158 28.746 5.194 ;
      RECT 28.694 6.358 28.746 6.394 ;
      RECT 28.694 7.558 28.746 7.594 ;
      RECT 28.694 8.758 28.746 8.794 ;
      RECT 28.694 9.958 28.746 9.994 ;
      RECT 28.694 11.158 28.746 11.194 ;
      RECT 28.694 12.358 28.746 12.394 ;
      RECT 28.694 13.558 28.746 13.594 ;
      RECT 28.694 14.758 28.746 14.794 ;
      RECT 28.694 15.958 28.746 15.994 ;
      RECT 28.694 17.158 28.746 17.194 ;
      RECT 28.694 18.358 28.746 18.394 ;
      RECT 28.694 19.558 28.746 19.594 ;
      RECT 28.694 20.758 28.746 20.794 ;
      RECT 28.694 21.958 28.746 21.994 ;
      RECT 28.694 23.158 28.746 23.194 ;
      RECT 28.694 24.358 28.746 24.394 ;
      RECT 28.694 25.558 28.746 25.594 ;
      RECT 28.694 26.758 28.746 26.794 ;
      RECT 28.694 27.958 28.746 27.994 ;
      RECT 28.694 29.158 28.746 29.194 ;
      RECT 28.694 30.358 28.746 30.394 ;
      RECT 28.694 31.558 28.746 31.594 ;
      RECT 28.694 33.342 28.746 33.378 ;
      RECT 28.694 33.582 28.746 33.618 ;
      RECT 28.694 37.902 28.746 37.938 ;
      RECT 28.694 38.142 28.746 38.178 ;
      RECT 28.694 40.678 28.746 40.714 ;
      RECT 28.694 41.878 28.746 41.914 ;
      RECT 28.694 43.078 28.746 43.114 ;
      RECT 28.694 44.278 28.746 44.314 ;
      RECT 28.694 45.478 28.746 45.514 ;
      RECT 28.694 46.678 28.746 46.714 ;
      RECT 28.694 47.878 28.746 47.914 ;
      RECT 28.694 49.078 28.746 49.114 ;
      RECT 28.694 50.278 28.746 50.314 ;
      RECT 28.694 51.478 28.746 51.514 ;
      RECT 28.694 52.678 28.746 52.714 ;
      RECT 28.694 53.878 28.746 53.914 ;
      RECT 28.694 55.078 28.746 55.114 ;
      RECT 28.694 56.278 28.746 56.314 ;
      RECT 28.694 57.478 28.746 57.514 ;
      RECT 28.694 58.678 28.746 58.714 ;
      RECT 28.694 59.878 28.746 59.914 ;
      RECT 28.694 61.078 28.746 61.114 ;
      RECT 28.694 62.278 28.746 62.314 ;
      RECT 28.694 63.478 28.746 63.514 ;
      RECT 28.694 64.678 28.746 64.714 ;
      RECT 28.694 65.878 28.746 65.914 ;
      RECT 28.694 67.078 28.746 67.114 ;
      RECT 28.694 68.278 28.746 68.314 ;
      RECT 28.694 69.478 28.746 69.514 ;
      RECT 28.694 70.678 28.746 70.714 ;
      RECT 28.694 71.878 28.746 71.914 ;
      RECT 28.774 0.281 28.826 0.317 ;
      RECT 28.774 72.403 28.826 72.439 ;
      RECT 28.854 0.806 28.906 0.842 ;
      RECT 28.854 2.006 28.906 2.042 ;
      RECT 28.854 3.206 28.906 3.242 ;
      RECT 28.854 4.406 28.906 4.442 ;
      RECT 28.854 5.606 28.906 5.642 ;
      RECT 28.854 6.806 28.906 6.842 ;
      RECT 28.854 8.006 28.906 8.042 ;
      RECT 28.854 9.206 28.906 9.242 ;
      RECT 28.854 10.406 28.906 10.442 ;
      RECT 28.854 11.606 28.906 11.642 ;
      RECT 28.854 12.806 28.906 12.842 ;
      RECT 28.854 14.006 28.906 14.042 ;
      RECT 28.854 15.206 28.906 15.242 ;
      RECT 28.854 16.406 28.906 16.442 ;
      RECT 28.854 17.606 28.906 17.642 ;
      RECT 28.854 18.806 28.906 18.842 ;
      RECT 28.854 20.006 28.906 20.042 ;
      RECT 28.854 21.206 28.906 21.242 ;
      RECT 28.854 22.406 28.906 22.442 ;
      RECT 28.854 23.606 28.906 23.642 ;
      RECT 28.854 24.806 28.906 24.842 ;
      RECT 28.854 26.006 28.906 26.042 ;
      RECT 28.854 27.206 28.906 27.242 ;
      RECT 28.854 28.406 28.906 28.442 ;
      RECT 28.854 29.606 28.906 29.642 ;
      RECT 28.854 30.806 28.906 30.842 ;
      RECT 28.854 32.622 28.906 32.658 ;
      RECT 28.854 32.862 28.906 32.898 ;
      RECT 28.854 34.302 28.906 34.338 ;
      RECT 28.854 34.782 28.906 34.818 ;
      RECT 28.854 36.702 28.906 36.738 ;
      RECT 28.854 37.182 28.906 37.218 ;
      RECT 28.854 38.622 28.906 38.658 ;
      RECT 28.854 38.862 28.906 38.898 ;
      RECT 28.854 39.926 28.906 39.962 ;
      RECT 28.854 41.126 28.906 41.162 ;
      RECT 28.854 42.326 28.906 42.362 ;
      RECT 28.854 43.526 28.906 43.562 ;
      RECT 28.854 44.726 28.906 44.762 ;
      RECT 28.854 45.926 28.906 45.962 ;
      RECT 28.854 47.126 28.906 47.162 ;
      RECT 28.854 48.326 28.906 48.362 ;
      RECT 28.854 49.526 28.906 49.562 ;
      RECT 28.854 50.726 28.906 50.762 ;
      RECT 28.854 51.926 28.906 51.962 ;
      RECT 28.854 53.126 28.906 53.162 ;
      RECT 28.854 54.326 28.906 54.362 ;
      RECT 28.854 55.526 28.906 55.562 ;
      RECT 28.854 56.726 28.906 56.762 ;
      RECT 28.854 57.926 28.906 57.962 ;
      RECT 28.854 59.126 28.906 59.162 ;
      RECT 28.854 60.326 28.906 60.362 ;
      RECT 28.854 61.526 28.906 61.562 ;
      RECT 28.854 62.726 28.906 62.762 ;
      RECT 28.854 63.926 28.906 63.962 ;
      RECT 28.854 65.126 28.906 65.162 ;
      RECT 28.854 66.326 28.906 66.362 ;
      RECT 28.854 67.526 28.906 67.562 ;
      RECT 28.854 68.726 28.906 68.762 ;
      RECT 28.854 69.926 28.906 69.962 ;
      RECT 28.854 71.126 28.906 71.162 ;
      RECT 28.934 1.558 28.986 1.594 ;
      RECT 28.934 2.758 28.986 2.794 ;
      RECT 28.934 3.958 28.986 3.994 ;
      RECT 28.934 5.158 28.986 5.194 ;
      RECT 28.934 6.358 28.986 6.394 ;
      RECT 28.934 7.558 28.986 7.594 ;
      RECT 28.934 8.758 28.986 8.794 ;
      RECT 28.934 9.958 28.986 9.994 ;
      RECT 28.934 11.158 28.986 11.194 ;
      RECT 28.934 12.358 28.986 12.394 ;
      RECT 28.934 13.558 28.986 13.594 ;
      RECT 28.934 14.758 28.986 14.794 ;
      RECT 28.934 15.958 28.986 15.994 ;
      RECT 28.934 17.158 28.986 17.194 ;
      RECT 28.934 18.358 28.986 18.394 ;
      RECT 28.934 19.558 28.986 19.594 ;
      RECT 28.934 20.758 28.986 20.794 ;
      RECT 28.934 21.958 28.986 21.994 ;
      RECT 28.934 23.158 28.986 23.194 ;
      RECT 28.934 24.358 28.986 24.394 ;
      RECT 28.934 25.558 28.986 25.594 ;
      RECT 28.934 26.758 28.986 26.794 ;
      RECT 28.934 27.958 28.986 27.994 ;
      RECT 28.934 29.158 28.986 29.194 ;
      RECT 28.934 30.358 28.986 30.394 ;
      RECT 28.934 31.558 28.986 31.594 ;
      RECT 28.934 33.342 28.986 33.378 ;
      RECT 28.934 33.582 28.986 33.618 ;
      RECT 28.934 37.902 28.986 37.938 ;
      RECT 28.934 38.142 28.986 38.178 ;
      RECT 28.934 40.678 28.986 40.714 ;
      RECT 28.934 41.878 28.986 41.914 ;
      RECT 28.934 43.078 28.986 43.114 ;
      RECT 28.934 44.278 28.986 44.314 ;
      RECT 28.934 45.478 28.986 45.514 ;
      RECT 28.934 46.678 28.986 46.714 ;
      RECT 28.934 47.878 28.986 47.914 ;
      RECT 28.934 49.078 28.986 49.114 ;
      RECT 28.934 50.278 28.986 50.314 ;
      RECT 28.934 51.478 28.986 51.514 ;
      RECT 28.934 52.678 28.986 52.714 ;
      RECT 28.934 53.878 28.986 53.914 ;
      RECT 28.934 55.078 28.986 55.114 ;
      RECT 28.934 56.278 28.986 56.314 ;
      RECT 28.934 57.478 28.986 57.514 ;
      RECT 28.934 58.678 28.986 58.714 ;
      RECT 28.934 59.878 28.986 59.914 ;
      RECT 28.934 61.078 28.986 61.114 ;
      RECT 28.934 62.278 28.986 62.314 ;
      RECT 28.934 63.478 28.986 63.514 ;
      RECT 28.934 64.678 28.986 64.714 ;
      RECT 28.934 65.878 28.986 65.914 ;
      RECT 28.934 67.078 28.986 67.114 ;
      RECT 28.934 68.278 28.986 68.314 ;
      RECT 28.934 69.478 28.986 69.514 ;
      RECT 28.934 70.678 28.986 70.714 ;
      RECT 28.934 71.878 28.986 71.914 ;
      RECT 29.014 0.806 29.066 0.842 ;
      RECT 29.014 2.006 29.066 2.042 ;
      RECT 29.014 3.206 29.066 3.242 ;
      RECT 29.014 4.406 29.066 4.442 ;
      RECT 29.014 5.606 29.066 5.642 ;
      RECT 29.014 6.806 29.066 6.842 ;
      RECT 29.014 8.006 29.066 8.042 ;
      RECT 29.014 9.206 29.066 9.242 ;
      RECT 29.014 10.406 29.066 10.442 ;
      RECT 29.014 11.606 29.066 11.642 ;
      RECT 29.014 12.806 29.066 12.842 ;
      RECT 29.014 14.006 29.066 14.042 ;
      RECT 29.014 15.206 29.066 15.242 ;
      RECT 29.014 16.406 29.066 16.442 ;
      RECT 29.014 17.606 29.066 17.642 ;
      RECT 29.014 18.806 29.066 18.842 ;
      RECT 29.014 20.006 29.066 20.042 ;
      RECT 29.014 21.206 29.066 21.242 ;
      RECT 29.014 22.406 29.066 22.442 ;
      RECT 29.014 23.606 29.066 23.642 ;
      RECT 29.014 24.806 29.066 24.842 ;
      RECT 29.014 26.006 29.066 26.042 ;
      RECT 29.014 27.206 29.066 27.242 ;
      RECT 29.014 28.406 29.066 28.442 ;
      RECT 29.014 29.606 29.066 29.642 ;
      RECT 29.014 30.806 29.066 30.842 ;
      RECT 29.014 32.622 29.066 32.658 ;
      RECT 29.014 32.862 29.066 32.898 ;
      RECT 29.014 38.622 29.066 38.658 ;
      RECT 29.014 38.862 29.066 38.898 ;
      RECT 29.014 39.926 29.066 39.962 ;
      RECT 29.014 41.126 29.066 41.162 ;
      RECT 29.014 42.326 29.066 42.362 ;
      RECT 29.014 43.526 29.066 43.562 ;
      RECT 29.014 44.726 29.066 44.762 ;
      RECT 29.014 45.926 29.066 45.962 ;
      RECT 29.014 47.126 29.066 47.162 ;
      RECT 29.014 48.326 29.066 48.362 ;
      RECT 29.014 49.526 29.066 49.562 ;
      RECT 29.014 50.726 29.066 50.762 ;
      RECT 29.014 51.926 29.066 51.962 ;
      RECT 29.014 53.126 29.066 53.162 ;
      RECT 29.014 54.326 29.066 54.362 ;
      RECT 29.014 55.526 29.066 55.562 ;
      RECT 29.014 56.726 29.066 56.762 ;
      RECT 29.014 57.926 29.066 57.962 ;
      RECT 29.014 59.126 29.066 59.162 ;
      RECT 29.014 60.326 29.066 60.362 ;
      RECT 29.014 61.526 29.066 61.562 ;
      RECT 29.014 62.726 29.066 62.762 ;
      RECT 29.014 63.926 29.066 63.962 ;
      RECT 29.014 65.126 29.066 65.162 ;
      RECT 29.014 66.326 29.066 66.362 ;
      RECT 29.014 67.526 29.066 67.562 ;
      RECT 29.014 68.726 29.066 68.762 ;
      RECT 29.014 69.926 29.066 69.962 ;
      RECT 29.014 71.126 29.066 71.162 ;
      RECT 29.094 1.558 29.146 1.594 ;
      RECT 29.094 2.758 29.146 2.794 ;
      RECT 29.094 3.958 29.146 3.994 ;
      RECT 29.094 5.158 29.146 5.194 ;
      RECT 29.094 6.358 29.146 6.394 ;
      RECT 29.094 7.558 29.146 7.594 ;
      RECT 29.094 8.758 29.146 8.794 ;
      RECT 29.094 9.958 29.146 9.994 ;
      RECT 29.094 11.158 29.146 11.194 ;
      RECT 29.094 12.358 29.146 12.394 ;
      RECT 29.094 13.558 29.146 13.594 ;
      RECT 29.094 14.758 29.146 14.794 ;
      RECT 29.094 15.958 29.146 15.994 ;
      RECT 29.094 17.158 29.146 17.194 ;
      RECT 29.094 18.358 29.146 18.394 ;
      RECT 29.094 19.558 29.146 19.594 ;
      RECT 29.094 20.758 29.146 20.794 ;
      RECT 29.094 21.958 29.146 21.994 ;
      RECT 29.094 23.158 29.146 23.194 ;
      RECT 29.094 24.358 29.146 24.394 ;
      RECT 29.094 25.558 29.146 25.594 ;
      RECT 29.094 26.758 29.146 26.794 ;
      RECT 29.094 27.958 29.146 27.994 ;
      RECT 29.094 29.158 29.146 29.194 ;
      RECT 29.094 30.358 29.146 30.394 ;
      RECT 29.094 31.558 29.146 31.594 ;
      RECT 29.094 33.342 29.146 33.378 ;
      RECT 29.094 33.582 29.146 33.618 ;
      RECT 29.094 37.902 29.146 37.938 ;
      RECT 29.094 38.142 29.146 38.178 ;
      RECT 29.094 40.678 29.146 40.714 ;
      RECT 29.094 41.878 29.146 41.914 ;
      RECT 29.094 43.078 29.146 43.114 ;
      RECT 29.094 44.278 29.146 44.314 ;
      RECT 29.094 45.478 29.146 45.514 ;
      RECT 29.094 46.678 29.146 46.714 ;
      RECT 29.094 47.878 29.146 47.914 ;
      RECT 29.094 49.078 29.146 49.114 ;
      RECT 29.094 50.278 29.146 50.314 ;
      RECT 29.094 51.478 29.146 51.514 ;
      RECT 29.094 52.678 29.146 52.714 ;
      RECT 29.094 53.878 29.146 53.914 ;
      RECT 29.094 55.078 29.146 55.114 ;
      RECT 29.094 56.278 29.146 56.314 ;
      RECT 29.094 57.478 29.146 57.514 ;
      RECT 29.094 58.678 29.146 58.714 ;
      RECT 29.094 59.878 29.146 59.914 ;
      RECT 29.094 61.078 29.146 61.114 ;
      RECT 29.094 62.278 29.146 62.314 ;
      RECT 29.094 63.478 29.146 63.514 ;
      RECT 29.094 64.678 29.146 64.714 ;
      RECT 29.094 65.878 29.146 65.914 ;
      RECT 29.094 67.078 29.146 67.114 ;
      RECT 29.094 68.278 29.146 68.314 ;
      RECT 29.094 69.478 29.146 69.514 ;
      RECT 29.094 70.678 29.146 70.714 ;
      RECT 29.094 71.878 29.146 71.914 ;
      RECT 29.174 0.281 29.226 0.317 ;
      RECT 29.174 72.403 29.226 72.439 ;
      RECT 29.254 0.806 29.306 0.842 ;
      RECT 29.254 2.006 29.306 2.042 ;
      RECT 29.254 3.206 29.306 3.242 ;
      RECT 29.254 4.406 29.306 4.442 ;
      RECT 29.254 5.606 29.306 5.642 ;
      RECT 29.254 6.806 29.306 6.842 ;
      RECT 29.254 8.006 29.306 8.042 ;
      RECT 29.254 9.206 29.306 9.242 ;
      RECT 29.254 10.406 29.306 10.442 ;
      RECT 29.254 11.606 29.306 11.642 ;
      RECT 29.254 12.806 29.306 12.842 ;
      RECT 29.254 14.006 29.306 14.042 ;
      RECT 29.254 15.206 29.306 15.242 ;
      RECT 29.254 16.406 29.306 16.442 ;
      RECT 29.254 17.606 29.306 17.642 ;
      RECT 29.254 18.806 29.306 18.842 ;
      RECT 29.254 20.006 29.306 20.042 ;
      RECT 29.254 21.206 29.306 21.242 ;
      RECT 29.254 22.406 29.306 22.442 ;
      RECT 29.254 23.606 29.306 23.642 ;
      RECT 29.254 24.806 29.306 24.842 ;
      RECT 29.254 26.006 29.306 26.042 ;
      RECT 29.254 27.206 29.306 27.242 ;
      RECT 29.254 28.406 29.306 28.442 ;
      RECT 29.254 29.606 29.306 29.642 ;
      RECT 29.254 30.806 29.306 30.842 ;
      RECT 29.254 32.622 29.306 32.658 ;
      RECT 29.254 32.862 29.306 32.898 ;
      RECT 29.254 38.622 29.306 38.658 ;
      RECT 29.254 38.862 29.306 38.898 ;
      RECT 29.254 39.926 29.306 39.962 ;
      RECT 29.254 41.126 29.306 41.162 ;
      RECT 29.254 42.326 29.306 42.362 ;
      RECT 29.254 43.526 29.306 43.562 ;
      RECT 29.254 44.726 29.306 44.762 ;
      RECT 29.254 45.926 29.306 45.962 ;
      RECT 29.254 47.126 29.306 47.162 ;
      RECT 29.254 48.326 29.306 48.362 ;
      RECT 29.254 49.526 29.306 49.562 ;
      RECT 29.254 50.726 29.306 50.762 ;
      RECT 29.254 51.926 29.306 51.962 ;
      RECT 29.254 53.126 29.306 53.162 ;
      RECT 29.254 54.326 29.306 54.362 ;
      RECT 29.254 55.526 29.306 55.562 ;
      RECT 29.254 56.726 29.306 56.762 ;
      RECT 29.254 57.926 29.306 57.962 ;
      RECT 29.254 59.126 29.306 59.162 ;
      RECT 29.254 60.326 29.306 60.362 ;
      RECT 29.254 61.526 29.306 61.562 ;
      RECT 29.254 62.726 29.306 62.762 ;
      RECT 29.254 63.926 29.306 63.962 ;
      RECT 29.254 65.126 29.306 65.162 ;
      RECT 29.254 66.326 29.306 66.362 ;
      RECT 29.254 67.526 29.306 67.562 ;
      RECT 29.254 68.726 29.306 68.762 ;
      RECT 29.254 69.926 29.306 69.962 ;
      RECT 29.254 71.126 29.306 71.162 ;
      RECT 29.334 1.558 29.386 1.594 ;
      RECT 29.334 2.758 29.386 2.794 ;
      RECT 29.334 3.958 29.386 3.994 ;
      RECT 29.334 5.158 29.386 5.194 ;
      RECT 29.334 6.358 29.386 6.394 ;
      RECT 29.334 7.558 29.386 7.594 ;
      RECT 29.334 8.758 29.386 8.794 ;
      RECT 29.334 9.958 29.386 9.994 ;
      RECT 29.334 11.158 29.386 11.194 ;
      RECT 29.334 12.358 29.386 12.394 ;
      RECT 29.334 13.558 29.386 13.594 ;
      RECT 29.334 14.758 29.386 14.794 ;
      RECT 29.334 15.958 29.386 15.994 ;
      RECT 29.334 17.158 29.386 17.194 ;
      RECT 29.334 18.358 29.386 18.394 ;
      RECT 29.334 19.558 29.386 19.594 ;
      RECT 29.334 20.758 29.386 20.794 ;
      RECT 29.334 21.958 29.386 21.994 ;
      RECT 29.334 23.158 29.386 23.194 ;
      RECT 29.334 24.358 29.386 24.394 ;
      RECT 29.334 25.558 29.386 25.594 ;
      RECT 29.334 26.758 29.386 26.794 ;
      RECT 29.334 27.958 29.386 27.994 ;
      RECT 29.334 29.158 29.386 29.194 ;
      RECT 29.334 30.358 29.386 30.394 ;
      RECT 29.334 31.558 29.386 31.594 ;
      RECT 29.334 33.342 29.386 33.378 ;
      RECT 29.334 33.582 29.386 33.618 ;
      RECT 29.334 37.902 29.386 37.938 ;
      RECT 29.334 38.142 29.386 38.178 ;
      RECT 29.334 40.678 29.386 40.714 ;
      RECT 29.334 41.878 29.386 41.914 ;
      RECT 29.334 43.078 29.386 43.114 ;
      RECT 29.334 44.278 29.386 44.314 ;
      RECT 29.334 45.478 29.386 45.514 ;
      RECT 29.334 46.678 29.386 46.714 ;
      RECT 29.334 47.878 29.386 47.914 ;
      RECT 29.334 49.078 29.386 49.114 ;
      RECT 29.334 50.278 29.386 50.314 ;
      RECT 29.334 51.478 29.386 51.514 ;
      RECT 29.334 52.678 29.386 52.714 ;
      RECT 29.334 53.878 29.386 53.914 ;
      RECT 29.334 55.078 29.386 55.114 ;
      RECT 29.334 56.278 29.386 56.314 ;
      RECT 29.334 57.478 29.386 57.514 ;
      RECT 29.334 58.678 29.386 58.714 ;
      RECT 29.334 59.878 29.386 59.914 ;
      RECT 29.334 61.078 29.386 61.114 ;
      RECT 29.334 62.278 29.386 62.314 ;
      RECT 29.334 63.478 29.386 63.514 ;
      RECT 29.334 64.678 29.386 64.714 ;
      RECT 29.334 65.878 29.386 65.914 ;
      RECT 29.334 67.078 29.386 67.114 ;
      RECT 29.334 68.278 29.386 68.314 ;
      RECT 29.334 69.478 29.386 69.514 ;
      RECT 29.334 70.678 29.386 70.714 ;
      RECT 29.334 71.878 29.386 71.914 ;
      RECT 29.414 0.806 29.466 0.842 ;
      RECT 29.414 2.006 29.466 2.042 ;
      RECT 29.414 3.206 29.466 3.242 ;
      RECT 29.414 4.406 29.466 4.442 ;
      RECT 29.414 5.606 29.466 5.642 ;
      RECT 29.414 6.806 29.466 6.842 ;
      RECT 29.414 8.006 29.466 8.042 ;
      RECT 29.414 9.206 29.466 9.242 ;
      RECT 29.414 10.406 29.466 10.442 ;
      RECT 29.414 11.606 29.466 11.642 ;
      RECT 29.414 12.806 29.466 12.842 ;
      RECT 29.414 14.006 29.466 14.042 ;
      RECT 29.414 15.206 29.466 15.242 ;
      RECT 29.414 16.406 29.466 16.442 ;
      RECT 29.414 17.606 29.466 17.642 ;
      RECT 29.414 18.806 29.466 18.842 ;
      RECT 29.414 20.006 29.466 20.042 ;
      RECT 29.414 21.206 29.466 21.242 ;
      RECT 29.414 22.406 29.466 22.442 ;
      RECT 29.414 23.606 29.466 23.642 ;
      RECT 29.414 24.806 29.466 24.842 ;
      RECT 29.414 26.006 29.466 26.042 ;
      RECT 29.414 27.206 29.466 27.242 ;
      RECT 29.414 28.406 29.466 28.442 ;
      RECT 29.414 29.606 29.466 29.642 ;
      RECT 29.414 30.806 29.466 30.842 ;
      RECT 29.414 32.622 29.466 32.658 ;
      RECT 29.414 32.862 29.466 32.898 ;
      RECT 29.414 38.622 29.466 38.658 ;
      RECT 29.414 38.862 29.466 38.898 ;
      RECT 29.414 39.926 29.466 39.962 ;
      RECT 29.414 41.126 29.466 41.162 ;
      RECT 29.414 42.326 29.466 42.362 ;
      RECT 29.414 43.526 29.466 43.562 ;
      RECT 29.414 44.726 29.466 44.762 ;
      RECT 29.414 45.926 29.466 45.962 ;
      RECT 29.414 47.126 29.466 47.162 ;
      RECT 29.414 48.326 29.466 48.362 ;
      RECT 29.414 49.526 29.466 49.562 ;
      RECT 29.414 50.726 29.466 50.762 ;
      RECT 29.414 51.926 29.466 51.962 ;
      RECT 29.414 53.126 29.466 53.162 ;
      RECT 29.414 54.326 29.466 54.362 ;
      RECT 29.414 55.526 29.466 55.562 ;
      RECT 29.414 56.726 29.466 56.762 ;
      RECT 29.414 57.926 29.466 57.962 ;
      RECT 29.414 59.126 29.466 59.162 ;
      RECT 29.414 60.326 29.466 60.362 ;
      RECT 29.414 61.526 29.466 61.562 ;
      RECT 29.414 62.726 29.466 62.762 ;
      RECT 29.414 63.926 29.466 63.962 ;
      RECT 29.414 65.126 29.466 65.162 ;
      RECT 29.414 66.326 29.466 66.362 ;
      RECT 29.414 67.526 29.466 67.562 ;
      RECT 29.414 68.726 29.466 68.762 ;
      RECT 29.414 69.926 29.466 69.962 ;
      RECT 29.414 71.126 29.466 71.162 ;
      RECT 29.494 1.558 29.546 1.594 ;
      RECT 29.494 2.758 29.546 2.794 ;
      RECT 29.494 3.958 29.546 3.994 ;
      RECT 29.494 5.158 29.546 5.194 ;
      RECT 29.494 6.358 29.546 6.394 ;
      RECT 29.494 7.558 29.546 7.594 ;
      RECT 29.494 8.758 29.546 8.794 ;
      RECT 29.494 9.958 29.546 9.994 ;
      RECT 29.494 11.158 29.546 11.194 ;
      RECT 29.494 12.358 29.546 12.394 ;
      RECT 29.494 13.558 29.546 13.594 ;
      RECT 29.494 14.758 29.546 14.794 ;
      RECT 29.494 15.958 29.546 15.994 ;
      RECT 29.494 17.158 29.546 17.194 ;
      RECT 29.494 18.358 29.546 18.394 ;
      RECT 29.494 19.558 29.546 19.594 ;
      RECT 29.494 20.758 29.546 20.794 ;
      RECT 29.494 21.958 29.546 21.994 ;
      RECT 29.494 23.158 29.546 23.194 ;
      RECT 29.494 24.358 29.546 24.394 ;
      RECT 29.494 25.558 29.546 25.594 ;
      RECT 29.494 26.758 29.546 26.794 ;
      RECT 29.494 27.958 29.546 27.994 ;
      RECT 29.494 29.158 29.546 29.194 ;
      RECT 29.494 30.358 29.546 30.394 ;
      RECT 29.494 31.558 29.546 31.594 ;
      RECT 29.494 33.342 29.546 33.378 ;
      RECT 29.494 33.582 29.546 33.618 ;
      RECT 29.494 37.902 29.546 37.938 ;
      RECT 29.494 38.142 29.546 38.178 ;
      RECT 29.494 40.678 29.546 40.714 ;
      RECT 29.494 41.878 29.546 41.914 ;
      RECT 29.494 43.078 29.546 43.114 ;
      RECT 29.494 44.278 29.546 44.314 ;
      RECT 29.494 45.478 29.546 45.514 ;
      RECT 29.494 46.678 29.546 46.714 ;
      RECT 29.494 47.878 29.546 47.914 ;
      RECT 29.494 49.078 29.546 49.114 ;
      RECT 29.494 50.278 29.546 50.314 ;
      RECT 29.494 51.478 29.546 51.514 ;
      RECT 29.494 52.678 29.546 52.714 ;
      RECT 29.494 53.878 29.546 53.914 ;
      RECT 29.494 55.078 29.546 55.114 ;
      RECT 29.494 56.278 29.546 56.314 ;
      RECT 29.494 57.478 29.546 57.514 ;
      RECT 29.494 58.678 29.546 58.714 ;
      RECT 29.494 59.878 29.546 59.914 ;
      RECT 29.494 61.078 29.546 61.114 ;
      RECT 29.494 62.278 29.546 62.314 ;
      RECT 29.494 63.478 29.546 63.514 ;
      RECT 29.494 64.678 29.546 64.714 ;
      RECT 29.494 65.878 29.546 65.914 ;
      RECT 29.494 67.078 29.546 67.114 ;
      RECT 29.494 68.278 29.546 68.314 ;
      RECT 29.494 69.478 29.546 69.514 ;
      RECT 29.494 70.678 29.546 70.714 ;
      RECT 29.494 71.878 29.546 71.914 ;
      RECT 29.574 0.281 29.626 0.317 ;
      RECT 29.574 72.403 29.626 72.439 ;
      RECT 29.654 0.806 29.706 0.842 ;
      RECT 29.654 2.006 29.706 2.042 ;
      RECT 29.654 3.206 29.706 3.242 ;
      RECT 29.654 4.406 29.706 4.442 ;
      RECT 29.654 5.606 29.706 5.642 ;
      RECT 29.654 6.806 29.706 6.842 ;
      RECT 29.654 8.006 29.706 8.042 ;
      RECT 29.654 9.206 29.706 9.242 ;
      RECT 29.654 10.406 29.706 10.442 ;
      RECT 29.654 11.606 29.706 11.642 ;
      RECT 29.654 12.806 29.706 12.842 ;
      RECT 29.654 14.006 29.706 14.042 ;
      RECT 29.654 15.206 29.706 15.242 ;
      RECT 29.654 16.406 29.706 16.442 ;
      RECT 29.654 17.606 29.706 17.642 ;
      RECT 29.654 18.806 29.706 18.842 ;
      RECT 29.654 20.006 29.706 20.042 ;
      RECT 29.654 21.206 29.706 21.242 ;
      RECT 29.654 22.406 29.706 22.442 ;
      RECT 29.654 23.606 29.706 23.642 ;
      RECT 29.654 24.806 29.706 24.842 ;
      RECT 29.654 26.006 29.706 26.042 ;
      RECT 29.654 27.206 29.706 27.242 ;
      RECT 29.654 28.406 29.706 28.442 ;
      RECT 29.654 29.606 29.706 29.642 ;
      RECT 29.654 30.806 29.706 30.842 ;
      RECT 29.654 32.622 29.706 32.658 ;
      RECT 29.654 32.862 29.706 32.898 ;
      RECT 29.654 34.302 29.706 34.338 ;
      RECT 29.654 34.782 29.706 34.818 ;
      RECT 29.654 36.702 29.706 36.738 ;
      RECT 29.654 37.182 29.706 37.218 ;
      RECT 29.654 38.622 29.706 38.658 ;
      RECT 29.654 38.862 29.706 38.898 ;
      RECT 29.654 39.926 29.706 39.962 ;
      RECT 29.654 41.126 29.706 41.162 ;
      RECT 29.654 42.326 29.706 42.362 ;
      RECT 29.654 43.526 29.706 43.562 ;
      RECT 29.654 44.726 29.706 44.762 ;
      RECT 29.654 45.926 29.706 45.962 ;
      RECT 29.654 47.126 29.706 47.162 ;
      RECT 29.654 48.326 29.706 48.362 ;
      RECT 29.654 49.526 29.706 49.562 ;
      RECT 29.654 50.726 29.706 50.762 ;
      RECT 29.654 51.926 29.706 51.962 ;
      RECT 29.654 53.126 29.706 53.162 ;
      RECT 29.654 54.326 29.706 54.362 ;
      RECT 29.654 55.526 29.706 55.562 ;
      RECT 29.654 56.726 29.706 56.762 ;
      RECT 29.654 57.926 29.706 57.962 ;
      RECT 29.654 59.126 29.706 59.162 ;
      RECT 29.654 60.326 29.706 60.362 ;
      RECT 29.654 61.526 29.706 61.562 ;
      RECT 29.654 62.726 29.706 62.762 ;
      RECT 29.654 63.926 29.706 63.962 ;
      RECT 29.654 65.126 29.706 65.162 ;
      RECT 29.654 66.326 29.706 66.362 ;
      RECT 29.654 67.526 29.706 67.562 ;
      RECT 29.654 68.726 29.706 68.762 ;
      RECT 29.654 69.926 29.706 69.962 ;
      RECT 29.654 71.126 29.706 71.162 ;
      RECT 29.734 1.558 29.786 1.594 ;
      RECT 29.734 2.758 29.786 2.794 ;
      RECT 29.734 3.958 29.786 3.994 ;
      RECT 29.734 5.158 29.786 5.194 ;
      RECT 29.734 6.358 29.786 6.394 ;
      RECT 29.734 7.558 29.786 7.594 ;
      RECT 29.734 8.758 29.786 8.794 ;
      RECT 29.734 9.958 29.786 9.994 ;
      RECT 29.734 11.158 29.786 11.194 ;
      RECT 29.734 12.358 29.786 12.394 ;
      RECT 29.734 13.558 29.786 13.594 ;
      RECT 29.734 14.758 29.786 14.794 ;
      RECT 29.734 15.958 29.786 15.994 ;
      RECT 29.734 17.158 29.786 17.194 ;
      RECT 29.734 18.358 29.786 18.394 ;
      RECT 29.734 19.558 29.786 19.594 ;
      RECT 29.734 20.758 29.786 20.794 ;
      RECT 29.734 21.958 29.786 21.994 ;
      RECT 29.734 23.158 29.786 23.194 ;
      RECT 29.734 24.358 29.786 24.394 ;
      RECT 29.734 25.558 29.786 25.594 ;
      RECT 29.734 26.758 29.786 26.794 ;
      RECT 29.734 27.958 29.786 27.994 ;
      RECT 29.734 29.158 29.786 29.194 ;
      RECT 29.734 30.358 29.786 30.394 ;
      RECT 29.734 31.558 29.786 31.594 ;
      RECT 29.734 33.342 29.786 33.378 ;
      RECT 29.734 33.582 29.786 33.618 ;
      RECT 29.734 37.902 29.786 37.938 ;
      RECT 29.734 38.142 29.786 38.178 ;
      RECT 29.734 40.678 29.786 40.714 ;
      RECT 29.734 41.878 29.786 41.914 ;
      RECT 29.734 43.078 29.786 43.114 ;
      RECT 29.734 44.278 29.786 44.314 ;
      RECT 29.734 45.478 29.786 45.514 ;
      RECT 29.734 46.678 29.786 46.714 ;
      RECT 29.734 47.878 29.786 47.914 ;
      RECT 29.734 49.078 29.786 49.114 ;
      RECT 29.734 50.278 29.786 50.314 ;
      RECT 29.734 51.478 29.786 51.514 ;
      RECT 29.734 52.678 29.786 52.714 ;
      RECT 29.734 53.878 29.786 53.914 ;
      RECT 29.734 55.078 29.786 55.114 ;
      RECT 29.734 56.278 29.786 56.314 ;
      RECT 29.734 57.478 29.786 57.514 ;
      RECT 29.734 58.678 29.786 58.714 ;
      RECT 29.734 59.878 29.786 59.914 ;
      RECT 29.734 61.078 29.786 61.114 ;
      RECT 29.734 62.278 29.786 62.314 ;
      RECT 29.734 63.478 29.786 63.514 ;
      RECT 29.734 64.678 29.786 64.714 ;
      RECT 29.734 65.878 29.786 65.914 ;
      RECT 29.734 67.078 29.786 67.114 ;
      RECT 29.734 68.278 29.786 68.314 ;
      RECT 29.734 69.478 29.786 69.514 ;
      RECT 29.734 70.678 29.786 70.714 ;
      RECT 29.734 71.878 29.786 71.914 ;
      RECT 29.814 0.806 29.866 0.842 ;
      RECT 29.814 2.006 29.866 2.042 ;
      RECT 29.814 3.206 29.866 3.242 ;
      RECT 29.814 4.406 29.866 4.442 ;
      RECT 29.814 5.606 29.866 5.642 ;
      RECT 29.814 6.806 29.866 6.842 ;
      RECT 29.814 8.006 29.866 8.042 ;
      RECT 29.814 9.206 29.866 9.242 ;
      RECT 29.814 10.406 29.866 10.442 ;
      RECT 29.814 11.606 29.866 11.642 ;
      RECT 29.814 12.806 29.866 12.842 ;
      RECT 29.814 14.006 29.866 14.042 ;
      RECT 29.814 15.206 29.866 15.242 ;
      RECT 29.814 16.406 29.866 16.442 ;
      RECT 29.814 17.606 29.866 17.642 ;
      RECT 29.814 18.806 29.866 18.842 ;
      RECT 29.814 20.006 29.866 20.042 ;
      RECT 29.814 21.206 29.866 21.242 ;
      RECT 29.814 22.406 29.866 22.442 ;
      RECT 29.814 23.606 29.866 23.642 ;
      RECT 29.814 24.806 29.866 24.842 ;
      RECT 29.814 26.006 29.866 26.042 ;
      RECT 29.814 27.206 29.866 27.242 ;
      RECT 29.814 28.406 29.866 28.442 ;
      RECT 29.814 29.606 29.866 29.642 ;
      RECT 29.814 30.806 29.866 30.842 ;
      RECT 29.814 32.622 29.866 32.658 ;
      RECT 29.814 32.862 29.866 32.898 ;
      RECT 29.814 38.622 29.866 38.658 ;
      RECT 29.814 38.862 29.866 38.898 ;
      RECT 29.814 39.926 29.866 39.962 ;
      RECT 29.814 41.126 29.866 41.162 ;
      RECT 29.814 42.326 29.866 42.362 ;
      RECT 29.814 43.526 29.866 43.562 ;
      RECT 29.814 44.726 29.866 44.762 ;
      RECT 29.814 45.926 29.866 45.962 ;
      RECT 29.814 47.126 29.866 47.162 ;
      RECT 29.814 48.326 29.866 48.362 ;
      RECT 29.814 49.526 29.866 49.562 ;
      RECT 29.814 50.726 29.866 50.762 ;
      RECT 29.814 51.926 29.866 51.962 ;
      RECT 29.814 53.126 29.866 53.162 ;
      RECT 29.814 54.326 29.866 54.362 ;
      RECT 29.814 55.526 29.866 55.562 ;
      RECT 29.814 56.726 29.866 56.762 ;
      RECT 29.814 57.926 29.866 57.962 ;
      RECT 29.814 59.126 29.866 59.162 ;
      RECT 29.814 60.326 29.866 60.362 ;
      RECT 29.814 61.526 29.866 61.562 ;
      RECT 29.814 62.726 29.866 62.762 ;
      RECT 29.814 63.926 29.866 63.962 ;
      RECT 29.814 65.126 29.866 65.162 ;
      RECT 29.814 66.326 29.866 66.362 ;
      RECT 29.814 67.526 29.866 67.562 ;
      RECT 29.814 68.726 29.866 68.762 ;
      RECT 29.814 69.926 29.866 69.962 ;
      RECT 29.814 71.126 29.866 71.162 ;
      RECT 29.894 1.558 29.946 1.594 ;
      RECT 29.894 2.758 29.946 2.794 ;
      RECT 29.894 3.958 29.946 3.994 ;
      RECT 29.894 5.158 29.946 5.194 ;
      RECT 29.894 6.358 29.946 6.394 ;
      RECT 29.894 7.558 29.946 7.594 ;
      RECT 29.894 8.758 29.946 8.794 ;
      RECT 29.894 9.958 29.946 9.994 ;
      RECT 29.894 11.158 29.946 11.194 ;
      RECT 29.894 12.358 29.946 12.394 ;
      RECT 29.894 13.558 29.946 13.594 ;
      RECT 29.894 14.758 29.946 14.794 ;
      RECT 29.894 15.958 29.946 15.994 ;
      RECT 29.894 17.158 29.946 17.194 ;
      RECT 29.894 18.358 29.946 18.394 ;
      RECT 29.894 19.558 29.946 19.594 ;
      RECT 29.894 20.758 29.946 20.794 ;
      RECT 29.894 21.958 29.946 21.994 ;
      RECT 29.894 23.158 29.946 23.194 ;
      RECT 29.894 24.358 29.946 24.394 ;
      RECT 29.894 25.558 29.946 25.594 ;
      RECT 29.894 26.758 29.946 26.794 ;
      RECT 29.894 27.958 29.946 27.994 ;
      RECT 29.894 29.158 29.946 29.194 ;
      RECT 29.894 30.358 29.946 30.394 ;
      RECT 29.894 31.558 29.946 31.594 ;
      RECT 29.894 33.342 29.946 33.378 ;
      RECT 29.894 33.582 29.946 33.618 ;
      RECT 29.894 37.902 29.946 37.938 ;
      RECT 29.894 38.142 29.946 38.178 ;
      RECT 29.894 40.678 29.946 40.714 ;
      RECT 29.894 41.878 29.946 41.914 ;
      RECT 29.894 43.078 29.946 43.114 ;
      RECT 29.894 44.278 29.946 44.314 ;
      RECT 29.894 45.478 29.946 45.514 ;
      RECT 29.894 46.678 29.946 46.714 ;
      RECT 29.894 47.878 29.946 47.914 ;
      RECT 29.894 49.078 29.946 49.114 ;
      RECT 29.894 50.278 29.946 50.314 ;
      RECT 29.894 51.478 29.946 51.514 ;
      RECT 29.894 52.678 29.946 52.714 ;
      RECT 29.894 53.878 29.946 53.914 ;
      RECT 29.894 55.078 29.946 55.114 ;
      RECT 29.894 56.278 29.946 56.314 ;
      RECT 29.894 57.478 29.946 57.514 ;
      RECT 29.894 58.678 29.946 58.714 ;
      RECT 29.894 59.878 29.946 59.914 ;
      RECT 29.894 61.078 29.946 61.114 ;
      RECT 29.894 62.278 29.946 62.314 ;
      RECT 29.894 63.478 29.946 63.514 ;
      RECT 29.894 64.678 29.946 64.714 ;
      RECT 29.894 65.878 29.946 65.914 ;
      RECT 29.894 67.078 29.946 67.114 ;
      RECT 29.894 68.278 29.946 68.314 ;
      RECT 29.894 69.478 29.946 69.514 ;
      RECT 29.894 70.678 29.946 70.714 ;
      RECT 29.894 71.878 29.946 71.914 ;
      RECT 29.974 0.281 30.026 0.317 ;
      RECT 29.974 72.403 30.026 72.439 ;
      RECT 30.054 0.806 30.106 0.842 ;
      RECT 30.054 2.006 30.106 2.042 ;
      RECT 30.054 3.206 30.106 3.242 ;
      RECT 30.054 4.406 30.106 4.442 ;
      RECT 30.054 5.606 30.106 5.642 ;
      RECT 30.054 6.806 30.106 6.842 ;
      RECT 30.054 8.006 30.106 8.042 ;
      RECT 30.054 9.206 30.106 9.242 ;
      RECT 30.054 10.406 30.106 10.442 ;
      RECT 30.054 11.606 30.106 11.642 ;
      RECT 30.054 12.806 30.106 12.842 ;
      RECT 30.054 14.006 30.106 14.042 ;
      RECT 30.054 15.206 30.106 15.242 ;
      RECT 30.054 16.406 30.106 16.442 ;
      RECT 30.054 17.606 30.106 17.642 ;
      RECT 30.054 18.806 30.106 18.842 ;
      RECT 30.054 20.006 30.106 20.042 ;
      RECT 30.054 21.206 30.106 21.242 ;
      RECT 30.054 22.406 30.106 22.442 ;
      RECT 30.054 23.606 30.106 23.642 ;
      RECT 30.054 24.806 30.106 24.842 ;
      RECT 30.054 26.006 30.106 26.042 ;
      RECT 30.054 27.206 30.106 27.242 ;
      RECT 30.054 28.406 30.106 28.442 ;
      RECT 30.054 29.606 30.106 29.642 ;
      RECT 30.054 30.806 30.106 30.842 ;
      RECT 30.054 32.622 30.106 32.658 ;
      RECT 30.054 32.862 30.106 32.898 ;
      RECT 30.054 38.622 30.106 38.658 ;
      RECT 30.054 38.862 30.106 38.898 ;
      RECT 30.054 39.926 30.106 39.962 ;
      RECT 30.054 41.126 30.106 41.162 ;
      RECT 30.054 42.326 30.106 42.362 ;
      RECT 30.054 43.526 30.106 43.562 ;
      RECT 30.054 44.726 30.106 44.762 ;
      RECT 30.054 45.926 30.106 45.962 ;
      RECT 30.054 47.126 30.106 47.162 ;
      RECT 30.054 48.326 30.106 48.362 ;
      RECT 30.054 49.526 30.106 49.562 ;
      RECT 30.054 50.726 30.106 50.762 ;
      RECT 30.054 51.926 30.106 51.962 ;
      RECT 30.054 53.126 30.106 53.162 ;
      RECT 30.054 54.326 30.106 54.362 ;
      RECT 30.054 55.526 30.106 55.562 ;
      RECT 30.054 56.726 30.106 56.762 ;
      RECT 30.054 57.926 30.106 57.962 ;
      RECT 30.054 59.126 30.106 59.162 ;
      RECT 30.054 60.326 30.106 60.362 ;
      RECT 30.054 61.526 30.106 61.562 ;
      RECT 30.054 62.726 30.106 62.762 ;
      RECT 30.054 63.926 30.106 63.962 ;
      RECT 30.054 65.126 30.106 65.162 ;
      RECT 30.054 66.326 30.106 66.362 ;
      RECT 30.054 67.526 30.106 67.562 ;
      RECT 30.054 68.726 30.106 68.762 ;
      RECT 30.054 69.926 30.106 69.962 ;
      RECT 30.054 71.126 30.106 71.162 ;
      RECT 30.134 1.558 30.186 1.594 ;
      RECT 30.134 2.758 30.186 2.794 ;
      RECT 30.134 3.958 30.186 3.994 ;
      RECT 30.134 5.158 30.186 5.194 ;
      RECT 30.134 6.358 30.186 6.394 ;
      RECT 30.134 7.558 30.186 7.594 ;
      RECT 30.134 8.758 30.186 8.794 ;
      RECT 30.134 9.958 30.186 9.994 ;
      RECT 30.134 11.158 30.186 11.194 ;
      RECT 30.134 12.358 30.186 12.394 ;
      RECT 30.134 13.558 30.186 13.594 ;
      RECT 30.134 14.758 30.186 14.794 ;
      RECT 30.134 15.958 30.186 15.994 ;
      RECT 30.134 17.158 30.186 17.194 ;
      RECT 30.134 18.358 30.186 18.394 ;
      RECT 30.134 19.558 30.186 19.594 ;
      RECT 30.134 20.758 30.186 20.794 ;
      RECT 30.134 21.958 30.186 21.994 ;
      RECT 30.134 23.158 30.186 23.194 ;
      RECT 30.134 24.358 30.186 24.394 ;
      RECT 30.134 25.558 30.186 25.594 ;
      RECT 30.134 26.758 30.186 26.794 ;
      RECT 30.134 27.958 30.186 27.994 ;
      RECT 30.134 29.158 30.186 29.194 ;
      RECT 30.134 30.358 30.186 30.394 ;
      RECT 30.134 31.558 30.186 31.594 ;
      RECT 30.134 33.342 30.186 33.378 ;
      RECT 30.134 33.582 30.186 33.618 ;
      RECT 30.134 37.902 30.186 37.938 ;
      RECT 30.134 38.142 30.186 38.178 ;
      RECT 30.134 40.678 30.186 40.714 ;
      RECT 30.134 41.878 30.186 41.914 ;
      RECT 30.134 43.078 30.186 43.114 ;
      RECT 30.134 44.278 30.186 44.314 ;
      RECT 30.134 45.478 30.186 45.514 ;
      RECT 30.134 46.678 30.186 46.714 ;
      RECT 30.134 47.878 30.186 47.914 ;
      RECT 30.134 49.078 30.186 49.114 ;
      RECT 30.134 50.278 30.186 50.314 ;
      RECT 30.134 51.478 30.186 51.514 ;
      RECT 30.134 52.678 30.186 52.714 ;
      RECT 30.134 53.878 30.186 53.914 ;
      RECT 30.134 55.078 30.186 55.114 ;
      RECT 30.134 56.278 30.186 56.314 ;
      RECT 30.134 57.478 30.186 57.514 ;
      RECT 30.134 58.678 30.186 58.714 ;
      RECT 30.134 59.878 30.186 59.914 ;
      RECT 30.134 61.078 30.186 61.114 ;
      RECT 30.134 62.278 30.186 62.314 ;
      RECT 30.134 63.478 30.186 63.514 ;
      RECT 30.134 64.678 30.186 64.714 ;
      RECT 30.134 65.878 30.186 65.914 ;
      RECT 30.134 67.078 30.186 67.114 ;
      RECT 30.134 68.278 30.186 68.314 ;
      RECT 30.134 69.478 30.186 69.514 ;
      RECT 30.134 70.678 30.186 70.714 ;
      RECT 30.134 71.878 30.186 71.914 ;
      RECT 30.214 0.806 30.266 0.842 ;
      RECT 30.214 2.006 30.266 2.042 ;
      RECT 30.214 3.206 30.266 3.242 ;
      RECT 30.214 4.406 30.266 4.442 ;
      RECT 30.214 5.606 30.266 5.642 ;
      RECT 30.214 6.806 30.266 6.842 ;
      RECT 30.214 8.006 30.266 8.042 ;
      RECT 30.214 9.206 30.266 9.242 ;
      RECT 30.214 10.406 30.266 10.442 ;
      RECT 30.214 11.606 30.266 11.642 ;
      RECT 30.214 12.806 30.266 12.842 ;
      RECT 30.214 14.006 30.266 14.042 ;
      RECT 30.214 15.206 30.266 15.242 ;
      RECT 30.214 16.406 30.266 16.442 ;
      RECT 30.214 17.606 30.266 17.642 ;
      RECT 30.214 18.806 30.266 18.842 ;
      RECT 30.214 20.006 30.266 20.042 ;
      RECT 30.214 21.206 30.266 21.242 ;
      RECT 30.214 22.406 30.266 22.442 ;
      RECT 30.214 23.606 30.266 23.642 ;
      RECT 30.214 24.806 30.266 24.842 ;
      RECT 30.214 26.006 30.266 26.042 ;
      RECT 30.214 27.206 30.266 27.242 ;
      RECT 30.214 28.406 30.266 28.442 ;
      RECT 30.214 29.606 30.266 29.642 ;
      RECT 30.214 30.806 30.266 30.842 ;
      RECT 30.214 32.622 30.266 32.658 ;
      RECT 30.214 32.862 30.266 32.898 ;
      RECT 30.214 38.622 30.266 38.658 ;
      RECT 30.214 38.862 30.266 38.898 ;
      RECT 30.214 39.926 30.266 39.962 ;
      RECT 30.214 41.126 30.266 41.162 ;
      RECT 30.214 42.326 30.266 42.362 ;
      RECT 30.214 43.526 30.266 43.562 ;
      RECT 30.214 44.726 30.266 44.762 ;
      RECT 30.214 45.926 30.266 45.962 ;
      RECT 30.214 47.126 30.266 47.162 ;
      RECT 30.214 48.326 30.266 48.362 ;
      RECT 30.214 49.526 30.266 49.562 ;
      RECT 30.214 50.726 30.266 50.762 ;
      RECT 30.214 51.926 30.266 51.962 ;
      RECT 30.214 53.126 30.266 53.162 ;
      RECT 30.214 54.326 30.266 54.362 ;
      RECT 30.214 55.526 30.266 55.562 ;
      RECT 30.214 56.726 30.266 56.762 ;
      RECT 30.214 57.926 30.266 57.962 ;
      RECT 30.214 59.126 30.266 59.162 ;
      RECT 30.214 60.326 30.266 60.362 ;
      RECT 30.214 61.526 30.266 61.562 ;
      RECT 30.214 62.726 30.266 62.762 ;
      RECT 30.214 63.926 30.266 63.962 ;
      RECT 30.214 65.126 30.266 65.162 ;
      RECT 30.214 66.326 30.266 66.362 ;
      RECT 30.214 67.526 30.266 67.562 ;
      RECT 30.214 68.726 30.266 68.762 ;
      RECT 30.214 69.926 30.266 69.962 ;
      RECT 30.214 71.126 30.266 71.162 ;
      RECT 30.294 1.558 30.346 1.594 ;
      RECT 30.294 2.758 30.346 2.794 ;
      RECT 30.294 3.958 30.346 3.994 ;
      RECT 30.294 5.158 30.346 5.194 ;
      RECT 30.294 6.358 30.346 6.394 ;
      RECT 30.294 7.558 30.346 7.594 ;
      RECT 30.294 8.758 30.346 8.794 ;
      RECT 30.294 9.958 30.346 9.994 ;
      RECT 30.294 11.158 30.346 11.194 ;
      RECT 30.294 12.358 30.346 12.394 ;
      RECT 30.294 13.558 30.346 13.594 ;
      RECT 30.294 14.758 30.346 14.794 ;
      RECT 30.294 15.958 30.346 15.994 ;
      RECT 30.294 17.158 30.346 17.194 ;
      RECT 30.294 18.358 30.346 18.394 ;
      RECT 30.294 19.558 30.346 19.594 ;
      RECT 30.294 20.758 30.346 20.794 ;
      RECT 30.294 21.958 30.346 21.994 ;
      RECT 30.294 23.158 30.346 23.194 ;
      RECT 30.294 24.358 30.346 24.394 ;
      RECT 30.294 25.558 30.346 25.594 ;
      RECT 30.294 26.758 30.346 26.794 ;
      RECT 30.294 27.958 30.346 27.994 ;
      RECT 30.294 29.158 30.346 29.194 ;
      RECT 30.294 30.358 30.346 30.394 ;
      RECT 30.294 31.558 30.346 31.594 ;
      RECT 30.294 33.342 30.346 33.378 ;
      RECT 30.294 33.582 30.346 33.618 ;
      RECT 30.294 37.902 30.346 37.938 ;
      RECT 30.294 38.142 30.346 38.178 ;
      RECT 30.294 40.678 30.346 40.714 ;
      RECT 30.294 41.878 30.346 41.914 ;
      RECT 30.294 43.078 30.346 43.114 ;
      RECT 30.294 44.278 30.346 44.314 ;
      RECT 30.294 45.478 30.346 45.514 ;
      RECT 30.294 46.678 30.346 46.714 ;
      RECT 30.294 47.878 30.346 47.914 ;
      RECT 30.294 49.078 30.346 49.114 ;
      RECT 30.294 50.278 30.346 50.314 ;
      RECT 30.294 51.478 30.346 51.514 ;
      RECT 30.294 52.678 30.346 52.714 ;
      RECT 30.294 53.878 30.346 53.914 ;
      RECT 30.294 55.078 30.346 55.114 ;
      RECT 30.294 56.278 30.346 56.314 ;
      RECT 30.294 57.478 30.346 57.514 ;
      RECT 30.294 58.678 30.346 58.714 ;
      RECT 30.294 59.878 30.346 59.914 ;
      RECT 30.294 61.078 30.346 61.114 ;
      RECT 30.294 62.278 30.346 62.314 ;
      RECT 30.294 63.478 30.346 63.514 ;
      RECT 30.294 64.678 30.346 64.714 ;
      RECT 30.294 65.878 30.346 65.914 ;
      RECT 30.294 67.078 30.346 67.114 ;
      RECT 30.294 68.278 30.346 68.314 ;
      RECT 30.294 69.478 30.346 69.514 ;
      RECT 30.294 70.678 30.346 70.714 ;
      RECT 30.294 71.878 30.346 71.914 ;
      RECT 30.374 0.281 30.426 0.317 ;
      RECT 30.374 72.403 30.426 72.439 ;
      RECT 30.454 0.806 30.506 0.842 ;
      RECT 30.454 2.006 30.506 2.042 ;
      RECT 30.454 3.206 30.506 3.242 ;
      RECT 30.454 4.406 30.506 4.442 ;
      RECT 30.454 5.606 30.506 5.642 ;
      RECT 30.454 6.806 30.506 6.842 ;
      RECT 30.454 8.006 30.506 8.042 ;
      RECT 30.454 9.206 30.506 9.242 ;
      RECT 30.454 10.406 30.506 10.442 ;
      RECT 30.454 11.606 30.506 11.642 ;
      RECT 30.454 12.806 30.506 12.842 ;
      RECT 30.454 14.006 30.506 14.042 ;
      RECT 30.454 15.206 30.506 15.242 ;
      RECT 30.454 16.406 30.506 16.442 ;
      RECT 30.454 17.606 30.506 17.642 ;
      RECT 30.454 18.806 30.506 18.842 ;
      RECT 30.454 20.006 30.506 20.042 ;
      RECT 30.454 21.206 30.506 21.242 ;
      RECT 30.454 22.406 30.506 22.442 ;
      RECT 30.454 23.606 30.506 23.642 ;
      RECT 30.454 24.806 30.506 24.842 ;
      RECT 30.454 26.006 30.506 26.042 ;
      RECT 30.454 27.206 30.506 27.242 ;
      RECT 30.454 28.406 30.506 28.442 ;
      RECT 30.454 29.606 30.506 29.642 ;
      RECT 30.454 30.806 30.506 30.842 ;
      RECT 30.454 32.622 30.506 32.658 ;
      RECT 30.454 32.862 30.506 32.898 ;
      RECT 30.454 34.302 30.506 34.338 ;
      RECT 30.454 34.782 30.506 34.818 ;
      RECT 30.454 36.702 30.506 36.738 ;
      RECT 30.454 37.182 30.506 37.218 ;
      RECT 30.454 38.622 30.506 38.658 ;
      RECT 30.454 38.862 30.506 38.898 ;
      RECT 30.454 39.926 30.506 39.962 ;
      RECT 30.454 41.126 30.506 41.162 ;
      RECT 30.454 42.326 30.506 42.362 ;
      RECT 30.454 43.526 30.506 43.562 ;
      RECT 30.454 44.726 30.506 44.762 ;
      RECT 30.454 45.926 30.506 45.962 ;
      RECT 30.454 47.126 30.506 47.162 ;
      RECT 30.454 48.326 30.506 48.362 ;
      RECT 30.454 49.526 30.506 49.562 ;
      RECT 30.454 50.726 30.506 50.762 ;
      RECT 30.454 51.926 30.506 51.962 ;
      RECT 30.454 53.126 30.506 53.162 ;
      RECT 30.454 54.326 30.506 54.362 ;
      RECT 30.454 55.526 30.506 55.562 ;
      RECT 30.454 56.726 30.506 56.762 ;
      RECT 30.454 57.926 30.506 57.962 ;
      RECT 30.454 59.126 30.506 59.162 ;
      RECT 30.454 60.326 30.506 60.362 ;
      RECT 30.454 61.526 30.506 61.562 ;
      RECT 30.454 62.726 30.506 62.762 ;
      RECT 30.454 63.926 30.506 63.962 ;
      RECT 30.454 65.126 30.506 65.162 ;
      RECT 30.454 66.326 30.506 66.362 ;
      RECT 30.454 67.526 30.506 67.562 ;
      RECT 30.454 68.726 30.506 68.762 ;
      RECT 30.454 69.926 30.506 69.962 ;
      RECT 30.454 71.126 30.506 71.162 ;
      RECT 30.534 1.558 30.586 1.594 ;
      RECT 30.534 2.758 30.586 2.794 ;
      RECT 30.534 3.958 30.586 3.994 ;
      RECT 30.534 5.158 30.586 5.194 ;
      RECT 30.534 6.358 30.586 6.394 ;
      RECT 30.534 7.558 30.586 7.594 ;
      RECT 30.534 8.758 30.586 8.794 ;
      RECT 30.534 9.958 30.586 9.994 ;
      RECT 30.534 11.158 30.586 11.194 ;
      RECT 30.534 12.358 30.586 12.394 ;
      RECT 30.534 13.558 30.586 13.594 ;
      RECT 30.534 14.758 30.586 14.794 ;
      RECT 30.534 15.958 30.586 15.994 ;
      RECT 30.534 17.158 30.586 17.194 ;
      RECT 30.534 18.358 30.586 18.394 ;
      RECT 30.534 19.558 30.586 19.594 ;
      RECT 30.534 20.758 30.586 20.794 ;
      RECT 30.534 21.958 30.586 21.994 ;
      RECT 30.534 23.158 30.586 23.194 ;
      RECT 30.534 24.358 30.586 24.394 ;
      RECT 30.534 25.558 30.586 25.594 ;
      RECT 30.534 26.758 30.586 26.794 ;
      RECT 30.534 27.958 30.586 27.994 ;
      RECT 30.534 29.158 30.586 29.194 ;
      RECT 30.534 30.358 30.586 30.394 ;
      RECT 30.534 31.558 30.586 31.594 ;
      RECT 30.534 33.342 30.586 33.378 ;
      RECT 30.534 33.582 30.586 33.618 ;
      RECT 30.534 37.902 30.586 37.938 ;
      RECT 30.534 38.142 30.586 38.178 ;
      RECT 30.534 40.678 30.586 40.714 ;
      RECT 30.534 41.878 30.586 41.914 ;
      RECT 30.534 43.078 30.586 43.114 ;
      RECT 30.534 44.278 30.586 44.314 ;
      RECT 30.534 45.478 30.586 45.514 ;
      RECT 30.534 46.678 30.586 46.714 ;
      RECT 30.534 47.878 30.586 47.914 ;
      RECT 30.534 49.078 30.586 49.114 ;
      RECT 30.534 50.278 30.586 50.314 ;
      RECT 30.534 51.478 30.586 51.514 ;
      RECT 30.534 52.678 30.586 52.714 ;
      RECT 30.534 53.878 30.586 53.914 ;
      RECT 30.534 55.078 30.586 55.114 ;
      RECT 30.534 56.278 30.586 56.314 ;
      RECT 30.534 57.478 30.586 57.514 ;
      RECT 30.534 58.678 30.586 58.714 ;
      RECT 30.534 59.878 30.586 59.914 ;
      RECT 30.534 61.078 30.586 61.114 ;
      RECT 30.534 62.278 30.586 62.314 ;
      RECT 30.534 63.478 30.586 63.514 ;
      RECT 30.534 64.678 30.586 64.714 ;
      RECT 30.534 65.878 30.586 65.914 ;
      RECT 30.534 67.078 30.586 67.114 ;
      RECT 30.534 68.278 30.586 68.314 ;
      RECT 30.534 69.478 30.586 69.514 ;
      RECT 30.534 70.678 30.586 70.714 ;
      RECT 30.534 71.878 30.586 71.914 ;
      RECT 30.614 0.806 30.666 0.842 ;
      RECT 30.614 2.006 30.666 2.042 ;
      RECT 30.614 3.206 30.666 3.242 ;
      RECT 30.614 4.406 30.666 4.442 ;
      RECT 30.614 5.606 30.666 5.642 ;
      RECT 30.614 6.806 30.666 6.842 ;
      RECT 30.614 8.006 30.666 8.042 ;
      RECT 30.614 9.206 30.666 9.242 ;
      RECT 30.614 10.406 30.666 10.442 ;
      RECT 30.614 11.606 30.666 11.642 ;
      RECT 30.614 12.806 30.666 12.842 ;
      RECT 30.614 14.006 30.666 14.042 ;
      RECT 30.614 15.206 30.666 15.242 ;
      RECT 30.614 16.406 30.666 16.442 ;
      RECT 30.614 17.606 30.666 17.642 ;
      RECT 30.614 18.806 30.666 18.842 ;
      RECT 30.614 20.006 30.666 20.042 ;
      RECT 30.614 21.206 30.666 21.242 ;
      RECT 30.614 22.406 30.666 22.442 ;
      RECT 30.614 23.606 30.666 23.642 ;
      RECT 30.614 24.806 30.666 24.842 ;
      RECT 30.614 26.006 30.666 26.042 ;
      RECT 30.614 27.206 30.666 27.242 ;
      RECT 30.614 28.406 30.666 28.442 ;
      RECT 30.614 29.606 30.666 29.642 ;
      RECT 30.614 30.806 30.666 30.842 ;
      RECT 30.614 32.622 30.666 32.658 ;
      RECT 30.614 32.862 30.666 32.898 ;
      RECT 30.614 38.622 30.666 38.658 ;
      RECT 30.614 38.862 30.666 38.898 ;
      RECT 30.614 39.926 30.666 39.962 ;
      RECT 30.614 41.126 30.666 41.162 ;
      RECT 30.614 42.326 30.666 42.362 ;
      RECT 30.614 43.526 30.666 43.562 ;
      RECT 30.614 44.726 30.666 44.762 ;
      RECT 30.614 45.926 30.666 45.962 ;
      RECT 30.614 47.126 30.666 47.162 ;
      RECT 30.614 48.326 30.666 48.362 ;
      RECT 30.614 49.526 30.666 49.562 ;
      RECT 30.614 50.726 30.666 50.762 ;
      RECT 30.614 51.926 30.666 51.962 ;
      RECT 30.614 53.126 30.666 53.162 ;
      RECT 30.614 54.326 30.666 54.362 ;
      RECT 30.614 55.526 30.666 55.562 ;
      RECT 30.614 56.726 30.666 56.762 ;
      RECT 30.614 57.926 30.666 57.962 ;
      RECT 30.614 59.126 30.666 59.162 ;
      RECT 30.614 60.326 30.666 60.362 ;
      RECT 30.614 61.526 30.666 61.562 ;
      RECT 30.614 62.726 30.666 62.762 ;
      RECT 30.614 63.926 30.666 63.962 ;
      RECT 30.614 65.126 30.666 65.162 ;
      RECT 30.614 66.326 30.666 66.362 ;
      RECT 30.614 67.526 30.666 67.562 ;
      RECT 30.614 68.726 30.666 68.762 ;
      RECT 30.614 69.926 30.666 69.962 ;
      RECT 30.614 71.126 30.666 71.162 ;
      RECT 30.694 1.558 30.746 1.594 ;
      RECT 30.694 2.758 30.746 2.794 ;
      RECT 30.694 3.958 30.746 3.994 ;
      RECT 30.694 5.158 30.746 5.194 ;
      RECT 30.694 6.358 30.746 6.394 ;
      RECT 30.694 7.558 30.746 7.594 ;
      RECT 30.694 8.758 30.746 8.794 ;
      RECT 30.694 9.958 30.746 9.994 ;
      RECT 30.694 11.158 30.746 11.194 ;
      RECT 30.694 12.358 30.746 12.394 ;
      RECT 30.694 13.558 30.746 13.594 ;
      RECT 30.694 14.758 30.746 14.794 ;
      RECT 30.694 15.958 30.746 15.994 ;
      RECT 30.694 17.158 30.746 17.194 ;
      RECT 30.694 18.358 30.746 18.394 ;
      RECT 30.694 19.558 30.746 19.594 ;
      RECT 30.694 20.758 30.746 20.794 ;
      RECT 30.694 21.958 30.746 21.994 ;
      RECT 30.694 23.158 30.746 23.194 ;
      RECT 30.694 24.358 30.746 24.394 ;
      RECT 30.694 25.558 30.746 25.594 ;
      RECT 30.694 26.758 30.746 26.794 ;
      RECT 30.694 27.958 30.746 27.994 ;
      RECT 30.694 29.158 30.746 29.194 ;
      RECT 30.694 30.358 30.746 30.394 ;
      RECT 30.694 31.558 30.746 31.594 ;
      RECT 30.694 33.342 30.746 33.378 ;
      RECT 30.694 33.582 30.746 33.618 ;
      RECT 30.694 37.902 30.746 37.938 ;
      RECT 30.694 38.142 30.746 38.178 ;
      RECT 30.694 40.678 30.746 40.714 ;
      RECT 30.694 41.878 30.746 41.914 ;
      RECT 30.694 43.078 30.746 43.114 ;
      RECT 30.694 44.278 30.746 44.314 ;
      RECT 30.694 45.478 30.746 45.514 ;
      RECT 30.694 46.678 30.746 46.714 ;
      RECT 30.694 47.878 30.746 47.914 ;
      RECT 30.694 49.078 30.746 49.114 ;
      RECT 30.694 50.278 30.746 50.314 ;
      RECT 30.694 51.478 30.746 51.514 ;
      RECT 30.694 52.678 30.746 52.714 ;
      RECT 30.694 53.878 30.746 53.914 ;
      RECT 30.694 55.078 30.746 55.114 ;
      RECT 30.694 56.278 30.746 56.314 ;
      RECT 30.694 57.478 30.746 57.514 ;
      RECT 30.694 58.678 30.746 58.714 ;
      RECT 30.694 59.878 30.746 59.914 ;
      RECT 30.694 61.078 30.746 61.114 ;
      RECT 30.694 62.278 30.746 62.314 ;
      RECT 30.694 63.478 30.746 63.514 ;
      RECT 30.694 64.678 30.746 64.714 ;
      RECT 30.694 65.878 30.746 65.914 ;
      RECT 30.694 67.078 30.746 67.114 ;
      RECT 30.694 68.278 30.746 68.314 ;
      RECT 30.694 69.478 30.746 69.514 ;
      RECT 30.694 70.678 30.746 70.714 ;
      RECT 30.694 71.878 30.746 71.914 ;
      RECT 30.774 0.281 30.826 0.317 ;
      RECT 30.774 72.403 30.826 72.439 ;
      RECT 30.854 0.806 30.906 0.842 ;
      RECT 30.854 2.006 30.906 2.042 ;
      RECT 30.854 3.206 30.906 3.242 ;
      RECT 30.854 4.406 30.906 4.442 ;
      RECT 30.854 5.606 30.906 5.642 ;
      RECT 30.854 6.806 30.906 6.842 ;
      RECT 30.854 8.006 30.906 8.042 ;
      RECT 30.854 9.206 30.906 9.242 ;
      RECT 30.854 10.406 30.906 10.442 ;
      RECT 30.854 11.606 30.906 11.642 ;
      RECT 30.854 12.806 30.906 12.842 ;
      RECT 30.854 14.006 30.906 14.042 ;
      RECT 30.854 15.206 30.906 15.242 ;
      RECT 30.854 16.406 30.906 16.442 ;
      RECT 30.854 17.606 30.906 17.642 ;
      RECT 30.854 18.806 30.906 18.842 ;
      RECT 30.854 20.006 30.906 20.042 ;
      RECT 30.854 21.206 30.906 21.242 ;
      RECT 30.854 22.406 30.906 22.442 ;
      RECT 30.854 23.606 30.906 23.642 ;
      RECT 30.854 24.806 30.906 24.842 ;
      RECT 30.854 26.006 30.906 26.042 ;
      RECT 30.854 27.206 30.906 27.242 ;
      RECT 30.854 28.406 30.906 28.442 ;
      RECT 30.854 29.606 30.906 29.642 ;
      RECT 30.854 30.806 30.906 30.842 ;
      RECT 30.854 32.622 30.906 32.658 ;
      RECT 30.854 32.862 30.906 32.898 ;
      RECT 30.854 38.622 30.906 38.658 ;
      RECT 30.854 38.862 30.906 38.898 ;
      RECT 30.854 39.926 30.906 39.962 ;
      RECT 30.854 41.126 30.906 41.162 ;
      RECT 30.854 42.326 30.906 42.362 ;
      RECT 30.854 43.526 30.906 43.562 ;
      RECT 30.854 44.726 30.906 44.762 ;
      RECT 30.854 45.926 30.906 45.962 ;
      RECT 30.854 47.126 30.906 47.162 ;
      RECT 30.854 48.326 30.906 48.362 ;
      RECT 30.854 49.526 30.906 49.562 ;
      RECT 30.854 50.726 30.906 50.762 ;
      RECT 30.854 51.926 30.906 51.962 ;
      RECT 30.854 53.126 30.906 53.162 ;
      RECT 30.854 54.326 30.906 54.362 ;
      RECT 30.854 55.526 30.906 55.562 ;
      RECT 30.854 56.726 30.906 56.762 ;
      RECT 30.854 57.926 30.906 57.962 ;
      RECT 30.854 59.126 30.906 59.162 ;
      RECT 30.854 60.326 30.906 60.362 ;
      RECT 30.854 61.526 30.906 61.562 ;
      RECT 30.854 62.726 30.906 62.762 ;
      RECT 30.854 63.926 30.906 63.962 ;
      RECT 30.854 65.126 30.906 65.162 ;
      RECT 30.854 66.326 30.906 66.362 ;
      RECT 30.854 67.526 30.906 67.562 ;
      RECT 30.854 68.726 30.906 68.762 ;
      RECT 30.854 69.926 30.906 69.962 ;
      RECT 30.854 71.126 30.906 71.162 ;
      RECT 30.934 1.558 30.986 1.594 ;
      RECT 30.934 2.758 30.986 2.794 ;
      RECT 30.934 3.958 30.986 3.994 ;
      RECT 30.934 5.158 30.986 5.194 ;
      RECT 30.934 6.358 30.986 6.394 ;
      RECT 30.934 7.558 30.986 7.594 ;
      RECT 30.934 8.758 30.986 8.794 ;
      RECT 30.934 9.958 30.986 9.994 ;
      RECT 30.934 11.158 30.986 11.194 ;
      RECT 30.934 12.358 30.986 12.394 ;
      RECT 30.934 13.558 30.986 13.594 ;
      RECT 30.934 14.758 30.986 14.794 ;
      RECT 30.934 15.958 30.986 15.994 ;
      RECT 30.934 17.158 30.986 17.194 ;
      RECT 30.934 18.358 30.986 18.394 ;
      RECT 30.934 19.558 30.986 19.594 ;
      RECT 30.934 20.758 30.986 20.794 ;
      RECT 30.934 21.958 30.986 21.994 ;
      RECT 30.934 23.158 30.986 23.194 ;
      RECT 30.934 24.358 30.986 24.394 ;
      RECT 30.934 25.558 30.986 25.594 ;
      RECT 30.934 26.758 30.986 26.794 ;
      RECT 30.934 27.958 30.986 27.994 ;
      RECT 30.934 29.158 30.986 29.194 ;
      RECT 30.934 30.358 30.986 30.394 ;
      RECT 30.934 31.558 30.986 31.594 ;
      RECT 30.934 33.342 30.986 33.378 ;
      RECT 30.934 33.582 30.986 33.618 ;
      RECT 30.934 37.902 30.986 37.938 ;
      RECT 30.934 38.142 30.986 38.178 ;
      RECT 30.934 40.678 30.986 40.714 ;
      RECT 30.934 41.878 30.986 41.914 ;
      RECT 30.934 43.078 30.986 43.114 ;
      RECT 30.934 44.278 30.986 44.314 ;
      RECT 30.934 45.478 30.986 45.514 ;
      RECT 30.934 46.678 30.986 46.714 ;
      RECT 30.934 47.878 30.986 47.914 ;
      RECT 30.934 49.078 30.986 49.114 ;
      RECT 30.934 50.278 30.986 50.314 ;
      RECT 30.934 51.478 30.986 51.514 ;
      RECT 30.934 52.678 30.986 52.714 ;
      RECT 30.934 53.878 30.986 53.914 ;
      RECT 30.934 55.078 30.986 55.114 ;
      RECT 30.934 56.278 30.986 56.314 ;
      RECT 30.934 57.478 30.986 57.514 ;
      RECT 30.934 58.678 30.986 58.714 ;
      RECT 30.934 59.878 30.986 59.914 ;
      RECT 30.934 61.078 30.986 61.114 ;
      RECT 30.934 62.278 30.986 62.314 ;
      RECT 30.934 63.478 30.986 63.514 ;
      RECT 30.934 64.678 30.986 64.714 ;
      RECT 30.934 65.878 30.986 65.914 ;
      RECT 30.934 67.078 30.986 67.114 ;
      RECT 30.934 68.278 30.986 68.314 ;
      RECT 30.934 69.478 30.986 69.514 ;
      RECT 30.934 70.678 30.986 70.714 ;
      RECT 30.934 71.878 30.986 71.914 ;
      RECT 31.014 0.806 31.066 0.842 ;
      RECT 31.014 2.006 31.066 2.042 ;
      RECT 31.014 3.206 31.066 3.242 ;
      RECT 31.014 4.406 31.066 4.442 ;
      RECT 31.014 5.606 31.066 5.642 ;
      RECT 31.014 6.806 31.066 6.842 ;
      RECT 31.014 8.006 31.066 8.042 ;
      RECT 31.014 9.206 31.066 9.242 ;
      RECT 31.014 10.406 31.066 10.442 ;
      RECT 31.014 11.606 31.066 11.642 ;
      RECT 31.014 12.806 31.066 12.842 ;
      RECT 31.014 14.006 31.066 14.042 ;
      RECT 31.014 15.206 31.066 15.242 ;
      RECT 31.014 16.406 31.066 16.442 ;
      RECT 31.014 17.606 31.066 17.642 ;
      RECT 31.014 18.806 31.066 18.842 ;
      RECT 31.014 20.006 31.066 20.042 ;
      RECT 31.014 21.206 31.066 21.242 ;
      RECT 31.014 22.406 31.066 22.442 ;
      RECT 31.014 23.606 31.066 23.642 ;
      RECT 31.014 24.806 31.066 24.842 ;
      RECT 31.014 26.006 31.066 26.042 ;
      RECT 31.014 27.206 31.066 27.242 ;
      RECT 31.014 28.406 31.066 28.442 ;
      RECT 31.014 29.606 31.066 29.642 ;
      RECT 31.014 30.806 31.066 30.842 ;
      RECT 31.014 32.622 31.066 32.658 ;
      RECT 31.014 32.862 31.066 32.898 ;
      RECT 31.014 38.622 31.066 38.658 ;
      RECT 31.014 38.862 31.066 38.898 ;
      RECT 31.014 39.926 31.066 39.962 ;
      RECT 31.014 41.126 31.066 41.162 ;
      RECT 31.014 42.326 31.066 42.362 ;
      RECT 31.014 43.526 31.066 43.562 ;
      RECT 31.014 44.726 31.066 44.762 ;
      RECT 31.014 45.926 31.066 45.962 ;
      RECT 31.014 47.126 31.066 47.162 ;
      RECT 31.014 48.326 31.066 48.362 ;
      RECT 31.014 49.526 31.066 49.562 ;
      RECT 31.014 50.726 31.066 50.762 ;
      RECT 31.014 51.926 31.066 51.962 ;
      RECT 31.014 53.126 31.066 53.162 ;
      RECT 31.014 54.326 31.066 54.362 ;
      RECT 31.014 55.526 31.066 55.562 ;
      RECT 31.014 56.726 31.066 56.762 ;
      RECT 31.014 57.926 31.066 57.962 ;
      RECT 31.014 59.126 31.066 59.162 ;
      RECT 31.014 60.326 31.066 60.362 ;
      RECT 31.014 61.526 31.066 61.562 ;
      RECT 31.014 62.726 31.066 62.762 ;
      RECT 31.014 63.926 31.066 63.962 ;
      RECT 31.014 65.126 31.066 65.162 ;
      RECT 31.014 66.326 31.066 66.362 ;
      RECT 31.014 67.526 31.066 67.562 ;
      RECT 31.014 68.726 31.066 68.762 ;
      RECT 31.014 69.926 31.066 69.962 ;
      RECT 31.014 71.126 31.066 71.162 ;
      RECT 31.094 1.558 31.146 1.594 ;
      RECT 31.094 2.758 31.146 2.794 ;
      RECT 31.094 3.958 31.146 3.994 ;
      RECT 31.094 5.158 31.146 5.194 ;
      RECT 31.094 6.358 31.146 6.394 ;
      RECT 31.094 7.558 31.146 7.594 ;
      RECT 31.094 8.758 31.146 8.794 ;
      RECT 31.094 9.958 31.146 9.994 ;
      RECT 31.094 11.158 31.146 11.194 ;
      RECT 31.094 12.358 31.146 12.394 ;
      RECT 31.094 13.558 31.146 13.594 ;
      RECT 31.094 14.758 31.146 14.794 ;
      RECT 31.094 15.958 31.146 15.994 ;
      RECT 31.094 17.158 31.146 17.194 ;
      RECT 31.094 18.358 31.146 18.394 ;
      RECT 31.094 19.558 31.146 19.594 ;
      RECT 31.094 20.758 31.146 20.794 ;
      RECT 31.094 21.958 31.146 21.994 ;
      RECT 31.094 23.158 31.146 23.194 ;
      RECT 31.094 24.358 31.146 24.394 ;
      RECT 31.094 25.558 31.146 25.594 ;
      RECT 31.094 26.758 31.146 26.794 ;
      RECT 31.094 27.958 31.146 27.994 ;
      RECT 31.094 29.158 31.146 29.194 ;
      RECT 31.094 30.358 31.146 30.394 ;
      RECT 31.094 31.558 31.146 31.594 ;
      RECT 31.094 33.342 31.146 33.378 ;
      RECT 31.094 33.582 31.146 33.618 ;
      RECT 31.094 37.902 31.146 37.938 ;
      RECT 31.094 38.142 31.146 38.178 ;
      RECT 31.094 40.678 31.146 40.714 ;
      RECT 31.094 41.878 31.146 41.914 ;
      RECT 31.094 43.078 31.146 43.114 ;
      RECT 31.094 44.278 31.146 44.314 ;
      RECT 31.094 45.478 31.146 45.514 ;
      RECT 31.094 46.678 31.146 46.714 ;
      RECT 31.094 47.878 31.146 47.914 ;
      RECT 31.094 49.078 31.146 49.114 ;
      RECT 31.094 50.278 31.146 50.314 ;
      RECT 31.094 51.478 31.146 51.514 ;
      RECT 31.094 52.678 31.146 52.714 ;
      RECT 31.094 53.878 31.146 53.914 ;
      RECT 31.094 55.078 31.146 55.114 ;
      RECT 31.094 56.278 31.146 56.314 ;
      RECT 31.094 57.478 31.146 57.514 ;
      RECT 31.094 58.678 31.146 58.714 ;
      RECT 31.094 59.878 31.146 59.914 ;
      RECT 31.094 61.078 31.146 61.114 ;
      RECT 31.094 62.278 31.146 62.314 ;
      RECT 31.094 63.478 31.146 63.514 ;
      RECT 31.094 64.678 31.146 64.714 ;
      RECT 31.094 65.878 31.146 65.914 ;
      RECT 31.094 67.078 31.146 67.114 ;
      RECT 31.094 68.278 31.146 68.314 ;
      RECT 31.094 69.478 31.146 69.514 ;
      RECT 31.094 70.678 31.146 70.714 ;
      RECT 31.094 71.878 31.146 71.914 ;
      RECT 31.174 0.281 31.226 0.317 ;
      RECT 31.174 72.403 31.226 72.439 ;
      RECT 31.254 0.806 31.306 0.842 ;
      RECT 31.254 2.006 31.306 2.042 ;
      RECT 31.254 3.206 31.306 3.242 ;
      RECT 31.254 4.406 31.306 4.442 ;
      RECT 31.254 5.606 31.306 5.642 ;
      RECT 31.254 6.806 31.306 6.842 ;
      RECT 31.254 8.006 31.306 8.042 ;
      RECT 31.254 9.206 31.306 9.242 ;
      RECT 31.254 10.406 31.306 10.442 ;
      RECT 31.254 11.606 31.306 11.642 ;
      RECT 31.254 12.806 31.306 12.842 ;
      RECT 31.254 14.006 31.306 14.042 ;
      RECT 31.254 15.206 31.306 15.242 ;
      RECT 31.254 16.406 31.306 16.442 ;
      RECT 31.254 17.606 31.306 17.642 ;
      RECT 31.254 18.806 31.306 18.842 ;
      RECT 31.254 20.006 31.306 20.042 ;
      RECT 31.254 21.206 31.306 21.242 ;
      RECT 31.254 22.406 31.306 22.442 ;
      RECT 31.254 23.606 31.306 23.642 ;
      RECT 31.254 24.806 31.306 24.842 ;
      RECT 31.254 26.006 31.306 26.042 ;
      RECT 31.254 27.206 31.306 27.242 ;
      RECT 31.254 28.406 31.306 28.442 ;
      RECT 31.254 29.606 31.306 29.642 ;
      RECT 31.254 30.806 31.306 30.842 ;
      RECT 31.254 32.622 31.306 32.658 ;
      RECT 31.254 32.862 31.306 32.898 ;
      RECT 31.254 34.302 31.306 34.338 ;
      RECT 31.254 34.782 31.306 34.818 ;
      RECT 31.254 36.702 31.306 36.738 ;
      RECT 31.254 37.182 31.306 37.218 ;
      RECT 31.254 38.622 31.306 38.658 ;
      RECT 31.254 38.862 31.306 38.898 ;
      RECT 31.254 39.926 31.306 39.962 ;
      RECT 31.254 41.126 31.306 41.162 ;
      RECT 31.254 42.326 31.306 42.362 ;
      RECT 31.254 43.526 31.306 43.562 ;
      RECT 31.254 44.726 31.306 44.762 ;
      RECT 31.254 45.926 31.306 45.962 ;
      RECT 31.254 47.126 31.306 47.162 ;
      RECT 31.254 48.326 31.306 48.362 ;
      RECT 31.254 49.526 31.306 49.562 ;
      RECT 31.254 50.726 31.306 50.762 ;
      RECT 31.254 51.926 31.306 51.962 ;
      RECT 31.254 53.126 31.306 53.162 ;
      RECT 31.254 54.326 31.306 54.362 ;
      RECT 31.254 55.526 31.306 55.562 ;
      RECT 31.254 56.726 31.306 56.762 ;
      RECT 31.254 57.926 31.306 57.962 ;
      RECT 31.254 59.126 31.306 59.162 ;
      RECT 31.254 60.326 31.306 60.362 ;
      RECT 31.254 61.526 31.306 61.562 ;
      RECT 31.254 62.726 31.306 62.762 ;
      RECT 31.254 63.926 31.306 63.962 ;
      RECT 31.254 65.126 31.306 65.162 ;
      RECT 31.254 66.326 31.306 66.362 ;
      RECT 31.254 67.526 31.306 67.562 ;
      RECT 31.254 68.726 31.306 68.762 ;
      RECT 31.254 69.926 31.306 69.962 ;
      RECT 31.254 71.126 31.306 71.162 ;
      RECT 31.334 1.558 31.386 1.594 ;
      RECT 31.334 2.758 31.386 2.794 ;
      RECT 31.334 3.958 31.386 3.994 ;
      RECT 31.334 5.158 31.386 5.194 ;
      RECT 31.334 6.358 31.386 6.394 ;
      RECT 31.334 7.558 31.386 7.594 ;
      RECT 31.334 8.758 31.386 8.794 ;
      RECT 31.334 9.958 31.386 9.994 ;
      RECT 31.334 11.158 31.386 11.194 ;
      RECT 31.334 12.358 31.386 12.394 ;
      RECT 31.334 13.558 31.386 13.594 ;
      RECT 31.334 14.758 31.386 14.794 ;
      RECT 31.334 15.958 31.386 15.994 ;
      RECT 31.334 17.158 31.386 17.194 ;
      RECT 31.334 18.358 31.386 18.394 ;
      RECT 31.334 19.558 31.386 19.594 ;
      RECT 31.334 20.758 31.386 20.794 ;
      RECT 31.334 21.958 31.386 21.994 ;
      RECT 31.334 23.158 31.386 23.194 ;
      RECT 31.334 24.358 31.386 24.394 ;
      RECT 31.334 25.558 31.386 25.594 ;
      RECT 31.334 26.758 31.386 26.794 ;
      RECT 31.334 27.958 31.386 27.994 ;
      RECT 31.334 29.158 31.386 29.194 ;
      RECT 31.334 30.358 31.386 30.394 ;
      RECT 31.334 31.558 31.386 31.594 ;
      RECT 31.334 33.342 31.386 33.378 ;
      RECT 31.334 33.582 31.386 33.618 ;
      RECT 31.334 37.902 31.386 37.938 ;
      RECT 31.334 38.142 31.386 38.178 ;
      RECT 31.334 40.678 31.386 40.714 ;
      RECT 31.334 41.878 31.386 41.914 ;
      RECT 31.334 43.078 31.386 43.114 ;
      RECT 31.334 44.278 31.386 44.314 ;
      RECT 31.334 45.478 31.386 45.514 ;
      RECT 31.334 46.678 31.386 46.714 ;
      RECT 31.334 47.878 31.386 47.914 ;
      RECT 31.334 49.078 31.386 49.114 ;
      RECT 31.334 50.278 31.386 50.314 ;
      RECT 31.334 51.478 31.386 51.514 ;
      RECT 31.334 52.678 31.386 52.714 ;
      RECT 31.334 53.878 31.386 53.914 ;
      RECT 31.334 55.078 31.386 55.114 ;
      RECT 31.334 56.278 31.386 56.314 ;
      RECT 31.334 57.478 31.386 57.514 ;
      RECT 31.334 58.678 31.386 58.714 ;
      RECT 31.334 59.878 31.386 59.914 ;
      RECT 31.334 61.078 31.386 61.114 ;
      RECT 31.334 62.278 31.386 62.314 ;
      RECT 31.334 63.478 31.386 63.514 ;
      RECT 31.334 64.678 31.386 64.714 ;
      RECT 31.334 65.878 31.386 65.914 ;
      RECT 31.334 67.078 31.386 67.114 ;
      RECT 31.334 68.278 31.386 68.314 ;
      RECT 31.334 69.478 31.386 69.514 ;
      RECT 31.334 70.678 31.386 70.714 ;
      RECT 31.334 71.878 31.386 71.914 ;
      RECT 31.414 0.806 31.466 0.842 ;
      RECT 31.414 2.006 31.466 2.042 ;
      RECT 31.414 3.206 31.466 3.242 ;
      RECT 31.414 4.406 31.466 4.442 ;
      RECT 31.414 5.606 31.466 5.642 ;
      RECT 31.414 6.806 31.466 6.842 ;
      RECT 31.414 8.006 31.466 8.042 ;
      RECT 31.414 9.206 31.466 9.242 ;
      RECT 31.414 10.406 31.466 10.442 ;
      RECT 31.414 11.606 31.466 11.642 ;
      RECT 31.414 12.806 31.466 12.842 ;
      RECT 31.414 14.006 31.466 14.042 ;
      RECT 31.414 15.206 31.466 15.242 ;
      RECT 31.414 16.406 31.466 16.442 ;
      RECT 31.414 17.606 31.466 17.642 ;
      RECT 31.414 18.806 31.466 18.842 ;
      RECT 31.414 20.006 31.466 20.042 ;
      RECT 31.414 21.206 31.466 21.242 ;
      RECT 31.414 22.406 31.466 22.442 ;
      RECT 31.414 23.606 31.466 23.642 ;
      RECT 31.414 24.806 31.466 24.842 ;
      RECT 31.414 26.006 31.466 26.042 ;
      RECT 31.414 27.206 31.466 27.242 ;
      RECT 31.414 28.406 31.466 28.442 ;
      RECT 31.414 29.606 31.466 29.642 ;
      RECT 31.414 30.806 31.466 30.842 ;
      RECT 31.414 32.622 31.466 32.658 ;
      RECT 31.414 32.862 31.466 32.898 ;
      RECT 31.414 38.622 31.466 38.658 ;
      RECT 31.414 38.862 31.466 38.898 ;
      RECT 31.414 39.926 31.466 39.962 ;
      RECT 31.414 41.126 31.466 41.162 ;
      RECT 31.414 42.326 31.466 42.362 ;
      RECT 31.414 43.526 31.466 43.562 ;
      RECT 31.414 44.726 31.466 44.762 ;
      RECT 31.414 45.926 31.466 45.962 ;
      RECT 31.414 47.126 31.466 47.162 ;
      RECT 31.414 48.326 31.466 48.362 ;
      RECT 31.414 49.526 31.466 49.562 ;
      RECT 31.414 50.726 31.466 50.762 ;
      RECT 31.414 51.926 31.466 51.962 ;
      RECT 31.414 53.126 31.466 53.162 ;
      RECT 31.414 54.326 31.466 54.362 ;
      RECT 31.414 55.526 31.466 55.562 ;
      RECT 31.414 56.726 31.466 56.762 ;
      RECT 31.414 57.926 31.466 57.962 ;
      RECT 31.414 59.126 31.466 59.162 ;
      RECT 31.414 60.326 31.466 60.362 ;
      RECT 31.414 61.526 31.466 61.562 ;
      RECT 31.414 62.726 31.466 62.762 ;
      RECT 31.414 63.926 31.466 63.962 ;
      RECT 31.414 65.126 31.466 65.162 ;
      RECT 31.414 66.326 31.466 66.362 ;
      RECT 31.414 67.526 31.466 67.562 ;
      RECT 31.414 68.726 31.466 68.762 ;
      RECT 31.414 69.926 31.466 69.962 ;
      RECT 31.414 71.126 31.466 71.162 ;
      RECT 31.494 1.558 31.546 1.594 ;
      RECT 31.494 2.758 31.546 2.794 ;
      RECT 31.494 3.958 31.546 3.994 ;
      RECT 31.494 5.158 31.546 5.194 ;
      RECT 31.494 6.358 31.546 6.394 ;
      RECT 31.494 7.558 31.546 7.594 ;
      RECT 31.494 8.758 31.546 8.794 ;
      RECT 31.494 9.958 31.546 9.994 ;
      RECT 31.494 11.158 31.546 11.194 ;
      RECT 31.494 12.358 31.546 12.394 ;
      RECT 31.494 13.558 31.546 13.594 ;
      RECT 31.494 14.758 31.546 14.794 ;
      RECT 31.494 15.958 31.546 15.994 ;
      RECT 31.494 17.158 31.546 17.194 ;
      RECT 31.494 18.358 31.546 18.394 ;
      RECT 31.494 19.558 31.546 19.594 ;
      RECT 31.494 20.758 31.546 20.794 ;
      RECT 31.494 21.958 31.546 21.994 ;
      RECT 31.494 23.158 31.546 23.194 ;
      RECT 31.494 24.358 31.546 24.394 ;
      RECT 31.494 25.558 31.546 25.594 ;
      RECT 31.494 26.758 31.546 26.794 ;
      RECT 31.494 27.958 31.546 27.994 ;
      RECT 31.494 29.158 31.546 29.194 ;
      RECT 31.494 30.358 31.546 30.394 ;
      RECT 31.494 31.558 31.546 31.594 ;
      RECT 31.494 33.342 31.546 33.378 ;
      RECT 31.494 33.582 31.546 33.618 ;
      RECT 31.494 37.902 31.546 37.938 ;
      RECT 31.494 38.142 31.546 38.178 ;
      RECT 31.494 40.678 31.546 40.714 ;
      RECT 31.494 41.878 31.546 41.914 ;
      RECT 31.494 43.078 31.546 43.114 ;
      RECT 31.494 44.278 31.546 44.314 ;
      RECT 31.494 45.478 31.546 45.514 ;
      RECT 31.494 46.678 31.546 46.714 ;
      RECT 31.494 47.878 31.546 47.914 ;
      RECT 31.494 49.078 31.546 49.114 ;
      RECT 31.494 50.278 31.546 50.314 ;
      RECT 31.494 51.478 31.546 51.514 ;
      RECT 31.494 52.678 31.546 52.714 ;
      RECT 31.494 53.878 31.546 53.914 ;
      RECT 31.494 55.078 31.546 55.114 ;
      RECT 31.494 56.278 31.546 56.314 ;
      RECT 31.494 57.478 31.546 57.514 ;
      RECT 31.494 58.678 31.546 58.714 ;
      RECT 31.494 59.878 31.546 59.914 ;
      RECT 31.494 61.078 31.546 61.114 ;
      RECT 31.494 62.278 31.546 62.314 ;
      RECT 31.494 63.478 31.546 63.514 ;
      RECT 31.494 64.678 31.546 64.714 ;
      RECT 31.494 65.878 31.546 65.914 ;
      RECT 31.494 67.078 31.546 67.114 ;
      RECT 31.494 68.278 31.546 68.314 ;
      RECT 31.494 69.478 31.546 69.514 ;
      RECT 31.494 70.678 31.546 70.714 ;
      RECT 31.494 71.878 31.546 71.914 ;
      RECT 31.574 0.281 31.626 0.317 ;
      RECT 31.574 72.403 31.626 72.439 ;
      RECT 31.654 0.806 31.706 0.842 ;
      RECT 31.654 2.006 31.706 2.042 ;
      RECT 31.654 3.206 31.706 3.242 ;
      RECT 31.654 4.406 31.706 4.442 ;
      RECT 31.654 5.606 31.706 5.642 ;
      RECT 31.654 6.806 31.706 6.842 ;
      RECT 31.654 8.006 31.706 8.042 ;
      RECT 31.654 9.206 31.706 9.242 ;
      RECT 31.654 10.406 31.706 10.442 ;
      RECT 31.654 11.606 31.706 11.642 ;
      RECT 31.654 12.806 31.706 12.842 ;
      RECT 31.654 14.006 31.706 14.042 ;
      RECT 31.654 15.206 31.706 15.242 ;
      RECT 31.654 16.406 31.706 16.442 ;
      RECT 31.654 17.606 31.706 17.642 ;
      RECT 31.654 18.806 31.706 18.842 ;
      RECT 31.654 20.006 31.706 20.042 ;
      RECT 31.654 21.206 31.706 21.242 ;
      RECT 31.654 22.406 31.706 22.442 ;
      RECT 31.654 23.606 31.706 23.642 ;
      RECT 31.654 24.806 31.706 24.842 ;
      RECT 31.654 26.006 31.706 26.042 ;
      RECT 31.654 27.206 31.706 27.242 ;
      RECT 31.654 28.406 31.706 28.442 ;
      RECT 31.654 29.606 31.706 29.642 ;
      RECT 31.654 30.806 31.706 30.842 ;
      RECT 31.654 32.622 31.706 32.658 ;
      RECT 31.654 32.862 31.706 32.898 ;
      RECT 31.654 38.622 31.706 38.658 ;
      RECT 31.654 38.862 31.706 38.898 ;
      RECT 31.654 39.926 31.706 39.962 ;
      RECT 31.654 41.126 31.706 41.162 ;
      RECT 31.654 42.326 31.706 42.362 ;
      RECT 31.654 43.526 31.706 43.562 ;
      RECT 31.654 44.726 31.706 44.762 ;
      RECT 31.654 45.926 31.706 45.962 ;
      RECT 31.654 47.126 31.706 47.162 ;
      RECT 31.654 48.326 31.706 48.362 ;
      RECT 31.654 49.526 31.706 49.562 ;
      RECT 31.654 50.726 31.706 50.762 ;
      RECT 31.654 51.926 31.706 51.962 ;
      RECT 31.654 53.126 31.706 53.162 ;
      RECT 31.654 54.326 31.706 54.362 ;
      RECT 31.654 55.526 31.706 55.562 ;
      RECT 31.654 56.726 31.706 56.762 ;
      RECT 31.654 57.926 31.706 57.962 ;
      RECT 31.654 59.126 31.706 59.162 ;
      RECT 31.654 60.326 31.706 60.362 ;
      RECT 31.654 61.526 31.706 61.562 ;
      RECT 31.654 62.726 31.706 62.762 ;
      RECT 31.654 63.926 31.706 63.962 ;
      RECT 31.654 65.126 31.706 65.162 ;
      RECT 31.654 66.326 31.706 66.362 ;
      RECT 31.654 67.526 31.706 67.562 ;
      RECT 31.654 68.726 31.706 68.762 ;
      RECT 31.654 69.926 31.706 69.962 ;
      RECT 31.654 71.126 31.706 71.162 ;
      RECT 31.734 1.558 31.786 1.594 ;
      RECT 31.734 2.758 31.786 2.794 ;
      RECT 31.734 3.958 31.786 3.994 ;
      RECT 31.734 5.158 31.786 5.194 ;
      RECT 31.734 6.358 31.786 6.394 ;
      RECT 31.734 7.558 31.786 7.594 ;
      RECT 31.734 8.758 31.786 8.794 ;
      RECT 31.734 9.958 31.786 9.994 ;
      RECT 31.734 11.158 31.786 11.194 ;
      RECT 31.734 12.358 31.786 12.394 ;
      RECT 31.734 13.558 31.786 13.594 ;
      RECT 31.734 14.758 31.786 14.794 ;
      RECT 31.734 15.958 31.786 15.994 ;
      RECT 31.734 17.158 31.786 17.194 ;
      RECT 31.734 18.358 31.786 18.394 ;
      RECT 31.734 19.558 31.786 19.594 ;
      RECT 31.734 20.758 31.786 20.794 ;
      RECT 31.734 21.958 31.786 21.994 ;
      RECT 31.734 23.158 31.786 23.194 ;
      RECT 31.734 24.358 31.786 24.394 ;
      RECT 31.734 25.558 31.786 25.594 ;
      RECT 31.734 26.758 31.786 26.794 ;
      RECT 31.734 27.958 31.786 27.994 ;
      RECT 31.734 29.158 31.786 29.194 ;
      RECT 31.734 30.358 31.786 30.394 ;
      RECT 31.734 31.558 31.786 31.594 ;
      RECT 31.734 33.342 31.786 33.378 ;
      RECT 31.734 33.582 31.786 33.618 ;
      RECT 31.734 37.902 31.786 37.938 ;
      RECT 31.734 38.142 31.786 38.178 ;
      RECT 31.734 40.678 31.786 40.714 ;
      RECT 31.734 41.878 31.786 41.914 ;
      RECT 31.734 43.078 31.786 43.114 ;
      RECT 31.734 44.278 31.786 44.314 ;
      RECT 31.734 45.478 31.786 45.514 ;
      RECT 31.734 46.678 31.786 46.714 ;
      RECT 31.734 47.878 31.786 47.914 ;
      RECT 31.734 49.078 31.786 49.114 ;
      RECT 31.734 50.278 31.786 50.314 ;
      RECT 31.734 51.478 31.786 51.514 ;
      RECT 31.734 52.678 31.786 52.714 ;
      RECT 31.734 53.878 31.786 53.914 ;
      RECT 31.734 55.078 31.786 55.114 ;
      RECT 31.734 56.278 31.786 56.314 ;
      RECT 31.734 57.478 31.786 57.514 ;
      RECT 31.734 58.678 31.786 58.714 ;
      RECT 31.734 59.878 31.786 59.914 ;
      RECT 31.734 61.078 31.786 61.114 ;
      RECT 31.734 62.278 31.786 62.314 ;
      RECT 31.734 63.478 31.786 63.514 ;
      RECT 31.734 64.678 31.786 64.714 ;
      RECT 31.734 65.878 31.786 65.914 ;
      RECT 31.734 67.078 31.786 67.114 ;
      RECT 31.734 68.278 31.786 68.314 ;
      RECT 31.734 69.478 31.786 69.514 ;
      RECT 31.734 70.678 31.786 70.714 ;
      RECT 31.734 71.878 31.786 71.914 ;
      RECT 31.814 0.806 31.866 0.842 ;
      RECT 31.814 2.006 31.866 2.042 ;
      RECT 31.814 3.206 31.866 3.242 ;
      RECT 31.814 4.406 31.866 4.442 ;
      RECT 31.814 5.606 31.866 5.642 ;
      RECT 31.814 6.806 31.866 6.842 ;
      RECT 31.814 8.006 31.866 8.042 ;
      RECT 31.814 9.206 31.866 9.242 ;
      RECT 31.814 10.406 31.866 10.442 ;
      RECT 31.814 11.606 31.866 11.642 ;
      RECT 31.814 12.806 31.866 12.842 ;
      RECT 31.814 14.006 31.866 14.042 ;
      RECT 31.814 15.206 31.866 15.242 ;
      RECT 31.814 16.406 31.866 16.442 ;
      RECT 31.814 17.606 31.866 17.642 ;
      RECT 31.814 18.806 31.866 18.842 ;
      RECT 31.814 20.006 31.866 20.042 ;
      RECT 31.814 21.206 31.866 21.242 ;
      RECT 31.814 22.406 31.866 22.442 ;
      RECT 31.814 23.606 31.866 23.642 ;
      RECT 31.814 24.806 31.866 24.842 ;
      RECT 31.814 26.006 31.866 26.042 ;
      RECT 31.814 27.206 31.866 27.242 ;
      RECT 31.814 28.406 31.866 28.442 ;
      RECT 31.814 29.606 31.866 29.642 ;
      RECT 31.814 30.806 31.866 30.842 ;
      RECT 31.814 32.622 31.866 32.658 ;
      RECT 31.814 32.862 31.866 32.898 ;
      RECT 31.814 38.622 31.866 38.658 ;
      RECT 31.814 38.862 31.866 38.898 ;
      RECT 31.814 39.926 31.866 39.962 ;
      RECT 31.814 41.126 31.866 41.162 ;
      RECT 31.814 42.326 31.866 42.362 ;
      RECT 31.814 43.526 31.866 43.562 ;
      RECT 31.814 44.726 31.866 44.762 ;
      RECT 31.814 45.926 31.866 45.962 ;
      RECT 31.814 47.126 31.866 47.162 ;
      RECT 31.814 48.326 31.866 48.362 ;
      RECT 31.814 49.526 31.866 49.562 ;
      RECT 31.814 50.726 31.866 50.762 ;
      RECT 31.814 51.926 31.866 51.962 ;
      RECT 31.814 53.126 31.866 53.162 ;
      RECT 31.814 54.326 31.866 54.362 ;
      RECT 31.814 55.526 31.866 55.562 ;
      RECT 31.814 56.726 31.866 56.762 ;
      RECT 31.814 57.926 31.866 57.962 ;
      RECT 31.814 59.126 31.866 59.162 ;
      RECT 31.814 60.326 31.866 60.362 ;
      RECT 31.814 61.526 31.866 61.562 ;
      RECT 31.814 62.726 31.866 62.762 ;
      RECT 31.814 63.926 31.866 63.962 ;
      RECT 31.814 65.126 31.866 65.162 ;
      RECT 31.814 66.326 31.866 66.362 ;
      RECT 31.814 67.526 31.866 67.562 ;
      RECT 31.814 68.726 31.866 68.762 ;
      RECT 31.814 69.926 31.866 69.962 ;
      RECT 31.814 71.126 31.866 71.162 ;
      RECT 31.894 1.558 31.946 1.594 ;
      RECT 31.894 2.758 31.946 2.794 ;
      RECT 31.894 3.958 31.946 3.994 ;
      RECT 31.894 5.158 31.946 5.194 ;
      RECT 31.894 6.358 31.946 6.394 ;
      RECT 31.894 7.558 31.946 7.594 ;
      RECT 31.894 8.758 31.946 8.794 ;
      RECT 31.894 9.958 31.946 9.994 ;
      RECT 31.894 11.158 31.946 11.194 ;
      RECT 31.894 12.358 31.946 12.394 ;
      RECT 31.894 13.558 31.946 13.594 ;
      RECT 31.894 14.758 31.946 14.794 ;
      RECT 31.894 15.958 31.946 15.994 ;
      RECT 31.894 17.158 31.946 17.194 ;
      RECT 31.894 18.358 31.946 18.394 ;
      RECT 31.894 19.558 31.946 19.594 ;
      RECT 31.894 20.758 31.946 20.794 ;
      RECT 31.894 21.958 31.946 21.994 ;
      RECT 31.894 23.158 31.946 23.194 ;
      RECT 31.894 24.358 31.946 24.394 ;
      RECT 31.894 25.558 31.946 25.594 ;
      RECT 31.894 26.758 31.946 26.794 ;
      RECT 31.894 27.958 31.946 27.994 ;
      RECT 31.894 29.158 31.946 29.194 ;
      RECT 31.894 30.358 31.946 30.394 ;
      RECT 31.894 31.558 31.946 31.594 ;
      RECT 31.894 33.342 31.946 33.378 ;
      RECT 31.894 33.582 31.946 33.618 ;
      RECT 31.894 37.902 31.946 37.938 ;
      RECT 31.894 38.142 31.946 38.178 ;
      RECT 31.894 40.678 31.946 40.714 ;
      RECT 31.894 41.878 31.946 41.914 ;
      RECT 31.894 43.078 31.946 43.114 ;
      RECT 31.894 44.278 31.946 44.314 ;
      RECT 31.894 45.478 31.946 45.514 ;
      RECT 31.894 46.678 31.946 46.714 ;
      RECT 31.894 47.878 31.946 47.914 ;
      RECT 31.894 49.078 31.946 49.114 ;
      RECT 31.894 50.278 31.946 50.314 ;
      RECT 31.894 51.478 31.946 51.514 ;
      RECT 31.894 52.678 31.946 52.714 ;
      RECT 31.894 53.878 31.946 53.914 ;
      RECT 31.894 55.078 31.946 55.114 ;
      RECT 31.894 56.278 31.946 56.314 ;
      RECT 31.894 57.478 31.946 57.514 ;
      RECT 31.894 58.678 31.946 58.714 ;
      RECT 31.894 59.878 31.946 59.914 ;
      RECT 31.894 61.078 31.946 61.114 ;
      RECT 31.894 62.278 31.946 62.314 ;
      RECT 31.894 63.478 31.946 63.514 ;
      RECT 31.894 64.678 31.946 64.714 ;
      RECT 31.894 65.878 31.946 65.914 ;
      RECT 31.894 67.078 31.946 67.114 ;
      RECT 31.894 68.278 31.946 68.314 ;
      RECT 31.894 69.478 31.946 69.514 ;
      RECT 31.894 70.678 31.946 70.714 ;
      RECT 31.894 71.878 31.946 71.914 ;
      RECT 31.974 0.281 32.026 0.317 ;
      RECT 31.974 72.403 32.026 72.439 ;
      RECT 32.054 0.806 32.106 0.842 ;
      RECT 32.054 2.006 32.106 2.042 ;
      RECT 32.054 3.206 32.106 3.242 ;
      RECT 32.054 4.406 32.106 4.442 ;
      RECT 32.054 5.606 32.106 5.642 ;
      RECT 32.054 6.806 32.106 6.842 ;
      RECT 32.054 8.006 32.106 8.042 ;
      RECT 32.054 9.206 32.106 9.242 ;
      RECT 32.054 10.406 32.106 10.442 ;
      RECT 32.054 11.606 32.106 11.642 ;
      RECT 32.054 12.806 32.106 12.842 ;
      RECT 32.054 14.006 32.106 14.042 ;
      RECT 32.054 15.206 32.106 15.242 ;
      RECT 32.054 16.406 32.106 16.442 ;
      RECT 32.054 17.606 32.106 17.642 ;
      RECT 32.054 18.806 32.106 18.842 ;
      RECT 32.054 20.006 32.106 20.042 ;
      RECT 32.054 21.206 32.106 21.242 ;
      RECT 32.054 22.406 32.106 22.442 ;
      RECT 32.054 23.606 32.106 23.642 ;
      RECT 32.054 24.806 32.106 24.842 ;
      RECT 32.054 26.006 32.106 26.042 ;
      RECT 32.054 27.206 32.106 27.242 ;
      RECT 32.054 28.406 32.106 28.442 ;
      RECT 32.054 29.606 32.106 29.642 ;
      RECT 32.054 30.806 32.106 30.842 ;
      RECT 32.054 32.622 32.106 32.658 ;
      RECT 32.054 32.862 32.106 32.898 ;
      RECT 32.054 34.302 32.106 34.338 ;
      RECT 32.054 34.782 32.106 34.818 ;
      RECT 32.054 36.702 32.106 36.738 ;
      RECT 32.054 37.182 32.106 37.218 ;
      RECT 32.054 38.622 32.106 38.658 ;
      RECT 32.054 38.862 32.106 38.898 ;
      RECT 32.054 39.926 32.106 39.962 ;
      RECT 32.054 41.126 32.106 41.162 ;
      RECT 32.054 42.326 32.106 42.362 ;
      RECT 32.054 43.526 32.106 43.562 ;
      RECT 32.054 44.726 32.106 44.762 ;
      RECT 32.054 45.926 32.106 45.962 ;
      RECT 32.054 47.126 32.106 47.162 ;
      RECT 32.054 48.326 32.106 48.362 ;
      RECT 32.054 49.526 32.106 49.562 ;
      RECT 32.054 50.726 32.106 50.762 ;
      RECT 32.054 51.926 32.106 51.962 ;
      RECT 32.054 53.126 32.106 53.162 ;
      RECT 32.054 54.326 32.106 54.362 ;
      RECT 32.054 55.526 32.106 55.562 ;
      RECT 32.054 56.726 32.106 56.762 ;
      RECT 32.054 57.926 32.106 57.962 ;
      RECT 32.054 59.126 32.106 59.162 ;
      RECT 32.054 60.326 32.106 60.362 ;
      RECT 32.054 61.526 32.106 61.562 ;
      RECT 32.054 62.726 32.106 62.762 ;
      RECT 32.054 63.926 32.106 63.962 ;
      RECT 32.054 65.126 32.106 65.162 ;
      RECT 32.054 66.326 32.106 66.362 ;
      RECT 32.054 67.526 32.106 67.562 ;
      RECT 32.054 68.726 32.106 68.762 ;
      RECT 32.054 69.926 32.106 69.962 ;
      RECT 32.054 71.126 32.106 71.162 ;
      RECT 32.134 1.558 32.186 1.594 ;
      RECT 32.134 2.758 32.186 2.794 ;
      RECT 32.134 3.958 32.186 3.994 ;
      RECT 32.134 5.158 32.186 5.194 ;
      RECT 32.134 6.358 32.186 6.394 ;
      RECT 32.134 7.558 32.186 7.594 ;
      RECT 32.134 8.758 32.186 8.794 ;
      RECT 32.134 9.958 32.186 9.994 ;
      RECT 32.134 11.158 32.186 11.194 ;
      RECT 32.134 12.358 32.186 12.394 ;
      RECT 32.134 13.558 32.186 13.594 ;
      RECT 32.134 14.758 32.186 14.794 ;
      RECT 32.134 15.958 32.186 15.994 ;
      RECT 32.134 17.158 32.186 17.194 ;
      RECT 32.134 18.358 32.186 18.394 ;
      RECT 32.134 19.558 32.186 19.594 ;
      RECT 32.134 20.758 32.186 20.794 ;
      RECT 32.134 21.958 32.186 21.994 ;
      RECT 32.134 23.158 32.186 23.194 ;
      RECT 32.134 24.358 32.186 24.394 ;
      RECT 32.134 25.558 32.186 25.594 ;
      RECT 32.134 26.758 32.186 26.794 ;
      RECT 32.134 27.958 32.186 27.994 ;
      RECT 32.134 29.158 32.186 29.194 ;
      RECT 32.134 30.358 32.186 30.394 ;
      RECT 32.134 31.558 32.186 31.594 ;
      RECT 32.134 33.342 32.186 33.378 ;
      RECT 32.134 33.582 32.186 33.618 ;
      RECT 32.134 37.902 32.186 37.938 ;
      RECT 32.134 38.142 32.186 38.178 ;
      RECT 32.134 40.678 32.186 40.714 ;
      RECT 32.134 41.878 32.186 41.914 ;
      RECT 32.134 43.078 32.186 43.114 ;
      RECT 32.134 44.278 32.186 44.314 ;
      RECT 32.134 45.478 32.186 45.514 ;
      RECT 32.134 46.678 32.186 46.714 ;
      RECT 32.134 47.878 32.186 47.914 ;
      RECT 32.134 49.078 32.186 49.114 ;
      RECT 32.134 50.278 32.186 50.314 ;
      RECT 32.134 51.478 32.186 51.514 ;
      RECT 32.134 52.678 32.186 52.714 ;
      RECT 32.134 53.878 32.186 53.914 ;
      RECT 32.134 55.078 32.186 55.114 ;
      RECT 32.134 56.278 32.186 56.314 ;
      RECT 32.134 57.478 32.186 57.514 ;
      RECT 32.134 58.678 32.186 58.714 ;
      RECT 32.134 59.878 32.186 59.914 ;
      RECT 32.134 61.078 32.186 61.114 ;
      RECT 32.134 62.278 32.186 62.314 ;
      RECT 32.134 63.478 32.186 63.514 ;
      RECT 32.134 64.678 32.186 64.714 ;
      RECT 32.134 65.878 32.186 65.914 ;
      RECT 32.134 67.078 32.186 67.114 ;
      RECT 32.134 68.278 32.186 68.314 ;
      RECT 32.134 69.478 32.186 69.514 ;
      RECT 32.134 70.678 32.186 70.714 ;
      RECT 32.134 71.878 32.186 71.914 ;
      RECT 32.214 0.806 32.266 0.842 ;
      RECT 32.214 2.006 32.266 2.042 ;
      RECT 32.214 3.206 32.266 3.242 ;
      RECT 32.214 4.406 32.266 4.442 ;
      RECT 32.214 5.606 32.266 5.642 ;
      RECT 32.214 6.806 32.266 6.842 ;
      RECT 32.214 8.006 32.266 8.042 ;
      RECT 32.214 9.206 32.266 9.242 ;
      RECT 32.214 10.406 32.266 10.442 ;
      RECT 32.214 11.606 32.266 11.642 ;
      RECT 32.214 12.806 32.266 12.842 ;
      RECT 32.214 14.006 32.266 14.042 ;
      RECT 32.214 15.206 32.266 15.242 ;
      RECT 32.214 16.406 32.266 16.442 ;
      RECT 32.214 17.606 32.266 17.642 ;
      RECT 32.214 18.806 32.266 18.842 ;
      RECT 32.214 20.006 32.266 20.042 ;
      RECT 32.214 21.206 32.266 21.242 ;
      RECT 32.214 22.406 32.266 22.442 ;
      RECT 32.214 23.606 32.266 23.642 ;
      RECT 32.214 24.806 32.266 24.842 ;
      RECT 32.214 26.006 32.266 26.042 ;
      RECT 32.214 27.206 32.266 27.242 ;
      RECT 32.214 28.406 32.266 28.442 ;
      RECT 32.214 29.606 32.266 29.642 ;
      RECT 32.214 30.806 32.266 30.842 ;
      RECT 32.214 32.622 32.266 32.658 ;
      RECT 32.214 32.862 32.266 32.898 ;
      RECT 32.214 38.622 32.266 38.658 ;
      RECT 32.214 38.862 32.266 38.898 ;
      RECT 32.214 39.926 32.266 39.962 ;
      RECT 32.214 41.126 32.266 41.162 ;
      RECT 32.214 42.326 32.266 42.362 ;
      RECT 32.214 43.526 32.266 43.562 ;
      RECT 32.214 44.726 32.266 44.762 ;
      RECT 32.214 45.926 32.266 45.962 ;
      RECT 32.214 47.126 32.266 47.162 ;
      RECT 32.214 48.326 32.266 48.362 ;
      RECT 32.214 49.526 32.266 49.562 ;
      RECT 32.214 50.726 32.266 50.762 ;
      RECT 32.214 51.926 32.266 51.962 ;
      RECT 32.214 53.126 32.266 53.162 ;
      RECT 32.214 54.326 32.266 54.362 ;
      RECT 32.214 55.526 32.266 55.562 ;
      RECT 32.214 56.726 32.266 56.762 ;
      RECT 32.214 57.926 32.266 57.962 ;
      RECT 32.214 59.126 32.266 59.162 ;
      RECT 32.214 60.326 32.266 60.362 ;
      RECT 32.214 61.526 32.266 61.562 ;
      RECT 32.214 62.726 32.266 62.762 ;
      RECT 32.214 63.926 32.266 63.962 ;
      RECT 32.214 65.126 32.266 65.162 ;
      RECT 32.214 66.326 32.266 66.362 ;
      RECT 32.214 67.526 32.266 67.562 ;
      RECT 32.214 68.726 32.266 68.762 ;
      RECT 32.214 69.926 32.266 69.962 ;
      RECT 32.214 71.126 32.266 71.162 ;
      RECT 32.294 1.558 32.346 1.594 ;
      RECT 32.294 2.758 32.346 2.794 ;
      RECT 32.294 3.958 32.346 3.994 ;
      RECT 32.294 5.158 32.346 5.194 ;
      RECT 32.294 6.358 32.346 6.394 ;
      RECT 32.294 7.558 32.346 7.594 ;
      RECT 32.294 8.758 32.346 8.794 ;
      RECT 32.294 9.958 32.346 9.994 ;
      RECT 32.294 11.158 32.346 11.194 ;
      RECT 32.294 12.358 32.346 12.394 ;
      RECT 32.294 13.558 32.346 13.594 ;
      RECT 32.294 14.758 32.346 14.794 ;
      RECT 32.294 15.958 32.346 15.994 ;
      RECT 32.294 17.158 32.346 17.194 ;
      RECT 32.294 18.358 32.346 18.394 ;
      RECT 32.294 19.558 32.346 19.594 ;
      RECT 32.294 20.758 32.346 20.794 ;
      RECT 32.294 21.958 32.346 21.994 ;
      RECT 32.294 23.158 32.346 23.194 ;
      RECT 32.294 24.358 32.346 24.394 ;
      RECT 32.294 25.558 32.346 25.594 ;
      RECT 32.294 26.758 32.346 26.794 ;
      RECT 32.294 27.958 32.346 27.994 ;
      RECT 32.294 29.158 32.346 29.194 ;
      RECT 32.294 30.358 32.346 30.394 ;
      RECT 32.294 31.558 32.346 31.594 ;
      RECT 32.294 33.342 32.346 33.378 ;
      RECT 32.294 33.582 32.346 33.618 ;
      RECT 32.294 37.902 32.346 37.938 ;
      RECT 32.294 38.142 32.346 38.178 ;
      RECT 32.294 40.678 32.346 40.714 ;
      RECT 32.294 41.878 32.346 41.914 ;
      RECT 32.294 43.078 32.346 43.114 ;
      RECT 32.294 44.278 32.346 44.314 ;
      RECT 32.294 45.478 32.346 45.514 ;
      RECT 32.294 46.678 32.346 46.714 ;
      RECT 32.294 47.878 32.346 47.914 ;
      RECT 32.294 49.078 32.346 49.114 ;
      RECT 32.294 50.278 32.346 50.314 ;
      RECT 32.294 51.478 32.346 51.514 ;
      RECT 32.294 52.678 32.346 52.714 ;
      RECT 32.294 53.878 32.346 53.914 ;
      RECT 32.294 55.078 32.346 55.114 ;
      RECT 32.294 56.278 32.346 56.314 ;
      RECT 32.294 57.478 32.346 57.514 ;
      RECT 32.294 58.678 32.346 58.714 ;
      RECT 32.294 59.878 32.346 59.914 ;
      RECT 32.294 61.078 32.346 61.114 ;
      RECT 32.294 62.278 32.346 62.314 ;
      RECT 32.294 63.478 32.346 63.514 ;
      RECT 32.294 64.678 32.346 64.714 ;
      RECT 32.294 65.878 32.346 65.914 ;
      RECT 32.294 67.078 32.346 67.114 ;
      RECT 32.294 68.278 32.346 68.314 ;
      RECT 32.294 69.478 32.346 69.514 ;
      RECT 32.294 70.678 32.346 70.714 ;
      RECT 32.294 71.878 32.346 71.914 ;
      RECT 32.374 0.281 32.426 0.317 ;
      RECT 32.374 72.403 32.426 72.439 ;
      RECT 32.454 0.806 32.506 0.842 ;
      RECT 32.454 2.006 32.506 2.042 ;
      RECT 32.454 3.206 32.506 3.242 ;
      RECT 32.454 4.406 32.506 4.442 ;
      RECT 32.454 5.606 32.506 5.642 ;
      RECT 32.454 6.806 32.506 6.842 ;
      RECT 32.454 8.006 32.506 8.042 ;
      RECT 32.454 9.206 32.506 9.242 ;
      RECT 32.454 10.406 32.506 10.442 ;
      RECT 32.454 11.606 32.506 11.642 ;
      RECT 32.454 12.806 32.506 12.842 ;
      RECT 32.454 14.006 32.506 14.042 ;
      RECT 32.454 15.206 32.506 15.242 ;
      RECT 32.454 16.406 32.506 16.442 ;
      RECT 32.454 17.606 32.506 17.642 ;
      RECT 32.454 18.806 32.506 18.842 ;
      RECT 32.454 20.006 32.506 20.042 ;
      RECT 32.454 21.206 32.506 21.242 ;
      RECT 32.454 22.406 32.506 22.442 ;
      RECT 32.454 23.606 32.506 23.642 ;
      RECT 32.454 24.806 32.506 24.842 ;
      RECT 32.454 26.006 32.506 26.042 ;
      RECT 32.454 27.206 32.506 27.242 ;
      RECT 32.454 28.406 32.506 28.442 ;
      RECT 32.454 29.606 32.506 29.642 ;
      RECT 32.454 30.806 32.506 30.842 ;
      RECT 32.454 32.622 32.506 32.658 ;
      RECT 32.454 32.862 32.506 32.898 ;
      RECT 32.454 38.622 32.506 38.658 ;
      RECT 32.454 38.862 32.506 38.898 ;
      RECT 32.454 39.926 32.506 39.962 ;
      RECT 32.454 41.126 32.506 41.162 ;
      RECT 32.454 42.326 32.506 42.362 ;
      RECT 32.454 43.526 32.506 43.562 ;
      RECT 32.454 44.726 32.506 44.762 ;
      RECT 32.454 45.926 32.506 45.962 ;
      RECT 32.454 47.126 32.506 47.162 ;
      RECT 32.454 48.326 32.506 48.362 ;
      RECT 32.454 49.526 32.506 49.562 ;
      RECT 32.454 50.726 32.506 50.762 ;
      RECT 32.454 51.926 32.506 51.962 ;
      RECT 32.454 53.126 32.506 53.162 ;
      RECT 32.454 54.326 32.506 54.362 ;
      RECT 32.454 55.526 32.506 55.562 ;
      RECT 32.454 56.726 32.506 56.762 ;
      RECT 32.454 57.926 32.506 57.962 ;
      RECT 32.454 59.126 32.506 59.162 ;
      RECT 32.454 60.326 32.506 60.362 ;
      RECT 32.454 61.526 32.506 61.562 ;
      RECT 32.454 62.726 32.506 62.762 ;
      RECT 32.454 63.926 32.506 63.962 ;
      RECT 32.454 65.126 32.506 65.162 ;
      RECT 32.454 66.326 32.506 66.362 ;
      RECT 32.454 67.526 32.506 67.562 ;
      RECT 32.454 68.726 32.506 68.762 ;
      RECT 32.454 69.926 32.506 69.962 ;
      RECT 32.454 71.126 32.506 71.162 ;
      RECT 32.534 1.558 32.586 1.594 ;
      RECT 32.534 2.758 32.586 2.794 ;
      RECT 32.534 3.958 32.586 3.994 ;
      RECT 32.534 5.158 32.586 5.194 ;
      RECT 32.534 6.358 32.586 6.394 ;
      RECT 32.534 7.558 32.586 7.594 ;
      RECT 32.534 8.758 32.586 8.794 ;
      RECT 32.534 9.958 32.586 9.994 ;
      RECT 32.534 11.158 32.586 11.194 ;
      RECT 32.534 12.358 32.586 12.394 ;
      RECT 32.534 13.558 32.586 13.594 ;
      RECT 32.534 14.758 32.586 14.794 ;
      RECT 32.534 15.958 32.586 15.994 ;
      RECT 32.534 17.158 32.586 17.194 ;
      RECT 32.534 18.358 32.586 18.394 ;
      RECT 32.534 19.558 32.586 19.594 ;
      RECT 32.534 20.758 32.586 20.794 ;
      RECT 32.534 21.958 32.586 21.994 ;
      RECT 32.534 23.158 32.586 23.194 ;
      RECT 32.534 24.358 32.586 24.394 ;
      RECT 32.534 25.558 32.586 25.594 ;
      RECT 32.534 26.758 32.586 26.794 ;
      RECT 32.534 27.958 32.586 27.994 ;
      RECT 32.534 29.158 32.586 29.194 ;
      RECT 32.534 30.358 32.586 30.394 ;
      RECT 32.534 31.558 32.586 31.594 ;
      RECT 32.534 33.342 32.586 33.378 ;
      RECT 32.534 33.582 32.586 33.618 ;
      RECT 32.534 37.902 32.586 37.938 ;
      RECT 32.534 38.142 32.586 38.178 ;
      RECT 32.534 40.678 32.586 40.714 ;
      RECT 32.534 41.878 32.586 41.914 ;
      RECT 32.534 43.078 32.586 43.114 ;
      RECT 32.534 44.278 32.586 44.314 ;
      RECT 32.534 45.478 32.586 45.514 ;
      RECT 32.534 46.678 32.586 46.714 ;
      RECT 32.534 47.878 32.586 47.914 ;
      RECT 32.534 49.078 32.586 49.114 ;
      RECT 32.534 50.278 32.586 50.314 ;
      RECT 32.534 51.478 32.586 51.514 ;
      RECT 32.534 52.678 32.586 52.714 ;
      RECT 32.534 53.878 32.586 53.914 ;
      RECT 32.534 55.078 32.586 55.114 ;
      RECT 32.534 56.278 32.586 56.314 ;
      RECT 32.534 57.478 32.586 57.514 ;
      RECT 32.534 58.678 32.586 58.714 ;
      RECT 32.534 59.878 32.586 59.914 ;
      RECT 32.534 61.078 32.586 61.114 ;
      RECT 32.534 62.278 32.586 62.314 ;
      RECT 32.534 63.478 32.586 63.514 ;
      RECT 32.534 64.678 32.586 64.714 ;
      RECT 32.534 65.878 32.586 65.914 ;
      RECT 32.534 67.078 32.586 67.114 ;
      RECT 32.534 68.278 32.586 68.314 ;
      RECT 32.534 69.478 32.586 69.514 ;
      RECT 32.534 70.678 32.586 70.714 ;
      RECT 32.534 71.878 32.586 71.914 ;
      RECT 32.614 0.806 32.666 0.842 ;
      RECT 32.614 2.006 32.666 2.042 ;
      RECT 32.614 3.206 32.666 3.242 ;
      RECT 32.614 4.406 32.666 4.442 ;
      RECT 32.614 5.606 32.666 5.642 ;
      RECT 32.614 6.806 32.666 6.842 ;
      RECT 32.614 8.006 32.666 8.042 ;
      RECT 32.614 9.206 32.666 9.242 ;
      RECT 32.614 10.406 32.666 10.442 ;
      RECT 32.614 11.606 32.666 11.642 ;
      RECT 32.614 12.806 32.666 12.842 ;
      RECT 32.614 14.006 32.666 14.042 ;
      RECT 32.614 15.206 32.666 15.242 ;
      RECT 32.614 16.406 32.666 16.442 ;
      RECT 32.614 17.606 32.666 17.642 ;
      RECT 32.614 18.806 32.666 18.842 ;
      RECT 32.614 20.006 32.666 20.042 ;
      RECT 32.614 21.206 32.666 21.242 ;
      RECT 32.614 22.406 32.666 22.442 ;
      RECT 32.614 23.606 32.666 23.642 ;
      RECT 32.614 24.806 32.666 24.842 ;
      RECT 32.614 26.006 32.666 26.042 ;
      RECT 32.614 27.206 32.666 27.242 ;
      RECT 32.614 28.406 32.666 28.442 ;
      RECT 32.614 29.606 32.666 29.642 ;
      RECT 32.614 30.806 32.666 30.842 ;
      RECT 32.614 32.622 32.666 32.658 ;
      RECT 32.614 32.862 32.666 32.898 ;
      RECT 32.614 38.622 32.666 38.658 ;
      RECT 32.614 38.862 32.666 38.898 ;
      RECT 32.614 39.926 32.666 39.962 ;
      RECT 32.614 41.126 32.666 41.162 ;
      RECT 32.614 42.326 32.666 42.362 ;
      RECT 32.614 43.526 32.666 43.562 ;
      RECT 32.614 44.726 32.666 44.762 ;
      RECT 32.614 45.926 32.666 45.962 ;
      RECT 32.614 47.126 32.666 47.162 ;
      RECT 32.614 48.326 32.666 48.362 ;
      RECT 32.614 49.526 32.666 49.562 ;
      RECT 32.614 50.726 32.666 50.762 ;
      RECT 32.614 51.926 32.666 51.962 ;
      RECT 32.614 53.126 32.666 53.162 ;
      RECT 32.614 54.326 32.666 54.362 ;
      RECT 32.614 55.526 32.666 55.562 ;
      RECT 32.614 56.726 32.666 56.762 ;
      RECT 32.614 57.926 32.666 57.962 ;
      RECT 32.614 59.126 32.666 59.162 ;
      RECT 32.614 60.326 32.666 60.362 ;
      RECT 32.614 61.526 32.666 61.562 ;
      RECT 32.614 62.726 32.666 62.762 ;
      RECT 32.614 63.926 32.666 63.962 ;
      RECT 32.614 65.126 32.666 65.162 ;
      RECT 32.614 66.326 32.666 66.362 ;
      RECT 32.614 67.526 32.666 67.562 ;
      RECT 32.614 68.726 32.666 68.762 ;
      RECT 32.614 69.926 32.666 69.962 ;
      RECT 32.614 71.126 32.666 71.162 ;
      RECT 32.694 1.558 32.746 1.594 ;
      RECT 32.694 2.758 32.746 2.794 ;
      RECT 32.694 3.958 32.746 3.994 ;
      RECT 32.694 5.158 32.746 5.194 ;
      RECT 32.694 6.358 32.746 6.394 ;
      RECT 32.694 7.558 32.746 7.594 ;
      RECT 32.694 8.758 32.746 8.794 ;
      RECT 32.694 9.958 32.746 9.994 ;
      RECT 32.694 11.158 32.746 11.194 ;
      RECT 32.694 12.358 32.746 12.394 ;
      RECT 32.694 13.558 32.746 13.594 ;
      RECT 32.694 14.758 32.746 14.794 ;
      RECT 32.694 15.958 32.746 15.994 ;
      RECT 32.694 17.158 32.746 17.194 ;
      RECT 32.694 18.358 32.746 18.394 ;
      RECT 32.694 19.558 32.746 19.594 ;
      RECT 32.694 20.758 32.746 20.794 ;
      RECT 32.694 21.958 32.746 21.994 ;
      RECT 32.694 23.158 32.746 23.194 ;
      RECT 32.694 24.358 32.746 24.394 ;
      RECT 32.694 25.558 32.746 25.594 ;
      RECT 32.694 26.758 32.746 26.794 ;
      RECT 32.694 27.958 32.746 27.994 ;
      RECT 32.694 29.158 32.746 29.194 ;
      RECT 32.694 30.358 32.746 30.394 ;
      RECT 32.694 31.558 32.746 31.594 ;
      RECT 32.694 33.342 32.746 33.378 ;
      RECT 32.694 33.582 32.746 33.618 ;
      RECT 32.694 37.902 32.746 37.938 ;
      RECT 32.694 38.142 32.746 38.178 ;
      RECT 32.694 40.678 32.746 40.714 ;
      RECT 32.694 41.878 32.746 41.914 ;
      RECT 32.694 43.078 32.746 43.114 ;
      RECT 32.694 44.278 32.746 44.314 ;
      RECT 32.694 45.478 32.746 45.514 ;
      RECT 32.694 46.678 32.746 46.714 ;
      RECT 32.694 47.878 32.746 47.914 ;
      RECT 32.694 49.078 32.746 49.114 ;
      RECT 32.694 50.278 32.746 50.314 ;
      RECT 32.694 51.478 32.746 51.514 ;
      RECT 32.694 52.678 32.746 52.714 ;
      RECT 32.694 53.878 32.746 53.914 ;
      RECT 32.694 55.078 32.746 55.114 ;
      RECT 32.694 56.278 32.746 56.314 ;
      RECT 32.694 57.478 32.746 57.514 ;
      RECT 32.694 58.678 32.746 58.714 ;
      RECT 32.694 59.878 32.746 59.914 ;
      RECT 32.694 61.078 32.746 61.114 ;
      RECT 32.694 62.278 32.746 62.314 ;
      RECT 32.694 63.478 32.746 63.514 ;
      RECT 32.694 64.678 32.746 64.714 ;
      RECT 32.694 65.878 32.746 65.914 ;
      RECT 32.694 67.078 32.746 67.114 ;
      RECT 32.694 68.278 32.746 68.314 ;
      RECT 32.694 69.478 32.746 69.514 ;
      RECT 32.694 70.678 32.746 70.714 ;
      RECT 32.694 71.878 32.746 71.914 ;
      RECT 32.774 0.281 32.826 0.317 ;
      RECT 32.774 72.403 32.826 72.439 ;
      RECT 32.854 0.806 32.906 0.842 ;
      RECT 32.854 2.006 32.906 2.042 ;
      RECT 32.854 3.206 32.906 3.242 ;
      RECT 32.854 4.406 32.906 4.442 ;
      RECT 32.854 5.606 32.906 5.642 ;
      RECT 32.854 6.806 32.906 6.842 ;
      RECT 32.854 8.006 32.906 8.042 ;
      RECT 32.854 9.206 32.906 9.242 ;
      RECT 32.854 10.406 32.906 10.442 ;
      RECT 32.854 11.606 32.906 11.642 ;
      RECT 32.854 12.806 32.906 12.842 ;
      RECT 32.854 14.006 32.906 14.042 ;
      RECT 32.854 15.206 32.906 15.242 ;
      RECT 32.854 16.406 32.906 16.442 ;
      RECT 32.854 17.606 32.906 17.642 ;
      RECT 32.854 18.806 32.906 18.842 ;
      RECT 32.854 20.006 32.906 20.042 ;
      RECT 32.854 21.206 32.906 21.242 ;
      RECT 32.854 22.406 32.906 22.442 ;
      RECT 32.854 23.606 32.906 23.642 ;
      RECT 32.854 24.806 32.906 24.842 ;
      RECT 32.854 26.006 32.906 26.042 ;
      RECT 32.854 27.206 32.906 27.242 ;
      RECT 32.854 28.406 32.906 28.442 ;
      RECT 32.854 29.606 32.906 29.642 ;
      RECT 32.854 30.806 32.906 30.842 ;
      RECT 32.854 32.622 32.906 32.658 ;
      RECT 32.854 32.862 32.906 32.898 ;
      RECT 32.854 34.302 32.906 34.338 ;
      RECT 32.854 34.782 32.906 34.818 ;
      RECT 32.854 36.702 32.906 36.738 ;
      RECT 32.854 37.182 32.906 37.218 ;
      RECT 32.854 38.622 32.906 38.658 ;
      RECT 32.854 38.862 32.906 38.898 ;
      RECT 32.854 39.926 32.906 39.962 ;
      RECT 32.854 41.126 32.906 41.162 ;
      RECT 32.854 42.326 32.906 42.362 ;
      RECT 32.854 43.526 32.906 43.562 ;
      RECT 32.854 44.726 32.906 44.762 ;
      RECT 32.854 45.926 32.906 45.962 ;
      RECT 32.854 47.126 32.906 47.162 ;
      RECT 32.854 48.326 32.906 48.362 ;
      RECT 32.854 49.526 32.906 49.562 ;
      RECT 32.854 50.726 32.906 50.762 ;
      RECT 32.854 51.926 32.906 51.962 ;
      RECT 32.854 53.126 32.906 53.162 ;
      RECT 32.854 54.326 32.906 54.362 ;
      RECT 32.854 55.526 32.906 55.562 ;
      RECT 32.854 56.726 32.906 56.762 ;
      RECT 32.854 57.926 32.906 57.962 ;
      RECT 32.854 59.126 32.906 59.162 ;
      RECT 32.854 60.326 32.906 60.362 ;
      RECT 32.854 61.526 32.906 61.562 ;
      RECT 32.854 62.726 32.906 62.762 ;
      RECT 32.854 63.926 32.906 63.962 ;
      RECT 32.854 65.126 32.906 65.162 ;
      RECT 32.854 66.326 32.906 66.362 ;
      RECT 32.854 67.526 32.906 67.562 ;
      RECT 32.854 68.726 32.906 68.762 ;
      RECT 32.854 69.926 32.906 69.962 ;
      RECT 32.854 71.126 32.906 71.162 ;
      RECT 32.934 1.558 32.986 1.594 ;
      RECT 32.934 2.758 32.986 2.794 ;
      RECT 32.934 3.958 32.986 3.994 ;
      RECT 32.934 5.158 32.986 5.194 ;
      RECT 32.934 6.358 32.986 6.394 ;
      RECT 32.934 7.558 32.986 7.594 ;
      RECT 32.934 8.758 32.986 8.794 ;
      RECT 32.934 9.958 32.986 9.994 ;
      RECT 32.934 11.158 32.986 11.194 ;
      RECT 32.934 12.358 32.986 12.394 ;
      RECT 32.934 13.558 32.986 13.594 ;
      RECT 32.934 14.758 32.986 14.794 ;
      RECT 32.934 15.958 32.986 15.994 ;
      RECT 32.934 17.158 32.986 17.194 ;
      RECT 32.934 18.358 32.986 18.394 ;
      RECT 32.934 19.558 32.986 19.594 ;
      RECT 32.934 20.758 32.986 20.794 ;
      RECT 32.934 21.958 32.986 21.994 ;
      RECT 32.934 23.158 32.986 23.194 ;
      RECT 32.934 24.358 32.986 24.394 ;
      RECT 32.934 25.558 32.986 25.594 ;
      RECT 32.934 26.758 32.986 26.794 ;
      RECT 32.934 27.958 32.986 27.994 ;
      RECT 32.934 29.158 32.986 29.194 ;
      RECT 32.934 30.358 32.986 30.394 ;
      RECT 32.934 31.558 32.986 31.594 ;
      RECT 32.934 33.342 32.986 33.378 ;
      RECT 32.934 33.582 32.986 33.618 ;
      RECT 32.934 37.902 32.986 37.938 ;
      RECT 32.934 38.142 32.986 38.178 ;
      RECT 32.934 40.678 32.986 40.714 ;
      RECT 32.934 41.878 32.986 41.914 ;
      RECT 32.934 43.078 32.986 43.114 ;
      RECT 32.934 44.278 32.986 44.314 ;
      RECT 32.934 45.478 32.986 45.514 ;
      RECT 32.934 46.678 32.986 46.714 ;
      RECT 32.934 47.878 32.986 47.914 ;
      RECT 32.934 49.078 32.986 49.114 ;
      RECT 32.934 50.278 32.986 50.314 ;
      RECT 32.934 51.478 32.986 51.514 ;
      RECT 32.934 52.678 32.986 52.714 ;
      RECT 32.934 53.878 32.986 53.914 ;
      RECT 32.934 55.078 32.986 55.114 ;
      RECT 32.934 56.278 32.986 56.314 ;
      RECT 32.934 57.478 32.986 57.514 ;
      RECT 32.934 58.678 32.986 58.714 ;
      RECT 32.934 59.878 32.986 59.914 ;
      RECT 32.934 61.078 32.986 61.114 ;
      RECT 32.934 62.278 32.986 62.314 ;
      RECT 32.934 63.478 32.986 63.514 ;
      RECT 32.934 64.678 32.986 64.714 ;
      RECT 32.934 65.878 32.986 65.914 ;
      RECT 32.934 67.078 32.986 67.114 ;
      RECT 32.934 68.278 32.986 68.314 ;
      RECT 32.934 69.478 32.986 69.514 ;
      RECT 32.934 70.678 32.986 70.714 ;
      RECT 32.934 71.878 32.986 71.914 ;
      RECT 33.014 0.806 33.066 0.842 ;
      RECT 33.014 2.006 33.066 2.042 ;
      RECT 33.014 3.206 33.066 3.242 ;
      RECT 33.014 4.406 33.066 4.442 ;
      RECT 33.014 5.606 33.066 5.642 ;
      RECT 33.014 6.806 33.066 6.842 ;
      RECT 33.014 8.006 33.066 8.042 ;
      RECT 33.014 9.206 33.066 9.242 ;
      RECT 33.014 10.406 33.066 10.442 ;
      RECT 33.014 11.606 33.066 11.642 ;
      RECT 33.014 12.806 33.066 12.842 ;
      RECT 33.014 14.006 33.066 14.042 ;
      RECT 33.014 15.206 33.066 15.242 ;
      RECT 33.014 16.406 33.066 16.442 ;
      RECT 33.014 17.606 33.066 17.642 ;
      RECT 33.014 18.806 33.066 18.842 ;
      RECT 33.014 20.006 33.066 20.042 ;
      RECT 33.014 21.206 33.066 21.242 ;
      RECT 33.014 22.406 33.066 22.442 ;
      RECT 33.014 23.606 33.066 23.642 ;
      RECT 33.014 24.806 33.066 24.842 ;
      RECT 33.014 26.006 33.066 26.042 ;
      RECT 33.014 27.206 33.066 27.242 ;
      RECT 33.014 28.406 33.066 28.442 ;
      RECT 33.014 29.606 33.066 29.642 ;
      RECT 33.014 30.806 33.066 30.842 ;
      RECT 33.014 32.622 33.066 32.658 ;
      RECT 33.014 32.862 33.066 32.898 ;
      RECT 33.014 38.622 33.066 38.658 ;
      RECT 33.014 38.862 33.066 38.898 ;
      RECT 33.014 39.926 33.066 39.962 ;
      RECT 33.014 41.126 33.066 41.162 ;
      RECT 33.014 42.326 33.066 42.362 ;
      RECT 33.014 43.526 33.066 43.562 ;
      RECT 33.014 44.726 33.066 44.762 ;
      RECT 33.014 45.926 33.066 45.962 ;
      RECT 33.014 47.126 33.066 47.162 ;
      RECT 33.014 48.326 33.066 48.362 ;
      RECT 33.014 49.526 33.066 49.562 ;
      RECT 33.014 50.726 33.066 50.762 ;
      RECT 33.014 51.926 33.066 51.962 ;
      RECT 33.014 53.126 33.066 53.162 ;
      RECT 33.014 54.326 33.066 54.362 ;
      RECT 33.014 55.526 33.066 55.562 ;
      RECT 33.014 56.726 33.066 56.762 ;
      RECT 33.014 57.926 33.066 57.962 ;
      RECT 33.014 59.126 33.066 59.162 ;
      RECT 33.014 60.326 33.066 60.362 ;
      RECT 33.014 61.526 33.066 61.562 ;
      RECT 33.014 62.726 33.066 62.762 ;
      RECT 33.014 63.926 33.066 63.962 ;
      RECT 33.014 65.126 33.066 65.162 ;
      RECT 33.014 66.326 33.066 66.362 ;
      RECT 33.014 67.526 33.066 67.562 ;
      RECT 33.014 68.726 33.066 68.762 ;
      RECT 33.014 69.926 33.066 69.962 ;
      RECT 33.014 71.126 33.066 71.162 ;
      RECT 33.094 1.558 33.146 1.594 ;
      RECT 33.094 2.758 33.146 2.794 ;
      RECT 33.094 3.958 33.146 3.994 ;
      RECT 33.094 5.158 33.146 5.194 ;
      RECT 33.094 6.358 33.146 6.394 ;
      RECT 33.094 7.558 33.146 7.594 ;
      RECT 33.094 8.758 33.146 8.794 ;
      RECT 33.094 9.958 33.146 9.994 ;
      RECT 33.094 11.158 33.146 11.194 ;
      RECT 33.094 12.358 33.146 12.394 ;
      RECT 33.094 13.558 33.146 13.594 ;
      RECT 33.094 14.758 33.146 14.794 ;
      RECT 33.094 15.958 33.146 15.994 ;
      RECT 33.094 17.158 33.146 17.194 ;
      RECT 33.094 18.358 33.146 18.394 ;
      RECT 33.094 19.558 33.146 19.594 ;
      RECT 33.094 20.758 33.146 20.794 ;
      RECT 33.094 21.958 33.146 21.994 ;
      RECT 33.094 23.158 33.146 23.194 ;
      RECT 33.094 24.358 33.146 24.394 ;
      RECT 33.094 25.558 33.146 25.594 ;
      RECT 33.094 26.758 33.146 26.794 ;
      RECT 33.094 27.958 33.146 27.994 ;
      RECT 33.094 29.158 33.146 29.194 ;
      RECT 33.094 30.358 33.146 30.394 ;
      RECT 33.094 31.558 33.146 31.594 ;
      RECT 33.094 33.342 33.146 33.378 ;
      RECT 33.094 33.582 33.146 33.618 ;
      RECT 33.094 37.902 33.146 37.938 ;
      RECT 33.094 38.142 33.146 38.178 ;
      RECT 33.094 40.678 33.146 40.714 ;
      RECT 33.094 41.878 33.146 41.914 ;
      RECT 33.094 43.078 33.146 43.114 ;
      RECT 33.094 44.278 33.146 44.314 ;
      RECT 33.094 45.478 33.146 45.514 ;
      RECT 33.094 46.678 33.146 46.714 ;
      RECT 33.094 47.878 33.146 47.914 ;
      RECT 33.094 49.078 33.146 49.114 ;
      RECT 33.094 50.278 33.146 50.314 ;
      RECT 33.094 51.478 33.146 51.514 ;
      RECT 33.094 52.678 33.146 52.714 ;
      RECT 33.094 53.878 33.146 53.914 ;
      RECT 33.094 55.078 33.146 55.114 ;
      RECT 33.094 56.278 33.146 56.314 ;
      RECT 33.094 57.478 33.146 57.514 ;
      RECT 33.094 58.678 33.146 58.714 ;
      RECT 33.094 59.878 33.146 59.914 ;
      RECT 33.094 61.078 33.146 61.114 ;
      RECT 33.094 62.278 33.146 62.314 ;
      RECT 33.094 63.478 33.146 63.514 ;
      RECT 33.094 64.678 33.146 64.714 ;
      RECT 33.094 65.878 33.146 65.914 ;
      RECT 33.094 67.078 33.146 67.114 ;
      RECT 33.094 68.278 33.146 68.314 ;
      RECT 33.094 69.478 33.146 69.514 ;
      RECT 33.094 70.678 33.146 70.714 ;
      RECT 33.094 71.878 33.146 71.914 ;
      RECT 33.174 0.281 33.226 0.317 ;
      RECT 33.174 72.403 33.226 72.439 ;
      RECT 33.254 0.806 33.306 0.842 ;
      RECT 33.254 2.006 33.306 2.042 ;
      RECT 33.254 3.206 33.306 3.242 ;
      RECT 33.254 4.406 33.306 4.442 ;
      RECT 33.254 5.606 33.306 5.642 ;
      RECT 33.254 6.806 33.306 6.842 ;
      RECT 33.254 8.006 33.306 8.042 ;
      RECT 33.254 9.206 33.306 9.242 ;
      RECT 33.254 10.406 33.306 10.442 ;
      RECT 33.254 11.606 33.306 11.642 ;
      RECT 33.254 12.806 33.306 12.842 ;
      RECT 33.254 14.006 33.306 14.042 ;
      RECT 33.254 15.206 33.306 15.242 ;
      RECT 33.254 16.406 33.306 16.442 ;
      RECT 33.254 17.606 33.306 17.642 ;
      RECT 33.254 18.806 33.306 18.842 ;
      RECT 33.254 20.006 33.306 20.042 ;
      RECT 33.254 21.206 33.306 21.242 ;
      RECT 33.254 22.406 33.306 22.442 ;
      RECT 33.254 23.606 33.306 23.642 ;
      RECT 33.254 24.806 33.306 24.842 ;
      RECT 33.254 26.006 33.306 26.042 ;
      RECT 33.254 27.206 33.306 27.242 ;
      RECT 33.254 28.406 33.306 28.442 ;
      RECT 33.254 29.606 33.306 29.642 ;
      RECT 33.254 30.806 33.306 30.842 ;
      RECT 33.254 32.622 33.306 32.658 ;
      RECT 33.254 32.862 33.306 32.898 ;
      RECT 33.254 38.622 33.306 38.658 ;
      RECT 33.254 38.862 33.306 38.898 ;
      RECT 33.254 39.926 33.306 39.962 ;
      RECT 33.254 41.126 33.306 41.162 ;
      RECT 33.254 42.326 33.306 42.362 ;
      RECT 33.254 43.526 33.306 43.562 ;
      RECT 33.254 44.726 33.306 44.762 ;
      RECT 33.254 45.926 33.306 45.962 ;
      RECT 33.254 47.126 33.306 47.162 ;
      RECT 33.254 48.326 33.306 48.362 ;
      RECT 33.254 49.526 33.306 49.562 ;
      RECT 33.254 50.726 33.306 50.762 ;
      RECT 33.254 51.926 33.306 51.962 ;
      RECT 33.254 53.126 33.306 53.162 ;
      RECT 33.254 54.326 33.306 54.362 ;
      RECT 33.254 55.526 33.306 55.562 ;
      RECT 33.254 56.726 33.306 56.762 ;
      RECT 33.254 57.926 33.306 57.962 ;
      RECT 33.254 59.126 33.306 59.162 ;
      RECT 33.254 60.326 33.306 60.362 ;
      RECT 33.254 61.526 33.306 61.562 ;
      RECT 33.254 62.726 33.306 62.762 ;
      RECT 33.254 63.926 33.306 63.962 ;
      RECT 33.254 65.126 33.306 65.162 ;
      RECT 33.254 66.326 33.306 66.362 ;
      RECT 33.254 67.526 33.306 67.562 ;
      RECT 33.254 68.726 33.306 68.762 ;
      RECT 33.254 69.926 33.306 69.962 ;
      RECT 33.254 71.126 33.306 71.162 ;
      RECT 33.334 1.558 33.386 1.594 ;
      RECT 33.334 2.758 33.386 2.794 ;
      RECT 33.334 3.958 33.386 3.994 ;
      RECT 33.334 5.158 33.386 5.194 ;
      RECT 33.334 6.358 33.386 6.394 ;
      RECT 33.334 7.558 33.386 7.594 ;
      RECT 33.334 8.758 33.386 8.794 ;
      RECT 33.334 9.958 33.386 9.994 ;
      RECT 33.334 11.158 33.386 11.194 ;
      RECT 33.334 12.358 33.386 12.394 ;
      RECT 33.334 13.558 33.386 13.594 ;
      RECT 33.334 14.758 33.386 14.794 ;
      RECT 33.334 15.958 33.386 15.994 ;
      RECT 33.334 17.158 33.386 17.194 ;
      RECT 33.334 18.358 33.386 18.394 ;
      RECT 33.334 19.558 33.386 19.594 ;
      RECT 33.334 20.758 33.386 20.794 ;
      RECT 33.334 21.958 33.386 21.994 ;
      RECT 33.334 23.158 33.386 23.194 ;
      RECT 33.334 24.358 33.386 24.394 ;
      RECT 33.334 25.558 33.386 25.594 ;
      RECT 33.334 26.758 33.386 26.794 ;
      RECT 33.334 27.958 33.386 27.994 ;
      RECT 33.334 29.158 33.386 29.194 ;
      RECT 33.334 30.358 33.386 30.394 ;
      RECT 33.334 31.558 33.386 31.594 ;
      RECT 33.334 33.342 33.386 33.378 ;
      RECT 33.334 33.582 33.386 33.618 ;
      RECT 33.334 37.902 33.386 37.938 ;
      RECT 33.334 38.142 33.386 38.178 ;
      RECT 33.334 40.678 33.386 40.714 ;
      RECT 33.334 41.878 33.386 41.914 ;
      RECT 33.334 43.078 33.386 43.114 ;
      RECT 33.334 44.278 33.386 44.314 ;
      RECT 33.334 45.478 33.386 45.514 ;
      RECT 33.334 46.678 33.386 46.714 ;
      RECT 33.334 47.878 33.386 47.914 ;
      RECT 33.334 49.078 33.386 49.114 ;
      RECT 33.334 50.278 33.386 50.314 ;
      RECT 33.334 51.478 33.386 51.514 ;
      RECT 33.334 52.678 33.386 52.714 ;
      RECT 33.334 53.878 33.386 53.914 ;
      RECT 33.334 55.078 33.386 55.114 ;
      RECT 33.334 56.278 33.386 56.314 ;
      RECT 33.334 57.478 33.386 57.514 ;
      RECT 33.334 58.678 33.386 58.714 ;
      RECT 33.334 59.878 33.386 59.914 ;
      RECT 33.334 61.078 33.386 61.114 ;
      RECT 33.334 62.278 33.386 62.314 ;
      RECT 33.334 63.478 33.386 63.514 ;
      RECT 33.334 64.678 33.386 64.714 ;
      RECT 33.334 65.878 33.386 65.914 ;
      RECT 33.334 67.078 33.386 67.114 ;
      RECT 33.334 68.278 33.386 68.314 ;
      RECT 33.334 69.478 33.386 69.514 ;
      RECT 33.334 70.678 33.386 70.714 ;
      RECT 33.334 71.878 33.386 71.914 ;
      RECT 33.414 0.806 33.466 0.842 ;
      RECT 33.414 2.006 33.466 2.042 ;
      RECT 33.414 3.206 33.466 3.242 ;
      RECT 33.414 4.406 33.466 4.442 ;
      RECT 33.414 5.606 33.466 5.642 ;
      RECT 33.414 6.806 33.466 6.842 ;
      RECT 33.414 8.006 33.466 8.042 ;
      RECT 33.414 9.206 33.466 9.242 ;
      RECT 33.414 10.406 33.466 10.442 ;
      RECT 33.414 11.606 33.466 11.642 ;
      RECT 33.414 12.806 33.466 12.842 ;
      RECT 33.414 14.006 33.466 14.042 ;
      RECT 33.414 15.206 33.466 15.242 ;
      RECT 33.414 16.406 33.466 16.442 ;
      RECT 33.414 17.606 33.466 17.642 ;
      RECT 33.414 18.806 33.466 18.842 ;
      RECT 33.414 20.006 33.466 20.042 ;
      RECT 33.414 21.206 33.466 21.242 ;
      RECT 33.414 22.406 33.466 22.442 ;
      RECT 33.414 23.606 33.466 23.642 ;
      RECT 33.414 24.806 33.466 24.842 ;
      RECT 33.414 26.006 33.466 26.042 ;
      RECT 33.414 27.206 33.466 27.242 ;
      RECT 33.414 28.406 33.466 28.442 ;
      RECT 33.414 29.606 33.466 29.642 ;
      RECT 33.414 30.806 33.466 30.842 ;
      RECT 33.414 32.622 33.466 32.658 ;
      RECT 33.414 32.862 33.466 32.898 ;
      RECT 33.414 38.622 33.466 38.658 ;
      RECT 33.414 38.862 33.466 38.898 ;
      RECT 33.414 39.926 33.466 39.962 ;
      RECT 33.414 41.126 33.466 41.162 ;
      RECT 33.414 42.326 33.466 42.362 ;
      RECT 33.414 43.526 33.466 43.562 ;
      RECT 33.414 44.726 33.466 44.762 ;
      RECT 33.414 45.926 33.466 45.962 ;
      RECT 33.414 47.126 33.466 47.162 ;
      RECT 33.414 48.326 33.466 48.362 ;
      RECT 33.414 49.526 33.466 49.562 ;
      RECT 33.414 50.726 33.466 50.762 ;
      RECT 33.414 51.926 33.466 51.962 ;
      RECT 33.414 53.126 33.466 53.162 ;
      RECT 33.414 54.326 33.466 54.362 ;
      RECT 33.414 55.526 33.466 55.562 ;
      RECT 33.414 56.726 33.466 56.762 ;
      RECT 33.414 57.926 33.466 57.962 ;
      RECT 33.414 59.126 33.466 59.162 ;
      RECT 33.414 60.326 33.466 60.362 ;
      RECT 33.414 61.526 33.466 61.562 ;
      RECT 33.414 62.726 33.466 62.762 ;
      RECT 33.414 63.926 33.466 63.962 ;
      RECT 33.414 65.126 33.466 65.162 ;
      RECT 33.414 66.326 33.466 66.362 ;
      RECT 33.414 67.526 33.466 67.562 ;
      RECT 33.414 68.726 33.466 68.762 ;
      RECT 33.414 69.926 33.466 69.962 ;
      RECT 33.414 71.126 33.466 71.162 ;
      RECT 33.494 1.558 33.546 1.594 ;
      RECT 33.494 2.758 33.546 2.794 ;
      RECT 33.494 3.958 33.546 3.994 ;
      RECT 33.494 5.158 33.546 5.194 ;
      RECT 33.494 6.358 33.546 6.394 ;
      RECT 33.494 7.558 33.546 7.594 ;
      RECT 33.494 8.758 33.546 8.794 ;
      RECT 33.494 9.958 33.546 9.994 ;
      RECT 33.494 11.158 33.546 11.194 ;
      RECT 33.494 12.358 33.546 12.394 ;
      RECT 33.494 13.558 33.546 13.594 ;
      RECT 33.494 14.758 33.546 14.794 ;
      RECT 33.494 15.958 33.546 15.994 ;
      RECT 33.494 17.158 33.546 17.194 ;
      RECT 33.494 18.358 33.546 18.394 ;
      RECT 33.494 19.558 33.546 19.594 ;
      RECT 33.494 20.758 33.546 20.794 ;
      RECT 33.494 21.958 33.546 21.994 ;
      RECT 33.494 23.158 33.546 23.194 ;
      RECT 33.494 24.358 33.546 24.394 ;
      RECT 33.494 25.558 33.546 25.594 ;
      RECT 33.494 26.758 33.546 26.794 ;
      RECT 33.494 27.958 33.546 27.994 ;
      RECT 33.494 29.158 33.546 29.194 ;
      RECT 33.494 30.358 33.546 30.394 ;
      RECT 33.494 31.558 33.546 31.594 ;
      RECT 33.494 33.342 33.546 33.378 ;
      RECT 33.494 33.582 33.546 33.618 ;
      RECT 33.494 37.902 33.546 37.938 ;
      RECT 33.494 38.142 33.546 38.178 ;
      RECT 33.494 40.678 33.546 40.714 ;
      RECT 33.494 41.878 33.546 41.914 ;
      RECT 33.494 43.078 33.546 43.114 ;
      RECT 33.494 44.278 33.546 44.314 ;
      RECT 33.494 45.478 33.546 45.514 ;
      RECT 33.494 46.678 33.546 46.714 ;
      RECT 33.494 47.878 33.546 47.914 ;
      RECT 33.494 49.078 33.546 49.114 ;
      RECT 33.494 50.278 33.546 50.314 ;
      RECT 33.494 51.478 33.546 51.514 ;
      RECT 33.494 52.678 33.546 52.714 ;
      RECT 33.494 53.878 33.546 53.914 ;
      RECT 33.494 55.078 33.546 55.114 ;
      RECT 33.494 56.278 33.546 56.314 ;
      RECT 33.494 57.478 33.546 57.514 ;
      RECT 33.494 58.678 33.546 58.714 ;
      RECT 33.494 59.878 33.546 59.914 ;
      RECT 33.494 61.078 33.546 61.114 ;
      RECT 33.494 62.278 33.546 62.314 ;
      RECT 33.494 63.478 33.546 63.514 ;
      RECT 33.494 64.678 33.546 64.714 ;
      RECT 33.494 65.878 33.546 65.914 ;
      RECT 33.494 67.078 33.546 67.114 ;
      RECT 33.494 68.278 33.546 68.314 ;
      RECT 33.494 69.478 33.546 69.514 ;
      RECT 33.494 70.678 33.546 70.714 ;
      RECT 33.494 71.878 33.546 71.914 ;
      RECT 33.574 0.281 33.626 0.317 ;
      RECT 33.574 72.403 33.626 72.439 ;
      RECT 33.654 0.806 33.706 0.842 ;
      RECT 33.654 2.006 33.706 2.042 ;
      RECT 33.654 3.206 33.706 3.242 ;
      RECT 33.654 4.406 33.706 4.442 ;
      RECT 33.654 5.606 33.706 5.642 ;
      RECT 33.654 6.806 33.706 6.842 ;
      RECT 33.654 8.006 33.706 8.042 ;
      RECT 33.654 9.206 33.706 9.242 ;
      RECT 33.654 10.406 33.706 10.442 ;
      RECT 33.654 11.606 33.706 11.642 ;
      RECT 33.654 12.806 33.706 12.842 ;
      RECT 33.654 14.006 33.706 14.042 ;
      RECT 33.654 15.206 33.706 15.242 ;
      RECT 33.654 16.406 33.706 16.442 ;
      RECT 33.654 17.606 33.706 17.642 ;
      RECT 33.654 18.806 33.706 18.842 ;
      RECT 33.654 20.006 33.706 20.042 ;
      RECT 33.654 21.206 33.706 21.242 ;
      RECT 33.654 22.406 33.706 22.442 ;
      RECT 33.654 23.606 33.706 23.642 ;
      RECT 33.654 24.806 33.706 24.842 ;
      RECT 33.654 26.006 33.706 26.042 ;
      RECT 33.654 27.206 33.706 27.242 ;
      RECT 33.654 28.406 33.706 28.442 ;
      RECT 33.654 29.606 33.706 29.642 ;
      RECT 33.654 30.806 33.706 30.842 ;
      RECT 33.654 32.622 33.706 32.658 ;
      RECT 33.654 32.862 33.706 32.898 ;
      RECT 33.654 34.302 33.706 34.338 ;
      RECT 33.654 34.782 33.706 34.818 ;
      RECT 33.654 36.702 33.706 36.738 ;
      RECT 33.654 37.182 33.706 37.218 ;
      RECT 33.654 38.622 33.706 38.658 ;
      RECT 33.654 38.862 33.706 38.898 ;
      RECT 33.654 39.926 33.706 39.962 ;
      RECT 33.654 41.126 33.706 41.162 ;
      RECT 33.654 42.326 33.706 42.362 ;
      RECT 33.654 43.526 33.706 43.562 ;
      RECT 33.654 44.726 33.706 44.762 ;
      RECT 33.654 45.926 33.706 45.962 ;
      RECT 33.654 47.126 33.706 47.162 ;
      RECT 33.654 48.326 33.706 48.362 ;
      RECT 33.654 49.526 33.706 49.562 ;
      RECT 33.654 50.726 33.706 50.762 ;
      RECT 33.654 51.926 33.706 51.962 ;
      RECT 33.654 53.126 33.706 53.162 ;
      RECT 33.654 54.326 33.706 54.362 ;
      RECT 33.654 55.526 33.706 55.562 ;
      RECT 33.654 56.726 33.706 56.762 ;
      RECT 33.654 57.926 33.706 57.962 ;
      RECT 33.654 59.126 33.706 59.162 ;
      RECT 33.654 60.326 33.706 60.362 ;
      RECT 33.654 61.526 33.706 61.562 ;
      RECT 33.654 62.726 33.706 62.762 ;
      RECT 33.654 63.926 33.706 63.962 ;
      RECT 33.654 65.126 33.706 65.162 ;
      RECT 33.654 66.326 33.706 66.362 ;
      RECT 33.654 67.526 33.706 67.562 ;
      RECT 33.654 68.726 33.706 68.762 ;
      RECT 33.654 69.926 33.706 69.962 ;
      RECT 33.654 71.126 33.706 71.162 ;
      RECT 33.734 1.558 33.786 1.594 ;
      RECT 33.734 2.758 33.786 2.794 ;
      RECT 33.734 3.958 33.786 3.994 ;
      RECT 33.734 5.158 33.786 5.194 ;
      RECT 33.734 6.358 33.786 6.394 ;
      RECT 33.734 7.558 33.786 7.594 ;
      RECT 33.734 8.758 33.786 8.794 ;
      RECT 33.734 9.958 33.786 9.994 ;
      RECT 33.734 11.158 33.786 11.194 ;
      RECT 33.734 12.358 33.786 12.394 ;
      RECT 33.734 13.558 33.786 13.594 ;
      RECT 33.734 14.758 33.786 14.794 ;
      RECT 33.734 15.958 33.786 15.994 ;
      RECT 33.734 17.158 33.786 17.194 ;
      RECT 33.734 18.358 33.786 18.394 ;
      RECT 33.734 19.558 33.786 19.594 ;
      RECT 33.734 20.758 33.786 20.794 ;
      RECT 33.734 21.958 33.786 21.994 ;
      RECT 33.734 23.158 33.786 23.194 ;
      RECT 33.734 24.358 33.786 24.394 ;
      RECT 33.734 25.558 33.786 25.594 ;
      RECT 33.734 26.758 33.786 26.794 ;
      RECT 33.734 27.958 33.786 27.994 ;
      RECT 33.734 29.158 33.786 29.194 ;
      RECT 33.734 30.358 33.786 30.394 ;
      RECT 33.734 31.558 33.786 31.594 ;
      RECT 33.734 33.342 33.786 33.378 ;
      RECT 33.734 33.582 33.786 33.618 ;
      RECT 33.734 37.902 33.786 37.938 ;
      RECT 33.734 38.142 33.786 38.178 ;
      RECT 33.734 40.678 33.786 40.714 ;
      RECT 33.734 41.878 33.786 41.914 ;
      RECT 33.734 43.078 33.786 43.114 ;
      RECT 33.734 44.278 33.786 44.314 ;
      RECT 33.734 45.478 33.786 45.514 ;
      RECT 33.734 46.678 33.786 46.714 ;
      RECT 33.734 47.878 33.786 47.914 ;
      RECT 33.734 49.078 33.786 49.114 ;
      RECT 33.734 50.278 33.786 50.314 ;
      RECT 33.734 51.478 33.786 51.514 ;
      RECT 33.734 52.678 33.786 52.714 ;
      RECT 33.734 53.878 33.786 53.914 ;
      RECT 33.734 55.078 33.786 55.114 ;
      RECT 33.734 56.278 33.786 56.314 ;
      RECT 33.734 57.478 33.786 57.514 ;
      RECT 33.734 58.678 33.786 58.714 ;
      RECT 33.734 59.878 33.786 59.914 ;
      RECT 33.734 61.078 33.786 61.114 ;
      RECT 33.734 62.278 33.786 62.314 ;
      RECT 33.734 63.478 33.786 63.514 ;
      RECT 33.734 64.678 33.786 64.714 ;
      RECT 33.734 65.878 33.786 65.914 ;
      RECT 33.734 67.078 33.786 67.114 ;
      RECT 33.734 68.278 33.786 68.314 ;
      RECT 33.734 69.478 33.786 69.514 ;
      RECT 33.734 70.678 33.786 70.714 ;
      RECT 33.734 71.878 33.786 71.914 ;
      RECT 33.814 0.806 33.866 0.842 ;
      RECT 33.814 2.006 33.866 2.042 ;
      RECT 33.814 3.206 33.866 3.242 ;
      RECT 33.814 4.406 33.866 4.442 ;
      RECT 33.814 5.606 33.866 5.642 ;
      RECT 33.814 6.806 33.866 6.842 ;
      RECT 33.814 8.006 33.866 8.042 ;
      RECT 33.814 9.206 33.866 9.242 ;
      RECT 33.814 10.406 33.866 10.442 ;
      RECT 33.814 11.606 33.866 11.642 ;
      RECT 33.814 12.806 33.866 12.842 ;
      RECT 33.814 14.006 33.866 14.042 ;
      RECT 33.814 15.206 33.866 15.242 ;
      RECT 33.814 16.406 33.866 16.442 ;
      RECT 33.814 17.606 33.866 17.642 ;
      RECT 33.814 18.806 33.866 18.842 ;
      RECT 33.814 20.006 33.866 20.042 ;
      RECT 33.814 21.206 33.866 21.242 ;
      RECT 33.814 22.406 33.866 22.442 ;
      RECT 33.814 23.606 33.866 23.642 ;
      RECT 33.814 24.806 33.866 24.842 ;
      RECT 33.814 26.006 33.866 26.042 ;
      RECT 33.814 27.206 33.866 27.242 ;
      RECT 33.814 28.406 33.866 28.442 ;
      RECT 33.814 29.606 33.866 29.642 ;
      RECT 33.814 30.806 33.866 30.842 ;
      RECT 33.814 32.622 33.866 32.658 ;
      RECT 33.814 32.862 33.866 32.898 ;
      RECT 33.814 38.622 33.866 38.658 ;
      RECT 33.814 38.862 33.866 38.898 ;
      RECT 33.814 39.926 33.866 39.962 ;
      RECT 33.814 41.126 33.866 41.162 ;
      RECT 33.814 42.326 33.866 42.362 ;
      RECT 33.814 43.526 33.866 43.562 ;
      RECT 33.814 44.726 33.866 44.762 ;
      RECT 33.814 45.926 33.866 45.962 ;
      RECT 33.814 47.126 33.866 47.162 ;
      RECT 33.814 48.326 33.866 48.362 ;
      RECT 33.814 49.526 33.866 49.562 ;
      RECT 33.814 50.726 33.866 50.762 ;
      RECT 33.814 51.926 33.866 51.962 ;
      RECT 33.814 53.126 33.866 53.162 ;
      RECT 33.814 54.326 33.866 54.362 ;
      RECT 33.814 55.526 33.866 55.562 ;
      RECT 33.814 56.726 33.866 56.762 ;
      RECT 33.814 57.926 33.866 57.962 ;
      RECT 33.814 59.126 33.866 59.162 ;
      RECT 33.814 60.326 33.866 60.362 ;
      RECT 33.814 61.526 33.866 61.562 ;
      RECT 33.814 62.726 33.866 62.762 ;
      RECT 33.814 63.926 33.866 63.962 ;
      RECT 33.814 65.126 33.866 65.162 ;
      RECT 33.814 66.326 33.866 66.362 ;
      RECT 33.814 67.526 33.866 67.562 ;
      RECT 33.814 68.726 33.866 68.762 ;
      RECT 33.814 69.926 33.866 69.962 ;
      RECT 33.814 71.126 33.866 71.162 ;
      RECT 33.894 1.558 33.946 1.594 ;
      RECT 33.894 2.758 33.946 2.794 ;
      RECT 33.894 3.958 33.946 3.994 ;
      RECT 33.894 5.158 33.946 5.194 ;
      RECT 33.894 6.358 33.946 6.394 ;
      RECT 33.894 7.558 33.946 7.594 ;
      RECT 33.894 8.758 33.946 8.794 ;
      RECT 33.894 9.958 33.946 9.994 ;
      RECT 33.894 11.158 33.946 11.194 ;
      RECT 33.894 12.358 33.946 12.394 ;
      RECT 33.894 13.558 33.946 13.594 ;
      RECT 33.894 14.758 33.946 14.794 ;
      RECT 33.894 15.958 33.946 15.994 ;
      RECT 33.894 17.158 33.946 17.194 ;
      RECT 33.894 18.358 33.946 18.394 ;
      RECT 33.894 19.558 33.946 19.594 ;
      RECT 33.894 20.758 33.946 20.794 ;
      RECT 33.894 21.958 33.946 21.994 ;
      RECT 33.894 23.158 33.946 23.194 ;
      RECT 33.894 24.358 33.946 24.394 ;
      RECT 33.894 25.558 33.946 25.594 ;
      RECT 33.894 26.758 33.946 26.794 ;
      RECT 33.894 27.958 33.946 27.994 ;
      RECT 33.894 29.158 33.946 29.194 ;
      RECT 33.894 30.358 33.946 30.394 ;
      RECT 33.894 31.558 33.946 31.594 ;
      RECT 33.894 33.342 33.946 33.378 ;
      RECT 33.894 33.582 33.946 33.618 ;
      RECT 33.894 37.902 33.946 37.938 ;
      RECT 33.894 38.142 33.946 38.178 ;
      RECT 33.894 40.678 33.946 40.714 ;
      RECT 33.894 41.878 33.946 41.914 ;
      RECT 33.894 43.078 33.946 43.114 ;
      RECT 33.894 44.278 33.946 44.314 ;
      RECT 33.894 45.478 33.946 45.514 ;
      RECT 33.894 46.678 33.946 46.714 ;
      RECT 33.894 47.878 33.946 47.914 ;
      RECT 33.894 49.078 33.946 49.114 ;
      RECT 33.894 50.278 33.946 50.314 ;
      RECT 33.894 51.478 33.946 51.514 ;
      RECT 33.894 52.678 33.946 52.714 ;
      RECT 33.894 53.878 33.946 53.914 ;
      RECT 33.894 55.078 33.946 55.114 ;
      RECT 33.894 56.278 33.946 56.314 ;
      RECT 33.894 57.478 33.946 57.514 ;
      RECT 33.894 58.678 33.946 58.714 ;
      RECT 33.894 59.878 33.946 59.914 ;
      RECT 33.894 61.078 33.946 61.114 ;
      RECT 33.894 62.278 33.946 62.314 ;
      RECT 33.894 63.478 33.946 63.514 ;
      RECT 33.894 64.678 33.946 64.714 ;
      RECT 33.894 65.878 33.946 65.914 ;
      RECT 33.894 67.078 33.946 67.114 ;
      RECT 33.894 68.278 33.946 68.314 ;
      RECT 33.894 69.478 33.946 69.514 ;
      RECT 33.894 70.678 33.946 70.714 ;
      RECT 33.894 71.878 33.946 71.914 ;
      RECT 33.974 0.281 34.026 0.317 ;
      RECT 33.974 72.403 34.026 72.439 ;
      RECT 34.054 0.806 34.106 0.842 ;
      RECT 34.054 2.006 34.106 2.042 ;
      RECT 34.054 3.206 34.106 3.242 ;
      RECT 34.054 4.406 34.106 4.442 ;
      RECT 34.054 5.606 34.106 5.642 ;
      RECT 34.054 6.806 34.106 6.842 ;
      RECT 34.054 8.006 34.106 8.042 ;
      RECT 34.054 9.206 34.106 9.242 ;
      RECT 34.054 10.406 34.106 10.442 ;
      RECT 34.054 11.606 34.106 11.642 ;
      RECT 34.054 12.806 34.106 12.842 ;
      RECT 34.054 14.006 34.106 14.042 ;
      RECT 34.054 15.206 34.106 15.242 ;
      RECT 34.054 16.406 34.106 16.442 ;
      RECT 34.054 17.606 34.106 17.642 ;
      RECT 34.054 18.806 34.106 18.842 ;
      RECT 34.054 20.006 34.106 20.042 ;
      RECT 34.054 21.206 34.106 21.242 ;
      RECT 34.054 22.406 34.106 22.442 ;
      RECT 34.054 23.606 34.106 23.642 ;
      RECT 34.054 24.806 34.106 24.842 ;
      RECT 34.054 26.006 34.106 26.042 ;
      RECT 34.054 27.206 34.106 27.242 ;
      RECT 34.054 28.406 34.106 28.442 ;
      RECT 34.054 29.606 34.106 29.642 ;
      RECT 34.054 30.806 34.106 30.842 ;
      RECT 34.054 32.622 34.106 32.658 ;
      RECT 34.054 32.862 34.106 32.898 ;
      RECT 34.054 38.622 34.106 38.658 ;
      RECT 34.054 38.862 34.106 38.898 ;
      RECT 34.054 39.926 34.106 39.962 ;
      RECT 34.054 41.126 34.106 41.162 ;
      RECT 34.054 42.326 34.106 42.362 ;
      RECT 34.054 43.526 34.106 43.562 ;
      RECT 34.054 44.726 34.106 44.762 ;
      RECT 34.054 45.926 34.106 45.962 ;
      RECT 34.054 47.126 34.106 47.162 ;
      RECT 34.054 48.326 34.106 48.362 ;
      RECT 34.054 49.526 34.106 49.562 ;
      RECT 34.054 50.726 34.106 50.762 ;
      RECT 34.054 51.926 34.106 51.962 ;
      RECT 34.054 53.126 34.106 53.162 ;
      RECT 34.054 54.326 34.106 54.362 ;
      RECT 34.054 55.526 34.106 55.562 ;
      RECT 34.054 56.726 34.106 56.762 ;
      RECT 34.054 57.926 34.106 57.962 ;
      RECT 34.054 59.126 34.106 59.162 ;
      RECT 34.054 60.326 34.106 60.362 ;
      RECT 34.054 61.526 34.106 61.562 ;
      RECT 34.054 62.726 34.106 62.762 ;
      RECT 34.054 63.926 34.106 63.962 ;
      RECT 34.054 65.126 34.106 65.162 ;
      RECT 34.054 66.326 34.106 66.362 ;
      RECT 34.054 67.526 34.106 67.562 ;
      RECT 34.054 68.726 34.106 68.762 ;
      RECT 34.054 69.926 34.106 69.962 ;
      RECT 34.054 71.126 34.106 71.162 ;
      RECT 34.134 1.558 34.186 1.594 ;
      RECT 34.134 2.758 34.186 2.794 ;
      RECT 34.134 3.958 34.186 3.994 ;
      RECT 34.134 5.158 34.186 5.194 ;
      RECT 34.134 6.358 34.186 6.394 ;
      RECT 34.134 7.558 34.186 7.594 ;
      RECT 34.134 8.758 34.186 8.794 ;
      RECT 34.134 9.958 34.186 9.994 ;
      RECT 34.134 11.158 34.186 11.194 ;
      RECT 34.134 12.358 34.186 12.394 ;
      RECT 34.134 13.558 34.186 13.594 ;
      RECT 34.134 14.758 34.186 14.794 ;
      RECT 34.134 15.958 34.186 15.994 ;
      RECT 34.134 17.158 34.186 17.194 ;
      RECT 34.134 18.358 34.186 18.394 ;
      RECT 34.134 19.558 34.186 19.594 ;
      RECT 34.134 20.758 34.186 20.794 ;
      RECT 34.134 21.958 34.186 21.994 ;
      RECT 34.134 23.158 34.186 23.194 ;
      RECT 34.134 24.358 34.186 24.394 ;
      RECT 34.134 25.558 34.186 25.594 ;
      RECT 34.134 26.758 34.186 26.794 ;
      RECT 34.134 27.958 34.186 27.994 ;
      RECT 34.134 29.158 34.186 29.194 ;
      RECT 34.134 30.358 34.186 30.394 ;
      RECT 34.134 31.558 34.186 31.594 ;
      RECT 34.134 33.342 34.186 33.378 ;
      RECT 34.134 33.582 34.186 33.618 ;
      RECT 34.134 37.902 34.186 37.938 ;
      RECT 34.134 38.142 34.186 38.178 ;
      RECT 34.134 40.678 34.186 40.714 ;
      RECT 34.134 41.878 34.186 41.914 ;
      RECT 34.134 43.078 34.186 43.114 ;
      RECT 34.134 44.278 34.186 44.314 ;
      RECT 34.134 45.478 34.186 45.514 ;
      RECT 34.134 46.678 34.186 46.714 ;
      RECT 34.134 47.878 34.186 47.914 ;
      RECT 34.134 49.078 34.186 49.114 ;
      RECT 34.134 50.278 34.186 50.314 ;
      RECT 34.134 51.478 34.186 51.514 ;
      RECT 34.134 52.678 34.186 52.714 ;
      RECT 34.134 53.878 34.186 53.914 ;
      RECT 34.134 55.078 34.186 55.114 ;
      RECT 34.134 56.278 34.186 56.314 ;
      RECT 34.134 57.478 34.186 57.514 ;
      RECT 34.134 58.678 34.186 58.714 ;
      RECT 34.134 59.878 34.186 59.914 ;
      RECT 34.134 61.078 34.186 61.114 ;
      RECT 34.134 62.278 34.186 62.314 ;
      RECT 34.134 63.478 34.186 63.514 ;
      RECT 34.134 64.678 34.186 64.714 ;
      RECT 34.134 65.878 34.186 65.914 ;
      RECT 34.134 67.078 34.186 67.114 ;
      RECT 34.134 68.278 34.186 68.314 ;
      RECT 34.134 69.478 34.186 69.514 ;
      RECT 34.134 70.678 34.186 70.714 ;
      RECT 34.134 71.878 34.186 71.914 ;
      RECT 34.214 0.806 34.266 0.842 ;
      RECT 34.214 2.006 34.266 2.042 ;
      RECT 34.214 3.206 34.266 3.242 ;
      RECT 34.214 4.406 34.266 4.442 ;
      RECT 34.214 5.606 34.266 5.642 ;
      RECT 34.214 6.806 34.266 6.842 ;
      RECT 34.214 8.006 34.266 8.042 ;
      RECT 34.214 9.206 34.266 9.242 ;
      RECT 34.214 10.406 34.266 10.442 ;
      RECT 34.214 11.606 34.266 11.642 ;
      RECT 34.214 12.806 34.266 12.842 ;
      RECT 34.214 14.006 34.266 14.042 ;
      RECT 34.214 15.206 34.266 15.242 ;
      RECT 34.214 16.406 34.266 16.442 ;
      RECT 34.214 17.606 34.266 17.642 ;
      RECT 34.214 18.806 34.266 18.842 ;
      RECT 34.214 20.006 34.266 20.042 ;
      RECT 34.214 21.206 34.266 21.242 ;
      RECT 34.214 22.406 34.266 22.442 ;
      RECT 34.214 23.606 34.266 23.642 ;
      RECT 34.214 24.806 34.266 24.842 ;
      RECT 34.214 26.006 34.266 26.042 ;
      RECT 34.214 27.206 34.266 27.242 ;
      RECT 34.214 28.406 34.266 28.442 ;
      RECT 34.214 29.606 34.266 29.642 ;
      RECT 34.214 30.806 34.266 30.842 ;
      RECT 34.214 32.622 34.266 32.658 ;
      RECT 34.214 32.862 34.266 32.898 ;
      RECT 34.214 38.622 34.266 38.658 ;
      RECT 34.214 38.862 34.266 38.898 ;
      RECT 34.214 39.926 34.266 39.962 ;
      RECT 34.214 41.126 34.266 41.162 ;
      RECT 34.214 42.326 34.266 42.362 ;
      RECT 34.214 43.526 34.266 43.562 ;
      RECT 34.214 44.726 34.266 44.762 ;
      RECT 34.214 45.926 34.266 45.962 ;
      RECT 34.214 47.126 34.266 47.162 ;
      RECT 34.214 48.326 34.266 48.362 ;
      RECT 34.214 49.526 34.266 49.562 ;
      RECT 34.214 50.726 34.266 50.762 ;
      RECT 34.214 51.926 34.266 51.962 ;
      RECT 34.214 53.126 34.266 53.162 ;
      RECT 34.214 54.326 34.266 54.362 ;
      RECT 34.214 55.526 34.266 55.562 ;
      RECT 34.214 56.726 34.266 56.762 ;
      RECT 34.214 57.926 34.266 57.962 ;
      RECT 34.214 59.126 34.266 59.162 ;
      RECT 34.214 60.326 34.266 60.362 ;
      RECT 34.214 61.526 34.266 61.562 ;
      RECT 34.214 62.726 34.266 62.762 ;
      RECT 34.214 63.926 34.266 63.962 ;
      RECT 34.214 65.126 34.266 65.162 ;
      RECT 34.214 66.326 34.266 66.362 ;
      RECT 34.214 67.526 34.266 67.562 ;
      RECT 34.214 68.726 34.266 68.762 ;
      RECT 34.214 69.926 34.266 69.962 ;
      RECT 34.214 71.126 34.266 71.162 ;
      RECT 34.294 1.558 34.346 1.594 ;
      RECT 34.294 2.758 34.346 2.794 ;
      RECT 34.294 3.958 34.346 3.994 ;
      RECT 34.294 5.158 34.346 5.194 ;
      RECT 34.294 6.358 34.346 6.394 ;
      RECT 34.294 7.558 34.346 7.594 ;
      RECT 34.294 8.758 34.346 8.794 ;
      RECT 34.294 9.958 34.346 9.994 ;
      RECT 34.294 11.158 34.346 11.194 ;
      RECT 34.294 12.358 34.346 12.394 ;
      RECT 34.294 13.558 34.346 13.594 ;
      RECT 34.294 14.758 34.346 14.794 ;
      RECT 34.294 15.958 34.346 15.994 ;
      RECT 34.294 17.158 34.346 17.194 ;
      RECT 34.294 18.358 34.346 18.394 ;
      RECT 34.294 19.558 34.346 19.594 ;
      RECT 34.294 20.758 34.346 20.794 ;
      RECT 34.294 21.958 34.346 21.994 ;
      RECT 34.294 23.158 34.346 23.194 ;
      RECT 34.294 24.358 34.346 24.394 ;
      RECT 34.294 25.558 34.346 25.594 ;
      RECT 34.294 26.758 34.346 26.794 ;
      RECT 34.294 27.958 34.346 27.994 ;
      RECT 34.294 29.158 34.346 29.194 ;
      RECT 34.294 30.358 34.346 30.394 ;
      RECT 34.294 31.558 34.346 31.594 ;
      RECT 34.294 33.342 34.346 33.378 ;
      RECT 34.294 33.582 34.346 33.618 ;
      RECT 34.294 37.902 34.346 37.938 ;
      RECT 34.294 38.142 34.346 38.178 ;
      RECT 34.294 40.678 34.346 40.714 ;
      RECT 34.294 41.878 34.346 41.914 ;
      RECT 34.294 43.078 34.346 43.114 ;
      RECT 34.294 44.278 34.346 44.314 ;
      RECT 34.294 45.478 34.346 45.514 ;
      RECT 34.294 46.678 34.346 46.714 ;
      RECT 34.294 47.878 34.346 47.914 ;
      RECT 34.294 49.078 34.346 49.114 ;
      RECT 34.294 50.278 34.346 50.314 ;
      RECT 34.294 51.478 34.346 51.514 ;
      RECT 34.294 52.678 34.346 52.714 ;
      RECT 34.294 53.878 34.346 53.914 ;
      RECT 34.294 55.078 34.346 55.114 ;
      RECT 34.294 56.278 34.346 56.314 ;
      RECT 34.294 57.478 34.346 57.514 ;
      RECT 34.294 58.678 34.346 58.714 ;
      RECT 34.294 59.878 34.346 59.914 ;
      RECT 34.294 61.078 34.346 61.114 ;
      RECT 34.294 62.278 34.346 62.314 ;
      RECT 34.294 63.478 34.346 63.514 ;
      RECT 34.294 64.678 34.346 64.714 ;
      RECT 34.294 65.878 34.346 65.914 ;
      RECT 34.294 67.078 34.346 67.114 ;
      RECT 34.294 68.278 34.346 68.314 ;
      RECT 34.294 69.478 34.346 69.514 ;
      RECT 34.294 70.678 34.346 70.714 ;
      RECT 34.294 71.878 34.346 71.914 ;
      RECT 34.374 0.281 34.426 0.317 ;
      RECT 34.374 72.403 34.426 72.439 ;
      RECT 34.454 0.806 34.506 0.842 ;
      RECT 34.454 2.006 34.506 2.042 ;
      RECT 34.454 3.206 34.506 3.242 ;
      RECT 34.454 4.406 34.506 4.442 ;
      RECT 34.454 5.606 34.506 5.642 ;
      RECT 34.454 6.806 34.506 6.842 ;
      RECT 34.454 8.006 34.506 8.042 ;
      RECT 34.454 9.206 34.506 9.242 ;
      RECT 34.454 10.406 34.506 10.442 ;
      RECT 34.454 11.606 34.506 11.642 ;
      RECT 34.454 12.806 34.506 12.842 ;
      RECT 34.454 14.006 34.506 14.042 ;
      RECT 34.454 15.206 34.506 15.242 ;
      RECT 34.454 16.406 34.506 16.442 ;
      RECT 34.454 17.606 34.506 17.642 ;
      RECT 34.454 18.806 34.506 18.842 ;
      RECT 34.454 20.006 34.506 20.042 ;
      RECT 34.454 21.206 34.506 21.242 ;
      RECT 34.454 22.406 34.506 22.442 ;
      RECT 34.454 23.606 34.506 23.642 ;
      RECT 34.454 24.806 34.506 24.842 ;
      RECT 34.454 26.006 34.506 26.042 ;
      RECT 34.454 27.206 34.506 27.242 ;
      RECT 34.454 28.406 34.506 28.442 ;
      RECT 34.454 29.606 34.506 29.642 ;
      RECT 34.454 30.806 34.506 30.842 ;
      RECT 34.454 32.622 34.506 32.658 ;
      RECT 34.454 32.862 34.506 32.898 ;
      RECT 34.454 34.302 34.506 34.338 ;
      RECT 34.454 34.782 34.506 34.818 ;
      RECT 34.454 36.702 34.506 36.738 ;
      RECT 34.454 37.182 34.506 37.218 ;
      RECT 34.454 38.622 34.506 38.658 ;
      RECT 34.454 38.862 34.506 38.898 ;
      RECT 34.454 39.926 34.506 39.962 ;
      RECT 34.454 41.126 34.506 41.162 ;
      RECT 34.454 42.326 34.506 42.362 ;
      RECT 34.454 43.526 34.506 43.562 ;
      RECT 34.454 44.726 34.506 44.762 ;
      RECT 34.454 45.926 34.506 45.962 ;
      RECT 34.454 47.126 34.506 47.162 ;
      RECT 34.454 48.326 34.506 48.362 ;
      RECT 34.454 49.526 34.506 49.562 ;
      RECT 34.454 50.726 34.506 50.762 ;
      RECT 34.454 51.926 34.506 51.962 ;
      RECT 34.454 53.126 34.506 53.162 ;
      RECT 34.454 54.326 34.506 54.362 ;
      RECT 34.454 55.526 34.506 55.562 ;
      RECT 34.454 56.726 34.506 56.762 ;
      RECT 34.454 57.926 34.506 57.962 ;
      RECT 34.454 59.126 34.506 59.162 ;
      RECT 34.454 60.326 34.506 60.362 ;
      RECT 34.454 61.526 34.506 61.562 ;
      RECT 34.454 62.726 34.506 62.762 ;
      RECT 34.454 63.926 34.506 63.962 ;
      RECT 34.454 65.126 34.506 65.162 ;
      RECT 34.454 66.326 34.506 66.362 ;
      RECT 34.454 67.526 34.506 67.562 ;
      RECT 34.454 68.726 34.506 68.762 ;
      RECT 34.454 69.926 34.506 69.962 ;
      RECT 34.454 71.126 34.506 71.162 ;
      RECT 34.534 1.558 34.586 1.594 ;
      RECT 34.534 2.758 34.586 2.794 ;
      RECT 34.534 3.958 34.586 3.994 ;
      RECT 34.534 5.158 34.586 5.194 ;
      RECT 34.534 6.358 34.586 6.394 ;
      RECT 34.534 7.558 34.586 7.594 ;
      RECT 34.534 8.758 34.586 8.794 ;
      RECT 34.534 9.958 34.586 9.994 ;
      RECT 34.534 11.158 34.586 11.194 ;
      RECT 34.534 12.358 34.586 12.394 ;
      RECT 34.534 13.558 34.586 13.594 ;
      RECT 34.534 14.758 34.586 14.794 ;
      RECT 34.534 15.958 34.586 15.994 ;
      RECT 34.534 17.158 34.586 17.194 ;
      RECT 34.534 18.358 34.586 18.394 ;
      RECT 34.534 19.558 34.586 19.594 ;
      RECT 34.534 20.758 34.586 20.794 ;
      RECT 34.534 21.958 34.586 21.994 ;
      RECT 34.534 23.158 34.586 23.194 ;
      RECT 34.534 24.358 34.586 24.394 ;
      RECT 34.534 25.558 34.586 25.594 ;
      RECT 34.534 26.758 34.586 26.794 ;
      RECT 34.534 27.958 34.586 27.994 ;
      RECT 34.534 29.158 34.586 29.194 ;
      RECT 34.534 30.358 34.586 30.394 ;
      RECT 34.534 31.558 34.586 31.594 ;
      RECT 34.534 33.342 34.586 33.378 ;
      RECT 34.534 33.582 34.586 33.618 ;
      RECT 34.534 37.902 34.586 37.938 ;
      RECT 34.534 38.142 34.586 38.178 ;
      RECT 34.534 40.678 34.586 40.714 ;
      RECT 34.534 41.878 34.586 41.914 ;
      RECT 34.534 43.078 34.586 43.114 ;
      RECT 34.534 44.278 34.586 44.314 ;
      RECT 34.534 45.478 34.586 45.514 ;
      RECT 34.534 46.678 34.586 46.714 ;
      RECT 34.534 47.878 34.586 47.914 ;
      RECT 34.534 49.078 34.586 49.114 ;
      RECT 34.534 50.278 34.586 50.314 ;
      RECT 34.534 51.478 34.586 51.514 ;
      RECT 34.534 52.678 34.586 52.714 ;
      RECT 34.534 53.878 34.586 53.914 ;
      RECT 34.534 55.078 34.586 55.114 ;
      RECT 34.534 56.278 34.586 56.314 ;
      RECT 34.534 57.478 34.586 57.514 ;
      RECT 34.534 58.678 34.586 58.714 ;
      RECT 34.534 59.878 34.586 59.914 ;
      RECT 34.534 61.078 34.586 61.114 ;
      RECT 34.534 62.278 34.586 62.314 ;
      RECT 34.534 63.478 34.586 63.514 ;
      RECT 34.534 64.678 34.586 64.714 ;
      RECT 34.534 65.878 34.586 65.914 ;
      RECT 34.534 67.078 34.586 67.114 ;
      RECT 34.534 68.278 34.586 68.314 ;
      RECT 34.534 69.478 34.586 69.514 ;
      RECT 34.534 70.678 34.586 70.714 ;
      RECT 34.534 71.878 34.586 71.914 ;
      RECT 34.614 0.806 34.666 0.842 ;
      RECT 34.614 2.006 34.666 2.042 ;
      RECT 34.614 3.206 34.666 3.242 ;
      RECT 34.614 4.406 34.666 4.442 ;
      RECT 34.614 5.606 34.666 5.642 ;
      RECT 34.614 6.806 34.666 6.842 ;
      RECT 34.614 8.006 34.666 8.042 ;
      RECT 34.614 9.206 34.666 9.242 ;
      RECT 34.614 10.406 34.666 10.442 ;
      RECT 34.614 11.606 34.666 11.642 ;
      RECT 34.614 12.806 34.666 12.842 ;
      RECT 34.614 14.006 34.666 14.042 ;
      RECT 34.614 15.206 34.666 15.242 ;
      RECT 34.614 16.406 34.666 16.442 ;
      RECT 34.614 17.606 34.666 17.642 ;
      RECT 34.614 18.806 34.666 18.842 ;
      RECT 34.614 20.006 34.666 20.042 ;
      RECT 34.614 21.206 34.666 21.242 ;
      RECT 34.614 22.406 34.666 22.442 ;
      RECT 34.614 23.606 34.666 23.642 ;
      RECT 34.614 24.806 34.666 24.842 ;
      RECT 34.614 26.006 34.666 26.042 ;
      RECT 34.614 27.206 34.666 27.242 ;
      RECT 34.614 28.406 34.666 28.442 ;
      RECT 34.614 29.606 34.666 29.642 ;
      RECT 34.614 30.806 34.666 30.842 ;
      RECT 34.614 32.622 34.666 32.658 ;
      RECT 34.614 32.862 34.666 32.898 ;
      RECT 34.614 38.622 34.666 38.658 ;
      RECT 34.614 38.862 34.666 38.898 ;
      RECT 34.614 39.926 34.666 39.962 ;
      RECT 34.614 41.126 34.666 41.162 ;
      RECT 34.614 42.326 34.666 42.362 ;
      RECT 34.614 43.526 34.666 43.562 ;
      RECT 34.614 44.726 34.666 44.762 ;
      RECT 34.614 45.926 34.666 45.962 ;
      RECT 34.614 47.126 34.666 47.162 ;
      RECT 34.614 48.326 34.666 48.362 ;
      RECT 34.614 49.526 34.666 49.562 ;
      RECT 34.614 50.726 34.666 50.762 ;
      RECT 34.614 51.926 34.666 51.962 ;
      RECT 34.614 53.126 34.666 53.162 ;
      RECT 34.614 54.326 34.666 54.362 ;
      RECT 34.614 55.526 34.666 55.562 ;
      RECT 34.614 56.726 34.666 56.762 ;
      RECT 34.614 57.926 34.666 57.962 ;
      RECT 34.614 59.126 34.666 59.162 ;
      RECT 34.614 60.326 34.666 60.362 ;
      RECT 34.614 61.526 34.666 61.562 ;
      RECT 34.614 62.726 34.666 62.762 ;
      RECT 34.614 63.926 34.666 63.962 ;
      RECT 34.614 65.126 34.666 65.162 ;
      RECT 34.614 66.326 34.666 66.362 ;
      RECT 34.614 67.526 34.666 67.562 ;
      RECT 34.614 68.726 34.666 68.762 ;
      RECT 34.614 69.926 34.666 69.962 ;
      RECT 34.614 71.126 34.666 71.162 ;
      RECT 34.694 1.558 34.746 1.594 ;
      RECT 34.694 2.758 34.746 2.794 ;
      RECT 34.694 3.958 34.746 3.994 ;
      RECT 34.694 5.158 34.746 5.194 ;
      RECT 34.694 6.358 34.746 6.394 ;
      RECT 34.694 7.558 34.746 7.594 ;
      RECT 34.694 8.758 34.746 8.794 ;
      RECT 34.694 9.958 34.746 9.994 ;
      RECT 34.694 11.158 34.746 11.194 ;
      RECT 34.694 12.358 34.746 12.394 ;
      RECT 34.694 13.558 34.746 13.594 ;
      RECT 34.694 14.758 34.746 14.794 ;
      RECT 34.694 15.958 34.746 15.994 ;
      RECT 34.694 17.158 34.746 17.194 ;
      RECT 34.694 18.358 34.746 18.394 ;
      RECT 34.694 19.558 34.746 19.594 ;
      RECT 34.694 20.758 34.746 20.794 ;
      RECT 34.694 21.958 34.746 21.994 ;
      RECT 34.694 23.158 34.746 23.194 ;
      RECT 34.694 24.358 34.746 24.394 ;
      RECT 34.694 25.558 34.746 25.594 ;
      RECT 34.694 26.758 34.746 26.794 ;
      RECT 34.694 27.958 34.746 27.994 ;
      RECT 34.694 29.158 34.746 29.194 ;
      RECT 34.694 30.358 34.746 30.394 ;
      RECT 34.694 31.558 34.746 31.594 ;
      RECT 34.694 33.342 34.746 33.378 ;
      RECT 34.694 33.582 34.746 33.618 ;
      RECT 34.694 37.902 34.746 37.938 ;
      RECT 34.694 38.142 34.746 38.178 ;
      RECT 34.694 40.678 34.746 40.714 ;
      RECT 34.694 41.878 34.746 41.914 ;
      RECT 34.694 43.078 34.746 43.114 ;
      RECT 34.694 44.278 34.746 44.314 ;
      RECT 34.694 45.478 34.746 45.514 ;
      RECT 34.694 46.678 34.746 46.714 ;
      RECT 34.694 47.878 34.746 47.914 ;
      RECT 34.694 49.078 34.746 49.114 ;
      RECT 34.694 50.278 34.746 50.314 ;
      RECT 34.694 51.478 34.746 51.514 ;
      RECT 34.694 52.678 34.746 52.714 ;
      RECT 34.694 53.878 34.746 53.914 ;
      RECT 34.694 55.078 34.746 55.114 ;
      RECT 34.694 56.278 34.746 56.314 ;
      RECT 34.694 57.478 34.746 57.514 ;
      RECT 34.694 58.678 34.746 58.714 ;
      RECT 34.694 59.878 34.746 59.914 ;
      RECT 34.694 61.078 34.746 61.114 ;
      RECT 34.694 62.278 34.746 62.314 ;
      RECT 34.694 63.478 34.746 63.514 ;
      RECT 34.694 64.678 34.746 64.714 ;
      RECT 34.694 65.878 34.746 65.914 ;
      RECT 34.694 67.078 34.746 67.114 ;
      RECT 34.694 68.278 34.746 68.314 ;
      RECT 34.694 69.478 34.746 69.514 ;
      RECT 34.694 70.678 34.746 70.714 ;
      RECT 34.694 71.878 34.746 71.914 ;
      RECT 34.774 0.281 34.826 0.317 ;
      RECT 34.774 72.403 34.826 72.439 ;
      RECT 34.854 0.806 34.906 0.842 ;
      RECT 34.854 2.006 34.906 2.042 ;
      RECT 34.854 3.206 34.906 3.242 ;
      RECT 34.854 4.406 34.906 4.442 ;
      RECT 34.854 5.606 34.906 5.642 ;
      RECT 34.854 6.806 34.906 6.842 ;
      RECT 34.854 8.006 34.906 8.042 ;
      RECT 34.854 9.206 34.906 9.242 ;
      RECT 34.854 10.406 34.906 10.442 ;
      RECT 34.854 11.606 34.906 11.642 ;
      RECT 34.854 12.806 34.906 12.842 ;
      RECT 34.854 14.006 34.906 14.042 ;
      RECT 34.854 15.206 34.906 15.242 ;
      RECT 34.854 16.406 34.906 16.442 ;
      RECT 34.854 17.606 34.906 17.642 ;
      RECT 34.854 18.806 34.906 18.842 ;
      RECT 34.854 20.006 34.906 20.042 ;
      RECT 34.854 21.206 34.906 21.242 ;
      RECT 34.854 22.406 34.906 22.442 ;
      RECT 34.854 23.606 34.906 23.642 ;
      RECT 34.854 24.806 34.906 24.842 ;
      RECT 34.854 26.006 34.906 26.042 ;
      RECT 34.854 27.206 34.906 27.242 ;
      RECT 34.854 28.406 34.906 28.442 ;
      RECT 34.854 29.606 34.906 29.642 ;
      RECT 34.854 30.806 34.906 30.842 ;
      RECT 34.854 32.622 34.906 32.658 ;
      RECT 34.854 32.862 34.906 32.898 ;
      RECT 34.854 38.622 34.906 38.658 ;
      RECT 34.854 38.862 34.906 38.898 ;
      RECT 34.854 39.926 34.906 39.962 ;
      RECT 34.854 41.126 34.906 41.162 ;
      RECT 34.854 42.326 34.906 42.362 ;
      RECT 34.854 43.526 34.906 43.562 ;
      RECT 34.854 44.726 34.906 44.762 ;
      RECT 34.854 45.926 34.906 45.962 ;
      RECT 34.854 47.126 34.906 47.162 ;
      RECT 34.854 48.326 34.906 48.362 ;
      RECT 34.854 49.526 34.906 49.562 ;
      RECT 34.854 50.726 34.906 50.762 ;
      RECT 34.854 51.926 34.906 51.962 ;
      RECT 34.854 53.126 34.906 53.162 ;
      RECT 34.854 54.326 34.906 54.362 ;
      RECT 34.854 55.526 34.906 55.562 ;
      RECT 34.854 56.726 34.906 56.762 ;
      RECT 34.854 57.926 34.906 57.962 ;
      RECT 34.854 59.126 34.906 59.162 ;
      RECT 34.854 60.326 34.906 60.362 ;
      RECT 34.854 61.526 34.906 61.562 ;
      RECT 34.854 62.726 34.906 62.762 ;
      RECT 34.854 63.926 34.906 63.962 ;
      RECT 34.854 65.126 34.906 65.162 ;
      RECT 34.854 66.326 34.906 66.362 ;
      RECT 34.854 67.526 34.906 67.562 ;
      RECT 34.854 68.726 34.906 68.762 ;
      RECT 34.854 69.926 34.906 69.962 ;
      RECT 34.854 71.126 34.906 71.162 ;
      RECT 34.934 1.558 34.986 1.594 ;
      RECT 34.934 2.758 34.986 2.794 ;
      RECT 34.934 3.958 34.986 3.994 ;
      RECT 34.934 5.158 34.986 5.194 ;
      RECT 34.934 6.358 34.986 6.394 ;
      RECT 34.934 7.558 34.986 7.594 ;
      RECT 34.934 8.758 34.986 8.794 ;
      RECT 34.934 9.958 34.986 9.994 ;
      RECT 34.934 11.158 34.986 11.194 ;
      RECT 34.934 12.358 34.986 12.394 ;
      RECT 34.934 13.558 34.986 13.594 ;
      RECT 34.934 14.758 34.986 14.794 ;
      RECT 34.934 15.958 34.986 15.994 ;
      RECT 34.934 17.158 34.986 17.194 ;
      RECT 34.934 18.358 34.986 18.394 ;
      RECT 34.934 19.558 34.986 19.594 ;
      RECT 34.934 20.758 34.986 20.794 ;
      RECT 34.934 21.958 34.986 21.994 ;
      RECT 34.934 23.158 34.986 23.194 ;
      RECT 34.934 24.358 34.986 24.394 ;
      RECT 34.934 25.558 34.986 25.594 ;
      RECT 34.934 26.758 34.986 26.794 ;
      RECT 34.934 27.958 34.986 27.994 ;
      RECT 34.934 29.158 34.986 29.194 ;
      RECT 34.934 30.358 34.986 30.394 ;
      RECT 34.934 31.558 34.986 31.594 ;
      RECT 34.934 33.342 34.986 33.378 ;
      RECT 34.934 33.582 34.986 33.618 ;
      RECT 34.934 37.902 34.986 37.938 ;
      RECT 34.934 38.142 34.986 38.178 ;
      RECT 34.934 40.678 34.986 40.714 ;
      RECT 34.934 41.878 34.986 41.914 ;
      RECT 34.934 43.078 34.986 43.114 ;
      RECT 34.934 44.278 34.986 44.314 ;
      RECT 34.934 45.478 34.986 45.514 ;
      RECT 34.934 46.678 34.986 46.714 ;
      RECT 34.934 47.878 34.986 47.914 ;
      RECT 34.934 49.078 34.986 49.114 ;
      RECT 34.934 50.278 34.986 50.314 ;
      RECT 34.934 51.478 34.986 51.514 ;
      RECT 34.934 52.678 34.986 52.714 ;
      RECT 34.934 53.878 34.986 53.914 ;
      RECT 34.934 55.078 34.986 55.114 ;
      RECT 34.934 56.278 34.986 56.314 ;
      RECT 34.934 57.478 34.986 57.514 ;
      RECT 34.934 58.678 34.986 58.714 ;
      RECT 34.934 59.878 34.986 59.914 ;
      RECT 34.934 61.078 34.986 61.114 ;
      RECT 34.934 62.278 34.986 62.314 ;
      RECT 34.934 63.478 34.986 63.514 ;
      RECT 34.934 64.678 34.986 64.714 ;
      RECT 34.934 65.878 34.986 65.914 ;
      RECT 34.934 67.078 34.986 67.114 ;
      RECT 34.934 68.278 34.986 68.314 ;
      RECT 34.934 69.478 34.986 69.514 ;
      RECT 34.934 70.678 34.986 70.714 ;
      RECT 34.934 71.878 34.986 71.914 ;
      RECT 35.014 0.806 35.066 0.842 ;
      RECT 35.014 2.006 35.066 2.042 ;
      RECT 35.014 3.206 35.066 3.242 ;
      RECT 35.014 4.406 35.066 4.442 ;
      RECT 35.014 5.606 35.066 5.642 ;
      RECT 35.014 6.806 35.066 6.842 ;
      RECT 35.014 8.006 35.066 8.042 ;
      RECT 35.014 9.206 35.066 9.242 ;
      RECT 35.014 10.406 35.066 10.442 ;
      RECT 35.014 11.606 35.066 11.642 ;
      RECT 35.014 12.806 35.066 12.842 ;
      RECT 35.014 14.006 35.066 14.042 ;
      RECT 35.014 15.206 35.066 15.242 ;
      RECT 35.014 16.406 35.066 16.442 ;
      RECT 35.014 17.606 35.066 17.642 ;
      RECT 35.014 18.806 35.066 18.842 ;
      RECT 35.014 20.006 35.066 20.042 ;
      RECT 35.014 21.206 35.066 21.242 ;
      RECT 35.014 22.406 35.066 22.442 ;
      RECT 35.014 23.606 35.066 23.642 ;
      RECT 35.014 24.806 35.066 24.842 ;
      RECT 35.014 26.006 35.066 26.042 ;
      RECT 35.014 27.206 35.066 27.242 ;
      RECT 35.014 28.406 35.066 28.442 ;
      RECT 35.014 29.606 35.066 29.642 ;
      RECT 35.014 30.806 35.066 30.842 ;
      RECT 35.014 32.622 35.066 32.658 ;
      RECT 35.014 32.862 35.066 32.898 ;
      RECT 35.014 38.622 35.066 38.658 ;
      RECT 35.014 38.862 35.066 38.898 ;
      RECT 35.014 39.926 35.066 39.962 ;
      RECT 35.014 41.126 35.066 41.162 ;
      RECT 35.014 42.326 35.066 42.362 ;
      RECT 35.014 43.526 35.066 43.562 ;
      RECT 35.014 44.726 35.066 44.762 ;
      RECT 35.014 45.926 35.066 45.962 ;
      RECT 35.014 47.126 35.066 47.162 ;
      RECT 35.014 48.326 35.066 48.362 ;
      RECT 35.014 49.526 35.066 49.562 ;
      RECT 35.014 50.726 35.066 50.762 ;
      RECT 35.014 51.926 35.066 51.962 ;
      RECT 35.014 53.126 35.066 53.162 ;
      RECT 35.014 54.326 35.066 54.362 ;
      RECT 35.014 55.526 35.066 55.562 ;
      RECT 35.014 56.726 35.066 56.762 ;
      RECT 35.014 57.926 35.066 57.962 ;
      RECT 35.014 59.126 35.066 59.162 ;
      RECT 35.014 60.326 35.066 60.362 ;
      RECT 35.014 61.526 35.066 61.562 ;
      RECT 35.014 62.726 35.066 62.762 ;
      RECT 35.014 63.926 35.066 63.962 ;
      RECT 35.014 65.126 35.066 65.162 ;
      RECT 35.014 66.326 35.066 66.362 ;
      RECT 35.014 67.526 35.066 67.562 ;
      RECT 35.014 68.726 35.066 68.762 ;
      RECT 35.014 69.926 35.066 69.962 ;
      RECT 35.014 71.126 35.066 71.162 ;
      RECT 35.094 1.558 35.146 1.594 ;
      RECT 35.094 2.758 35.146 2.794 ;
      RECT 35.094 3.958 35.146 3.994 ;
      RECT 35.094 5.158 35.146 5.194 ;
      RECT 35.094 6.358 35.146 6.394 ;
      RECT 35.094 7.558 35.146 7.594 ;
      RECT 35.094 8.758 35.146 8.794 ;
      RECT 35.094 9.958 35.146 9.994 ;
      RECT 35.094 11.158 35.146 11.194 ;
      RECT 35.094 12.358 35.146 12.394 ;
      RECT 35.094 13.558 35.146 13.594 ;
      RECT 35.094 14.758 35.146 14.794 ;
      RECT 35.094 15.958 35.146 15.994 ;
      RECT 35.094 17.158 35.146 17.194 ;
      RECT 35.094 18.358 35.146 18.394 ;
      RECT 35.094 19.558 35.146 19.594 ;
      RECT 35.094 20.758 35.146 20.794 ;
      RECT 35.094 21.958 35.146 21.994 ;
      RECT 35.094 23.158 35.146 23.194 ;
      RECT 35.094 24.358 35.146 24.394 ;
      RECT 35.094 25.558 35.146 25.594 ;
      RECT 35.094 26.758 35.146 26.794 ;
      RECT 35.094 27.958 35.146 27.994 ;
      RECT 35.094 29.158 35.146 29.194 ;
      RECT 35.094 30.358 35.146 30.394 ;
      RECT 35.094 31.558 35.146 31.594 ;
      RECT 35.094 33.342 35.146 33.378 ;
      RECT 35.094 33.582 35.146 33.618 ;
      RECT 35.094 37.902 35.146 37.938 ;
      RECT 35.094 38.142 35.146 38.178 ;
      RECT 35.094 40.678 35.146 40.714 ;
      RECT 35.094 41.878 35.146 41.914 ;
      RECT 35.094 43.078 35.146 43.114 ;
      RECT 35.094 44.278 35.146 44.314 ;
      RECT 35.094 45.478 35.146 45.514 ;
      RECT 35.094 46.678 35.146 46.714 ;
      RECT 35.094 47.878 35.146 47.914 ;
      RECT 35.094 49.078 35.146 49.114 ;
      RECT 35.094 50.278 35.146 50.314 ;
      RECT 35.094 51.478 35.146 51.514 ;
      RECT 35.094 52.678 35.146 52.714 ;
      RECT 35.094 53.878 35.146 53.914 ;
      RECT 35.094 55.078 35.146 55.114 ;
      RECT 35.094 56.278 35.146 56.314 ;
      RECT 35.094 57.478 35.146 57.514 ;
      RECT 35.094 58.678 35.146 58.714 ;
      RECT 35.094 59.878 35.146 59.914 ;
      RECT 35.094 61.078 35.146 61.114 ;
      RECT 35.094 62.278 35.146 62.314 ;
      RECT 35.094 63.478 35.146 63.514 ;
      RECT 35.094 64.678 35.146 64.714 ;
      RECT 35.094 65.878 35.146 65.914 ;
      RECT 35.094 67.078 35.146 67.114 ;
      RECT 35.094 68.278 35.146 68.314 ;
      RECT 35.094 69.478 35.146 69.514 ;
      RECT 35.094 70.678 35.146 70.714 ;
      RECT 35.094 71.878 35.146 71.914 ;
      RECT 35.174 0.281 35.226 0.317 ;
      RECT 35.174 72.403 35.226 72.439 ;
      RECT 35.254 0.806 35.306 0.842 ;
      RECT 35.254 2.006 35.306 2.042 ;
      RECT 35.254 3.206 35.306 3.242 ;
      RECT 35.254 4.406 35.306 4.442 ;
      RECT 35.254 5.606 35.306 5.642 ;
      RECT 35.254 6.806 35.306 6.842 ;
      RECT 35.254 8.006 35.306 8.042 ;
      RECT 35.254 9.206 35.306 9.242 ;
      RECT 35.254 10.406 35.306 10.442 ;
      RECT 35.254 11.606 35.306 11.642 ;
      RECT 35.254 12.806 35.306 12.842 ;
      RECT 35.254 14.006 35.306 14.042 ;
      RECT 35.254 15.206 35.306 15.242 ;
      RECT 35.254 16.406 35.306 16.442 ;
      RECT 35.254 17.606 35.306 17.642 ;
      RECT 35.254 18.806 35.306 18.842 ;
      RECT 35.254 20.006 35.306 20.042 ;
      RECT 35.254 21.206 35.306 21.242 ;
      RECT 35.254 22.406 35.306 22.442 ;
      RECT 35.254 23.606 35.306 23.642 ;
      RECT 35.254 24.806 35.306 24.842 ;
      RECT 35.254 26.006 35.306 26.042 ;
      RECT 35.254 27.206 35.306 27.242 ;
      RECT 35.254 28.406 35.306 28.442 ;
      RECT 35.254 29.606 35.306 29.642 ;
      RECT 35.254 30.806 35.306 30.842 ;
      RECT 35.254 32.622 35.306 32.658 ;
      RECT 35.254 32.862 35.306 32.898 ;
      RECT 35.254 34.302 35.306 34.338 ;
      RECT 35.254 34.782 35.306 34.818 ;
      RECT 35.254 36.702 35.306 36.738 ;
      RECT 35.254 37.182 35.306 37.218 ;
      RECT 35.254 38.622 35.306 38.658 ;
      RECT 35.254 38.862 35.306 38.898 ;
      RECT 35.254 39.926 35.306 39.962 ;
      RECT 35.254 41.126 35.306 41.162 ;
      RECT 35.254 42.326 35.306 42.362 ;
      RECT 35.254 43.526 35.306 43.562 ;
      RECT 35.254 44.726 35.306 44.762 ;
      RECT 35.254 45.926 35.306 45.962 ;
      RECT 35.254 47.126 35.306 47.162 ;
      RECT 35.254 48.326 35.306 48.362 ;
      RECT 35.254 49.526 35.306 49.562 ;
      RECT 35.254 50.726 35.306 50.762 ;
      RECT 35.254 51.926 35.306 51.962 ;
      RECT 35.254 53.126 35.306 53.162 ;
      RECT 35.254 54.326 35.306 54.362 ;
      RECT 35.254 55.526 35.306 55.562 ;
      RECT 35.254 56.726 35.306 56.762 ;
      RECT 35.254 57.926 35.306 57.962 ;
      RECT 35.254 59.126 35.306 59.162 ;
      RECT 35.254 60.326 35.306 60.362 ;
      RECT 35.254 61.526 35.306 61.562 ;
      RECT 35.254 62.726 35.306 62.762 ;
      RECT 35.254 63.926 35.306 63.962 ;
      RECT 35.254 65.126 35.306 65.162 ;
      RECT 35.254 66.326 35.306 66.362 ;
      RECT 35.254 67.526 35.306 67.562 ;
      RECT 35.254 68.726 35.306 68.762 ;
      RECT 35.254 69.926 35.306 69.962 ;
      RECT 35.254 71.126 35.306 71.162 ;
      RECT 35.334 1.558 35.386 1.594 ;
      RECT 35.334 2.758 35.386 2.794 ;
      RECT 35.334 3.958 35.386 3.994 ;
      RECT 35.334 5.158 35.386 5.194 ;
      RECT 35.334 6.358 35.386 6.394 ;
      RECT 35.334 7.558 35.386 7.594 ;
      RECT 35.334 8.758 35.386 8.794 ;
      RECT 35.334 9.958 35.386 9.994 ;
      RECT 35.334 11.158 35.386 11.194 ;
      RECT 35.334 12.358 35.386 12.394 ;
      RECT 35.334 13.558 35.386 13.594 ;
      RECT 35.334 14.758 35.386 14.794 ;
      RECT 35.334 15.958 35.386 15.994 ;
      RECT 35.334 17.158 35.386 17.194 ;
      RECT 35.334 18.358 35.386 18.394 ;
      RECT 35.334 19.558 35.386 19.594 ;
      RECT 35.334 20.758 35.386 20.794 ;
      RECT 35.334 21.958 35.386 21.994 ;
      RECT 35.334 23.158 35.386 23.194 ;
      RECT 35.334 24.358 35.386 24.394 ;
      RECT 35.334 25.558 35.386 25.594 ;
      RECT 35.334 26.758 35.386 26.794 ;
      RECT 35.334 27.958 35.386 27.994 ;
      RECT 35.334 29.158 35.386 29.194 ;
      RECT 35.334 30.358 35.386 30.394 ;
      RECT 35.334 31.558 35.386 31.594 ;
      RECT 35.334 33.342 35.386 33.378 ;
      RECT 35.334 33.582 35.386 33.618 ;
      RECT 35.334 37.902 35.386 37.938 ;
      RECT 35.334 38.142 35.386 38.178 ;
      RECT 35.334 40.678 35.386 40.714 ;
      RECT 35.334 41.878 35.386 41.914 ;
      RECT 35.334 43.078 35.386 43.114 ;
      RECT 35.334 44.278 35.386 44.314 ;
      RECT 35.334 45.478 35.386 45.514 ;
      RECT 35.334 46.678 35.386 46.714 ;
      RECT 35.334 47.878 35.386 47.914 ;
      RECT 35.334 49.078 35.386 49.114 ;
      RECT 35.334 50.278 35.386 50.314 ;
      RECT 35.334 51.478 35.386 51.514 ;
      RECT 35.334 52.678 35.386 52.714 ;
      RECT 35.334 53.878 35.386 53.914 ;
      RECT 35.334 55.078 35.386 55.114 ;
      RECT 35.334 56.278 35.386 56.314 ;
      RECT 35.334 57.478 35.386 57.514 ;
      RECT 35.334 58.678 35.386 58.714 ;
      RECT 35.334 59.878 35.386 59.914 ;
      RECT 35.334 61.078 35.386 61.114 ;
      RECT 35.334 62.278 35.386 62.314 ;
      RECT 35.334 63.478 35.386 63.514 ;
      RECT 35.334 64.678 35.386 64.714 ;
      RECT 35.334 65.878 35.386 65.914 ;
      RECT 35.334 67.078 35.386 67.114 ;
      RECT 35.334 68.278 35.386 68.314 ;
      RECT 35.334 69.478 35.386 69.514 ;
      RECT 35.334 70.678 35.386 70.714 ;
      RECT 35.334 71.878 35.386 71.914 ;
      RECT 35.414 0.806 35.466 0.842 ;
      RECT 35.414 2.006 35.466 2.042 ;
      RECT 35.414 3.206 35.466 3.242 ;
      RECT 35.414 4.406 35.466 4.442 ;
      RECT 35.414 5.606 35.466 5.642 ;
      RECT 35.414 6.806 35.466 6.842 ;
      RECT 35.414 8.006 35.466 8.042 ;
      RECT 35.414 9.206 35.466 9.242 ;
      RECT 35.414 10.406 35.466 10.442 ;
      RECT 35.414 11.606 35.466 11.642 ;
      RECT 35.414 12.806 35.466 12.842 ;
      RECT 35.414 14.006 35.466 14.042 ;
      RECT 35.414 15.206 35.466 15.242 ;
      RECT 35.414 16.406 35.466 16.442 ;
      RECT 35.414 17.606 35.466 17.642 ;
      RECT 35.414 18.806 35.466 18.842 ;
      RECT 35.414 20.006 35.466 20.042 ;
      RECT 35.414 21.206 35.466 21.242 ;
      RECT 35.414 22.406 35.466 22.442 ;
      RECT 35.414 23.606 35.466 23.642 ;
      RECT 35.414 24.806 35.466 24.842 ;
      RECT 35.414 26.006 35.466 26.042 ;
      RECT 35.414 27.206 35.466 27.242 ;
      RECT 35.414 28.406 35.466 28.442 ;
      RECT 35.414 29.606 35.466 29.642 ;
      RECT 35.414 30.806 35.466 30.842 ;
      RECT 35.414 32.622 35.466 32.658 ;
      RECT 35.414 32.862 35.466 32.898 ;
      RECT 35.414 38.622 35.466 38.658 ;
      RECT 35.414 38.862 35.466 38.898 ;
      RECT 35.414 39.926 35.466 39.962 ;
      RECT 35.414 41.126 35.466 41.162 ;
      RECT 35.414 42.326 35.466 42.362 ;
      RECT 35.414 43.526 35.466 43.562 ;
      RECT 35.414 44.726 35.466 44.762 ;
      RECT 35.414 45.926 35.466 45.962 ;
      RECT 35.414 47.126 35.466 47.162 ;
      RECT 35.414 48.326 35.466 48.362 ;
      RECT 35.414 49.526 35.466 49.562 ;
      RECT 35.414 50.726 35.466 50.762 ;
      RECT 35.414 51.926 35.466 51.962 ;
      RECT 35.414 53.126 35.466 53.162 ;
      RECT 35.414 54.326 35.466 54.362 ;
      RECT 35.414 55.526 35.466 55.562 ;
      RECT 35.414 56.726 35.466 56.762 ;
      RECT 35.414 57.926 35.466 57.962 ;
      RECT 35.414 59.126 35.466 59.162 ;
      RECT 35.414 60.326 35.466 60.362 ;
      RECT 35.414 61.526 35.466 61.562 ;
      RECT 35.414 62.726 35.466 62.762 ;
      RECT 35.414 63.926 35.466 63.962 ;
      RECT 35.414 65.126 35.466 65.162 ;
      RECT 35.414 66.326 35.466 66.362 ;
      RECT 35.414 67.526 35.466 67.562 ;
      RECT 35.414 68.726 35.466 68.762 ;
      RECT 35.414 69.926 35.466 69.962 ;
      RECT 35.414 71.126 35.466 71.162 ;
      RECT 35.494 1.558 35.546 1.594 ;
      RECT 35.494 2.758 35.546 2.794 ;
      RECT 35.494 3.958 35.546 3.994 ;
      RECT 35.494 5.158 35.546 5.194 ;
      RECT 35.494 6.358 35.546 6.394 ;
      RECT 35.494 7.558 35.546 7.594 ;
      RECT 35.494 8.758 35.546 8.794 ;
      RECT 35.494 9.958 35.546 9.994 ;
      RECT 35.494 11.158 35.546 11.194 ;
      RECT 35.494 12.358 35.546 12.394 ;
      RECT 35.494 13.558 35.546 13.594 ;
      RECT 35.494 14.758 35.546 14.794 ;
      RECT 35.494 15.958 35.546 15.994 ;
      RECT 35.494 17.158 35.546 17.194 ;
      RECT 35.494 18.358 35.546 18.394 ;
      RECT 35.494 19.558 35.546 19.594 ;
      RECT 35.494 20.758 35.546 20.794 ;
      RECT 35.494 21.958 35.546 21.994 ;
      RECT 35.494 23.158 35.546 23.194 ;
      RECT 35.494 24.358 35.546 24.394 ;
      RECT 35.494 25.558 35.546 25.594 ;
      RECT 35.494 26.758 35.546 26.794 ;
      RECT 35.494 27.958 35.546 27.994 ;
      RECT 35.494 29.158 35.546 29.194 ;
      RECT 35.494 30.358 35.546 30.394 ;
      RECT 35.494 31.558 35.546 31.594 ;
      RECT 35.494 33.342 35.546 33.378 ;
      RECT 35.494 33.582 35.546 33.618 ;
      RECT 35.494 37.902 35.546 37.938 ;
      RECT 35.494 38.142 35.546 38.178 ;
      RECT 35.494 40.678 35.546 40.714 ;
      RECT 35.494 41.878 35.546 41.914 ;
      RECT 35.494 43.078 35.546 43.114 ;
      RECT 35.494 44.278 35.546 44.314 ;
      RECT 35.494 45.478 35.546 45.514 ;
      RECT 35.494 46.678 35.546 46.714 ;
      RECT 35.494 47.878 35.546 47.914 ;
      RECT 35.494 49.078 35.546 49.114 ;
      RECT 35.494 50.278 35.546 50.314 ;
      RECT 35.494 51.478 35.546 51.514 ;
      RECT 35.494 52.678 35.546 52.714 ;
      RECT 35.494 53.878 35.546 53.914 ;
      RECT 35.494 55.078 35.546 55.114 ;
      RECT 35.494 56.278 35.546 56.314 ;
      RECT 35.494 57.478 35.546 57.514 ;
      RECT 35.494 58.678 35.546 58.714 ;
      RECT 35.494 59.878 35.546 59.914 ;
      RECT 35.494 61.078 35.546 61.114 ;
      RECT 35.494 62.278 35.546 62.314 ;
      RECT 35.494 63.478 35.546 63.514 ;
      RECT 35.494 64.678 35.546 64.714 ;
      RECT 35.494 65.878 35.546 65.914 ;
      RECT 35.494 67.078 35.546 67.114 ;
      RECT 35.494 68.278 35.546 68.314 ;
      RECT 35.494 69.478 35.546 69.514 ;
      RECT 35.494 70.678 35.546 70.714 ;
      RECT 35.494 71.878 35.546 71.914 ;
      RECT 35.574 0.281 35.626 0.317 ;
      RECT 35.574 72.403 35.626 72.439 ;
      RECT 35.946 0.582 35.994 0.618 ;
      RECT 35.946 0.882 35.994 0.918 ;
      RECT 35.946 1.182 35.994 1.218 ;
      RECT 35.946 1.482 35.994 1.518 ;
      RECT 35.946 1.782 35.994 1.818 ;
      RECT 35.946 2.082 35.994 2.118 ;
      RECT 35.946 2.382 35.994 2.418 ;
      RECT 35.946 2.682 35.994 2.718 ;
      RECT 35.946 2.982 35.994 3.018 ;
      RECT 35.946 3.282 35.994 3.318 ;
      RECT 35.946 3.582 35.994 3.618 ;
      RECT 35.946 3.882 35.994 3.918 ;
      RECT 35.946 4.182 35.994 4.218 ;
      RECT 35.946 4.482 35.994 4.518 ;
      RECT 35.946 4.782 35.994 4.818 ;
      RECT 35.946 5.082 35.994 5.118 ;
      RECT 35.946 5.382 35.994 5.418 ;
      RECT 35.946 5.682 35.994 5.718 ;
      RECT 35.946 5.982 35.994 6.018 ;
      RECT 35.946 6.282 35.994 6.318 ;
      RECT 35.946 6.582 35.994 6.618 ;
      RECT 35.946 6.882 35.994 6.918 ;
      RECT 35.946 7.182 35.994 7.218 ;
      RECT 35.946 7.482 35.994 7.518 ;
      RECT 35.946 7.782 35.994 7.818 ;
      RECT 35.946 8.082 35.994 8.118 ;
      RECT 35.946 8.382 35.994 8.418 ;
      RECT 35.946 8.682 35.994 8.718 ;
      RECT 35.946 8.982 35.994 9.018 ;
      RECT 35.946 9.282 35.994 9.318 ;
      RECT 35.946 9.582 35.994 9.618 ;
      RECT 35.946 9.882 35.994 9.918 ;
      RECT 35.946 10.182 35.994 10.218 ;
      RECT 35.946 10.482 35.994 10.518 ;
      RECT 35.946 10.782 35.994 10.818 ;
      RECT 35.946 11.082 35.994 11.118 ;
      RECT 35.946 11.382 35.994 11.418 ;
      RECT 35.946 11.682 35.994 11.718 ;
      RECT 35.946 11.982 35.994 12.018 ;
      RECT 35.946 12.282 35.994 12.318 ;
      RECT 35.946 12.582 35.994 12.618 ;
      RECT 35.946 12.882 35.994 12.918 ;
      RECT 35.946 13.182 35.994 13.218 ;
      RECT 35.946 13.482 35.994 13.518 ;
      RECT 35.946 13.782 35.994 13.818 ;
      RECT 35.946 14.082 35.994 14.118 ;
      RECT 35.946 14.382 35.994 14.418 ;
      RECT 35.946 14.682 35.994 14.718 ;
      RECT 35.946 14.982 35.994 15.018 ;
      RECT 35.946 15.282 35.994 15.318 ;
      RECT 35.946 15.582 35.994 15.618 ;
      RECT 35.946 15.882 35.994 15.918 ;
      RECT 35.946 16.182 35.994 16.218 ;
      RECT 35.946 16.482 35.994 16.518 ;
      RECT 35.946 16.782 35.994 16.818 ;
      RECT 35.946 17.082 35.994 17.118 ;
      RECT 35.946 17.382 35.994 17.418 ;
      RECT 35.946 17.682 35.994 17.718 ;
      RECT 35.946 17.982 35.994 18.018 ;
      RECT 35.946 18.282 35.994 18.318 ;
      RECT 35.946 18.582 35.994 18.618 ;
      RECT 35.946 18.882 35.994 18.918 ;
      RECT 35.946 19.182 35.994 19.218 ;
      RECT 35.946 19.482 35.994 19.518 ;
      RECT 35.946 19.782 35.994 19.818 ;
      RECT 35.946 20.082 35.994 20.118 ;
      RECT 35.946 20.382 35.994 20.418 ;
      RECT 35.946 20.682 35.994 20.718 ;
      RECT 35.946 20.982 35.994 21.018 ;
      RECT 35.946 21.282 35.994 21.318 ;
      RECT 35.946 21.582 35.994 21.618 ;
      RECT 35.946 21.882 35.994 21.918 ;
      RECT 35.946 22.182 35.994 22.218 ;
      RECT 35.946 22.482 35.994 22.518 ;
      RECT 35.946 22.782 35.994 22.818 ;
      RECT 35.946 23.082 35.994 23.118 ;
      RECT 35.946 23.382 35.994 23.418 ;
      RECT 35.946 23.682 35.994 23.718 ;
      RECT 35.946 23.982 35.994 24.018 ;
      RECT 35.946 24.282 35.994 24.318 ;
      RECT 35.946 24.582 35.994 24.618 ;
      RECT 35.946 24.882 35.994 24.918 ;
      RECT 35.946 25.182 35.994 25.218 ;
      RECT 35.946 25.482 35.994 25.518 ;
      RECT 35.946 25.782 35.994 25.818 ;
      RECT 35.946 26.082 35.994 26.118 ;
      RECT 35.946 26.382 35.994 26.418 ;
      RECT 35.946 26.682 35.994 26.718 ;
      RECT 35.946 26.982 35.994 27.018 ;
      RECT 35.946 27.282 35.994 27.318 ;
      RECT 35.946 27.582 35.994 27.618 ;
      RECT 35.946 27.882 35.994 27.918 ;
      RECT 35.946 28.182 35.994 28.218 ;
      RECT 35.946 28.482 35.994 28.518 ;
      RECT 35.946 28.782 35.994 28.818 ;
      RECT 35.946 29.082 35.994 29.118 ;
      RECT 35.946 29.382 35.994 29.418 ;
      RECT 35.946 29.682 35.994 29.718 ;
      RECT 35.946 29.982 35.994 30.018 ;
      RECT 35.946 30.282 35.994 30.318 ;
      RECT 35.946 30.582 35.994 30.618 ;
      RECT 35.946 30.882 35.994 30.918 ;
      RECT 35.946 31.182 35.994 31.218 ;
      RECT 35.946 31.482 35.994 31.518 ;
      RECT 35.946 31.782 35.994 31.818 ;
      RECT 35.946 32.3235 35.994 32.3595 ;
      RECT 35.946 32.622 35.994 32.658 ;
      RECT 35.946 32.9205 35.994 32.9565 ;
      RECT 35.946 33.222 35.994 33.258 ;
      RECT 35.946 33.5235 35.994 33.5595 ;
      RECT 35.946 33.822 35.994 33.858 ;
      RECT 35.946 34.1205 35.994 34.1565 ;
      RECT 35.946 34.422 35.994 34.458 ;
      RECT 35.946 34.7235 35.994 34.7595 ;
      RECT 35.946 35.262 35.994 35.298 ;
      RECT 35.946 35.862 35.994 35.898 ;
      RECT 35.946 36.1635 35.994 36.1995 ;
      RECT 35.946 36.462 35.994 36.498 ;
      RECT 35.946 36.7605 35.994 36.7965 ;
      RECT 35.946 37.062 35.994 37.098 ;
      RECT 35.946 37.3635 35.994 37.3995 ;
      RECT 35.946 37.662 35.994 37.698 ;
      RECT 35.946 37.9605 35.994 37.9965 ;
      RECT 35.946 38.262 35.994 38.298 ;
      RECT 35.946 38.5635 35.994 38.5995 ;
      RECT 35.946 38.862 35.994 38.898 ;
      RECT 35.946 39.1605 35.994 39.1965 ;
      RECT 35.946 39.702 35.994 39.738 ;
      RECT 35.946 40.002 35.994 40.038 ;
      RECT 35.946 40.302 35.994 40.338 ;
      RECT 35.946 40.602 35.994 40.638 ;
      RECT 35.946 40.902 35.994 40.938 ;
      RECT 35.946 41.202 35.994 41.238 ;
      RECT 35.946 41.502 35.994 41.538 ;
      RECT 35.946 41.802 35.994 41.838 ;
      RECT 35.946 42.102 35.994 42.138 ;
      RECT 35.946 42.402 35.994 42.438 ;
      RECT 35.946 42.702 35.994 42.738 ;
      RECT 35.946 43.002 35.994 43.038 ;
      RECT 35.946 43.302 35.994 43.338 ;
      RECT 35.946 43.602 35.994 43.638 ;
      RECT 35.946 43.902 35.994 43.938 ;
      RECT 35.946 44.202 35.994 44.238 ;
      RECT 35.946 44.502 35.994 44.538 ;
      RECT 35.946 44.802 35.994 44.838 ;
      RECT 35.946 45.102 35.994 45.138 ;
      RECT 35.946 45.402 35.994 45.438 ;
      RECT 35.946 45.702 35.994 45.738 ;
      RECT 35.946 46.002 35.994 46.038 ;
      RECT 35.946 46.302 35.994 46.338 ;
      RECT 35.946 46.602 35.994 46.638 ;
      RECT 35.946 46.902 35.994 46.938 ;
      RECT 35.946 47.202 35.994 47.238 ;
      RECT 35.946 47.502 35.994 47.538 ;
      RECT 35.946 47.802 35.994 47.838 ;
      RECT 35.946 48.102 35.994 48.138 ;
      RECT 35.946 48.402 35.994 48.438 ;
      RECT 35.946 48.702 35.994 48.738 ;
      RECT 35.946 49.002 35.994 49.038 ;
      RECT 35.946 49.302 35.994 49.338 ;
      RECT 35.946 49.602 35.994 49.638 ;
      RECT 35.946 49.902 35.994 49.938 ;
      RECT 35.946 50.202 35.994 50.238 ;
      RECT 35.946 50.502 35.994 50.538 ;
      RECT 35.946 50.802 35.994 50.838 ;
      RECT 35.946 51.102 35.994 51.138 ;
      RECT 35.946 51.402 35.994 51.438 ;
      RECT 35.946 51.702 35.994 51.738 ;
      RECT 35.946 52.002 35.994 52.038 ;
      RECT 35.946 52.302 35.994 52.338 ;
      RECT 35.946 52.602 35.994 52.638 ;
      RECT 35.946 52.902 35.994 52.938 ;
      RECT 35.946 53.202 35.994 53.238 ;
      RECT 35.946 53.502 35.994 53.538 ;
      RECT 35.946 53.802 35.994 53.838 ;
      RECT 35.946 54.102 35.994 54.138 ;
      RECT 35.946 54.402 35.994 54.438 ;
      RECT 35.946 54.702 35.994 54.738 ;
      RECT 35.946 55.002 35.994 55.038 ;
      RECT 35.946 55.302 35.994 55.338 ;
      RECT 35.946 55.602 35.994 55.638 ;
      RECT 35.946 55.902 35.994 55.938 ;
      RECT 35.946 56.202 35.994 56.238 ;
      RECT 35.946 56.502 35.994 56.538 ;
      RECT 35.946 56.802 35.994 56.838 ;
      RECT 35.946 57.102 35.994 57.138 ;
      RECT 35.946 57.402 35.994 57.438 ;
      RECT 35.946 57.702 35.994 57.738 ;
      RECT 35.946 58.002 35.994 58.038 ;
      RECT 35.946 58.302 35.994 58.338 ;
      RECT 35.946 58.602 35.994 58.638 ;
      RECT 35.946 58.902 35.994 58.938 ;
      RECT 35.946 59.202 35.994 59.238 ;
      RECT 35.946 59.502 35.994 59.538 ;
      RECT 35.946 59.802 35.994 59.838 ;
      RECT 35.946 60.102 35.994 60.138 ;
      RECT 35.946 60.402 35.994 60.438 ;
      RECT 35.946 60.702 35.994 60.738 ;
      RECT 35.946 61.002 35.994 61.038 ;
      RECT 35.946 61.302 35.994 61.338 ;
      RECT 35.946 61.602 35.994 61.638 ;
      RECT 35.946 61.902 35.994 61.938 ;
      RECT 35.946 62.202 35.994 62.238 ;
      RECT 35.946 62.502 35.994 62.538 ;
      RECT 35.946 62.802 35.994 62.838 ;
      RECT 35.946 63.102 35.994 63.138 ;
      RECT 35.946 63.402 35.994 63.438 ;
      RECT 35.946 63.702 35.994 63.738 ;
      RECT 35.946 64.002 35.994 64.038 ;
      RECT 35.946 64.302 35.994 64.338 ;
      RECT 35.946 64.602 35.994 64.638 ;
      RECT 35.946 64.902 35.994 64.938 ;
      RECT 35.946 65.202 35.994 65.238 ;
      RECT 35.946 65.502 35.994 65.538 ;
      RECT 35.946 65.802 35.994 65.838 ;
      RECT 35.946 66.102 35.994 66.138 ;
      RECT 35.946 66.402 35.994 66.438 ;
      RECT 35.946 66.702 35.994 66.738 ;
      RECT 35.946 67.002 35.994 67.038 ;
      RECT 35.946 67.302 35.994 67.338 ;
      RECT 35.946 67.602 35.994 67.638 ;
      RECT 35.946 67.902 35.994 67.938 ;
      RECT 35.946 68.202 35.994 68.238 ;
      RECT 35.946 68.502 35.994 68.538 ;
      RECT 35.946 68.802 35.994 68.838 ;
      RECT 35.946 69.102 35.994 69.138 ;
      RECT 35.946 69.402 35.994 69.438 ;
      RECT 35.946 69.702 35.994 69.738 ;
      RECT 35.946 70.002 35.994 70.038 ;
      RECT 35.946 70.302 35.994 70.338 ;
      RECT 35.946 70.602 35.994 70.638 ;
      RECT 35.946 70.902 35.994 70.938 ;
      RECT 35.946 71.202 35.994 71.238 ;
      RECT 35.946 71.502 35.994 71.538 ;
      RECT 35.946 71.802 35.994 71.838 ;
      RECT 35.946 72.102 35.994 72.138 ;
    LAYER m5 ;
      RECT 0.012 72.1905 36.288 72.72 ;
      RECT 15.75 72.16 15.914 72.1905 ;
      RECT 20.086 72.16 20.25 72.1905 ;
      RECT 17.076 72.14 17.304 72.1905 ;
      RECT 17.424 72.14 17.644 72.1905 ;
      RECT 19.076 39.76 19.41 72.1905 ;
      RECT 18.228 39.74 18.316 72.1905 ;
      RECT 17.216 39.74 17.304 72.14 ;
      RECT 17.076 39.7 17.096 72.14 ;
      RECT 17.492 39.7 17.644 72.14 ;
      RECT 17.424 39.38 17.644 39.7 ;
      RECT 16.894 39.2325 16.924 72.1905 ;
      RECT 17.284 39.34 17.304 39.74 ;
      RECT 17.492 38.97 17.644 39.38 ;
      RECT 0.666 72.16 1.334 72.1905 ;
      RECT 1.466 72.16 2.134 72.1905 ;
      RECT 2.266 72.16 2.934 72.1905 ;
      RECT 3.066 72.16 3.734 72.1905 ;
      RECT 3.866 72.16 4.534 72.1905 ;
      RECT 4.666 72.16 5.334 72.1905 ;
      RECT 5.466 72.16 6.134 72.1905 ;
      RECT 6.266 72.16 6.934 72.1905 ;
      RECT 7.066 72.16 7.734 72.1905 ;
      RECT 7.866 72.16 8.534 72.1905 ;
      RECT 8.666 72.16 9.334 72.1905 ;
      RECT 9.466 72.16 10.134 72.1905 ;
      RECT 10.266 72.16 10.934 72.1905 ;
      RECT 11.066 72.16 11.734 72.1905 ;
      RECT 11.866 72.16 12.534 72.1905 ;
      RECT 12.666 72.16 13.334 72.1905 ;
      RECT 22.866 72.16 23.534 72.1905 ;
      RECT 23.666 72.16 24.334 72.1905 ;
      RECT 24.466 72.16 25.134 72.1905 ;
      RECT 25.266 72.16 25.934 72.1905 ;
      RECT 26.066 72.16 26.734 72.1905 ;
      RECT 27.666 72.16 28.334 72.1905 ;
      RECT 28.466 72.16 29.134 72.1905 ;
      RECT 29.266 72.16 29.934 72.1905 ;
      RECT 30.066 72.16 30.734 72.1905 ;
      RECT 30.866 72.16 31.534 72.1905 ;
      RECT 31.666 72.16 32.334 72.1905 ;
      RECT 32.466 72.16 33.134 72.1905 ;
      RECT 33.266 72.16 33.934 72.1905 ;
      RECT 34.066 72.16 34.734 72.1905 ;
      RECT 34.866 72.16 35.534 72.1905 ;
      RECT 19.076 39.72 19.27 39.76 ;
      RECT 20.382 38.159 20.43 72.1905 ;
      RECT 20.562 38.159 20.59 72.1905 ;
      RECT 17.956 37.85 18.108 72.1905 ;
      RECT 17.076 38.85 17.164 39.7 ;
      RECT 17.284 38.85 17.372 39.34 ;
      RECT 17.56 38.85 17.644 38.97 ;
      RECT 18.436 37.85 18.524 72.1905 ;
      RECT 17.492 36.81 17.508 36.93 ;
      RECT 17.076 35.81 17.096 38.85 ;
      RECT 17.284 35.81 17.304 38.85 ;
      RECT 17.492 35.81 17.576 36.81 ;
      RECT 17.076 35.3 17.164 35.81 ;
      RECT 17.492 35.3 17.644 35.81 ;
      RECT 17.956 35.18 18.108 36.81 ;
      RECT 17.284 35.18 17.372 35.81 ;
      RECT 17.076 35.18 17.096 35.3 ;
      RECT 17.56 35.18 17.644 35.3 ;
      RECT 17.956 34.18 17.972 35.18 ;
      RECT 17.56 34.14 17.576 35.18 ;
      RECT 17.076 33.26 17.096 34.14 ;
      RECT 17.56 33.26 17.644 34.14 ;
      RECT 17.492 33.18 17.644 33.26 ;
      RECT 0.666 38.6095 0.934 72.16 ;
      RECT 1.466 38.6095 1.734 72.16 ;
      RECT 2.266 38.6095 2.534 72.16 ;
      RECT 3.066 38.6095 3.334 72.16 ;
      RECT 3.866 38.6095 4.134 72.16 ;
      RECT 4.666 38.6095 4.934 72.16 ;
      RECT 5.466 38.6095 5.734 72.16 ;
      RECT 6.266 38.6095 6.534 72.16 ;
      RECT 7.066 38.6095 7.334 72.16 ;
      RECT 7.866 38.6095 8.134 72.16 ;
      RECT 8.666 38.6095 8.934 72.16 ;
      RECT 9.466 38.6095 9.734 72.16 ;
      RECT 10.266 38.6095 10.534 72.16 ;
      RECT 11.066 38.6095 11.334 72.16 ;
      RECT 11.866 38.6095 12.134 72.16 ;
      RECT 12.666 38.6095 12.934 72.16 ;
      RECT 22.866 38.6095 23.134 72.16 ;
      RECT 23.666 38.6095 23.934 72.16 ;
      RECT 24.466 38.6095 24.734 72.16 ;
      RECT 25.266 38.6095 25.534 72.16 ;
      RECT 26.066 38.6095 26.334 72.16 ;
      RECT 26.866 38.6095 27.134 72.16 ;
      RECT 27.666 38.6095 27.934 72.16 ;
      RECT 28.466 38.6095 28.734 72.16 ;
      RECT 29.266 38.6095 29.534 72.16 ;
      RECT 30.066 38.6095 30.334 72.16 ;
      RECT 30.866 38.6095 31.134 72.16 ;
      RECT 31.666 38.6095 31.934 72.16 ;
      RECT 32.466 38.6095 32.734 72.16 ;
      RECT 33.266 38.6095 33.534 72.16 ;
      RECT 34.066 38.6095 34.334 72.16 ;
      RECT 34.866 38.6095 35.134 72.16 ;
      RECT 15.41 38.159 15.438 72.1905 ;
      RECT 15.57 38.159 15.618 72.1905 ;
      RECT 18.296 35.18 18.316 39.74 ;
      RECT 18.504 36.81 18.524 37.85 ;
      RECT 18.092 33.14 18.108 35.18 ;
      RECT 20.382 32.8995 20.59 38.159 ;
      RECT 17.492 32.14 17.508 33.18 ;
      RECT 17.076 31.82 17.164 33.26 ;
      RECT 17.424 31.82 17.644 32.14 ;
      RECT 19.076 31.8 19.188 39.72 ;
      RECT 18.296 31.78 18.316 32.14 ;
      RECT 17.284 31.78 17.304 33.14 ;
      RECT 0.746 32.9105 0.934 38.6095 ;
      RECT 1.546 32.9105 1.734 38.6095 ;
      RECT 2.346 32.9105 2.534 38.6095 ;
      RECT 3.146 32.9105 3.334 38.6095 ;
      RECT 3.946 32.9105 4.134 38.6095 ;
      RECT 4.746 32.9105 4.934 38.6095 ;
      RECT 5.546 32.9105 5.734 38.6095 ;
      RECT 6.346 32.9105 6.534 38.6095 ;
      RECT 7.146 32.9105 7.334 38.6095 ;
      RECT 7.946 32.9105 8.134 38.6095 ;
      RECT 8.746 32.9105 8.934 38.6095 ;
      RECT 9.546 32.9105 9.734 38.6095 ;
      RECT 10.346 32.9105 10.534 38.6095 ;
      RECT 11.146 32.9105 11.334 38.6095 ;
      RECT 11.946 32.9105 12.134 38.6095 ;
      RECT 12.746 32.9105 12.934 38.6095 ;
      RECT 15.41 32.8995 15.618 38.159 ;
      RECT 19.39 31.76 19.41 39.76 ;
      RECT 19.076 31.76 19.27 31.8 ;
      RECT 22.946 32.9105 23.134 38.6095 ;
      RECT 23.746 32.9105 23.934 38.6095 ;
      RECT 24.546 32.9105 24.734 38.6095 ;
      RECT 25.346 32.9105 25.534 38.6095 ;
      RECT 26.146 32.9105 26.334 38.6095 ;
      RECT 26.946 32.9105 27.134 38.6095 ;
      RECT 27.746 32.9105 27.934 38.6095 ;
      RECT 28.546 32.9105 28.734 38.6095 ;
      RECT 29.346 32.9105 29.534 38.6095 ;
      RECT 30.146 32.9105 30.334 38.6095 ;
      RECT 30.946 32.9105 31.134 38.6095 ;
      RECT 31.746 32.9105 31.934 38.6095 ;
      RECT 32.546 32.9105 32.734 38.6095 ;
      RECT 33.346 32.9105 33.534 38.6095 ;
      RECT 34.146 32.9105 34.334 38.6095 ;
      RECT 34.946 32.9105 35.134 38.6095 ;
      RECT 26.866 72.16 27.534 72.1905 ;
      RECT 31.666 0.56 31.934 32.9105 ;
      RECT 32.066 0.56 32.334 72.16 ;
      RECT 32.866 0.56 33.134 72.16 ;
      RECT 33.666 0.56 33.934 72.16 ;
      RECT 34.466 0.56 34.734 72.16 ;
      RECT 35.266 0.56 35.534 72.16 ;
      RECT 32.466 0.56 32.734 32.9105 ;
      RECT 33.266 0.56 33.534 32.9105 ;
      RECT 34.066 0.56 34.334 32.9105 ;
      RECT 34.866 0.56 35.134 32.9105 ;
      RECT 27.266 0.56 27.534 72.16 ;
      RECT 28.066 0.56 28.334 72.16 ;
      RECT 28.866 0.56 29.134 72.16 ;
      RECT 29.666 0.56 29.934 72.16 ;
      RECT 30.466 0.56 30.734 72.16 ;
      RECT 31.266 0.56 31.534 72.16 ;
      RECT 27.666 0.56 27.934 32.9105 ;
      RECT 28.466 0.56 28.734 32.9105 ;
      RECT 29.266 0.56 29.534 32.9105 ;
      RECT 30.066 0.56 30.334 32.9105 ;
      RECT 30.866 0.56 31.134 32.9105 ;
      RECT 24.866 0.56 25.134 72.16 ;
      RECT 25.666 0.56 25.934 72.16 ;
      RECT 26.466 0.56 26.734 72.16 ;
      RECT 25.266 0.56 25.534 32.9105 ;
      RECT 26.066 0.56 26.334 32.9105 ;
      RECT 26.866 0.56 27.134 32.9105 ;
      RECT 23.266 0.56 23.534 72.16 ;
      RECT 24.066 0.56 24.334 72.16 ;
      RECT 22.866 0.56 23.134 32.9105 ;
      RECT 23.666 0.56 23.934 32.9105 ;
      RECT 24.466 0.56 24.734 32.9105 ;
      RECT 20.166 0.56 20.25 72.16 ;
      RECT 9.066 0.56 9.334 72.16 ;
      RECT 17.076 0.58 17.096 31.82 ;
      RECT 17.492 0.58 17.644 31.82 ;
      RECT 17.216 0.58 17.304 31.78 ;
      RECT 15.75 0.56 15.834 72.16 ;
      RECT 9.866 0.56 10.134 72.16 ;
      RECT 10.666 0.56 10.934 72.16 ;
      RECT 11.466 0.56 11.734 72.16 ;
      RECT 12.266 0.56 12.534 72.16 ;
      RECT 13.066 0.56 13.334 72.16 ;
      RECT 9.466 0.56 9.734 32.9105 ;
      RECT 10.266 0.56 10.534 32.9105 ;
      RECT 11.066 0.56 11.334 32.9105 ;
      RECT 11.866 0.56 12.134 32.9105 ;
      RECT 12.666 0.56 12.934 32.9105 ;
      RECT 6.666 0.56 6.934 72.16 ;
      RECT 7.466 0.56 7.734 72.16 ;
      RECT 8.266 0.56 8.534 72.16 ;
      RECT 7.066 0.56 7.334 32.9105 ;
      RECT 7.866 0.56 8.134 32.9105 ;
      RECT 8.666 0.56 8.934 32.9105 ;
      RECT 5.066 0.56 5.334 72.16 ;
      RECT 5.866 0.56 6.134 72.16 ;
      RECT 4.666 0.56 4.934 32.9105 ;
      RECT 5.466 0.56 5.734 32.9105 ;
      RECT 6.266 0.56 6.534 32.9105 ;
      RECT 1.066 0.56 1.334 72.16 ;
      RECT 1.866 0.56 2.134 72.16 ;
      RECT 2.666 0.56 2.934 72.16 ;
      RECT 3.466 0.56 3.734 72.16 ;
      RECT 4.266 0.56 4.534 72.16 ;
      RECT 0.666 0.56 0.934 32.9105 ;
      RECT 1.466 0.56 1.734 32.9105 ;
      RECT 2.266 0.56 2.534 32.9105 ;
      RECT 3.066 0.56 3.334 32.9105 ;
      RECT 3.866 0.56 4.134 32.9105 ;
      RECT 0.012 0 36.288 0.5295 ;
      RECT 26.866 0.5295 27.534 0.56 ;
      RECT 31.666 0.5295 32.334 0.56 ;
      RECT 35.666 0.5295 36.288 72.1905 ;
      RECT 32.466 0.5295 33.134 0.56 ;
      RECT 33.266 0.5295 33.934 0.56 ;
      RECT 34.066 0.5295 34.734 0.56 ;
      RECT 34.866 0.5295 35.534 0.56 ;
      RECT 27.666 0.5295 28.334 0.56 ;
      RECT 28.466 0.5295 29.134 0.56 ;
      RECT 29.266 0.5295 29.934 0.56 ;
      RECT 30.066 0.5295 30.734 0.56 ;
      RECT 30.866 0.5295 31.534 0.56 ;
      RECT 21.99 0.5295 22.734 72.1905 ;
      RECT 24.466 0.5295 25.134 0.56 ;
      RECT 25.266 0.5295 25.934 0.56 ;
      RECT 26.066 0.5295 26.734 0.56 ;
      RECT 22.866 0.5295 23.534 0.56 ;
      RECT 23.666 0.5295 24.334 0.56 ;
      RECT 18.776 0.5295 18.824 72.1905 ;
      RECT 19.542 0.5295 19.642 72.1905 ;
      RECT 19.774 0.5295 19.874 72.1905 ;
      RECT 20.722 0.5295 20.974 72.1905 ;
      RECT 21.108 0.5295 21.456 72.1905 ;
      RECT 21.59 0.5295 21.61 72.1905 ;
      RECT 21.744 0.5295 21.856 72.1905 ;
      RECT 18.436 0.5295 18.524 36.81 ;
      RECT 20.382 0.5295 20.43 32.8995 ;
      RECT 20.562 0.5295 20.59 32.8995 ;
      RECT 18.228 0.5295 18.316 31.78 ;
      RECT 19.076 0.5295 19.41 31.76 ;
      RECT 20.086 0.5295 20.25 0.56 ;
      RECT 8.666 0.5295 9.334 0.56 ;
      RECT 13.466 0.5295 14.01 72.1905 ;
      RECT 15.75 0.5295 15.914 0.56 ;
      RECT 16.126 0.5295 16.226 72.1905 ;
      RECT 16.358 0.5295 16.458 72.1905 ;
      RECT 16.59 0.5295 16.76 72.1905 ;
      RECT 17.776 0.5295 17.804 72.1905 ;
      RECT 17.956 0.5295 18.108 33.14 ;
      RECT 16.894 0.5295 16.924 32.313 ;
      RECT 17.076 0.5295 17.304 0.58 ;
      RECT 17.424 0.5295 17.644 0.58 ;
      RECT 14.144 0.5295 14.256 72.1905 ;
      RECT 14.39 0.5295 14.41 72.1905 ;
      RECT 14.544 0.5295 14.892 72.1905 ;
      RECT 15.026 0.5295 15.278 72.1905 ;
      RECT 15.41 0.5295 15.438 32.8995 ;
      RECT 15.57 0.5295 15.618 32.8995 ;
      RECT 9.466 0.5295 10.134 0.56 ;
      RECT 10.266 0.5295 10.934 0.56 ;
      RECT 11.066 0.5295 11.734 0.56 ;
      RECT 11.866 0.5295 12.534 0.56 ;
      RECT 12.666 0.5295 13.334 0.56 ;
      RECT 6.266 0.5295 6.934 0.56 ;
      RECT 7.066 0.5295 7.734 0.56 ;
      RECT 7.866 0.5295 8.534 0.56 ;
      RECT 4.666 0.5295 5.334 0.56 ;
      RECT 5.466 0.5295 6.134 0.56 ;
      RECT 0.012 0.5295 0.534 72.1905 ;
      RECT 0.666 0.5295 1.334 0.56 ;
      RECT 1.466 0.5295 2.134 0.56 ;
      RECT 2.266 0.5295 2.934 0.56 ;
      RECT 3.066 0.5295 3.734 0.56 ;
      RECT 3.866 0.5295 4.534 0.56 ;
      RECT 17.356 33.18 17.372 34.14 ;
    LAYER m0 ;
      RECT 0 0.002 36.3 72.718 ;
    LAYER m1 ;
      RECT 0 0 36.3 72.72 ;
    LAYER m2 ;
      RECT 0 0.015 36.3 72.705 ;
    LAYER m3 ;
      RECT 0.015 0 36.285 72.72 ;
    LAYER m4 ;
      RECT 0 0.02 36.3 72.7 ;
  END
  PROPERTY hpml_layer "5" ;
  PROPERTY heml_layer "5" ;
END ip764hduspsr1024x52m4b2s0r2p0d0

END LIBRARY
