VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf124b192e1r1w0cbbehcaa4acw
  CLASS BLOCK ;
  FOREIGN arf124b192e1r1w0cbbehcaa4acw ;
  ORIGIN 0 0 ;
  SIZE 70.2 BY 28.8 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.644 14.76 33.688 15.96 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.644 12.84 33.688 14.04 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.796 14.76 34.84 15.96 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.972 14.76 35.016 15.96 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.272 14.76 35.316 15.96 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.812 14.76 33.856 15.96 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.984 14.76 34.028 15.96 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.284 14.76 34.328 15.96 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.46 14.76 34.504 15.96 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.712 14.76 34.756 15.96 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.896 14.76 33.94 15.96 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.072 14.76 34.116 15.96 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.372 14.76 34.416 15.96 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.544 14.76 34.588 15.96 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.972 12.84 35.016 14.04 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.272 12.84 35.316 14.04 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.812 12.84 33.856 14.04 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.984 12.84 34.028 14.04 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.284 12.84 34.328 14.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.46 12.84 34.504 14.04 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.712 12.84 34.756 14.04 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.884 12.84 34.928 14.04 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.896 12.84 33.94 14.04 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.072 12.84 34.116 14.04 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 23.04 12.988 24.24 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 23.04 13.072 24.24 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 23.04 47.916 24.24 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.044 23.04 48.088 24.24 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 23.76 13.972 24.96 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 23.76 14.056 24.96 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 23.76 48.988 24.96 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 23.76 49.072 24.96 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 24.48 10.372 25.68 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 24.48 10.456 25.68 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 1.68 47.528 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.512 24.48 45.556 25.68 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 24.48 45.728 25.68 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 25.2 11.916 26.4 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 25.2 12.088 26.4 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 25.2 46.928 26.4 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 25.2 47.016 26.4 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 25.92 12.988 27.12 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 25.92 13.072 27.12 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 25.92 47.916 27.12 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.044 25.92 48.088 27.12 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 1.68 47.616 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 26.64 13.972 27.84 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 26.64 14.056 27.84 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 26.64 48.988 27.84 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 26.64 49.072 27.84 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 27.36 10.372 28.56 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 27.36 10.456 28.56 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.512 27.36 45.556 28.56 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 27.36 45.728 28.56 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 2.4 13.628 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 2.4 13.716 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 2.4 48.516 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 2.4 48.728 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.12 14.616 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 3.12 10.116 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 3.12 44.916 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 3.12 45.128 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 3.84 11.356 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 3.84 11.528 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.412 3.84 46.456 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 3.84 46.628 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 4.56 12.516 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 4.56 12.728 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 4.56 47.528 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 4.56 47.616 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 5.28 13.628 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 5.28 13.716 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 0.24 44.916 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 5.28 48.516 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 5.28 48.728 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6 14.616 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 6 10.116 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 6 44.916 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 6 45.128 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 6.72 11.356 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 6.72 11.528 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.412 6.72 46.456 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 6.72 46.628 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 0.24 45.128 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 7.44 12.516 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 7.44 12.728 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 7.44 47.528 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 7.44 47.616 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 8.16 13.628 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 8.16 13.716 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 8.16 48.516 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 8.16 48.728 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.88 14.616 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.88 10.116 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 0.96 11.528 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 8.88 44.916 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 8.88 45.128 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 9.6 11.356 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 9.6 11.528 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.412 9.6 46.456 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 9.6 46.628 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 10.32 12.516 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 10.32 12.728 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 10.32 47.528 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 10.32 47.616 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 0.96 11.616 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.04 13.628 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 11.04 13.716 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 11.04 48.516 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 11.04 48.728 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 16.56 11.356 17.76 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 16.56 11.528 17.76 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.328 16.56 46.372 17.76 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.412 16.56 46.456 17.76 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 17.28 12.988 18.48 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 17.28 13.072 18.48 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.412 0.96 46.456 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 17.28 47.916 18.48 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.044 17.28 48.088 18.48 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 18 13.972 19.2 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 18 14.056 19.2 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 18 48.988 19.2 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 18 49.072 19.2 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 18.72 10.372 19.92 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 18.72 10.456 19.92 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.512 18.72 45.556 19.92 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 18.72 45.728 19.92 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 0.96 46.628 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 19.44 11.916 20.64 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 19.44 12.088 20.64 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 19.44 46.928 20.64 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 19.44 47.016 20.64 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 20.16 12.988 21.36 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 20.16 13.072 21.36 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 20.16 47.916 21.36 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.044 20.16 48.088 21.36 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 20.88 13.972 22.08 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 20.88 14.056 22.08 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 1.68 12.516 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 20.88 48.988 22.08 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 20.88 49.072 22.08 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 21.6 10.372 22.8 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 21.6 10.456 22.8 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.512 21.6 45.556 22.8 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 21.6 45.728 22.8 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 22.32 11.916 23.52 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 22.32 12.088 23.52 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 22.32 46.928 23.52 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 22.32 47.016 23.52 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 1.68 12.728 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.544 12.84 34.588 14.04 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.796 12.84 34.84 14.04 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.372 12.84 34.416 14.04 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 0.24 10.288 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 23.04 13.156 24.24 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 23.04 13.328 24.24 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 23.04 48.172 24.24 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.212 23.04 48.256 24.24 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 23.76 14.228 24.96 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 23.76 14.316 24.96 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 23.76 44.572 24.96 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.612 23.76 44.656 24.96 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 24.48 10.628 25.68 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 24.48 10.716 25.68 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 1.68 47.828 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 24.48 45.816 25.68 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 24.48 46.028 25.68 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 25.2 12.172 26.4 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 25.2 12.256 26.4 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.144 25.2 47.188 26.4 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 25.2 47.272 26.4 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 25.92 13.156 27.12 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 25.92 13.328 27.12 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 25.92 48.172 27.12 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.212 25.92 48.256 27.12 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 1.68 47.916 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 26.64 14.228 27.84 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 26.64 14.316 27.84 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 26.64 44.572 27.84 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.612 26.64 44.656 27.84 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 27.36 10.628 28.56 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 27.36 10.716 28.56 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 27.36 45.816 28.56 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 27.36 46.028 28.56 ;
    END
  END rddatap0[127]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 2.4 13.888 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 2.4 13.972 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 2.4 48.816 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 2.4 48.988 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 3.12 10.288 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 3.12 10.372 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 3.12 45.216 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.344 3.12 45.388 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.24 10.372 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 3.84 11.616 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 3.84 11.828 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 3.84 46.716 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 3.84 46.928 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 4.56 12.816 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 4.56 12.988 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 4.56 47.828 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 4.56 47.916 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 5.28 13.888 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 5.28 13.972 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 0.24 45.216 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 5.28 48.816 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 5.28 48.988 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 6 10.288 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 6 10.372 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 6 45.216 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.344 6 45.388 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 6.72 11.616 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 6.72 11.828 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 6.72 46.716 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 6.72 46.928 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.344 0.24 45.388 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 7.44 12.816 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 7.44 12.988 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 7.44 47.828 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 7.44 47.916 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 8.16 13.888 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 8.16 13.972 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 8.16 48.816 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 8.16 48.988 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 8.88 10.288 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 8.88 10.372 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 0.96 11.828 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 8.88 45.216 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.344 8.88 45.388 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 9.6 11.616 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 9.6 11.828 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 9.6 46.716 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 9.6 46.928 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 10.32 12.816 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 10.32 12.988 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 10.32 47.828 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 10.32 47.916 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 0.96 11.916 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 11.04 13.888 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 11.04 13.972 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 11.04 48.816 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.944 11.04 48.988 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 16.56 11.616 17.76 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 16.56 11.828 17.76 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 16.56 46.628 17.76 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 16.56 46.716 17.76 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 17.28 13.156 18.48 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 17.28 13.328 18.48 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 0.96 46.716 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 17.28 48.172 18.48 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.212 17.28 48.256 18.48 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 18 14.228 19.2 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 18 14.316 19.2 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 18 44.572 19.2 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.612 18 44.656 19.2 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 18.72 10.628 19.92 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 18.72 10.716 19.92 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 18.72 45.816 19.92 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 18.72 46.028 19.92 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 0.96 46.928 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 19.44 12.172 20.64 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 19.44 12.256 20.64 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.144 19.44 47.188 20.64 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 19.44 47.272 20.64 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 20.16 13.156 21.36 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 20.16 13.328 21.36 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 20.16 48.172 21.36 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.212 20.16 48.256 21.36 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 20.88 14.228 22.08 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 20.88 14.316 22.08 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 1.68 12.816 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 20.88 44.572 22.08 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.612 20.88 44.656 22.08 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 21.6 10.628 22.8 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 21.6 10.716 22.8 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 21.6 45.816 22.8 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 21.6 46.028 22.8 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 22.32 12.172 23.52 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 22.32 12.256 23.52 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.144 22.32 47.188 23.52 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 22.32 47.272 23.52 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 1.68 12.988 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 28.74 ;
        RECT 2.662 0.06 2.738 28.74 ;
        RECT 4.462 0.06 4.538 28.74 ;
        RECT 6.262 0.06 6.338 28.74 ;
        RECT 8.062 0.06 8.138 28.74 ;
        RECT 9.862 0.06 9.938 28.74 ;
        RECT 11.662 0.06 11.738 28.74 ;
        RECT 13.462 0.06 13.538 28.74 ;
        RECT 15.262 0.06 15.338 28.74 ;
        RECT 17.062 0.06 17.138 28.74 ;
        RECT 18.862 0.06 18.938 28.74 ;
        RECT 20.662 0.06 20.738 28.74 ;
        RECT 22.462 0.06 22.538 28.74 ;
        RECT 24.262 0.06 24.338 28.74 ;
        RECT 26.062 0.06 26.138 28.74 ;
        RECT 27.862 0.06 27.938 28.74 ;
        RECT 29.662 0.06 29.738 28.74 ;
        RECT 31.462 0.06 31.538 28.74 ;
        RECT 33.262 0.06 33.338 28.74 ;
        RECT 35.062 0.06 35.138 28.74 ;
        RECT 36.862 0.06 36.938 28.74 ;
        RECT 38.662 0.06 38.738 28.74 ;
        RECT 40.462 0.06 40.538 28.74 ;
        RECT 42.262 0.06 42.338 28.74 ;
        RECT 44.062 0.06 44.138 28.74 ;
        RECT 45.862 0.06 45.938 28.74 ;
        RECT 47.662 0.06 47.738 28.74 ;
        RECT 49.462 0.06 49.538 28.74 ;
        RECT 51.262 0.06 51.338 28.74 ;
        RECT 53.062 0.06 53.138 28.74 ;
        RECT 54.862 0.06 54.938 28.74 ;
        RECT 56.662 0.06 56.738 28.74 ;
        RECT 58.462 0.06 58.538 28.74 ;
        RECT 60.262 0.06 60.338 28.74 ;
        RECT 62.062 0.06 62.138 28.74 ;
        RECT 63.862 0.06 63.938 28.74 ;
        RECT 65.662 0.06 65.738 28.74 ;
        RECT 67.462 0.06 67.538 28.74 ;
        RECT 69.262 0.06 69.338 28.74 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 28.74 ;
        RECT 3.562 0.06 3.638 28.74 ;
        RECT 5.362 0.06 5.438 28.74 ;
        RECT 7.162 0.06 7.238 28.74 ;
        RECT 8.962 0.06 9.038 28.74 ;
        RECT 10.762 0.06 10.838 28.74 ;
        RECT 12.562 0.06 12.638 28.74 ;
        RECT 14.362 0.06 14.438 28.74 ;
        RECT 16.162 0.06 16.238 28.74 ;
        RECT 17.962 0.06 18.038 28.74 ;
        RECT 19.762 0.06 19.838 28.74 ;
        RECT 21.562 0.06 21.638 28.74 ;
        RECT 23.362 0.06 23.438 28.74 ;
        RECT 25.162 0.06 25.238 28.74 ;
        RECT 26.962 0.06 27.038 28.74 ;
        RECT 28.762 0.06 28.838 28.74 ;
        RECT 30.562 0.06 30.638 28.74 ;
        RECT 32.362 0.06 32.438 28.74 ;
        RECT 34.162 0.06 34.238 28.74 ;
        RECT 35.962 0.06 36.038 28.74 ;
        RECT 37.762 0.06 37.838 28.74 ;
        RECT 39.562 0.06 39.638 28.74 ;
        RECT 41.362 0.06 41.438 28.74 ;
        RECT 43.162 0.06 43.238 28.74 ;
        RECT 44.962 0.06 45.038 28.74 ;
        RECT 46.762 0.06 46.838 28.74 ;
        RECT 48.562 0.06 48.638 28.74 ;
        RECT 50.362 0.06 50.438 28.74 ;
        RECT 52.162 0.06 52.238 28.74 ;
        RECT 53.962 0.06 54.038 28.74 ;
        RECT 55.762 0.06 55.838 28.74 ;
        RECT 57.562 0.06 57.638 28.74 ;
        RECT 59.362 0.06 59.438 28.74 ;
        RECT 61.162 0.06 61.238 28.74 ;
        RECT 62.962 0.06 63.038 28.74 ;
        RECT 64.762 0.06 64.838 28.74 ;
        RECT 66.562 0.06 66.638 28.74 ;
        RECT 68.362 0.06 68.438 28.74 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 70.216 28.814 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 70.22 28.82 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 70.2705 28.838 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 70.235 28.87 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 70.27 28.838 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 70.259 28.89 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 70.29 28.862 ;
    LAYER m7 SPACING 0 ;
      RECT 69.338 28.86 70.24 28.92 ;
      RECT 69.338 -0.06 70.292 28.86 ;
      RECT 69.338 -0.12 70.24 -0.06 ;
      RECT 68.438 -0.12 69.262 28.92 ;
      RECT 67.538 -0.12 68.362 28.92 ;
      RECT 66.638 -0.12 67.462 28.92 ;
      RECT 65.738 -0.12 66.562 28.92 ;
      RECT 64.838 -0.12 65.662 28.92 ;
      RECT 63.938 -0.12 64.762 28.92 ;
      RECT 63.038 -0.12 63.862 28.92 ;
      RECT 62.138 -0.12 62.962 28.92 ;
      RECT 61.238 -0.12 62.062 28.92 ;
      RECT 60.338 -0.12 61.162 28.92 ;
      RECT 59.438 -0.12 60.262 28.92 ;
      RECT 58.538 -0.12 59.362 28.92 ;
      RECT 57.638 -0.12 58.462 28.92 ;
      RECT 56.738 -0.12 57.562 28.92 ;
      RECT 55.838 -0.12 56.662 28.92 ;
      RECT 54.938 -0.12 55.762 28.92 ;
      RECT 54.038 -0.12 54.862 28.92 ;
      RECT 53.138 -0.12 53.962 28.92 ;
      RECT 52.238 -0.12 53.062 28.92 ;
      RECT 51.338 -0.12 52.162 28.92 ;
      RECT 50.438 -0.12 51.262 28.92 ;
      RECT 49.538 -0.12 50.362 28.92 ;
      RECT 48.638 27.84 49.462 28.92 ;
      RECT 48.638 26.64 48.944 27.84 ;
      RECT 48.988 26.64 49.028 27.84 ;
      RECT 49.072 26.64 49.462 27.84 ;
      RECT 48.638 24.96 49.462 26.64 ;
      RECT 48.638 23.76 48.944 24.96 ;
      RECT 48.988 23.76 49.028 24.96 ;
      RECT 49.072 23.76 49.462 24.96 ;
      RECT 48.638 22.08 49.462 23.76 ;
      RECT 48.638 20.88 48.944 22.08 ;
      RECT 48.988 20.88 49.028 22.08 ;
      RECT 49.072 20.88 49.462 22.08 ;
      RECT 48.638 19.2 49.462 20.88 ;
      RECT 48.638 18 48.944 19.2 ;
      RECT 48.988 18 49.028 19.2 ;
      RECT 49.072 18 49.462 19.2 ;
      RECT 48.638 12.24 49.462 18 ;
      RECT 48.638 11.04 48.684 12.24 ;
      RECT 48.728 11.04 48.772 12.24 ;
      RECT 48.816 11.04 48.944 12.24 ;
      RECT 48.988 11.04 49.462 12.24 ;
      RECT 48.638 9.36 49.462 11.04 ;
      RECT 48.638 8.16 48.684 9.36 ;
      RECT 48.728 8.16 48.772 9.36 ;
      RECT 48.816 8.16 48.944 9.36 ;
      RECT 48.988 8.16 49.462 9.36 ;
      RECT 48.638 6.48 49.462 8.16 ;
      RECT 48.638 5.28 48.684 6.48 ;
      RECT 48.728 5.28 48.772 6.48 ;
      RECT 48.816 5.28 48.944 6.48 ;
      RECT 48.988 5.28 49.462 6.48 ;
      RECT 48.638 3.6 49.462 5.28 ;
      RECT 48.638 2.4 48.684 3.6 ;
      RECT 48.728 2.4 48.772 3.6 ;
      RECT 48.816 2.4 48.944 3.6 ;
      RECT 48.988 2.4 49.462 3.6 ;
      RECT 48.638 -0.12 49.462 2.4 ;
      RECT 47.738 27.12 48.562 28.92 ;
      RECT 47.738 25.92 47.872 27.12 ;
      RECT 47.916 25.92 48.044 27.12 ;
      RECT 48.088 25.92 48.128 27.12 ;
      RECT 48.172 25.92 48.212 27.12 ;
      RECT 48.256 25.92 48.562 27.12 ;
      RECT 47.738 24.24 48.562 25.92 ;
      RECT 47.738 23.04 47.872 24.24 ;
      RECT 47.916 23.04 48.044 24.24 ;
      RECT 48.088 23.04 48.128 24.24 ;
      RECT 48.172 23.04 48.212 24.24 ;
      RECT 48.256 23.04 48.562 24.24 ;
      RECT 47.738 21.36 48.562 23.04 ;
      RECT 47.738 20.16 47.872 21.36 ;
      RECT 47.916 20.16 48.044 21.36 ;
      RECT 48.088 20.16 48.128 21.36 ;
      RECT 48.172 20.16 48.212 21.36 ;
      RECT 48.256 20.16 48.562 21.36 ;
      RECT 47.738 18.48 48.562 20.16 ;
      RECT 47.738 17.28 47.872 18.48 ;
      RECT 47.916 17.28 48.044 18.48 ;
      RECT 48.088 17.28 48.128 18.48 ;
      RECT 48.172 17.28 48.212 18.48 ;
      RECT 48.256 17.28 48.562 18.48 ;
      RECT 47.738 12.24 48.562 17.28 ;
      RECT 47.738 11.52 48.472 12.24 ;
      RECT 48.516 11.04 48.562 12.24 ;
      RECT 47.916 11.04 48.472 11.52 ;
      RECT 47.738 10.32 47.784 11.52 ;
      RECT 47.828 10.32 47.872 11.52 ;
      RECT 47.916 10.32 48.562 11.04 ;
      RECT 47.738 9.36 48.562 10.32 ;
      RECT 47.738 8.64 48.472 9.36 ;
      RECT 48.516 8.16 48.562 9.36 ;
      RECT 47.916 8.16 48.472 8.64 ;
      RECT 47.738 7.44 47.784 8.64 ;
      RECT 47.828 7.44 47.872 8.64 ;
      RECT 47.916 7.44 48.562 8.16 ;
      RECT 47.738 6.48 48.562 7.44 ;
      RECT 47.738 5.76 48.472 6.48 ;
      RECT 48.516 5.28 48.562 6.48 ;
      RECT 47.916 5.28 48.472 5.76 ;
      RECT 47.738 4.56 47.784 5.76 ;
      RECT 47.828 4.56 47.872 5.76 ;
      RECT 47.916 4.56 48.562 5.28 ;
      RECT 47.738 3.6 48.562 4.56 ;
      RECT 47.738 2.88 48.472 3.6 ;
      RECT 48.516 2.4 48.562 3.6 ;
      RECT 47.916 2.4 48.472 2.88 ;
      RECT 47.738 1.68 47.784 2.88 ;
      RECT 47.828 1.68 47.872 2.88 ;
      RECT 47.916 1.68 48.562 2.4 ;
      RECT 47.738 -0.12 48.562 1.68 ;
      RECT 46.838 26.4 47.662 28.92 ;
      RECT 46.838 25.2 46.884 26.4 ;
      RECT 46.928 25.2 46.972 26.4 ;
      RECT 47.016 25.2 47.144 26.4 ;
      RECT 47.188 25.2 47.228 26.4 ;
      RECT 47.272 25.2 47.662 26.4 ;
      RECT 46.838 23.52 47.662 25.2 ;
      RECT 46.838 22.32 46.884 23.52 ;
      RECT 46.928 22.32 46.972 23.52 ;
      RECT 47.016 22.32 47.144 23.52 ;
      RECT 47.188 22.32 47.228 23.52 ;
      RECT 47.272 22.32 47.662 23.52 ;
      RECT 46.838 20.64 47.662 22.32 ;
      RECT 46.838 19.44 46.884 20.64 ;
      RECT 46.928 19.44 46.972 20.64 ;
      RECT 47.016 19.44 47.144 20.64 ;
      RECT 47.188 19.44 47.228 20.64 ;
      RECT 47.272 19.44 47.662 20.64 ;
      RECT 46.838 11.52 47.662 19.44 ;
      RECT 46.838 10.8 47.484 11.52 ;
      RECT 47.528 10.32 47.572 11.52 ;
      RECT 47.616 10.32 47.662 11.52 ;
      RECT 46.928 10.32 47.484 10.8 ;
      RECT 46.838 9.6 46.884 10.8 ;
      RECT 46.928 9.6 47.662 10.32 ;
      RECT 46.838 8.64 47.662 9.6 ;
      RECT 46.838 7.92 47.484 8.64 ;
      RECT 47.528 7.44 47.572 8.64 ;
      RECT 47.616 7.44 47.662 8.64 ;
      RECT 46.928 7.44 47.484 7.92 ;
      RECT 46.838 6.72 46.884 7.92 ;
      RECT 46.928 6.72 47.662 7.44 ;
      RECT 46.838 5.76 47.662 6.72 ;
      RECT 46.838 5.04 47.484 5.76 ;
      RECT 47.528 4.56 47.572 5.76 ;
      RECT 47.616 4.56 47.662 5.76 ;
      RECT 46.928 4.56 47.484 5.04 ;
      RECT 46.838 3.84 46.884 5.04 ;
      RECT 46.928 3.84 47.662 4.56 ;
      RECT 46.838 2.88 47.662 3.84 ;
      RECT 46.838 2.16 47.484 2.88 ;
      RECT 47.528 1.68 47.572 2.88 ;
      RECT 47.616 1.68 47.662 2.88 ;
      RECT 46.928 1.68 47.484 2.16 ;
      RECT 46.838 0.96 46.884 2.16 ;
      RECT 46.928 0.96 47.662 1.68 ;
      RECT 46.838 -0.12 47.662 0.96 ;
      RECT 45.938 28.56 46.762 28.92 ;
      RECT 45.938 27.36 45.984 28.56 ;
      RECT 46.028 27.36 46.762 28.56 ;
      RECT 45.938 25.68 46.762 27.36 ;
      RECT 45.938 24.48 45.984 25.68 ;
      RECT 46.028 24.48 46.762 25.68 ;
      RECT 45.938 22.8 46.762 24.48 ;
      RECT 45.938 21.6 45.984 22.8 ;
      RECT 46.028 21.6 46.762 22.8 ;
      RECT 45.938 19.92 46.762 21.6 ;
      RECT 45.938 18.72 45.984 19.92 ;
      RECT 46.028 18.72 46.762 19.92 ;
      RECT 45.938 17.76 46.762 18.72 ;
      RECT 45.938 16.56 46.328 17.76 ;
      RECT 46.372 16.56 46.412 17.76 ;
      RECT 46.456 16.56 46.584 17.76 ;
      RECT 46.628 16.56 46.672 17.76 ;
      RECT 46.716 16.56 46.762 17.76 ;
      RECT 45.938 10.8 46.762 16.56 ;
      RECT 45.938 9.6 46.412 10.8 ;
      RECT 46.456 9.6 46.584 10.8 ;
      RECT 46.628 9.6 46.672 10.8 ;
      RECT 46.716 9.6 46.762 10.8 ;
      RECT 45.938 7.92 46.762 9.6 ;
      RECT 45.938 6.72 46.412 7.92 ;
      RECT 46.456 6.72 46.584 7.92 ;
      RECT 46.628 6.72 46.672 7.92 ;
      RECT 46.716 6.72 46.762 7.92 ;
      RECT 45.938 5.04 46.762 6.72 ;
      RECT 45.938 3.84 46.412 5.04 ;
      RECT 46.456 3.84 46.584 5.04 ;
      RECT 46.628 3.84 46.672 5.04 ;
      RECT 46.716 3.84 46.762 5.04 ;
      RECT 45.938 2.16 46.762 3.84 ;
      RECT 45.938 0.96 46.412 2.16 ;
      RECT 46.456 0.96 46.584 2.16 ;
      RECT 46.628 0.96 46.672 2.16 ;
      RECT 46.716 0.96 46.762 2.16 ;
      RECT 45.938 -0.12 46.762 0.96 ;
      RECT 45.038 28.56 45.862 28.92 ;
      RECT 45.038 27.36 45.512 28.56 ;
      RECT 45.556 27.36 45.684 28.56 ;
      RECT 45.728 27.36 45.772 28.56 ;
      RECT 45.816 27.36 45.862 28.56 ;
      RECT 45.038 25.68 45.862 27.36 ;
      RECT 45.038 24.48 45.512 25.68 ;
      RECT 45.556 24.48 45.684 25.68 ;
      RECT 45.728 24.48 45.772 25.68 ;
      RECT 45.816 24.48 45.862 25.68 ;
      RECT 45.038 22.8 45.862 24.48 ;
      RECT 45.038 21.6 45.512 22.8 ;
      RECT 45.556 21.6 45.684 22.8 ;
      RECT 45.728 21.6 45.772 22.8 ;
      RECT 45.816 21.6 45.862 22.8 ;
      RECT 45.038 19.92 45.862 21.6 ;
      RECT 45.038 18.72 45.512 19.92 ;
      RECT 45.556 18.72 45.684 19.92 ;
      RECT 45.728 18.72 45.772 19.92 ;
      RECT 45.816 18.72 45.862 19.92 ;
      RECT 45.038 10.08 45.862 18.72 ;
      RECT 45.038 8.88 45.084 10.08 ;
      RECT 45.128 8.88 45.172 10.08 ;
      RECT 45.216 8.88 45.344 10.08 ;
      RECT 45.388 8.88 45.862 10.08 ;
      RECT 45.038 7.2 45.862 8.88 ;
      RECT 45.038 6 45.084 7.2 ;
      RECT 45.128 6 45.172 7.2 ;
      RECT 45.216 6 45.344 7.2 ;
      RECT 45.388 6 45.862 7.2 ;
      RECT 45.038 4.32 45.862 6 ;
      RECT 45.038 3.12 45.084 4.32 ;
      RECT 45.128 3.12 45.172 4.32 ;
      RECT 45.216 3.12 45.344 4.32 ;
      RECT 45.388 3.12 45.862 4.32 ;
      RECT 45.038 1.44 45.862 3.12 ;
      RECT 45.038 0.24 45.084 1.44 ;
      RECT 45.128 0.24 45.172 1.44 ;
      RECT 45.216 0.24 45.344 1.44 ;
      RECT 45.388 0.24 45.862 1.44 ;
      RECT 45.038 -0.12 45.862 0.24 ;
      RECT 44.138 27.84 44.962 28.92 ;
      RECT 44.138 26.64 44.528 27.84 ;
      RECT 44.572 26.64 44.612 27.84 ;
      RECT 44.656 26.64 44.962 27.84 ;
      RECT 44.138 24.96 44.962 26.64 ;
      RECT 44.138 23.76 44.528 24.96 ;
      RECT 44.572 23.76 44.612 24.96 ;
      RECT 44.656 23.76 44.962 24.96 ;
      RECT 44.138 22.08 44.962 23.76 ;
      RECT 44.138 20.88 44.528 22.08 ;
      RECT 44.572 20.88 44.612 22.08 ;
      RECT 44.656 20.88 44.962 22.08 ;
      RECT 44.138 19.2 44.962 20.88 ;
      RECT 44.138 18 44.528 19.2 ;
      RECT 44.572 18 44.612 19.2 ;
      RECT 44.656 18 44.962 19.2 ;
      RECT 44.138 10.08 44.962 18 ;
      RECT 44.138 8.88 44.872 10.08 ;
      RECT 44.916 8.88 44.962 10.08 ;
      RECT 44.138 7.2 44.962 8.88 ;
      RECT 44.138 6 44.872 7.2 ;
      RECT 44.916 6 44.962 7.2 ;
      RECT 44.138 4.32 44.962 6 ;
      RECT 44.138 3.12 44.872 4.32 ;
      RECT 44.916 3.12 44.962 4.32 ;
      RECT 44.138 1.44 44.962 3.12 ;
      RECT 44.138 0.24 44.872 1.44 ;
      RECT 44.916 0.24 44.962 1.44 ;
      RECT 44.138 -0.12 44.962 0.24 ;
      RECT 43.238 -0.12 44.062 28.92 ;
      RECT 42.338 -0.12 43.162 28.92 ;
      RECT 41.438 -0.12 42.262 28.92 ;
      RECT 40.538 -0.12 41.362 28.92 ;
      RECT 39.638 -0.12 40.462 28.92 ;
      RECT 38.738 -0.12 39.562 28.92 ;
      RECT 37.838 -0.12 38.662 28.92 ;
      RECT 36.938 -0.12 37.762 28.92 ;
      RECT 36.038 -0.12 36.862 28.92 ;
      RECT 35.138 15.96 35.962 28.92 ;
      RECT 35.138 14.76 35.272 15.96 ;
      RECT 35.316 14.76 35.962 15.96 ;
      RECT 35.138 14.04 35.962 14.76 ;
      RECT 35.138 12.84 35.272 14.04 ;
      RECT 35.316 12.84 35.962 14.04 ;
      RECT 35.138 -0.12 35.962 12.84 ;
      RECT 34.238 15.96 35.062 28.92 ;
      RECT 34.238 14.76 34.284 15.96 ;
      RECT 34.328 14.76 34.372 15.96 ;
      RECT 34.416 14.76 34.46 15.96 ;
      RECT 34.504 14.76 34.544 15.96 ;
      RECT 34.588 14.76 34.712 15.96 ;
      RECT 34.756 14.76 34.796 15.96 ;
      RECT 34.84 14.76 34.972 15.96 ;
      RECT 35.016 14.76 35.062 15.96 ;
      RECT 34.238 14.04 35.062 14.76 ;
      RECT 34.238 12.84 34.284 14.04 ;
      RECT 34.328 12.84 34.372 14.04 ;
      RECT 34.416 12.84 34.46 14.04 ;
      RECT 34.504 12.84 34.544 14.04 ;
      RECT 34.588 12.84 34.712 14.04 ;
      RECT 34.756 12.84 34.796 14.04 ;
      RECT 34.84 12.84 34.884 14.04 ;
      RECT 34.928 12.84 34.972 14.04 ;
      RECT 35.016 12.84 35.062 14.04 ;
      RECT 34.238 -0.12 35.062 12.84 ;
      RECT 33.338 15.96 34.162 28.92 ;
      RECT 33.338 14.76 33.644 15.96 ;
      RECT 33.688 14.76 33.812 15.96 ;
      RECT 33.856 14.76 33.896 15.96 ;
      RECT 33.94 14.76 33.984 15.96 ;
      RECT 34.028 14.76 34.072 15.96 ;
      RECT 34.116 14.76 34.162 15.96 ;
      RECT 33.338 14.04 34.162 14.76 ;
      RECT 33.338 12.84 33.644 14.04 ;
      RECT 33.688 12.84 33.812 14.04 ;
      RECT 33.856 12.84 33.896 14.04 ;
      RECT 33.94 12.84 33.984 14.04 ;
      RECT 34.028 12.84 34.072 14.04 ;
      RECT 34.116 12.84 34.162 14.04 ;
      RECT 33.338 -0.12 34.162 12.84 ;
      RECT 32.438 -0.12 33.262 28.92 ;
      RECT 31.538 -0.12 32.362 28.92 ;
      RECT 30.638 -0.12 31.462 28.92 ;
      RECT 29.738 -0.12 30.562 28.92 ;
      RECT 28.838 -0.12 29.662 28.92 ;
      RECT 27.938 -0.12 28.762 28.92 ;
      RECT 27.038 -0.12 27.862 28.92 ;
      RECT 26.138 -0.12 26.962 28.92 ;
      RECT 25.238 -0.12 26.062 28.92 ;
      RECT 24.338 -0.12 25.162 28.92 ;
      RECT 23.438 -0.12 24.262 28.92 ;
      RECT 22.538 -0.12 23.362 28.92 ;
      RECT 21.638 -0.12 22.462 28.92 ;
      RECT 20.738 -0.12 21.562 28.92 ;
      RECT 19.838 -0.12 20.662 28.92 ;
      RECT 18.938 -0.12 19.762 28.92 ;
      RECT 18.038 -0.12 18.862 28.92 ;
      RECT 17.138 -0.12 17.962 28.92 ;
      RECT 16.238 -0.12 17.062 28.92 ;
      RECT 15.338 -0.12 16.162 28.92 ;
      RECT 14.438 10.08 15.262 28.92 ;
      RECT 14.438 8.88 14.572 10.08 ;
      RECT 14.616 8.88 15.262 10.08 ;
      RECT 14.438 7.2 15.262 8.88 ;
      RECT 14.438 6 14.572 7.2 ;
      RECT 14.616 6 15.262 7.2 ;
      RECT 14.438 4.32 15.262 6 ;
      RECT 14.438 3.12 14.572 4.32 ;
      RECT 14.616 3.12 15.262 4.32 ;
      RECT 14.438 -0.12 15.262 3.12 ;
      RECT 13.538 27.84 14.362 28.92 ;
      RECT 13.538 26.64 13.928 27.84 ;
      RECT 13.972 26.64 14.012 27.84 ;
      RECT 14.056 26.64 14.184 27.84 ;
      RECT 14.228 26.64 14.272 27.84 ;
      RECT 14.316 26.64 14.362 27.84 ;
      RECT 13.538 24.96 14.362 26.64 ;
      RECT 13.538 23.76 13.928 24.96 ;
      RECT 13.972 23.76 14.012 24.96 ;
      RECT 14.056 23.76 14.184 24.96 ;
      RECT 14.228 23.76 14.272 24.96 ;
      RECT 14.316 23.76 14.362 24.96 ;
      RECT 13.538 22.08 14.362 23.76 ;
      RECT 13.538 20.88 13.928 22.08 ;
      RECT 13.972 20.88 14.012 22.08 ;
      RECT 14.056 20.88 14.184 22.08 ;
      RECT 14.228 20.88 14.272 22.08 ;
      RECT 14.316 20.88 14.362 22.08 ;
      RECT 13.538 19.2 14.362 20.88 ;
      RECT 13.538 18 13.928 19.2 ;
      RECT 13.972 18 14.012 19.2 ;
      RECT 14.056 18 14.184 19.2 ;
      RECT 14.228 18 14.272 19.2 ;
      RECT 14.316 18 14.362 19.2 ;
      RECT 13.538 12.24 14.362 18 ;
      RECT 13.538 11.04 13.584 12.24 ;
      RECT 13.628 11.04 13.672 12.24 ;
      RECT 13.716 11.04 13.844 12.24 ;
      RECT 13.888 11.04 13.928 12.24 ;
      RECT 13.972 11.04 14.362 12.24 ;
      RECT 13.538 9.36 14.362 11.04 ;
      RECT 13.538 8.16 13.584 9.36 ;
      RECT 13.628 8.16 13.672 9.36 ;
      RECT 13.716 8.16 13.844 9.36 ;
      RECT 13.888 8.16 13.928 9.36 ;
      RECT 13.972 8.16 14.362 9.36 ;
      RECT 13.538 6.48 14.362 8.16 ;
      RECT 13.538 5.28 13.584 6.48 ;
      RECT 13.628 5.28 13.672 6.48 ;
      RECT 13.716 5.28 13.844 6.48 ;
      RECT 13.888 5.28 13.928 6.48 ;
      RECT 13.972 5.28 14.362 6.48 ;
      RECT 13.538 3.6 14.362 5.28 ;
      RECT 13.538 2.4 13.584 3.6 ;
      RECT 13.628 2.4 13.672 3.6 ;
      RECT 13.716 2.4 13.844 3.6 ;
      RECT 13.888 2.4 13.928 3.6 ;
      RECT 13.972 2.4 14.362 3.6 ;
      RECT 13.538 -0.12 14.362 2.4 ;
      RECT 12.638 27.12 13.462 28.92 ;
      RECT 12.638 25.92 12.944 27.12 ;
      RECT 12.988 25.92 13.028 27.12 ;
      RECT 13.072 25.92 13.112 27.12 ;
      RECT 13.156 25.92 13.284 27.12 ;
      RECT 13.328 25.92 13.462 27.12 ;
      RECT 12.638 24.24 13.462 25.92 ;
      RECT 12.638 23.04 12.944 24.24 ;
      RECT 12.988 23.04 13.028 24.24 ;
      RECT 13.072 23.04 13.112 24.24 ;
      RECT 13.156 23.04 13.284 24.24 ;
      RECT 13.328 23.04 13.462 24.24 ;
      RECT 12.638 21.36 13.462 23.04 ;
      RECT 12.638 20.16 12.944 21.36 ;
      RECT 12.988 20.16 13.028 21.36 ;
      RECT 13.072 20.16 13.112 21.36 ;
      RECT 13.156 20.16 13.284 21.36 ;
      RECT 13.328 20.16 13.462 21.36 ;
      RECT 12.638 18.48 13.462 20.16 ;
      RECT 12.638 17.28 12.944 18.48 ;
      RECT 12.988 17.28 13.028 18.48 ;
      RECT 13.072 17.28 13.112 18.48 ;
      RECT 13.156 17.28 13.284 18.48 ;
      RECT 13.328 17.28 13.462 18.48 ;
      RECT 12.638 11.52 13.462 17.28 ;
      RECT 12.638 10.32 12.684 11.52 ;
      RECT 12.728 10.32 12.772 11.52 ;
      RECT 12.816 10.32 12.944 11.52 ;
      RECT 12.988 10.32 13.462 11.52 ;
      RECT 12.638 8.64 13.462 10.32 ;
      RECT 12.638 7.44 12.684 8.64 ;
      RECT 12.728 7.44 12.772 8.64 ;
      RECT 12.816 7.44 12.944 8.64 ;
      RECT 12.988 7.44 13.462 8.64 ;
      RECT 12.638 5.76 13.462 7.44 ;
      RECT 12.638 4.56 12.684 5.76 ;
      RECT 12.728 4.56 12.772 5.76 ;
      RECT 12.816 4.56 12.944 5.76 ;
      RECT 12.988 4.56 13.462 5.76 ;
      RECT 12.638 2.88 13.462 4.56 ;
      RECT 12.638 1.68 12.684 2.88 ;
      RECT 12.728 1.68 12.772 2.88 ;
      RECT 12.816 1.68 12.944 2.88 ;
      RECT 12.988 1.68 13.462 2.88 ;
      RECT 12.638 -0.12 13.462 1.68 ;
      RECT 11.738 26.4 12.562 28.92 ;
      RECT 11.738 25.2 11.872 26.4 ;
      RECT 11.916 25.2 12.044 26.4 ;
      RECT 12.088 25.2 12.128 26.4 ;
      RECT 12.172 25.2 12.212 26.4 ;
      RECT 12.256 25.2 12.562 26.4 ;
      RECT 11.738 23.52 12.562 25.2 ;
      RECT 11.738 22.32 11.872 23.52 ;
      RECT 11.916 22.32 12.044 23.52 ;
      RECT 12.088 22.32 12.128 23.52 ;
      RECT 12.172 22.32 12.212 23.52 ;
      RECT 12.256 22.32 12.562 23.52 ;
      RECT 11.738 20.64 12.562 22.32 ;
      RECT 11.738 19.44 11.872 20.64 ;
      RECT 11.916 19.44 12.044 20.64 ;
      RECT 12.088 19.44 12.128 20.64 ;
      RECT 12.172 19.44 12.212 20.64 ;
      RECT 12.256 19.44 12.562 20.64 ;
      RECT 11.738 17.76 12.562 19.44 ;
      RECT 11.738 16.56 11.784 17.76 ;
      RECT 11.828 16.56 12.562 17.76 ;
      RECT 11.738 11.52 12.562 16.56 ;
      RECT 11.738 10.8 12.472 11.52 ;
      RECT 12.516 10.32 12.562 11.52 ;
      RECT 11.828 10.32 12.472 10.8 ;
      RECT 11.738 9.6 11.784 10.8 ;
      RECT 11.828 9.6 12.562 10.32 ;
      RECT 11.738 8.64 12.562 9.6 ;
      RECT 11.738 7.92 12.472 8.64 ;
      RECT 12.516 7.44 12.562 8.64 ;
      RECT 11.828 7.44 12.472 7.92 ;
      RECT 11.738 6.72 11.784 7.92 ;
      RECT 11.828 6.72 12.562 7.44 ;
      RECT 11.738 5.76 12.562 6.72 ;
      RECT 11.738 5.04 12.472 5.76 ;
      RECT 12.516 4.56 12.562 5.76 ;
      RECT 11.828 4.56 12.472 5.04 ;
      RECT 11.738 3.84 11.784 5.04 ;
      RECT 11.828 3.84 12.562 4.56 ;
      RECT 11.738 2.88 12.562 3.84 ;
      RECT 11.738 2.16 12.472 2.88 ;
      RECT 12.516 1.68 12.562 2.88 ;
      RECT 11.916 1.68 12.472 2.16 ;
      RECT 11.738 0.96 11.784 2.16 ;
      RECT 11.828 0.96 11.872 2.16 ;
      RECT 11.916 0.96 12.562 1.68 ;
      RECT 11.738 -0.12 12.562 0.96 ;
      RECT 10.838 17.76 11.662 28.92 ;
      RECT 10.838 16.56 11.312 17.76 ;
      RECT 11.356 16.56 11.484 17.76 ;
      RECT 11.528 16.56 11.572 17.76 ;
      RECT 11.616 16.56 11.662 17.76 ;
      RECT 10.838 10.8 11.662 16.56 ;
      RECT 10.838 9.6 11.312 10.8 ;
      RECT 11.356 9.6 11.484 10.8 ;
      RECT 11.528 9.6 11.572 10.8 ;
      RECT 11.616 9.6 11.662 10.8 ;
      RECT 10.838 7.92 11.662 9.6 ;
      RECT 10.838 6.72 11.312 7.92 ;
      RECT 11.356 6.72 11.484 7.92 ;
      RECT 11.528 6.72 11.572 7.92 ;
      RECT 11.616 6.72 11.662 7.92 ;
      RECT 10.838 5.04 11.662 6.72 ;
      RECT 10.838 3.84 11.312 5.04 ;
      RECT 11.356 3.84 11.484 5.04 ;
      RECT 11.528 3.84 11.572 5.04 ;
      RECT 11.616 3.84 11.662 5.04 ;
      RECT 10.838 2.16 11.662 3.84 ;
      RECT 10.838 0.96 11.484 2.16 ;
      RECT 11.528 0.96 11.572 2.16 ;
      RECT 11.616 0.96 11.662 2.16 ;
      RECT 10.838 -0.12 11.662 0.96 ;
      RECT 9.938 28.56 10.762 28.92 ;
      RECT 9.938 27.36 10.328 28.56 ;
      RECT 10.372 27.36 10.412 28.56 ;
      RECT 10.456 27.36 10.584 28.56 ;
      RECT 10.628 27.36 10.672 28.56 ;
      RECT 10.716 27.36 10.762 28.56 ;
      RECT 9.938 25.68 10.762 27.36 ;
      RECT 9.938 24.48 10.328 25.68 ;
      RECT 10.372 24.48 10.412 25.68 ;
      RECT 10.456 24.48 10.584 25.68 ;
      RECT 10.628 24.48 10.672 25.68 ;
      RECT 10.716 24.48 10.762 25.68 ;
      RECT 9.938 22.8 10.762 24.48 ;
      RECT 9.938 21.6 10.328 22.8 ;
      RECT 10.372 21.6 10.412 22.8 ;
      RECT 10.456 21.6 10.584 22.8 ;
      RECT 10.628 21.6 10.672 22.8 ;
      RECT 10.716 21.6 10.762 22.8 ;
      RECT 9.938 19.92 10.762 21.6 ;
      RECT 9.938 18.72 10.328 19.92 ;
      RECT 10.372 18.72 10.412 19.92 ;
      RECT 10.456 18.72 10.584 19.92 ;
      RECT 10.628 18.72 10.672 19.92 ;
      RECT 10.716 18.72 10.762 19.92 ;
      RECT 9.938 10.08 10.762 18.72 ;
      RECT 9.938 8.88 10.072 10.08 ;
      RECT 10.116 8.88 10.244 10.08 ;
      RECT 10.288 8.88 10.328 10.08 ;
      RECT 10.372 8.88 10.762 10.08 ;
      RECT 9.938 7.2 10.762 8.88 ;
      RECT 9.938 6 10.072 7.2 ;
      RECT 10.116 6 10.244 7.2 ;
      RECT 10.288 6 10.328 7.2 ;
      RECT 10.372 6 10.762 7.2 ;
      RECT 9.938 4.32 10.762 6 ;
      RECT 9.938 3.12 10.072 4.32 ;
      RECT 10.116 3.12 10.244 4.32 ;
      RECT 10.288 3.12 10.328 4.32 ;
      RECT 10.372 3.12 10.762 4.32 ;
      RECT 9.938 1.44 10.762 3.12 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.244 1.44 ;
      RECT 10.288 0.24 10.328 1.44 ;
      RECT 10.372 0.24 10.762 1.44 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 28.92 ;
      RECT 8.138 -0.12 8.962 28.92 ;
      RECT 7.238 -0.12 8.062 28.92 ;
      RECT 6.338 -0.12 7.162 28.92 ;
      RECT 5.438 -0.12 6.262 28.92 ;
      RECT 4.538 -0.12 5.362 28.92 ;
      RECT 3.638 -0.12 4.462 28.92 ;
      RECT 2.738 -0.12 3.562 28.92 ;
      RECT 1.838 -0.12 2.662 28.92 ;
      RECT 0.938 -0.12 1.762 28.92 ;
      RECT -0.04 28.86 0.862 28.92 ;
      RECT -0.092 -0.06 0.862 28.86 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 69.458 0 70.12 28.8 ;
      RECT 68.558 0 69.142 28.8 ;
      RECT 67.658 0 68.242 28.8 ;
      RECT 66.758 0 67.342 28.8 ;
      RECT 65.858 0 66.442 28.8 ;
      RECT 64.958 0 65.542 28.8 ;
      RECT 64.058 0 64.642 28.8 ;
      RECT 63.158 0 63.742 28.8 ;
      RECT 62.258 0 62.842 28.8 ;
      RECT 61.358 0 61.942 28.8 ;
      RECT 60.458 0 61.042 28.8 ;
      RECT 59.558 0 60.142 28.8 ;
      RECT 58.658 0 59.242 28.8 ;
      RECT 57.758 0 58.342 28.8 ;
      RECT 56.858 0 57.442 28.8 ;
      RECT 55.958 0 56.542 28.8 ;
      RECT 55.058 0 55.642 28.8 ;
      RECT 54.158 0 54.742 28.8 ;
      RECT 53.258 0 53.842 28.8 ;
      RECT 52.358 0 52.942 28.8 ;
      RECT 51.458 0 52.042 28.8 ;
      RECT 50.558 0 51.142 28.8 ;
      RECT 49.658 0 50.242 28.8 ;
      RECT 48.758 27.96 49.342 28.8 ;
      RECT 48.758 26.52 48.824 27.96 ;
      RECT 49.192 26.52 49.342 27.96 ;
      RECT 48.758 25.08 49.342 26.52 ;
      RECT 48.758 23.64 48.824 25.08 ;
      RECT 49.192 23.64 49.342 25.08 ;
      RECT 48.758 22.2 49.342 23.64 ;
      RECT 48.758 20.76 48.824 22.2 ;
      RECT 49.192 20.76 49.342 22.2 ;
      RECT 48.758 19.32 49.342 20.76 ;
      RECT 48.758 17.88 48.824 19.32 ;
      RECT 49.192 17.88 49.342 19.32 ;
      RECT 48.758 12.36 49.342 17.88 ;
      RECT 49.108 10.92 49.342 12.36 ;
      RECT 48.758 9.48 49.342 10.92 ;
      RECT 49.108 8.04 49.342 9.48 ;
      RECT 48.758 6.6 49.342 8.04 ;
      RECT 49.108 5.16 49.342 6.6 ;
      RECT 48.758 3.72 49.342 5.16 ;
      RECT 49.108 2.28 49.342 3.72 ;
      RECT 48.758 0 49.342 2.28 ;
      RECT 47.858 27.24 48.442 28.8 ;
      RECT 48.376 25.8 48.442 27.24 ;
      RECT 47.858 24.36 48.442 25.8 ;
      RECT 48.376 22.92 48.442 24.36 ;
      RECT 47.858 21.48 48.442 22.92 ;
      RECT 48.376 20.04 48.442 21.48 ;
      RECT 47.858 18.6 48.442 20.04 ;
      RECT 48.376 17.16 48.442 18.6 ;
      RECT 47.858 12.36 48.442 17.16 ;
      RECT 47.858 11.64 48.352 12.36 ;
      RECT 48.036 10.92 48.352 11.64 ;
      RECT 48.036 10.2 48.442 10.92 ;
      RECT 47.858 9.48 48.442 10.2 ;
      RECT 47.858 8.76 48.352 9.48 ;
      RECT 48.036 8.04 48.352 8.76 ;
      RECT 48.036 7.32 48.442 8.04 ;
      RECT 47.858 6.6 48.442 7.32 ;
      RECT 47.858 5.88 48.352 6.6 ;
      RECT 48.036 5.16 48.352 5.88 ;
      RECT 48.036 4.44 48.442 5.16 ;
      RECT 47.858 3.72 48.442 4.44 ;
      RECT 47.858 3 48.352 3.72 ;
      RECT 48.036 2.28 48.352 3 ;
      RECT 48.036 1.56 48.442 2.28 ;
      RECT 47.858 0 48.442 1.56 ;
      RECT 46.958 26.52 47.542 28.8 ;
      RECT 47.392 25.08 47.542 26.52 ;
      RECT 46.958 23.64 47.542 25.08 ;
      RECT 47.392 22.2 47.542 23.64 ;
      RECT 46.958 20.76 47.542 22.2 ;
      RECT 47.392 19.32 47.542 20.76 ;
      RECT 46.958 11.64 47.542 19.32 ;
      RECT 46.958 10.92 47.364 11.64 ;
      RECT 47.048 10.2 47.364 10.92 ;
      RECT 47.048 9.48 47.542 10.2 ;
      RECT 46.958 8.76 47.542 9.48 ;
      RECT 46.958 8.04 47.364 8.76 ;
      RECT 47.048 7.32 47.364 8.04 ;
      RECT 47.048 6.6 47.542 7.32 ;
      RECT 46.958 5.88 47.542 6.6 ;
      RECT 46.958 5.16 47.364 5.88 ;
      RECT 47.048 4.44 47.364 5.16 ;
      RECT 47.048 3.72 47.542 4.44 ;
      RECT 46.958 3 47.542 3.72 ;
      RECT 46.958 2.28 47.364 3 ;
      RECT 47.048 1.56 47.364 2.28 ;
      RECT 47.048 0.84 47.542 1.56 ;
      RECT 46.958 0 47.542 0.84 ;
      RECT 46.058 28.68 46.642 28.8 ;
      RECT 46.148 27.24 46.642 28.68 ;
      RECT 46.058 25.8 46.642 27.24 ;
      RECT 46.148 24.36 46.642 25.8 ;
      RECT 46.058 22.92 46.642 24.36 ;
      RECT 46.148 21.48 46.642 22.92 ;
      RECT 46.058 20.04 46.642 21.48 ;
      RECT 46.148 18.6 46.642 20.04 ;
      RECT 46.058 17.88 46.642 18.6 ;
      RECT 46.058 16.44 46.208 17.88 ;
      RECT 46.058 10.92 46.642 16.44 ;
      RECT 46.058 9.48 46.292 10.92 ;
      RECT 46.058 8.04 46.642 9.48 ;
      RECT 46.058 6.6 46.292 8.04 ;
      RECT 46.058 5.16 46.642 6.6 ;
      RECT 46.058 3.72 46.292 5.16 ;
      RECT 46.058 2.28 46.642 3.72 ;
      RECT 46.058 0.84 46.292 2.28 ;
      RECT 46.058 0 46.642 0.84 ;
      RECT 45.158 28.68 45.742 28.8 ;
      RECT 45.158 27.24 45.392 28.68 ;
      RECT 45.158 25.8 45.742 27.24 ;
      RECT 45.158 24.36 45.392 25.8 ;
      RECT 45.158 22.92 45.742 24.36 ;
      RECT 45.158 21.48 45.392 22.92 ;
      RECT 45.158 20.04 45.742 21.48 ;
      RECT 45.158 18.6 45.392 20.04 ;
      RECT 45.158 10.2 45.742 18.6 ;
      RECT 45.508 8.76 45.742 10.2 ;
      RECT 45.158 7.32 45.742 8.76 ;
      RECT 45.508 5.88 45.742 7.32 ;
      RECT 45.158 4.44 45.742 5.88 ;
      RECT 45.508 3 45.742 4.44 ;
      RECT 45.158 1.56 45.742 3 ;
      RECT 45.508 0.12 45.742 1.56 ;
      RECT 45.158 0 45.742 0.12 ;
      RECT 44.258 27.96 44.842 28.8 ;
      RECT 44.258 26.52 44.408 27.96 ;
      RECT 44.776 26.52 44.842 27.96 ;
      RECT 44.258 25.08 44.842 26.52 ;
      RECT 44.258 23.64 44.408 25.08 ;
      RECT 44.776 23.64 44.842 25.08 ;
      RECT 44.258 22.2 44.842 23.64 ;
      RECT 44.258 20.76 44.408 22.2 ;
      RECT 44.776 20.76 44.842 22.2 ;
      RECT 44.258 19.32 44.842 20.76 ;
      RECT 44.258 17.88 44.408 19.32 ;
      RECT 44.776 17.88 44.842 19.32 ;
      RECT 44.258 10.2 44.842 17.88 ;
      RECT 44.258 8.76 44.752 10.2 ;
      RECT 44.258 7.32 44.842 8.76 ;
      RECT 44.258 5.88 44.752 7.32 ;
      RECT 44.258 4.44 44.842 5.88 ;
      RECT 44.258 3 44.752 4.44 ;
      RECT 44.258 1.56 44.842 3 ;
      RECT 44.258 0.12 44.752 1.56 ;
      RECT 44.258 0 44.842 0.12 ;
      RECT 43.358 0 43.942 28.8 ;
      RECT 42.458 0 43.042 28.8 ;
      RECT 41.558 0 42.142 28.8 ;
      RECT 40.658 0 41.242 28.8 ;
      RECT 39.758 0 40.342 28.8 ;
      RECT 38.858 0 39.442 28.8 ;
      RECT 37.958 0 38.542 28.8 ;
      RECT 37.058 0 37.642 28.8 ;
      RECT 36.158 0 36.742 28.8 ;
      RECT 35.258 16.08 35.842 28.8 ;
      RECT 35.436 14.64 35.842 16.08 ;
      RECT 35.258 14.16 35.842 14.64 ;
      RECT 35.436 12.72 35.842 14.16 ;
      RECT 35.258 0 35.842 12.72 ;
      RECT 34.358 16.08 34.942 28.8 ;
      RECT 33.458 16.08 34.042 28.8 ;
      RECT 33.458 14.64 33.524 16.08 ;
      RECT 33.458 14.16 34.042 14.64 ;
      RECT 33.458 12.72 33.524 14.16 ;
      RECT 33.458 0 34.042 12.72 ;
      RECT 32.558 0 33.142 28.8 ;
      RECT 31.658 0 32.242 28.8 ;
      RECT 30.758 0 31.342 28.8 ;
      RECT 29.858 0 30.442 28.8 ;
      RECT 28.958 0 29.542 28.8 ;
      RECT 28.058 0 28.642 28.8 ;
      RECT 27.158 0 27.742 28.8 ;
      RECT 26.258 0 26.842 28.8 ;
      RECT 25.358 0 25.942 28.8 ;
      RECT 24.458 0 25.042 28.8 ;
      RECT 23.558 0 24.142 28.8 ;
      RECT 22.658 0 23.242 28.8 ;
      RECT 21.758 0 22.342 28.8 ;
      RECT 20.858 0 21.442 28.8 ;
      RECT 19.958 0 20.542 28.8 ;
      RECT 19.058 0 19.642 28.8 ;
      RECT 18.158 0 18.742 28.8 ;
      RECT 17.258 0 17.842 28.8 ;
      RECT 16.358 0 16.942 28.8 ;
      RECT 15.458 0 16.042 28.8 ;
      RECT 14.558 10.2 15.142 28.8 ;
      RECT 14.736 8.76 15.142 10.2 ;
      RECT 14.558 7.32 15.142 8.76 ;
      RECT 14.736 5.88 15.142 7.32 ;
      RECT 14.558 4.44 15.142 5.88 ;
      RECT 14.736 3 15.142 4.44 ;
      RECT 14.558 0 15.142 3 ;
      RECT 13.658 27.96 14.242 28.8 ;
      RECT 13.658 26.52 13.808 27.96 ;
      RECT 13.658 25.08 14.242 26.52 ;
      RECT 13.658 23.64 13.808 25.08 ;
      RECT 13.658 22.2 14.242 23.64 ;
      RECT 13.658 20.76 13.808 22.2 ;
      RECT 13.658 19.32 14.242 20.76 ;
      RECT 13.658 17.88 13.808 19.32 ;
      RECT 13.658 12.36 14.242 17.88 ;
      RECT 14.092 10.92 14.242 12.36 ;
      RECT 13.658 9.48 14.242 10.92 ;
      RECT 14.092 8.04 14.242 9.48 ;
      RECT 13.658 6.6 14.242 8.04 ;
      RECT 14.092 5.16 14.242 6.6 ;
      RECT 13.658 3.72 14.242 5.16 ;
      RECT 14.092 2.28 14.242 3.72 ;
      RECT 13.658 0 14.242 2.28 ;
      RECT 12.758 27.24 13.342 28.8 ;
      RECT 12.758 25.8 12.824 27.24 ;
      RECT 12.758 24.36 13.342 25.8 ;
      RECT 12.758 22.92 12.824 24.36 ;
      RECT 12.758 21.48 13.342 22.92 ;
      RECT 12.758 20.04 12.824 21.48 ;
      RECT 12.758 18.6 13.342 20.04 ;
      RECT 12.758 17.16 12.824 18.6 ;
      RECT 12.758 11.64 13.342 17.16 ;
      RECT 13.108 10.2 13.342 11.64 ;
      RECT 12.758 8.76 13.342 10.2 ;
      RECT 13.108 7.32 13.342 8.76 ;
      RECT 12.758 5.88 13.342 7.32 ;
      RECT 13.108 4.44 13.342 5.88 ;
      RECT 12.758 3 13.342 4.44 ;
      RECT 13.108 1.56 13.342 3 ;
      RECT 12.758 0 13.342 1.56 ;
      RECT 11.858 26.52 12.442 28.8 ;
      RECT 12.376 25.08 12.442 26.52 ;
      RECT 11.858 23.64 12.442 25.08 ;
      RECT 12.376 22.2 12.442 23.64 ;
      RECT 11.858 20.76 12.442 22.2 ;
      RECT 12.376 19.32 12.442 20.76 ;
      RECT 11.858 17.88 12.442 19.32 ;
      RECT 11.948 16.44 12.442 17.88 ;
      RECT 11.858 11.64 12.442 16.44 ;
      RECT 11.858 10.92 12.352 11.64 ;
      RECT 11.948 10.2 12.352 10.92 ;
      RECT 11.948 9.48 12.442 10.2 ;
      RECT 11.858 8.76 12.442 9.48 ;
      RECT 11.858 8.04 12.352 8.76 ;
      RECT 11.948 7.32 12.352 8.04 ;
      RECT 11.948 6.6 12.442 7.32 ;
      RECT 11.858 5.88 12.442 6.6 ;
      RECT 11.858 5.16 12.352 5.88 ;
      RECT 11.948 4.44 12.352 5.16 ;
      RECT 11.948 3.72 12.442 4.44 ;
      RECT 11.858 3 12.442 3.72 ;
      RECT 11.858 2.28 12.352 3 ;
      RECT 12.036 1.56 12.352 2.28 ;
      RECT 12.036 0.84 12.442 1.56 ;
      RECT 11.858 0 12.442 0.84 ;
      RECT 10.958 17.88 11.542 28.8 ;
      RECT 10.958 16.44 11.192 17.88 ;
      RECT 10.958 10.92 11.542 16.44 ;
      RECT 10.958 9.48 11.192 10.92 ;
      RECT 10.958 8.04 11.542 9.48 ;
      RECT 10.958 6.6 11.192 8.04 ;
      RECT 10.958 5.16 11.542 6.6 ;
      RECT 10.958 3.72 11.192 5.16 ;
      RECT 10.958 2.28 11.542 3.72 ;
      RECT 10.958 0.84 11.364 2.28 ;
      RECT 10.958 0 11.542 0.84 ;
      RECT 10.058 28.68 10.642 28.8 ;
      RECT 10.058 27.24 10.208 28.68 ;
      RECT 10.058 25.8 10.642 27.24 ;
      RECT 10.058 24.36 10.208 25.8 ;
      RECT 10.058 22.92 10.642 24.36 ;
      RECT 10.058 21.48 10.208 22.92 ;
      RECT 10.058 20.04 10.642 21.48 ;
      RECT 10.058 18.6 10.208 20.04 ;
      RECT 10.058 10.2 10.642 18.6 ;
      RECT 10.492 8.76 10.642 10.2 ;
      RECT 10.058 7.32 10.642 8.76 ;
      RECT 10.492 5.88 10.642 7.32 ;
      RECT 10.058 4.44 10.642 5.88 ;
      RECT 10.492 3 10.642 4.44 ;
      RECT 10.058 1.56 10.642 3 ;
      RECT 10.492 0.12 10.642 1.56 ;
      RECT 10.058 0 10.642 0.12 ;
      RECT 9.158 0 9.742 28.8 ;
      RECT 8.258 0 8.842 28.8 ;
      RECT 7.358 0 7.942 28.8 ;
      RECT 6.458 0 7.042 28.8 ;
      RECT 5.558 0 6.142 28.8 ;
      RECT 4.658 0 5.242 28.8 ;
      RECT 3.758 0 4.342 28.8 ;
      RECT 2.858 0 3.442 28.8 ;
      RECT 1.958 0 2.542 28.8 ;
      RECT 1.058 0 1.642 28.8 ;
      RECT 0.08 0 0.742 28.8 ;
      RECT 34.358 14.16 34.942 14.64 ;
      RECT 34.358 0 34.942 12.72 ;
    LAYER m0 ;
      RECT 0 0.002 70.2 28.798 ;
    LAYER m1 ;
      RECT 0 0 70.2 28.8 ;
    LAYER m2 ;
      RECT 0 0.015 70.2 28.785 ;
    LAYER m3 ;
      RECT 0.015 0 70.185 28.8 ;
    LAYER m4 ;
      RECT 0 0.02 70.2 28.78 ;
    LAYER m5 ;
      RECT 0.012 0 70.188 28.8 ;
    LAYER m6 ;
      RECT 0 0.012 70.2 28.788 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf124b192e1r1w0cbbehcaa4acw

END LIBRARY
