library ieee;
use ieee.std_logic_1164.all;
entity bogus_vhdl_module is 
port (bogus : in std_logic);
end bogus_vhdl_module;
architecture bogus_vhdl_module of bogus_vhdl_module is
begin
end bogus_vhdl_module;