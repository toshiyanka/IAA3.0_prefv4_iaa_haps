//----------------------------------------------------------------------
// ENUM DECLARATIONS
//------------------------------------------------------------------------
typedef enum int {
   IPLEVEL_STAP  =  'd0,
   NOTAP         =  'hFFFF_FFFF
} Tap_t;


