VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf074b064e1r1w0cbbehsaa4acw
  CLASS BLOCK ;
  FOREIGN arf074b064e1r1w0cbbehsaa4acw ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 32.64 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 16.68 3.172 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 14.76 0.728 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 16.68 0.472 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 16.68 0.728 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 16.68 0.816 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 16.68 1.028 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 16.68 1.116 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 16.68 1.372 17.88 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.68 3.516 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 16.68 3.728 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 16.68 3.816 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.68 4.072 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 14.76 1.716 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 14.76 1.928 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 14.76 2.016 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.76 2.616 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 14.76 2.828 15.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 14.76 2.916 15.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 14.76 0.816 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 14.76 1.028 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.24 1.928 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 3.84 1.928 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 3.84 2.272 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 4.56 2.916 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 4.56 2.016 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.28 2.616 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.28 2.828 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 6 2.272 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6 2.528 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 6.72 2.016 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 6.72 2.616 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 0.24 2.016 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 7.44 1.928 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 7.44 2.272 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 8.16 2.916 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 8.16 2.016 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 8.88 2.616 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 8.88 2.828 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 9.6 2.272 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 9.6 2.528 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 10.32 2.016 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 10.32 2.616 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.96 2.916 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 11.04 1.928 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 11.04 2.272 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 11.76 2.916 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 11.76 2.016 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 12.48 2.616 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12.48 2.828 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 13.2 2.272 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 13.2 2.528 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 18.24 2.916 19.44 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 18.24 1.928 19.44 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.96 2.272 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 18.96 2.272 20.16 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 18.96 2.528 20.16 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 19.68 1.928 20.88 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 19.68 2.016 20.88 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 20.4 2.916 21.6 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 20.4 2.272 21.6 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 21.12 2.616 22.32 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 21.12 2.828 22.32 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 21.84 2.272 23.04 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 21.84 2.528 23.04 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 1.68 2.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 22.56 2.016 23.76 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 22.56 2.616 23.76 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 23.28 1.928 24.48 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 23.28 2.272 24.48 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 24 2.916 25.2 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 24 2.016 25.2 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 24.72 2.616 25.92 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 24.72 2.828 25.92 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 25.44 2.272 26.64 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 25.44 2.528 26.64 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 1.68 2.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 26.16 2.016 27.36 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 26.16 2.616 27.36 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 26.88 1.928 28.08 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 26.88 2.272 28.08 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 27.6 2.916 28.8 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 27.6 2.016 28.8 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 28.32 2.616 29.52 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 28.32 2.828 29.52 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 29.04 2.272 30.24 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 29.04 2.528 30.24 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 2.4 2.272 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 29.76 2.016 30.96 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 29.76 2.616 30.96 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 30.48 1.928 31.68 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 30.48 2.272 31.68 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 31.2 2.916 32.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 31.2 2.016 32.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.4 2.528 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 3.12 2.016 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.12 2.616 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 14.76 1.372 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 14.76 1.628 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 14.76 1.116 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 0.24 3.516 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.84 3.516 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.84 3.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.56 3.428 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 4.56 3.816 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 5.28 3.172 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.28 3.516 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6 4.328 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6 3.428 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 6.72 3.816 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.72 4.072 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.24 3.728 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.44 3.516 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 7.44 3.728 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 8.16 3.428 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 8.16 3.816 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 8.88 3.172 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.88 3.516 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.6 4.328 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9.6 3.428 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 10.32 3.816 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 10.32 4.072 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.96 3.428 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.04 3.516 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 11.04 3.728 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 11.76 3.428 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 11.76 3.816 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 12.48 3.172 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.48 3.516 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 13.2 4.328 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 13.2 3.428 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 18.24 4.328 19.44 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 18.24 3.428 19.44 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 0.96 3.816 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 18.96 3.816 20.16 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 18.96 4.072 20.16 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.68 3.516 20.88 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 19.68 3.728 20.88 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.4 3.428 21.6 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 20.4 3.816 21.6 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 21.12 3.172 22.32 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 21.12 3.516 22.32 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 21.84 4.328 23.04 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 21.84 3.428 23.04 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 1.68 3.172 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 22.56 3.816 23.76 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 22.56 4.072 23.76 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 23.28 3.516 24.48 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 23.28 3.728 24.48 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 24 3.428 25.2 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 24 3.816 25.2 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 24.72 3.172 25.92 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 24.72 3.516 25.92 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 25.44 4.328 26.64 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 25.44 3.428 26.64 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 1.68 3.516 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 26.16 3.816 27.36 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 26.16 4.072 27.36 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 26.88 3.516 28.08 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 26.88 3.728 28.08 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 27.6 3.428 28.8 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 27.6 3.816 28.8 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 28.32 3.172 29.52 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 28.32 3.516 29.52 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 29.04 4.328 30.24 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 29.04 3.428 30.24 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 2.4 4.328 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 29.76 3.816 30.96 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 29.76 4.072 30.96 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 30.48 3.516 31.68 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 30.48 3.728 31.68 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 31.2 3.428 32.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 31.2 3.816 32.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.4 3.428 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 3.12 3.816 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 3.12 4.072 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 32.58 ;
        RECT 2.662 0.06 2.738 32.58 ;
        RECT 4.462 0.06 4.538 32.58 ;
        RECT 6.262 0.06 6.338 32.58 ;
        RECT 8.062 0.06 8.138 32.58 ;
        RECT 9.862 0.06 9.938 32.58 ;
        RECT 11.662 0.06 11.738 32.58 ;
        RECT 13.462 0.06 13.538 32.58 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 32.58 ;
        RECT 3.562 0.06 3.638 32.58 ;
        RECT 5.362 0.06 5.438 32.58 ;
        RECT 7.162 0.06 7.238 32.58 ;
        RECT 8.962 0.06 9.038 32.58 ;
        RECT 10.762 0.06 10.838 32.58 ;
        RECT 12.562 0.06 12.638 32.58 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 14.416 32.654 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 14.42 32.66 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 14.4705 32.678 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 14.435 32.71 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 14.47 32.678 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 14.459 32.73 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 14.49 32.702 ;
    LAYER m7 SPACING 0 ;
      RECT 13.538 32.7 14.44 32.76 ;
      RECT 13.538 -0.06 14.492 32.7 ;
      RECT 13.538 -0.12 14.44 -0.06 ;
      RECT 12.638 -0.12 13.462 32.76 ;
      RECT 11.738 -0.12 12.562 32.76 ;
      RECT 10.838 -0.12 11.662 32.76 ;
      RECT 9.938 -0.12 10.762 32.76 ;
      RECT 9.038 -0.12 9.862 32.76 ;
      RECT 8.138 -0.12 8.962 32.76 ;
      RECT 7.238 -0.12 8.062 32.76 ;
      RECT 6.338 -0.12 7.162 32.76 ;
      RECT 5.438 -0.12 6.262 32.76 ;
      RECT 4.538 -0.12 5.362 32.76 ;
      RECT 3.638 32.4 4.462 32.76 ;
      RECT 3.638 31.68 3.772 32.4 ;
      RECT 3.816 31.2 4.462 32.4 ;
      RECT 3.728 31.2 3.772 31.68 ;
      RECT 3.728 30.96 4.462 31.2 ;
      RECT 3.638 30.48 3.684 31.68 ;
      RECT 3.728 30.48 3.772 30.96 ;
      RECT 4.072 30.24 4.462 30.96 ;
      RECT 3.816 29.76 4.028 30.96 ;
      RECT 3.638 29.76 3.772 30.48 ;
      RECT 4.072 29.76 4.284 30.24 ;
      RECT 4.328 29.04 4.462 30.24 ;
      RECT 3.638 29.04 4.284 29.76 ;
      RECT 3.638 28.8 4.462 29.04 ;
      RECT 3.638 28.08 3.772 28.8 ;
      RECT 3.816 27.6 4.462 28.8 ;
      RECT 3.728 27.6 3.772 28.08 ;
      RECT 3.728 27.36 4.462 27.6 ;
      RECT 3.638 26.88 3.684 28.08 ;
      RECT 3.728 26.88 3.772 27.36 ;
      RECT 4.072 26.64 4.462 27.36 ;
      RECT 3.816 26.16 4.028 27.36 ;
      RECT 3.638 26.16 3.772 26.88 ;
      RECT 4.072 26.16 4.284 26.64 ;
      RECT 4.328 25.44 4.462 26.64 ;
      RECT 3.638 25.44 4.284 26.16 ;
      RECT 3.638 25.2 4.462 25.44 ;
      RECT 3.638 24.48 3.772 25.2 ;
      RECT 3.816 24 4.462 25.2 ;
      RECT 3.728 24 3.772 24.48 ;
      RECT 3.728 23.76 4.462 24 ;
      RECT 3.638 23.28 3.684 24.48 ;
      RECT 3.728 23.28 3.772 23.76 ;
      RECT 4.072 23.04 4.462 23.76 ;
      RECT 3.816 22.56 4.028 23.76 ;
      RECT 3.638 22.56 3.772 23.28 ;
      RECT 4.072 22.56 4.284 23.04 ;
      RECT 4.328 21.84 4.462 23.04 ;
      RECT 3.638 21.84 4.284 22.56 ;
      RECT 3.638 21.6 4.462 21.84 ;
      RECT 3.638 20.88 3.772 21.6 ;
      RECT 3.816 20.4 4.462 21.6 ;
      RECT 3.728 20.4 3.772 20.88 ;
      RECT 3.728 20.16 4.462 20.4 ;
      RECT 3.638 19.68 3.684 20.88 ;
      RECT 3.728 19.68 3.772 20.16 ;
      RECT 4.072 19.44 4.462 20.16 ;
      RECT 3.816 18.96 4.028 20.16 ;
      RECT 3.638 18.96 3.772 19.68 ;
      RECT 4.072 18.96 4.284 19.44 ;
      RECT 4.328 18.24 4.462 19.44 ;
      RECT 3.638 18.24 4.284 18.96 ;
      RECT 3.638 17.88 4.462 18.24 ;
      RECT 3.638 16.68 3.684 17.88 ;
      RECT 3.728 16.68 3.772 17.88 ;
      RECT 3.816 16.68 4.028 17.88 ;
      RECT 4.072 16.68 4.462 17.88 ;
      RECT 3.638 14.4 4.462 16.68 ;
      RECT 3.638 13.2 4.284 14.4 ;
      RECT 4.328 13.2 4.462 14.4 ;
      RECT 3.638 12.96 4.462 13.2 ;
      RECT 3.638 12.24 3.772 12.96 ;
      RECT 3.816 11.76 4.462 12.96 ;
      RECT 3.728 11.76 3.772 12.24 ;
      RECT 3.728 11.52 4.462 11.76 ;
      RECT 3.638 11.04 3.684 12.24 ;
      RECT 3.728 11.04 3.772 11.52 ;
      RECT 4.072 10.8 4.462 11.52 ;
      RECT 3.816 10.32 4.028 11.52 ;
      RECT 3.638 10.32 3.772 11.04 ;
      RECT 4.072 10.32 4.284 10.8 ;
      RECT 4.328 9.6 4.462 10.8 ;
      RECT 3.638 9.6 4.284 10.32 ;
      RECT 3.638 9.36 4.462 9.6 ;
      RECT 3.638 8.64 3.772 9.36 ;
      RECT 3.816 8.16 4.462 9.36 ;
      RECT 3.728 8.16 3.772 8.64 ;
      RECT 3.728 7.92 4.462 8.16 ;
      RECT 3.638 7.44 3.684 8.64 ;
      RECT 3.728 7.44 3.772 7.92 ;
      RECT 4.072 7.2 4.462 7.92 ;
      RECT 3.816 6.72 4.028 7.92 ;
      RECT 3.638 6.72 3.772 7.44 ;
      RECT 4.072 6.72 4.284 7.2 ;
      RECT 4.328 6 4.462 7.2 ;
      RECT 3.638 6 4.284 6.72 ;
      RECT 3.638 5.76 4.462 6 ;
      RECT 3.638 5.04 3.772 5.76 ;
      RECT 3.816 4.56 4.462 5.76 ;
      RECT 3.728 4.56 3.772 5.04 ;
      RECT 3.728 4.32 4.462 4.56 ;
      RECT 3.638 3.84 3.684 5.04 ;
      RECT 3.728 3.84 3.772 4.32 ;
      RECT 4.072 3.6 4.462 4.32 ;
      RECT 3.816 3.12 4.028 4.32 ;
      RECT 3.638 3.12 3.772 3.84 ;
      RECT 4.072 3.12 4.284 3.6 ;
      RECT 4.328 2.4 4.462 3.6 ;
      RECT 3.638 2.4 4.284 3.12 ;
      RECT 3.638 2.16 4.462 2.4 ;
      RECT 3.638 1.44 3.772 2.16 ;
      RECT 3.816 0.96 4.462 2.16 ;
      RECT 3.728 0.96 3.772 1.44 ;
      RECT 3.638 0.24 3.684 1.44 ;
      RECT 3.728 0.24 4.462 0.96 ;
      RECT 3.638 -0.12 4.462 0.24 ;
      RECT 2.738 32.4 3.562 32.76 ;
      RECT 3.428 31.68 3.562 32.4 ;
      RECT 2.738 31.2 2.872 32.4 ;
      RECT 2.916 31.2 3.384 32.4 ;
      RECT 3.428 31.2 3.472 31.68 ;
      RECT 3.516 30.48 3.562 31.68 ;
      RECT 2.738 30.48 3.472 31.2 ;
      RECT 2.738 30.24 3.562 30.48 ;
      RECT 2.738 29.52 3.384 30.24 ;
      RECT 3.428 29.52 3.562 30.24 ;
      RECT 3.172 29.04 3.384 29.52 ;
      RECT 3.428 29.04 3.472 29.52 ;
      RECT 2.828 28.8 3.128 29.52 ;
      RECT 3.172 28.8 3.472 29.04 ;
      RECT 2.738 28.32 2.784 29.52 ;
      RECT 3.516 28.32 3.562 29.52 ;
      RECT 2.828 28.32 2.872 28.8 ;
      RECT 2.916 28.32 3.128 28.8 ;
      RECT 3.172 28.32 3.384 28.8 ;
      RECT 3.428 28.32 3.472 28.8 ;
      RECT 3.428 28.08 3.562 28.32 ;
      RECT 2.738 27.6 2.872 28.32 ;
      RECT 2.916 27.6 3.384 28.32 ;
      RECT 3.428 27.6 3.472 28.08 ;
      RECT 3.516 26.88 3.562 28.08 ;
      RECT 2.738 26.88 3.472 27.6 ;
      RECT 2.738 26.64 3.562 26.88 ;
      RECT 2.738 25.92 3.384 26.64 ;
      RECT 3.428 25.92 3.562 26.64 ;
      RECT 3.172 25.44 3.384 25.92 ;
      RECT 3.428 25.44 3.472 25.92 ;
      RECT 2.828 25.2 3.128 25.92 ;
      RECT 3.172 25.2 3.472 25.44 ;
      RECT 2.738 24.72 2.784 25.92 ;
      RECT 3.516 24.72 3.562 25.92 ;
      RECT 2.828 24.72 2.872 25.2 ;
      RECT 2.916 24.72 3.128 25.2 ;
      RECT 3.172 24.72 3.384 25.2 ;
      RECT 3.428 24.72 3.472 25.2 ;
      RECT 3.428 24.48 3.562 24.72 ;
      RECT 2.738 24 2.872 24.72 ;
      RECT 2.916 24 3.384 24.72 ;
      RECT 3.428 24 3.472 24.48 ;
      RECT 3.516 23.28 3.562 24.48 ;
      RECT 2.738 23.28 3.472 24 ;
      RECT 2.738 23.04 3.562 23.28 ;
      RECT 2.738 22.32 3.384 23.04 ;
      RECT 3.428 22.32 3.562 23.04 ;
      RECT 3.172 21.84 3.384 22.32 ;
      RECT 3.428 21.84 3.472 22.32 ;
      RECT 2.828 21.6 3.128 22.32 ;
      RECT 3.172 21.6 3.472 21.84 ;
      RECT 2.738 21.12 2.784 22.32 ;
      RECT 3.516 21.12 3.562 22.32 ;
      RECT 2.828 21.12 2.872 21.6 ;
      RECT 2.916 21.12 3.128 21.6 ;
      RECT 3.172 21.12 3.384 21.6 ;
      RECT 3.428 21.12 3.472 21.6 ;
      RECT 3.428 20.88 3.562 21.12 ;
      RECT 2.738 20.4 2.872 21.12 ;
      RECT 2.916 20.4 3.384 21.12 ;
      RECT 3.428 20.4 3.472 20.88 ;
      RECT 3.516 19.68 3.562 20.88 ;
      RECT 2.738 19.68 3.472 20.4 ;
      RECT 2.738 19.44 3.562 19.68 ;
      RECT 2.738 18.24 2.872 19.44 ;
      RECT 2.916 18.24 3.384 19.44 ;
      RECT 3.428 18.24 3.562 19.44 ;
      RECT 2.738 17.88 3.562 18.24 ;
      RECT 2.738 16.68 3.128 17.88 ;
      RECT 3.172 16.68 3.472 17.88 ;
      RECT 3.516 16.68 3.562 17.88 ;
      RECT 2.738 15.96 3.562 16.68 ;
      RECT 2.738 14.76 2.784 15.96 ;
      RECT 2.828 14.76 2.872 15.96 ;
      RECT 2.916 14.76 3.562 15.96 ;
      RECT 2.738 14.4 3.562 14.76 ;
      RECT 2.738 13.68 3.384 14.4 ;
      RECT 3.428 13.68 3.562 14.4 ;
      RECT 3.172 13.2 3.384 13.68 ;
      RECT 3.428 13.2 3.472 13.68 ;
      RECT 2.828 12.96 3.128 13.68 ;
      RECT 3.172 12.96 3.472 13.2 ;
      RECT 2.738 12.48 2.784 13.68 ;
      RECT 3.516 12.48 3.562 13.68 ;
      RECT 2.828 12.48 2.872 12.96 ;
      RECT 2.916 12.48 3.128 12.96 ;
      RECT 3.172 12.48 3.384 12.96 ;
      RECT 3.428 12.48 3.472 12.96 ;
      RECT 3.428 12.24 3.562 12.48 ;
      RECT 2.738 11.76 2.872 12.48 ;
      RECT 2.916 11.76 3.384 12.48 ;
      RECT 3.428 11.76 3.472 12.24 ;
      RECT 3.516 11.04 3.562 12.24 ;
      RECT 2.738 11.04 3.472 11.76 ;
      RECT 2.738 10.8 3.562 11.04 ;
      RECT 2.738 10.08 3.384 10.8 ;
      RECT 3.428 10.08 3.562 10.8 ;
      RECT 3.172 9.6 3.384 10.08 ;
      RECT 3.428 9.6 3.472 10.08 ;
      RECT 2.828 9.36 3.128 10.08 ;
      RECT 3.172 9.36 3.472 9.6 ;
      RECT 2.738 8.88 2.784 10.08 ;
      RECT 3.516 8.88 3.562 10.08 ;
      RECT 2.828 8.88 2.872 9.36 ;
      RECT 2.916 8.88 3.128 9.36 ;
      RECT 3.172 8.88 3.384 9.36 ;
      RECT 3.428 8.88 3.472 9.36 ;
      RECT 3.428 8.64 3.562 8.88 ;
      RECT 2.738 8.16 2.872 8.88 ;
      RECT 2.916 8.16 3.384 8.88 ;
      RECT 3.428 8.16 3.472 8.64 ;
      RECT 3.516 7.44 3.562 8.64 ;
      RECT 2.738 7.44 3.472 8.16 ;
      RECT 2.738 7.2 3.562 7.44 ;
      RECT 2.738 6.48 3.384 7.2 ;
      RECT 3.428 6.48 3.562 7.2 ;
      RECT 3.172 6 3.384 6.48 ;
      RECT 3.428 6 3.472 6.48 ;
      RECT 2.828 5.76 3.128 6.48 ;
      RECT 3.172 5.76 3.472 6 ;
      RECT 2.738 5.28 2.784 6.48 ;
      RECT 3.516 5.28 3.562 6.48 ;
      RECT 2.828 5.28 2.872 5.76 ;
      RECT 2.916 5.28 3.128 5.76 ;
      RECT 3.172 5.28 3.384 5.76 ;
      RECT 3.428 5.28 3.472 5.76 ;
      RECT 3.428 5.04 3.562 5.28 ;
      RECT 2.738 4.56 2.872 5.28 ;
      RECT 2.916 4.56 3.384 5.28 ;
      RECT 3.428 4.56 3.472 5.04 ;
      RECT 3.516 3.84 3.562 5.04 ;
      RECT 2.738 3.84 3.472 4.56 ;
      RECT 2.738 3.6 3.562 3.84 ;
      RECT 2.738 2.88 3.384 3.6 ;
      RECT 3.428 2.88 3.562 3.6 ;
      RECT 3.172 2.4 3.384 2.88 ;
      RECT 3.428 2.4 3.472 2.88 ;
      RECT 2.828 2.16 3.128 2.88 ;
      RECT 3.172 2.16 3.472 2.4 ;
      RECT 2.738 1.68 2.784 2.88 ;
      RECT 3.516 1.68 3.562 2.88 ;
      RECT 2.828 1.68 2.872 2.16 ;
      RECT 2.916 1.68 3.128 2.16 ;
      RECT 3.172 1.68 3.384 2.16 ;
      RECT 3.428 1.68 3.472 2.16 ;
      RECT 3.428 1.44 3.562 1.68 ;
      RECT 2.738 0.96 2.872 1.68 ;
      RECT 2.916 0.96 3.384 1.68 ;
      RECT 3.428 0.96 3.472 1.44 ;
      RECT 3.516 0.24 3.562 1.44 ;
      RECT 2.738 0.24 3.472 0.96 ;
      RECT 2.738 -0.12 3.562 0.24 ;
      RECT 1.838 32.4 2.662 32.76 ;
      RECT 1.838 31.68 1.972 32.4 ;
      RECT 2.016 31.68 2.662 32.4 ;
      RECT 1.928 31.2 1.972 31.68 ;
      RECT 2.016 31.2 2.228 31.68 ;
      RECT 2.272 30.96 2.662 31.68 ;
      RECT 1.928 30.96 2.228 31.2 ;
      RECT 1.838 30.48 1.884 31.68 ;
      RECT 1.928 30.48 1.972 30.96 ;
      RECT 2.016 30.48 2.228 30.96 ;
      RECT 2.272 30.48 2.572 30.96 ;
      RECT 2.016 30.24 2.572 30.48 ;
      RECT 2.616 29.76 2.662 30.96 ;
      RECT 1.838 29.76 1.972 30.48 ;
      RECT 2.016 29.76 2.228 30.24 ;
      RECT 2.528 29.76 2.572 30.24 ;
      RECT 2.528 29.52 2.662 29.76 ;
      RECT 2.272 29.04 2.484 30.24 ;
      RECT 1.838 29.04 2.228 29.76 ;
      RECT 2.528 29.04 2.572 29.52 ;
      RECT 1.838 28.8 2.572 29.04 ;
      RECT 2.616 28.32 2.662 29.52 ;
      RECT 2.016 28.32 2.572 28.8 ;
      RECT 1.838 28.08 1.972 28.8 ;
      RECT 2.016 28.08 2.662 28.32 ;
      RECT 1.928 27.6 1.972 28.08 ;
      RECT 2.016 27.6 2.228 28.08 ;
      RECT 2.272 27.36 2.662 28.08 ;
      RECT 1.928 27.36 2.228 27.6 ;
      RECT 1.838 26.88 1.884 28.08 ;
      RECT 1.928 26.88 1.972 27.36 ;
      RECT 2.016 26.88 2.228 27.36 ;
      RECT 2.272 26.88 2.572 27.36 ;
      RECT 2.016 26.64 2.572 26.88 ;
      RECT 2.616 26.16 2.662 27.36 ;
      RECT 1.838 26.16 1.972 26.88 ;
      RECT 2.016 26.16 2.228 26.64 ;
      RECT 2.528 26.16 2.572 26.64 ;
      RECT 2.528 25.92 2.662 26.16 ;
      RECT 2.272 25.44 2.484 26.64 ;
      RECT 1.838 25.44 2.228 26.16 ;
      RECT 2.528 25.44 2.572 25.92 ;
      RECT 1.838 25.2 2.572 25.44 ;
      RECT 2.616 24.72 2.662 25.92 ;
      RECT 2.016 24.72 2.572 25.2 ;
      RECT 1.838 24.48 1.972 25.2 ;
      RECT 2.016 24.48 2.662 24.72 ;
      RECT 1.928 24 1.972 24.48 ;
      RECT 2.016 24 2.228 24.48 ;
      RECT 2.272 23.76 2.662 24.48 ;
      RECT 1.928 23.76 2.228 24 ;
      RECT 1.838 23.28 1.884 24.48 ;
      RECT 1.928 23.28 1.972 23.76 ;
      RECT 2.016 23.28 2.228 23.76 ;
      RECT 2.272 23.28 2.572 23.76 ;
      RECT 2.016 23.04 2.572 23.28 ;
      RECT 2.616 22.56 2.662 23.76 ;
      RECT 1.838 22.56 1.972 23.28 ;
      RECT 2.016 22.56 2.228 23.04 ;
      RECT 2.528 22.56 2.572 23.04 ;
      RECT 2.528 22.32 2.662 22.56 ;
      RECT 2.272 21.84 2.484 23.04 ;
      RECT 1.838 21.84 2.228 22.56 ;
      RECT 2.528 21.84 2.572 22.32 ;
      RECT 1.838 21.6 2.572 21.84 ;
      RECT 2.616 21.12 2.662 22.32 ;
      RECT 2.272 21.12 2.572 21.6 ;
      RECT 1.838 20.88 2.228 21.6 ;
      RECT 2.272 20.4 2.662 21.12 ;
      RECT 2.016 20.4 2.228 20.88 ;
      RECT 2.016 20.16 2.662 20.4 ;
      RECT 1.838 19.68 1.884 20.88 ;
      RECT 1.928 19.68 1.972 20.88 ;
      RECT 2.016 19.68 2.228 20.16 ;
      RECT 1.838 19.44 2.228 19.68 ;
      RECT 2.272 18.96 2.484 20.16 ;
      RECT 2.528 18.96 2.662 20.16 ;
      RECT 1.928 18.96 2.228 19.44 ;
      RECT 1.838 18.24 1.884 19.44 ;
      RECT 1.928 18.24 2.662 18.96 ;
      RECT 1.838 15.96 2.662 18.24 ;
      RECT 1.838 14.76 1.884 15.96 ;
      RECT 1.928 14.76 1.972 15.96 ;
      RECT 2.016 14.76 2.572 15.96 ;
      RECT 2.616 14.76 2.662 15.96 ;
      RECT 1.838 14.4 2.662 14.76 ;
      RECT 2.528 13.68 2.662 14.4 ;
      RECT 1.838 13.2 2.228 14.4 ;
      RECT 2.272 13.2 2.484 14.4 ;
      RECT 2.528 13.2 2.572 13.68 ;
      RECT 1.838 12.96 2.572 13.2 ;
      RECT 2.616 12.48 2.662 13.68 ;
      RECT 2.016 12.48 2.572 12.96 ;
      RECT 1.838 12.24 1.972 12.96 ;
      RECT 2.016 12.24 2.662 12.48 ;
      RECT 1.928 11.76 1.972 12.24 ;
      RECT 2.016 11.76 2.228 12.24 ;
      RECT 2.272 11.52 2.662 12.24 ;
      RECT 1.928 11.52 2.228 11.76 ;
      RECT 1.838 11.04 1.884 12.24 ;
      RECT 1.928 11.04 1.972 11.52 ;
      RECT 2.016 11.04 2.228 11.52 ;
      RECT 2.272 11.04 2.572 11.52 ;
      RECT 2.016 10.8 2.572 11.04 ;
      RECT 2.616 10.32 2.662 11.52 ;
      RECT 1.838 10.32 1.972 11.04 ;
      RECT 2.016 10.32 2.228 10.8 ;
      RECT 2.528 10.32 2.572 10.8 ;
      RECT 2.528 10.08 2.662 10.32 ;
      RECT 2.272 9.6 2.484 10.8 ;
      RECT 1.838 9.6 2.228 10.32 ;
      RECT 2.528 9.6 2.572 10.08 ;
      RECT 1.838 9.36 2.572 9.6 ;
      RECT 2.616 8.88 2.662 10.08 ;
      RECT 2.016 8.88 2.572 9.36 ;
      RECT 1.838 8.64 1.972 9.36 ;
      RECT 2.016 8.64 2.662 8.88 ;
      RECT 1.928 8.16 1.972 8.64 ;
      RECT 2.016 8.16 2.228 8.64 ;
      RECT 2.272 7.92 2.662 8.64 ;
      RECT 1.928 7.92 2.228 8.16 ;
      RECT 1.838 7.44 1.884 8.64 ;
      RECT 1.928 7.44 1.972 7.92 ;
      RECT 2.016 7.44 2.228 7.92 ;
      RECT 2.272 7.44 2.572 7.92 ;
      RECT 2.016 7.2 2.572 7.44 ;
      RECT 2.616 6.72 2.662 7.92 ;
      RECT 1.838 6.72 1.972 7.44 ;
      RECT 2.016 6.72 2.228 7.2 ;
      RECT 2.528 6.72 2.572 7.2 ;
      RECT 2.528 6.48 2.662 6.72 ;
      RECT 2.272 6 2.484 7.2 ;
      RECT 1.838 6 2.228 6.72 ;
      RECT 2.528 6 2.572 6.48 ;
      RECT 1.838 5.76 2.572 6 ;
      RECT 2.616 5.28 2.662 6.48 ;
      RECT 2.016 5.28 2.572 5.76 ;
      RECT 1.838 5.04 1.972 5.76 ;
      RECT 2.016 5.04 2.662 5.28 ;
      RECT 1.928 4.56 1.972 5.04 ;
      RECT 2.016 4.56 2.228 5.04 ;
      RECT 2.272 4.32 2.662 5.04 ;
      RECT 1.928 4.32 2.228 4.56 ;
      RECT 1.838 3.84 1.884 5.04 ;
      RECT 1.928 3.84 1.972 4.32 ;
      RECT 2.016 3.84 2.228 4.32 ;
      RECT 2.272 3.84 2.572 4.32 ;
      RECT 2.016 3.6 2.572 3.84 ;
      RECT 2.616 3.12 2.662 4.32 ;
      RECT 1.838 3.12 1.972 3.84 ;
      RECT 2.016 3.12 2.228 3.6 ;
      RECT 2.528 3.12 2.572 3.6 ;
      RECT 2.528 2.88 2.662 3.12 ;
      RECT 2.272 2.4 2.484 3.6 ;
      RECT 1.838 2.4 2.228 3.12 ;
      RECT 2.528 2.4 2.572 2.88 ;
      RECT 1.838 2.16 2.572 2.4 ;
      RECT 2.616 1.68 2.662 2.88 ;
      RECT 2.272 1.68 2.572 2.16 ;
      RECT 1.838 1.44 2.228 2.16 ;
      RECT 2.272 0.96 2.662 1.68 ;
      RECT 2.016 0.96 2.228 1.44 ;
      RECT 1.838 0.24 1.884 1.44 ;
      RECT 1.928 0.24 1.972 1.44 ;
      RECT 2.016 0.24 2.662 0.96 ;
      RECT 1.838 -0.12 2.662 0.24 ;
      RECT 0.938 17.88 1.762 32.76 ;
      RECT 0.938 16.68 0.984 17.88 ;
      RECT 1.028 16.68 1.072 17.88 ;
      RECT 1.116 16.68 1.328 17.88 ;
      RECT 1.372 16.68 1.762 17.88 ;
      RECT 0.938 15.96 1.762 16.68 ;
      RECT 0.938 14.76 0.984 15.96 ;
      RECT 1.028 14.76 1.072 15.96 ;
      RECT 1.116 14.76 1.328 15.96 ;
      RECT 1.372 14.76 1.584 15.96 ;
      RECT 1.628 14.76 1.672 15.96 ;
      RECT 1.716 14.76 1.762 15.96 ;
      RECT 0.938 -0.12 1.762 14.76 ;
      RECT -0.04 32.7 0.862 32.76 ;
      RECT -0.092 17.88 0.862 32.7 ;
      RECT -0.092 16.68 0.428 17.88 ;
      RECT 0.472 16.68 0.684 17.88 ;
      RECT 0.728 16.68 0.772 17.88 ;
      RECT 0.816 16.68 0.862 17.88 ;
      RECT -0.092 15.96 0.862 16.68 ;
      RECT -0.092 14.76 0.684 15.96 ;
      RECT 0.728 14.76 0.772 15.96 ;
      RECT 0.816 14.76 0.862 15.96 ;
      RECT -0.092 -0.06 0.862 14.76 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 13.658 0 14.32 32.64 ;
      RECT 12.758 0 13.342 32.64 ;
      RECT 11.858 0 12.442 32.64 ;
      RECT 10.958 0 11.542 32.64 ;
      RECT 10.058 0 10.642 32.64 ;
      RECT 9.158 0 9.742 32.64 ;
      RECT 8.258 0 8.842 32.64 ;
      RECT 7.358 0 7.942 32.64 ;
      RECT 6.458 0 7.042 32.64 ;
      RECT 5.558 0 6.142 32.64 ;
      RECT 4.658 0 5.242 32.64 ;
      RECT 3.758 32.52 4.342 32.64 ;
      RECT 3.936 31.08 4.342 32.52 ;
      RECT 4.192 30.36 4.342 31.08 ;
      RECT 2.858 32.52 3.442 32.64 ;
      RECT 3.036 31.08 3.264 32.52 ;
      RECT 2.858 30.36 3.352 31.08 ;
      RECT 2.858 29.64 3.264 30.36 ;
      RECT 2.948 28.92 3.008 29.64 ;
      RECT 1.958 32.52 2.542 32.64 ;
      RECT 2.136 31.8 2.542 32.52 ;
      RECT 2.392 31.08 2.542 31.8 ;
      RECT 2.392 30.36 2.452 31.08 ;
      RECT 1.058 18 1.642 32.64 ;
      RECT 1.492 16.56 1.642 18 ;
      RECT 1.058 16.08 1.642 16.56 ;
      RECT 0.08 18 0.742 32.64 ;
      RECT 0.08 16.56 0.308 18 ;
      RECT 0.08 16.08 0.742 16.56 ;
      RECT 0.08 14.64 0.564 16.08 ;
      RECT 0.08 0 0.742 14.64 ;
      RECT 3.758 28.92 4.164 29.64 ;
      RECT 3.936 27.48 4.342 28.92 ;
      RECT 4.192 26.76 4.342 27.48 ;
      RECT 1.958 28.92 2.108 29.64 ;
      RECT 2.136 28.2 2.452 28.92 ;
      RECT 2.392 27.48 2.542 28.2 ;
      RECT 2.392 26.76 2.452 27.48 ;
      RECT 3.036 27.48 3.264 28.2 ;
      RECT 2.858 26.76 3.352 27.48 ;
      RECT 2.858 26.04 3.264 26.76 ;
      RECT 2.948 25.32 3.008 26.04 ;
      RECT 3.758 25.32 4.164 26.04 ;
      RECT 3.936 23.88 4.342 25.32 ;
      RECT 4.192 23.16 4.342 23.88 ;
      RECT 1.958 25.32 2.108 26.04 ;
      RECT 2.136 24.6 2.452 25.32 ;
      RECT 2.392 23.88 2.542 24.6 ;
      RECT 2.392 23.16 2.452 23.88 ;
      RECT 3.036 23.88 3.264 24.6 ;
      RECT 2.858 23.16 3.352 23.88 ;
      RECT 2.858 22.44 3.264 23.16 ;
      RECT 2.948 21.72 3.008 22.44 ;
      RECT 3.758 21.72 4.164 22.44 ;
      RECT 3.936 20.28 4.342 21.72 ;
      RECT 4.192 19.56 4.342 20.28 ;
      RECT 1.958 21 2.108 22.44 ;
      RECT 2.392 21 2.452 21.72 ;
      RECT 2.392 20.28 2.542 21 ;
      RECT 3.036 20.28 3.264 21 ;
      RECT 2.858 19.56 3.352 20.28 ;
      RECT 3.036 18.12 3.264 19.56 ;
      RECT 2.858 18 3.442 18.12 ;
      RECT 2.858 16.56 3.008 18 ;
      RECT 3.292 16.56 3.352 18 ;
      RECT 2.858 16.08 3.442 16.56 ;
      RECT 3.036 14.64 3.442 16.08 ;
      RECT 2.858 14.52 3.442 14.64 ;
      RECT 2.858 13.8 3.264 14.52 ;
      RECT 2.948 13.08 3.008 13.8 ;
      RECT 2.048 18.84 2.108 19.56 ;
      RECT 2.048 18.12 2.542 18.84 ;
      RECT 1.958 16.08 2.542 18.12 ;
      RECT 2.136 14.64 2.452 16.08 ;
      RECT 1.958 14.52 2.542 14.64 ;
      RECT 1.958 13.08 2.108 14.52 ;
      RECT 3.758 18.12 4.164 18.84 ;
      RECT 3.758 18 4.342 18.12 ;
      RECT 4.192 16.56 4.342 18 ;
      RECT 3.758 14.52 4.342 16.56 ;
      RECT 3.758 13.08 4.164 14.52 ;
      RECT 3.936 11.64 4.342 13.08 ;
      RECT 4.192 10.92 4.342 11.64 ;
      RECT 1.058 0 1.642 14.64 ;
      RECT 2.136 12.36 2.452 13.08 ;
      RECT 2.392 11.64 2.542 12.36 ;
      RECT 2.392 10.92 2.452 11.64 ;
      RECT 3.036 11.64 3.264 12.36 ;
      RECT 2.858 10.92 3.352 11.64 ;
      RECT 2.858 10.2 3.264 10.92 ;
      RECT 2.948 9.48 3.008 10.2 ;
      RECT 3.758 9.48 4.164 10.2 ;
      RECT 3.936 8.04 4.342 9.48 ;
      RECT 4.192 7.32 4.342 8.04 ;
      RECT 1.958 9.48 2.108 10.2 ;
      RECT 2.136 8.76 2.452 9.48 ;
      RECT 2.392 8.04 2.542 8.76 ;
      RECT 2.392 7.32 2.452 8.04 ;
      RECT 3.036 8.04 3.264 8.76 ;
      RECT 2.858 7.32 3.352 8.04 ;
      RECT 2.858 6.6 3.264 7.32 ;
      RECT 2.948 5.88 3.008 6.6 ;
      RECT 3.758 5.88 4.164 6.6 ;
      RECT 3.936 4.44 4.342 5.88 ;
      RECT 4.192 3.72 4.342 4.44 ;
      RECT 1.958 5.88 2.108 6.6 ;
      RECT 2.136 5.16 2.452 5.88 ;
      RECT 2.392 4.44 2.542 5.16 ;
      RECT 2.392 3.72 2.452 4.44 ;
      RECT 3.036 4.44 3.264 5.16 ;
      RECT 2.858 3.72 3.352 4.44 ;
      RECT 2.858 3 3.264 3.72 ;
      RECT 2.948 2.28 3.008 3 ;
      RECT 3.758 2.28 4.164 3 ;
      RECT 3.936 0.84 4.342 2.28 ;
      RECT 3.848 0.12 4.342 0.84 ;
      RECT 3.758 0 4.342 0.12 ;
      RECT 1.958 1.56 2.108 3 ;
      RECT 2.392 1.56 2.452 2.28 ;
      RECT 2.392 0.84 2.542 1.56 ;
      RECT 2.136 0.12 2.542 0.84 ;
      RECT 1.958 0 2.542 0.12 ;
      RECT 3.036 0.84 3.264 1.56 ;
      RECT 2.858 0.12 3.352 0.84 ;
      RECT 2.858 0 3.442 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 14.4 32.638 ;
    LAYER m1 ;
      RECT 0 0 14.4 32.64 ;
    LAYER m2 ;
      RECT 0 0.015 14.4 32.625 ;
    LAYER m3 ;
      RECT 0.015 0 14.385 32.64 ;
    LAYER m4 ;
      RECT 0 0.02 14.4 32.62 ;
    LAYER m5 ;
      RECT 0.012 0 14.388 32.64 ;
    LAYER m6 ;
      RECT 0 0.012 14.4 32.628 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf074b064e1r1w0cbbehsaa4acw

END LIBRARY
