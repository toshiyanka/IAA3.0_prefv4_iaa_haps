package sip_vintf_pkg;

endpackage;
