VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf030b256e1r1w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf030b256e1r1w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 43.2 BY 17.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.484 9 23.528 10.2 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 7.08 20.916 8.28 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 9 18.816 10.2 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 9 19.028 10.2 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 9 19.116 10.2 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 9 19.372 10.2 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 9 19.628 10.2 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 9 19.716 10.2 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 9 19.928 10.2 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 9 20.016 10.2 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 9 23.616 10.2 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 9 23.872 10.2 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 9 18.472 10.2 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 9 18.728 10.2 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 7.08 22.072 8.28 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 7.08 22.328 8.28 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 7.08 22.416 8.28 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 7.08 22.628 8.28 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 7.08 22.716 8.28 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 7.08 22.972 8.28 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 7.08 23.228 8.28 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 7.08 23.316 8.28 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 7.08 21.172 8.28 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 7.08 21.428 8.28 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 3.84 22.716 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 3.84 22.972 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 4.56 19.116 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 4.56 19.372 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 5.28 20.272 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 5.28 20.528 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 10.8 22.072 12 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 10.8 22.328 12 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 11.52 20.916 12.72 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 11.52 21.172 12.72 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 12.24 22.416 13.44 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 12.24 22.628 13.44 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 12.96 18.472 14.16 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 12.96 18.728 14.16 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 13.68 19.928 14.88 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 13.68 20.016 14.88 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 14.4 20.616 15.6 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 14.4 20.828 15.6 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 15.12 21.428 16.32 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 15.12 21.516 16.32 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 0.96 19.928 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 15.84 22.072 17.04 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 15.84 22.328 17.04 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 0.96 20.016 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.68 20.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 1.68 20.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 2.4 21.428 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 2.4 21.516 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 3.12 22.072 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 3.12 22.328 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 7.08 21.728 8.28 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 7.08 21.816 8.28 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 7.08 21.516 8.28 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 3.84 18.472 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 3.84 18.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 4.56 19.628 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 4.56 19.716 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 5.28 20.616 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 5.28 20.828 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 10.8 22.416 12 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 10.8 22.628 12 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 11.52 21.428 12.72 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 11.52 21.516 12.72 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 12.24 22.716 13.44 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 12.24 22.972 13.44 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 12.96 18.816 14.16 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 12.96 19.028 14.16 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 13.68 20.272 14.88 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 13.68 20.528 14.88 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 14.4 20.916 15.6 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 14.4 21.172 15.6 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 15.12 21.728 16.32 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 15.12 21.816 16.32 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 0.96 20.272 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 15.84 22.416 17.04 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 15.84 22.628 17.04 ;
    END
  END rddatap0[31]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 0.96 20.528 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 1.68 20.916 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 1.68 21.172 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 2.4 21.728 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.4 21.816 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 3.12 22.416 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 3.12 22.628 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 17.22 ;
        RECT 2.662 0.06 2.738 17.22 ;
        RECT 4.462 0.06 4.538 17.22 ;
        RECT 6.262 0.06 6.338 17.22 ;
        RECT 8.062 0.06 8.138 17.22 ;
        RECT 9.862 0.06 9.938 17.22 ;
        RECT 11.662 0.06 11.738 17.22 ;
        RECT 13.462 0.06 13.538 17.22 ;
        RECT 15.262 0.06 15.338 17.22 ;
        RECT 17.062 0.06 17.138 17.22 ;
        RECT 18.862 0.06 18.938 17.22 ;
        RECT 20.662 0.06 20.738 17.22 ;
        RECT 22.462 0.06 22.538 17.22 ;
        RECT 24.262 0.06 24.338 17.22 ;
        RECT 26.062 0.06 26.138 17.22 ;
        RECT 27.862 0.06 27.938 17.22 ;
        RECT 29.662 0.06 29.738 17.22 ;
        RECT 31.462 0.06 31.538 17.22 ;
        RECT 33.262 0.06 33.338 17.22 ;
        RECT 35.062 0.06 35.138 17.22 ;
        RECT 36.862 0.06 36.938 17.22 ;
        RECT 38.662 0.06 38.738 17.22 ;
        RECT 40.462 0.06 40.538 17.22 ;
        RECT 42.262 0.06 42.338 17.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 17.22 ;
        RECT 3.562 0.06 3.638 17.22 ;
        RECT 5.362 0.06 5.438 17.22 ;
        RECT 7.162 0.06 7.238 17.22 ;
        RECT 8.962 0.06 9.038 17.22 ;
        RECT 10.762 0.06 10.838 17.22 ;
        RECT 12.562 0.06 12.638 17.22 ;
        RECT 14.362 0.06 14.438 17.22 ;
        RECT 16.162 0.06 16.238 17.22 ;
        RECT 17.962 0.06 18.038 17.22 ;
        RECT 19.762 0.06 19.838 17.22 ;
        RECT 21.562 0.06 21.638 17.22 ;
        RECT 23.362 0.06 23.438 17.22 ;
        RECT 25.162 0.06 25.238 17.22 ;
        RECT 26.962 0.06 27.038 17.22 ;
        RECT 28.762 0.06 28.838 17.22 ;
        RECT 30.562 0.06 30.638 17.22 ;
        RECT 32.362 0.06 32.438 17.22 ;
        RECT 34.162 0.06 34.238 17.22 ;
        RECT 35.962 0.06 36.038 17.22 ;
        RECT 37.762 0.06 37.838 17.22 ;
        RECT 39.562 0.06 39.638 17.22 ;
        RECT 41.362 0.06 41.438 17.22 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 43.216 17.294 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 43.22 17.3 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 43.2705 17.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 43.235 17.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 43.27 17.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 43.259 17.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 43.29 17.342 ;
    LAYER m7 SPACING 0 ;
      RECT 42.338 17.34 43.24 17.4 ;
      RECT 42.338 -0.06 43.292 17.34 ;
      RECT 42.338 -0.12 43.24 -0.06 ;
      RECT 41.438 -0.12 42.262 17.4 ;
      RECT 40.538 -0.12 41.362 17.4 ;
      RECT 39.638 -0.12 40.462 17.4 ;
      RECT 38.738 -0.12 39.562 17.4 ;
      RECT 37.838 -0.12 38.662 17.4 ;
      RECT 36.938 -0.12 37.762 17.4 ;
      RECT 36.038 -0.12 36.862 17.4 ;
      RECT 35.138 -0.12 35.962 17.4 ;
      RECT 34.238 -0.12 35.062 17.4 ;
      RECT 33.338 -0.12 34.162 17.4 ;
      RECT 32.438 -0.12 33.262 17.4 ;
      RECT 31.538 -0.12 32.362 17.4 ;
      RECT 30.638 -0.12 31.462 17.4 ;
      RECT 29.738 -0.12 30.562 17.4 ;
      RECT 28.838 -0.12 29.662 17.4 ;
      RECT 27.938 -0.12 28.762 17.4 ;
      RECT 27.038 -0.12 27.862 17.4 ;
      RECT 26.138 -0.12 26.962 17.4 ;
      RECT 25.238 -0.12 26.062 17.4 ;
      RECT 24.338 -0.12 25.162 17.4 ;
      RECT 23.438 10.2 24.262 17.4 ;
      RECT 23.438 9 23.484 10.2 ;
      RECT 23.528 9 23.572 10.2 ;
      RECT 23.616 9 23.828 10.2 ;
      RECT 23.872 9 24.262 10.2 ;
      RECT 23.438 -0.12 24.262 9 ;
      RECT 22.538 17.04 23.362 17.4 ;
      RECT 22.538 15.84 22.584 17.04 ;
      RECT 22.628 15.84 23.362 17.04 ;
      RECT 22.538 13.44 23.362 15.84 ;
      RECT 22.538 12.24 22.584 13.44 ;
      RECT 22.628 12.24 22.672 13.44 ;
      RECT 22.716 12.24 22.928 13.44 ;
      RECT 22.972 12.24 23.362 13.44 ;
      RECT 22.538 12 23.362 12.24 ;
      RECT 22.538 10.8 22.584 12 ;
      RECT 22.628 10.8 23.362 12 ;
      RECT 22.538 8.28 23.362 10.8 ;
      RECT 22.538 7.08 22.584 8.28 ;
      RECT 22.628 7.08 22.672 8.28 ;
      RECT 22.716 7.08 22.928 8.28 ;
      RECT 22.972 7.08 23.184 8.28 ;
      RECT 23.228 7.08 23.272 8.28 ;
      RECT 23.316 7.08 23.362 8.28 ;
      RECT 22.538 5.04 23.362 7.08 ;
      RECT 22.538 4.32 22.672 5.04 ;
      RECT 22.716 3.84 22.928 5.04 ;
      RECT 22.972 3.84 23.362 5.04 ;
      RECT 22.628 3.84 22.672 4.32 ;
      RECT 22.538 3.12 22.584 4.32 ;
      RECT 22.628 3.12 23.362 3.84 ;
      RECT 22.538 -0.12 23.362 3.12 ;
      RECT 21.638 17.04 22.462 17.4 ;
      RECT 21.638 16.32 22.028 17.04 ;
      RECT 22.072 15.84 22.284 17.04 ;
      RECT 22.328 15.84 22.372 17.04 ;
      RECT 22.416 15.84 22.462 17.04 ;
      RECT 21.816 15.84 22.028 16.32 ;
      RECT 21.638 15.12 21.684 16.32 ;
      RECT 21.728 15.12 21.772 16.32 ;
      RECT 21.816 15.12 22.462 15.84 ;
      RECT 21.638 13.44 22.462 15.12 ;
      RECT 21.638 12.24 22.372 13.44 ;
      RECT 22.416 12.24 22.462 13.44 ;
      RECT 21.638 12 22.462 12.24 ;
      RECT 21.638 10.8 22.028 12 ;
      RECT 22.072 10.8 22.284 12 ;
      RECT 22.328 10.8 22.372 12 ;
      RECT 22.416 10.8 22.462 12 ;
      RECT 21.638 8.28 22.462 10.8 ;
      RECT 21.638 7.08 21.684 8.28 ;
      RECT 21.728 7.08 21.772 8.28 ;
      RECT 21.816 7.08 22.028 8.28 ;
      RECT 22.072 7.08 22.284 8.28 ;
      RECT 22.328 7.08 22.372 8.28 ;
      RECT 22.416 7.08 22.462 8.28 ;
      RECT 21.638 4.32 22.462 7.08 ;
      RECT 21.638 3.6 22.028 4.32 ;
      RECT 22.072 3.12 22.284 4.32 ;
      RECT 22.328 3.12 22.372 4.32 ;
      RECT 22.416 3.12 22.462 4.32 ;
      RECT 21.816 3.12 22.028 3.6 ;
      RECT 21.638 2.4 21.684 3.6 ;
      RECT 21.728 2.4 21.772 3.6 ;
      RECT 21.816 2.4 22.462 3.12 ;
      RECT 21.638 -0.12 22.462 2.4 ;
      RECT 20.738 16.32 21.562 17.4 ;
      RECT 20.738 15.6 21.384 16.32 ;
      RECT 21.428 15.12 21.472 16.32 ;
      RECT 21.516 15.12 21.562 16.32 ;
      RECT 21.172 15.12 21.384 15.6 ;
      RECT 20.738 14.4 20.784 15.6 ;
      RECT 20.828 14.4 20.872 15.6 ;
      RECT 20.916 14.4 21.128 15.6 ;
      RECT 21.172 14.4 21.562 15.12 ;
      RECT 20.738 12.72 21.562 14.4 ;
      RECT 20.738 11.52 20.872 12.72 ;
      RECT 20.916 11.52 21.128 12.72 ;
      RECT 21.172 11.52 21.384 12.72 ;
      RECT 21.428 11.52 21.472 12.72 ;
      RECT 21.516 11.52 21.562 12.72 ;
      RECT 20.738 8.28 21.562 11.52 ;
      RECT 20.738 7.08 20.872 8.28 ;
      RECT 20.916 7.08 21.128 8.28 ;
      RECT 21.172 7.08 21.384 8.28 ;
      RECT 21.428 7.08 21.472 8.28 ;
      RECT 21.516 7.08 21.562 8.28 ;
      RECT 20.738 6.48 21.562 7.08 ;
      RECT 20.738 5.28 20.784 6.48 ;
      RECT 20.828 5.28 21.562 6.48 ;
      RECT 20.738 3.6 21.562 5.28 ;
      RECT 20.738 2.88 21.384 3.6 ;
      RECT 21.428 2.4 21.472 3.6 ;
      RECT 21.516 2.4 21.562 3.6 ;
      RECT 21.172 2.4 21.384 2.88 ;
      RECT 20.738 1.68 20.784 2.88 ;
      RECT 20.828 1.68 20.872 2.88 ;
      RECT 20.916 1.68 21.128 2.88 ;
      RECT 21.172 1.68 21.562 2.4 ;
      RECT 20.738 -0.12 21.562 1.68 ;
      RECT 19.838 15.6 20.662 17.4 ;
      RECT 19.838 14.88 20.572 15.6 ;
      RECT 20.616 14.4 20.662 15.6 ;
      RECT 20.528 14.4 20.572 14.88 ;
      RECT 19.838 13.68 19.884 14.88 ;
      RECT 19.928 13.68 19.972 14.88 ;
      RECT 20.016 13.68 20.228 14.88 ;
      RECT 20.272 13.68 20.484 14.88 ;
      RECT 20.528 13.68 20.662 14.4 ;
      RECT 19.838 10.2 20.662 13.68 ;
      RECT 19.838 9 19.884 10.2 ;
      RECT 19.928 9 19.972 10.2 ;
      RECT 20.016 9 20.662 10.2 ;
      RECT 19.838 6.48 20.662 9 ;
      RECT 19.838 5.28 20.228 6.48 ;
      RECT 20.272 5.28 20.484 6.48 ;
      RECT 20.528 5.28 20.572 6.48 ;
      RECT 20.616 5.28 20.662 6.48 ;
      RECT 19.838 2.88 20.662 5.28 ;
      RECT 19.838 2.16 20.572 2.88 ;
      RECT 20.616 1.68 20.662 2.88 ;
      RECT 20.528 1.68 20.572 2.16 ;
      RECT 19.838 0.96 19.884 2.16 ;
      RECT 19.928 0.96 19.972 2.16 ;
      RECT 20.016 0.96 20.228 2.16 ;
      RECT 20.272 0.96 20.484 2.16 ;
      RECT 20.528 0.96 20.662 1.68 ;
      RECT 19.838 -0.12 20.662 0.96 ;
      RECT 18.938 14.16 19.762 17.4 ;
      RECT 18.938 12.96 18.984 14.16 ;
      RECT 19.028 12.96 19.762 14.16 ;
      RECT 18.938 10.2 19.762 12.96 ;
      RECT 18.938 9 18.984 10.2 ;
      RECT 19.028 9 19.072 10.2 ;
      RECT 19.116 9 19.328 10.2 ;
      RECT 19.372 9 19.584 10.2 ;
      RECT 19.628 9 19.672 10.2 ;
      RECT 19.716 9 19.762 10.2 ;
      RECT 18.938 5.76 19.762 9 ;
      RECT 18.938 4.56 19.072 5.76 ;
      RECT 19.116 4.56 19.328 5.76 ;
      RECT 19.372 4.56 19.584 5.76 ;
      RECT 19.628 4.56 19.672 5.76 ;
      RECT 19.716 4.56 19.762 5.76 ;
      RECT 18.938 1.44 19.762 4.56 ;
      RECT 18.938 0.24 18.984 1.44 ;
      RECT 19.028 0.24 19.762 1.44 ;
      RECT 18.938 -0.12 19.762 0.24 ;
      RECT 18.038 14.16 18.862 17.4 ;
      RECT 18.038 12.96 18.428 14.16 ;
      RECT 18.472 12.96 18.684 14.16 ;
      RECT 18.728 12.96 18.772 14.16 ;
      RECT 18.816 12.96 18.862 14.16 ;
      RECT 18.038 10.2 18.862 12.96 ;
      RECT 18.038 9 18.428 10.2 ;
      RECT 18.472 9 18.684 10.2 ;
      RECT 18.728 9 18.772 10.2 ;
      RECT 18.816 9 18.862 10.2 ;
      RECT 18.038 5.04 18.862 9 ;
      RECT 18.038 3.84 18.428 5.04 ;
      RECT 18.472 3.84 18.684 5.04 ;
      RECT 18.728 3.84 18.862 5.04 ;
      RECT 18.038 1.44 18.862 3.84 ;
      RECT 18.038 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.772 1.44 ;
      RECT 18.816 0.24 18.862 1.44 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 17.4 ;
      RECT 16.238 -0.12 17.062 17.4 ;
      RECT 15.338 -0.12 16.162 17.4 ;
      RECT 14.438 -0.12 15.262 17.4 ;
      RECT 13.538 -0.12 14.362 17.4 ;
      RECT 12.638 -0.12 13.462 17.4 ;
      RECT 11.738 -0.12 12.562 17.4 ;
      RECT 10.838 -0.12 11.662 17.4 ;
      RECT 9.938 -0.12 10.762 17.4 ;
      RECT 9.038 -0.12 9.862 17.4 ;
      RECT 8.138 -0.12 8.962 17.4 ;
      RECT 7.238 -0.12 8.062 17.4 ;
      RECT 6.338 -0.12 7.162 17.4 ;
      RECT 5.438 -0.12 6.262 17.4 ;
      RECT 4.538 -0.12 5.362 17.4 ;
      RECT 3.638 -0.12 4.462 17.4 ;
      RECT 2.738 -0.12 3.562 17.4 ;
      RECT 1.838 -0.12 2.662 17.4 ;
      RECT 0.938 -0.12 1.762 17.4 ;
      RECT -0.04 17.34 0.862 17.4 ;
      RECT -0.092 -0.06 0.862 17.34 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 42.458 0 43.12 17.28 ;
      RECT 41.558 0 42.142 17.28 ;
      RECT 40.658 0 41.242 17.28 ;
      RECT 39.758 0 40.342 17.28 ;
      RECT 38.858 0 39.442 17.28 ;
      RECT 37.958 0 38.542 17.28 ;
      RECT 37.058 0 37.642 17.28 ;
      RECT 36.158 0 36.742 17.28 ;
      RECT 35.258 0 35.842 17.28 ;
      RECT 34.358 0 34.942 17.28 ;
      RECT 33.458 0 34.042 17.28 ;
      RECT 32.558 0 33.142 17.28 ;
      RECT 31.658 0 32.242 17.28 ;
      RECT 30.758 0 31.342 17.28 ;
      RECT 29.858 0 30.442 17.28 ;
      RECT 28.958 0 29.542 17.28 ;
      RECT 28.058 0 28.642 17.28 ;
      RECT 27.158 0 27.742 17.28 ;
      RECT 26.258 0 26.842 17.28 ;
      RECT 25.358 0 25.942 17.28 ;
      RECT 24.458 0 25.042 17.28 ;
      RECT 23.558 10.32 24.142 17.28 ;
      RECT 23.992 8.88 24.142 10.32 ;
      RECT 23.558 0 24.142 8.88 ;
      RECT 22.658 17.16 23.242 17.28 ;
      RECT 22.748 15.72 23.242 17.16 ;
      RECT 22.658 13.56 23.242 15.72 ;
      RECT 23.092 12.12 23.242 13.56 ;
      RECT 22.748 10.68 23.242 12.12 ;
      RECT 22.658 8.4 23.242 10.68 ;
      RECT 21.758 17.16 22.342 17.28 ;
      RECT 21.758 16.44 21.908 17.16 ;
      RECT 20.858 16.44 21.442 17.28 ;
      RECT 20.858 15.72 21.264 16.44 ;
      RECT 19.958 15.72 20.542 17.28 ;
      RECT 19.958 15 20.452 15.72 ;
      RECT 19.058 14.28 19.642 17.28 ;
      RECT 19.148 12.84 19.642 14.28 ;
      RECT 19.058 10.32 19.642 12.84 ;
      RECT 18.158 14.28 18.742 17.28 ;
      RECT 18.158 12.84 18.308 14.28 ;
      RECT 18.158 10.32 18.742 12.84 ;
      RECT 18.158 8.88 18.308 10.32 ;
      RECT 18.158 5.16 18.742 8.88 ;
      RECT 18.158 3.72 18.308 5.16 ;
      RECT 18.158 1.56 18.742 3.72 ;
      RECT 18.158 0.12 18.308 1.56 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 17.28 ;
      RECT 16.358 0 16.942 17.28 ;
      RECT 15.458 0 16.042 17.28 ;
      RECT 14.558 0 15.142 17.28 ;
      RECT 13.658 0 14.242 17.28 ;
      RECT 12.758 0 13.342 17.28 ;
      RECT 11.858 0 12.442 17.28 ;
      RECT 10.958 0 11.542 17.28 ;
      RECT 10.058 0 10.642 17.28 ;
      RECT 9.158 0 9.742 17.28 ;
      RECT 8.258 0 8.842 17.28 ;
      RECT 7.358 0 7.942 17.28 ;
      RECT 6.458 0 7.042 17.28 ;
      RECT 5.558 0 6.142 17.28 ;
      RECT 4.658 0 5.242 17.28 ;
      RECT 3.758 0 4.342 17.28 ;
      RECT 2.858 0 3.442 17.28 ;
      RECT 1.958 0 2.542 17.28 ;
      RECT 1.058 0 1.642 17.28 ;
      RECT 0.08 0 0.742 17.28 ;
      RECT 21.936 15 22.342 15.72 ;
      RECT 21.758 13.56 22.342 15 ;
      RECT 21.758 12.12 22.252 13.56 ;
      RECT 21.758 10.68 21.908 12.12 ;
      RECT 21.758 8.4 22.342 10.68 ;
      RECT 21.292 14.28 21.442 15 ;
      RECT 20.858 12.84 21.442 14.28 ;
      RECT 19.958 10.32 20.542 13.56 ;
      RECT 20.136 8.88 20.542 10.32 ;
      RECT 19.958 6.6 20.542 8.88 ;
      RECT 19.958 5.16 20.108 6.6 ;
      RECT 19.958 3 20.542 5.16 ;
      RECT 19.958 2.28 20.452 3 ;
      RECT 20.858 8.4 21.442 11.4 ;
      RECT 19.058 5.88 19.642 8.88 ;
      RECT 22.658 5.16 23.242 6.96 ;
      RECT 23.092 3.72 23.242 5.16 ;
      RECT 22.748 3 23.242 3.72 ;
      RECT 22.658 0 23.242 3 ;
      RECT 21.758 4.44 22.342 6.96 ;
      RECT 21.758 3.72 21.908 4.44 ;
      RECT 20.858 6.6 21.442 6.96 ;
      RECT 20.948 5.16 21.442 6.6 ;
      RECT 20.858 3.72 21.442 5.16 ;
      RECT 20.858 3 21.264 3.72 ;
      RECT 19.058 1.56 19.642 4.44 ;
      RECT 19.148 0.12 19.642 1.56 ;
      RECT 19.058 0 19.642 0.12 ;
      RECT 21.936 2.28 22.342 3 ;
      RECT 21.758 0 22.342 2.28 ;
      RECT 21.292 1.56 21.442 2.28 ;
      RECT 20.858 0 21.442 1.56 ;
      RECT 19.958 0 20.542 0.84 ;
    LAYER m0 ;
      RECT 0 0.002 43.2 17.278 ;
    LAYER m1 ;
      RECT 0 0 43.2 17.28 ;
    LAYER m2 ;
      RECT 0 0.015 43.2 17.265 ;
    LAYER m3 ;
      RECT 0.015 0 43.185 17.28 ;
    LAYER m4 ;
      RECT 0 0.02 43.2 17.26 ;
    LAYER m5 ;
      RECT 0.012 0 43.188 17.28 ;
    LAYER m6 ;
      RECT 0 0.012 43.2 17.268 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf030b256e1r1w0cbbeheaa4acw

END LIBRARY
