
//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2015 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
//-- Test
//-----------------------------------------------------------------------------------------------------
`ifndef VERIF_DOMAIN_BASE_TEST
`define VERIF_DOMAIN_BASE_TEST hqm_base_test;
`endif

import hqm_tb_cfg_sequences_pkg::*;

//-------------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------------
class hqm_visa_test extends `VERIF_DOMAIN_BASE_TEST;
   
  `ovm_component_utils(hqm_visa_test)

  function new(string name = "hqm_visa_test", ovm_component parent = null);
    super.new(name,parent);
  endfunction : new

  virtual function void build();
     super.build();
  endfunction : build
  

  virtual function void connect();
    super.connect();
    if ($test$plusargs("VISA_SKIP_INIT")) begin
        i_hqm_tb_env.skip_test_phase("PCIE_CONFIG_PHASE");
    end
       // i_hqm_tb_env.skip_test_phase("CONFIG_PHASE");
        i_hqm_tb_env.skip_test_phase("PCIE_FLUSH_PHASE");
        i_hqm_tb_env.skip_test_phase("FLUSH_PHASE");

        i_hqm_tb_env.set_test_phase_type("i_hqm_tb_env","CONFIG_PHASE","hqm_tb_cfg_file_mode_seq");

    if ($test$plusargs("VISA_SECURITY_TEST")) 
        i_hqm_tb_env.set_test_phase_type("i_hqm_tb_env", "USER_DATA_PHASE", "hqm_visa_security_seq"); 
    else
        i_hqm_tb_env.set_test_phase_type("i_hqm_tb_env", "USER_DATA_PHASE", "hqm_visa_seq"); 
  endfunction // void

   task run();
     ovm_report_info("hqm_visa_test", "hqm_visa_test run is executing\!");
   endtask

endclass : hqm_visa_test 
