VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf028b256e2r2w0cbbeheaa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf028b256e2r2w0cbbeheaa4acw 0 0 ;
  SIZE 81 BY 22.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 12.12 35.828 13.32 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 12.12 40.156 13.32 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 9.24 35.828 10.44 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 9.24 40.416 10.44 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 12.12 38.188 13.32 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 12.12 38.356 13.32 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 12.12 38.616 13.32 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 12.12 38.916 13.32 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 12.12 39.172 13.32 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 12.12 39.428 13.32 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 12.12 39.728 13.32 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 12.12 39.988 13.32 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.072 12.12 37.116 13.32 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.328 12.12 37.372 13.32 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 12.12 41.528 13.32 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 12.12 41.788 13.32 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 12.12 41.956 13.32 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 12.12 42.216 13.32 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 12.12 42.516 13.32 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 12.12 42.772 13.32 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 12.12 43.028 13.32 ;
    END
  END rdaddrp1[6]
  PIN rdaddrp1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 12.12 43.328 13.32 ;
    END
  END rdaddrp1[7]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 12.12 40.416 13.32 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 12.12 40.716 13.32 ;
    END
  END rdaddrp1_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 0.36 36.388 1.56 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 5.16 42.516 6.36 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.644 5.16 42.688 6.36 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 6.12 43.588 7.32 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 6.12 43.672 7.32 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 7.08 36.472 8.28 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 7.08 36.556 8.28 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 14.28 36.556 15.48 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 14.28 36.728 15.48 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.484 15.24 38.528 16.44 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 15.24 38.616 16.44 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 0.36 36.472 1.56 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 16.2 39.516 17.4 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 16.2 39.728 17.4 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.584 17.16 40.628 18.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 17.16 40.716 18.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.572 18.12 41.616 19.32 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 18.12 41.788 19.32 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.644 19.08 42.688 20.28 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 19.08 42.772 20.28 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.628 20.04 43.672 21.24 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 20.04 43.756 21.24 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 1.32 38.356 2.52 ;
    END
  END rddatap0[2]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.484 1.32 38.528 2.52 ;
    END
  END rddatap0[3]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 2.28 39.428 3.48 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.472 2.28 39.516 3.48 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 3.24 40.416 4.44 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.584 3.24 40.628 4.44 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 4.2 41.528 5.4 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.572 4.2 41.616 5.4 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.512 0.36 36.556 1.56 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 5.16 42.772 6.36 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.812 5.16 42.856 6.36 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 6.12 43.756 7.32 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.884 6.12 43.928 7.32 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 7.08 36.728 8.28 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.772 7.08 36.816 8.28 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.772 14.28 36.816 15.48 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.984 14.28 37.028 15.48 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 15.24 38.828 16.44 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 15.24 38.916 16.44 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.684 0.36 36.728 1.56 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 16.2 39.816 17.4 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 16.2 39.988 17.4 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.844 17.16 40.888 18.36 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 17.16 40.972 18.36 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.828 18.12 41.872 19.32 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 18.12 41.956 19.32 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.812 19.08 42.856 20.28 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 19.08 43.028 20.28 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.884 20.04 43.928 21.24 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 20.04 35.916 21.24 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 1.32 38.616 2.52 ;
    END
  END rddatap1[2]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.784 1.32 38.828 2.52 ;
    END
  END rddatap1[3]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 2.28 39.728 3.48 ;
    END
  END rddatap1[4]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.772 2.28 39.816 3.48 ;
    END
  END rddatap1[5]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 3.24 40.716 4.44 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.844 3.24 40.888 4.44 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 4.2 41.788 5.4 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.828 4.2 41.872 5.4 ;
    END
  END rddatap1[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.584 12.12 37.628 13.32 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 12.12 40.972 13.32 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 12.12 37.928 13.32 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 12.12 41.228 13.32 ;
    END
  END sdl_initp1
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 80.062 0.06 80.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 78.262 0.06 78.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 76.462 0.06 76.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 74.662 0.06 74.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 72.862 0.06 72.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 71.062 0.06 71.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 69.262 0.06 69.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 67.462 0.06 67.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 65.662 0.06 65.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 63.862 0.06 63.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 62.062 0.06 62.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 60.262 0.06 60.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 58.462 0.06 58.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 56.662 0.06 56.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 54.862 0.06 54.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 53.062 0.06 53.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 51.262 0.06 51.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 49.462 0.06 49.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 47.662 0.06 47.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 45.862 0.06 45.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 44.062 0.06 44.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 42.262 0.06 42.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 40.462 0.06 40.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 38.662 0.06 38.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 36.862 0.06 36.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.062 0.06 35.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 33.262 0.06 33.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.462 0.06 31.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.662 0.06 29.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 27.862 0.06 27.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.062 0.06 26.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.262 0.06 24.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 22.462 0.06 22.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.662 0.06 20.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.862 0.06 18.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.062 0.06 17.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.262 0.06 15.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 22.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 79.162 0.06 79.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 77.362 0.06 77.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 75.562 0.06 75.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 73.762 0.06 73.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 71.962 0.06 72.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 70.162 0.06 70.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 68.362 0.06 68.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 66.562 0.06 66.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 64.762 0.06 64.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 62.962 0.06 63.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 61.162 0.06 61.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 59.362 0.06 59.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 57.562 0.06 57.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 55.762 0.06 55.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 53.962 0.06 54.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 52.162 0.06 52.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 50.362 0.06 50.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 48.562 0.06 48.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 46.762 0.06 46.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 44.962 0.06 45.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 43.162 0.06 43.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 41.362 0.06 41.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 39.562 0.06 39.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 37.762 0.06 37.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.962 0.06 36.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 34.162 0.06 34.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 32.362 0.06 32.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.562 0.06 30.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 28.762 0.06 28.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.962 0.06 27.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.162 0.06 25.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.362 0.06 23.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 21.562 0.06 21.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 19.762 0.06 19.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.962 0.06 18.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 16.162 0.06 16.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.362 0.06 14.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 22.02 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 9.24 38.356 10.44 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.572 9.24 38.616 10.44 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 9.24 38.916 10.44 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 9.24 39.172 10.44 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 9.24 39.428 10.44 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.684 9.24 39.728 10.44 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 9.24 39.988 10.44 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 9.24 40.156 10.44 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.072 9.24 37.116 10.44 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.328 9.24 37.372 10.44 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 9.24 41.956 10.44 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 9.24 42.216 10.44 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 9.24 42.516 10.44 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.728 9.24 42.772 10.44 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 9.24 43.028 10.44 ;
    END
  END wraddrp1[4]
  PIN wraddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 9.24 43.328 10.44 ;
    END
  END wraddrp1[5]
  PIN wraddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 9.24 43.588 10.44 ;
    END
  END wraddrp1[6]
  PIN wraddrp1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.712 9.24 43.756 10.44 ;
    END
  END wraddrp1[7]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.672 9.24 40.716 10.44 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 9.24 40.972 10.44 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.784 0.36 35.828 1.56 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.912 5.16 41.956 6.36 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 5.16 42.128 6.36 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.984 6.12 43.028 7.32 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 6.12 43.116 7.32 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 7.08 35.916 8.28 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 7.08 36.128 8.28 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 14.28 36.128 15.48 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 14.28 36.216 15.48 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.972 15.24 38.016 16.44 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 15.24 38.188 16.44 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.872 0.36 35.916 1.56 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 16.2 39.088 17.4 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 16.2 39.172 17.4 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.028 17.16 40.072 18.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 17.16 40.156 18.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.012 18.12 41.056 19.32 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 18.12 41.228 19.32 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.084 19.08 42.128 20.28 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 19.08 42.216 20.28 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.072 20.04 43.116 21.24 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 20.04 43.328 21.24 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 1.32 37.928 2.52 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.972 1.32 38.016 2.52 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.872 2.28 38.916 3.48 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.044 2.28 39.088 3.48 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.944 3.24 39.988 4.44 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.028 3.24 40.072 4.44 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.928 4.2 40.972 5.4 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.012 4.2 41.056 5.4 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.884 9.24 37.928 10.44 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 9.24 38.188 10.44 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.084 0.36 36.128 1.56 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.172 5.16 42.216 6.36 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 5.16 42.428 6.36 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.284 6.12 43.328 7.32 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 6.12 43.416 7.32 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 7.08 36.216 8.28 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 7.08 36.388 8.28 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.344 14.28 36.388 15.48 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.428 14.28 36.472 15.48 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.228 15.24 38.272 16.44 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.312 15.24 38.356 16.44 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 36.172 0.36 36.216 1.56 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 16.2 39.256 17.4 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.384 16.2 39.428 17.4 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 17.16 40.328 18.36 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.372 17.16 40.416 18.36 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.272 18.12 41.316 19.32 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 18.12 41.528 19.32 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.384 19.08 42.428 20.28 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 42.472 19.08 42.516 20.28 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.372 20.04 43.416 21.24 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 43.544 20.04 43.588 21.24 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.144 1.32 38.188 2.52 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 38.228 1.32 38.272 2.52 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.128 2.28 39.172 3.48 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 39.212 2.28 39.256 3.48 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.112 3.24 40.156 4.44 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 40.284 3.24 40.328 4.44 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 4.2 41.228 5.4 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.272 4.2 41.316 5.4 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.484 9.24 41.528 10.44 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.744 9.24 41.788 10.44 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.584 9.24 37.628 10.44 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 41.184 9.24 41.228 10.44 ;
    END
  END wrenp1
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 81 22.08 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 81 22.08 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 81.0705 22.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 81.035 22.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 81.07 22.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 81.059 22.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 81.09 22.142 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 81.092 22.14 ;
  END
END arf028b256e2r2w0cbbeheaa4acw
END LIBRARY
