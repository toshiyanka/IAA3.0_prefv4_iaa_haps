//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr_c : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr_c
(
  // Synchronous Clock/Reset
  clk_100,
  rst_b_100,

  // Asynchronous Clock/Reset(s)
  clk_200,

  // Power Well Isolation Input Signals
  island0_pok,
  island2_pok,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  p3_fab_init_idle_exit,
  p3_fab_init_idle_exit_ack,
  p4_fab_init_idle_exit,
  p4_fab_init_idle_exit_ack,
  p5_fab_init_idle_exit,
  p5_fab_init_idle_exit_ack,
  p6_fab_init_idle_exit,
  p6_fab_init_idle_exit_ack,
  p7_fab_init_idle_exit,
  p7_fab_init_idle_exit_ack,
  p8_fab_init_idle_exit,
  p8_fab_init_idle_exit_ack,
  p9_fab_init_idle_exit,
  p9_fab_init_idle_exit_ack,
  p10_fab_init_idle_exit,
  p10_fab_init_idle_exit_ack,
  p11_fab_init_idle_exit,
  p11_fab_init_idle_exit_ack,
  p12_fab_init_idle_exit,
  p12_fab_init_idle_exit_ack,
  p13_fab_init_idle_exit,
  p13_fab_init_idle_exit_ack,
  p14_fab_init_idle_exit,
  p14_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_clk_100,
  visa_vp_clk_100,
  visa_p0_tier1_clk_100,
  visa_p0_tier2_clk_100,
  visa_p1_tier1_clk_100,
  visa_p1_tier2_clk_100,
  visa_p2_tier1_clk_200,
  visa_p2_tier2_clk_200,
  visa_p2_ififo_tier1_clk_100,
  visa_p2_ififo_tier2_clk_100,
  visa_p2_efifo_tier1_clk_100,
  visa_p2_efifo_tier2_clk_100,
  visa_p3_tier1_clk_200,
  visa_p3_tier2_clk_200,
  visa_p3_ififo_tier1_clk_100,
  visa_p3_ififo_tier2_clk_100,
  visa_p3_efifo_tier1_clk_100,
  visa_p3_efifo_tier2_clk_100,
  visa_p4_tier1_clk_200,
  visa_p4_tier2_clk_200,
  visa_p4_ififo_tier1_clk_100,
  visa_p4_ififo_tier2_clk_100,
  visa_p4_efifo_tier1_clk_100,
  visa_p4_efifo_tier2_clk_100,
  visa_p5_tier1_clk_200,
  visa_p5_tier2_clk_200,
  visa_p5_ififo_tier1_clk_100,
  visa_p5_ififo_tier2_clk_100,
  visa_p5_efifo_tier1_clk_100,
  visa_p5_efifo_tier2_clk_100,
  visa_p6_tier1_clk_100,
  visa_p6_tier2_clk_100,
  visa_p7_tier1_clk_100,
  visa_p7_tier2_clk_100,
  visa_p8_tier1_clk_100,
  visa_p8_tier2_clk_100,
  visa_p9_tier1_clk_100,
  visa_p9_tier2_clk_100,
  visa_p10_tier1_clk_100,
  visa_p10_tier2_clk_100,
  visa_p11_tier1_clk_100,
  visa_p11_tier2_clk_100,
  visa_p12_tier1_clk_200,
  visa_p12_tier2_clk_200,
  visa_p12_ififo_tier1_clk_100,
  visa_p12_ififo_tier2_clk_100,
  visa_p12_efifo_tier1_clk_100,
  visa_p12_efifo_tier2_clk_100,
  visa_p13_tier1_clk_100,
  visa_p13_tier2_clk_100,
  visa_p14_tier1_clk_100,
  visa_p14_tier2_clk_100,


  // Register wires
  cfg_sbr_c_cgovrd,
  cfg_sbr_c_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  sbr_a_sbr_c_side_ism_agent,
  sbr_c_sbr_a_side_ism_fabric,
  sbr_a_sbr_c_pccup,
  sbr_a_sbr_c_npcup,
  sbr_c_sbr_a_pcput,
  sbr_c_sbr_a_npput,
  sbr_c_sbr_a_eom,
  sbr_c_sbr_a_payload,
  sbr_c_sbr_a_pccup,
  sbr_c_sbr_a_npcup,
  sbr_a_sbr_c_pcput,
  sbr_a_sbr_c_npput,
  sbr_a_sbr_c_eom,
  sbr_a_sbr_c_payload,

  // Port 1 declarations
  sbr_d_sbr_c_side_ism_fabric,
  sbr_c_sbr_d_side_ism_agent,
  sbr_d_sbr_c_pccup,
  sbr_d_sbr_c_npcup,
  sbr_c_sbr_d_pcput,
  sbr_c_sbr_d_npput,
  sbr_c_sbr_d_eom,
  sbr_c_sbr_d_payload,
  sbr_c_sbr_d_pccup,
  sbr_c_sbr_d_npcup,
  sbr_d_sbr_c_pcput,
  sbr_d_sbr_c_npput,
  sbr_d_sbr_c_eom,
  sbr_d_sbr_c_payload,

  // Port 2 declarations
  vtunit_sbr_c_side_ism_agent,
  sbr_c_vtunit_side_ism_fabric,
  vtunit_sbr_c_pccup,
  vtunit_sbr_c_npcup,
  sbr_c_vtunit_pcput,
  sbr_c_vtunit_npput,
  sbr_c_vtunit_eom,
  sbr_c_vtunit_payload,
  sbr_c_vtunit_pccup,
  sbr_c_vtunit_npcup,
  vtunit_sbr_c_pcput,
  vtunit_sbr_c_npput,
  vtunit_sbr_c_eom,
  vtunit_sbr_c_payload,

  // Port 3 declarations
  hunit_sbr_c_side_ism_agent,
  sbr_c_hunit_side_ism_fabric,
  hunit_sbr_c_pccup,
  hunit_sbr_c_npcup,
  sbr_c_hunit_pcput,
  sbr_c_hunit_npput,
  sbr_c_hunit_eom,
  sbr_c_hunit_payload,
  sbr_c_hunit_pccup,
  sbr_c_hunit_npcup,
  hunit_sbr_c_pcput,
  hunit_sbr_c_npput,
  hunit_sbr_c_eom,
  hunit_sbr_c_payload,

  // Port 4 declarations
  bunit_sbr_c_side_ism_agent,
  sbr_c_bunit_side_ism_fabric,
  bunit_sbr_c_pccup,
  bunit_sbr_c_npcup,
  sbr_c_bunit_pcput,
  sbr_c_bunit_npput,
  sbr_c_bunit_eom,
  sbr_c_bunit_payload,
  sbr_c_bunit_pccup,
  sbr_c_bunit_npcup,
  bunit_sbr_c_pcput,
  bunit_sbr_c_npput,
  bunit_sbr_c_eom,
  bunit_sbr_c_payload,

  // Port 5 declarations
  cunit_sbr_c_side_ism_agent,
  sbr_c_cunit_side_ism_fabric,
  cunit_sbr_c_pccup,
  cunit_sbr_c_npcup,
  sbr_c_cunit_pcput,
  sbr_c_cunit_npput,
  sbr_c_cunit_eom,
  sbr_c_cunit_payload,
  sbr_c_cunit_pccup,
  sbr_c_cunit_npcup,
  cunit_sbr_c_pcput,
  cunit_sbr_c_npput,
  cunit_sbr_c_eom,
  cunit_sbr_c_payload,

  // Port 6 declarations
  cpunit_sbr_c_side_ism_agent,
  sbr_c_cpunit_side_ism_fabric,
  cpunit_sbr_c_pccup,
  cpunit_sbr_c_npcup,
  sbr_c_cpunit_pcput,
  sbr_c_cpunit_npput,
  sbr_c_cpunit_eom,
  sbr_c_cpunit_payload,
  sbr_c_cpunit_pccup,
  sbr_c_cpunit_npcup,
  cpunit_sbr_c_pcput,
  cpunit_sbr_c_npput,
  cpunit_sbr_c_eom,
  cpunit_sbr_c_payload,

  // Port 7 declarations
  legacy_sbr_c_side_ism_agent,
  sbr_c_legacy_side_ism_fabric,
  legacy_sbr_c_pccup,
  legacy_sbr_c_npcup,
  sbr_c_legacy_pcput,
  sbr_c_legacy_npput,
  sbr_c_legacy_eom,
  sbr_c_legacy_payload,
  sbr_c_legacy_pccup,
  sbr_c_legacy_npcup,
  legacy_sbr_c_pcput,
  legacy_sbr_c_npput,
  legacy_sbr_c_eom,
  legacy_sbr_c_payload,

  // Port 8 declarations
  dfx_lakemore_sbr_c_side_ism_agent,
  sbr_c_dfx_lakemore_side_ism_fabric,
  dfx_lakemore_sbr_c_pccup,
  dfx_lakemore_sbr_c_npcup,
  sbr_c_dfx_lakemore_pcput,
  sbr_c_dfx_lakemore_npput,
  sbr_c_dfx_lakemore_eom,
  sbr_c_dfx_lakemore_payload,
  sbr_c_dfx_lakemore_pccup,
  sbr_c_dfx_lakemore_npcup,
  dfx_lakemore_sbr_c_pcput,
  dfx_lakemore_sbr_c_npput,
  dfx_lakemore_sbr_c_eom,
  dfx_lakemore_sbr_c_payload,

  // Port 9 declarations
  dfx_omar_sbr_c_side_ism_agent,
  sbr_c_dfx_omar_side_ism_fabric,
  dfx_omar_sbr_c_pccup,
  dfx_omar_sbr_c_npcup,
  sbr_c_dfx_omar_pcput,
  sbr_c_dfx_omar_npput,
  sbr_c_dfx_omar_eom,
  sbr_c_dfx_omar_payload,
  sbr_c_dfx_omar_pccup,
  sbr_c_dfx_omar_npcup,
  dfx_omar_sbr_c_pcput,
  dfx_omar_sbr_c_npput,
  dfx_omar_sbr_c_eom,
  dfx_omar_sbr_c_payload,

  // Port 10 declarations
  dfx_jtag_sbr_c_side_ism_agent,
  sbr_c_dfx_jtag_side_ism_fabric,
  dfx_jtag_sbr_c_pccup,
  dfx_jtag_sbr_c_npcup,
  sbr_c_dfx_jtag_pcput,
  sbr_c_dfx_jtag_npput,
  sbr_c_dfx_jtag_eom,
  sbr_c_dfx_jtag_payload,
  sbr_c_dfx_jtag_pccup,
  sbr_c_dfx_jtag_npcup,
  dfx_jtag_sbr_c_pcput,
  dfx_jtag_sbr_c_npput,
  dfx_jtag_sbr_c_eom,
  dfx_jtag_sbr_c_payload,

  // Port 11 declarations
  itunit_sbr_c_side_ism_agent,
  sbr_c_itunit_side_ism_fabric,
  itunit_sbr_c_pccup,
  itunit_sbr_c_npcup,
  sbr_c_itunit_pcput,
  sbr_c_itunit_npput,
  sbr_c_itunit_eom,
  sbr_c_itunit_payload,
  sbr_c_itunit_pccup,
  sbr_c_itunit_npcup,
  itunit_sbr_c_pcput,
  itunit_sbr_c_npput,
  itunit_sbr_c_eom,
  itunit_sbr_c_payload,

  // Port 12 declarations
  psf_3_sbr_c_side_ism_agent,
  sbr_c_psf_3_side_ism_fabric,
  psf_3_sbr_c_pccup,
  psf_3_sbr_c_npcup,
  sbr_c_psf_3_pcput,
  sbr_c_psf_3_npput,
  sbr_c_psf_3_eom,
  sbr_c_psf_3_payload,
  sbr_c_psf_3_pccup,
  sbr_c_psf_3_npcup,
  psf_3_sbr_c_pcput,
  psf_3_sbr_c_npput,
  psf_3_sbr_c_eom,
  psf_3_sbr_c_payload,

  // Port 13 declarations
  SAPms_sbr_c_side_ism_agent,
  sbr_c_SAPms_side_ism_fabric,
  SAPms_sbr_c_pccup,
  SAPms_sbr_c_npcup,
  sbr_c_SAPms_pcput,
  sbr_c_SAPms_npput,
  sbr_c_SAPms_eom,
  sbr_c_SAPms_payload,
  sbr_c_SAPms_pccup,
  sbr_c_SAPms_npcup,
  SAPms_sbr_c_pcput,
  SAPms_sbr_c_npput,
  SAPms_sbr_c_eom,
  SAPms_sbr_c_payload,

  // Port 14 declarations
  itunit2_sbr_c_side_ism_agent,
  sbr_c_itunit2_side_ism_fabric,
  itunit2_sbr_c_pccup,
  itunit2_sbr_c_npcup,
  sbr_c_itunit2_pcput,
  sbr_c_itunit2_npput,
  sbr_c_itunit2_eom,
  sbr_c_itunit2_payload,
  sbr_c_itunit2_pccup,
  sbr_c_itunit2_npcup,
  itunit2_sbr_c_pcput,
  itunit2_sbr_c_npput,
  itunit2_sbr_c_eom,
  itunit2_sbr_c_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic clk_100;
  input logic rst_b_100;

  // Asynchronous Clock/Reset(s)
  input logic clk_200;

  // Power Well Isolation Input Signals
  input logic island0_pok;
  input logic island2_pok;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic p3_fab_init_idle_exit;
  input logic p3_fab_init_idle_exit_ack;
  output logic p4_fab_init_idle_exit;
  input logic p4_fab_init_idle_exit_ack;
  output logic p5_fab_init_idle_exit;
  input logic p5_fab_init_idle_exit_ack;
  output logic p6_fab_init_idle_exit;
  input logic p6_fab_init_idle_exit_ack;
  output logic p7_fab_init_idle_exit;
  input logic p7_fab_init_idle_exit_ack;
  output logic p8_fab_init_idle_exit;
  input logic p8_fab_init_idle_exit_ack;
  output logic p9_fab_init_idle_exit;
  input logic p9_fab_init_idle_exit_ack;
  output logic p10_fab_init_idle_exit;
  input logic p10_fab_init_idle_exit_ack;
  output logic p11_fab_init_idle_exit;
  input logic p11_fab_init_idle_exit_ack;
  output logic p12_fab_init_idle_exit;
  input logic p12_fab_init_idle_exit_ack;
  output logic p13_fab_init_idle_exit;
  input logic p13_fab_init_idle_exit_ack;
  output logic p14_fab_init_idle_exit;
  input logic p14_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_clk_100;
  output visa_vp  visa_vp_clk_100;
  output visa_port_tier1 visa_p0_tier1_clk_100;
  output visa_port_tier2 visa_p0_tier2_clk_100;
  output visa_port_tier1 visa_p1_tier1_clk_100;
  output visa_port_tier2 visa_p1_tier2_clk_100;
  output visa_port_tier1 visa_p2_tier1_clk_200;
  output visa_port_tier2 visa_p2_tier2_clk_200;
  output visa_ififo_tier1 visa_p2_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p2_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p2_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p2_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p3_tier1_clk_200;
  output visa_port_tier2 visa_p3_tier2_clk_200;
  output visa_ififo_tier1 visa_p3_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p3_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p3_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p3_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p4_tier1_clk_200;
  output visa_port_tier2 visa_p4_tier2_clk_200;
  output visa_ififo_tier1 visa_p4_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p4_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p4_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p4_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p5_tier1_clk_200;
  output visa_port_tier2 visa_p5_tier2_clk_200;
  output visa_ififo_tier1 visa_p5_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p5_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p5_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p5_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p6_tier1_clk_100;
  output visa_port_tier2 visa_p6_tier2_clk_100;
  output visa_port_tier1 visa_p7_tier1_clk_100;
  output visa_port_tier2 visa_p7_tier2_clk_100;
  output visa_port_tier1 visa_p8_tier1_clk_100;
  output visa_port_tier2 visa_p8_tier2_clk_100;
  output visa_port_tier1 visa_p9_tier1_clk_100;
  output visa_port_tier2 visa_p9_tier2_clk_100;
  output visa_port_tier1 visa_p10_tier1_clk_100;
  output visa_port_tier2 visa_p10_tier2_clk_100;
  output visa_port_tier1 visa_p11_tier1_clk_100;
  output visa_port_tier2 visa_p11_tier2_clk_100;
  output visa_port_tier1 visa_p12_tier1_clk_200;
  output visa_port_tier2 visa_p12_tier2_clk_200;
  output visa_ififo_tier1 visa_p12_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p12_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p12_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p12_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p13_tier1_clk_100;
  output visa_port_tier2 visa_p13_tier2_clk_100;
  output visa_port_tier1 visa_p14_tier1_clk_100;
  output visa_port_tier2 visa_p14_tier2_clk_100;

  // Register wires
  input logic [4:0]  cfg_sbr_c_cgovrd;
  input logic [15:0] cfg_sbr_c_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic fscan_rstbypen;
  input logic fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] sbr_a_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_sbr_a_side_ism_fabric;
  input logic sbr_a_sbr_c_pccup;
  input logic sbr_a_sbr_c_npcup;
  output logic sbr_c_sbr_a_pcput;
  output logic sbr_c_sbr_a_npput;
  output logic sbr_c_sbr_a_eom;
  output logic [7:0] sbr_c_sbr_a_payload;
  output logic sbr_c_sbr_a_pccup;
  output logic sbr_c_sbr_a_npcup;
  input logic sbr_a_sbr_c_pcput;
  input logic sbr_a_sbr_c_npput;
  input logic sbr_a_sbr_c_eom;
  input logic [7:0] sbr_a_sbr_c_payload;

  // Port 1 declarations
  input logic [2:0] sbr_d_sbr_c_side_ism_fabric;
  output logic [2:0] sbr_c_sbr_d_side_ism_agent;
  input logic sbr_d_sbr_c_pccup;
  input logic sbr_d_sbr_c_npcup;
  output logic sbr_c_sbr_d_pcput;
  output logic sbr_c_sbr_d_npput;
  output logic sbr_c_sbr_d_eom;
  output logic [7:0] sbr_c_sbr_d_payload;
  output logic sbr_c_sbr_d_pccup;
  output logic sbr_c_sbr_d_npcup;
  input logic sbr_d_sbr_c_pcput;
  input logic sbr_d_sbr_c_npput;
  input logic sbr_d_sbr_c_eom;
  input logic [7:0] sbr_d_sbr_c_payload;

  // Port 2 declarations
  input logic [2:0] vtunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_vtunit_side_ism_fabric;
  input logic vtunit_sbr_c_pccup;
  input logic vtunit_sbr_c_npcup;
  output logic sbr_c_vtunit_pcput;
  output logic sbr_c_vtunit_npput;
  output logic sbr_c_vtunit_eom;
  output logic [7:0] sbr_c_vtunit_payload;
  output logic sbr_c_vtunit_pccup;
  output logic sbr_c_vtunit_npcup;
  input logic vtunit_sbr_c_pcput;
  input logic vtunit_sbr_c_npput;
  input logic vtunit_sbr_c_eom;
  input logic [7:0] vtunit_sbr_c_payload;

  // Port 3 declarations
  input logic [2:0] hunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_hunit_side_ism_fabric;
  input logic hunit_sbr_c_pccup;
  input logic hunit_sbr_c_npcup;
  output logic sbr_c_hunit_pcput;
  output logic sbr_c_hunit_npput;
  output logic sbr_c_hunit_eom;
  output logic [7:0] sbr_c_hunit_payload;
  output logic sbr_c_hunit_pccup;
  output logic sbr_c_hunit_npcup;
  input logic hunit_sbr_c_pcput;
  input logic hunit_sbr_c_npput;
  input logic hunit_sbr_c_eom;
  input logic [7:0] hunit_sbr_c_payload;

  // Port 4 declarations
  input logic [2:0] bunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_bunit_side_ism_fabric;
  input logic bunit_sbr_c_pccup;
  input logic bunit_sbr_c_npcup;
  output logic sbr_c_bunit_pcput;
  output logic sbr_c_bunit_npput;
  output logic sbr_c_bunit_eom;
  output logic [7:0] sbr_c_bunit_payload;
  output logic sbr_c_bunit_pccup;
  output logic sbr_c_bunit_npcup;
  input logic bunit_sbr_c_pcput;
  input logic bunit_sbr_c_npput;
  input logic bunit_sbr_c_eom;
  input logic [7:0] bunit_sbr_c_payload;

  // Port 5 declarations
  input logic [2:0] cunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_cunit_side_ism_fabric;
  input logic cunit_sbr_c_pccup;
  input logic cunit_sbr_c_npcup;
  output logic sbr_c_cunit_pcput;
  output logic sbr_c_cunit_npput;
  output logic sbr_c_cunit_eom;
  output logic [7:0] sbr_c_cunit_payload;
  output logic sbr_c_cunit_pccup;
  output logic sbr_c_cunit_npcup;
  input logic cunit_sbr_c_pcput;
  input logic cunit_sbr_c_npput;
  input logic cunit_sbr_c_eom;
  input logic [7:0] cunit_sbr_c_payload;

  // Port 6 declarations
  input logic [2:0] cpunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_cpunit_side_ism_fabric;
  input logic cpunit_sbr_c_pccup;
  input logic cpunit_sbr_c_npcup;
  output logic sbr_c_cpunit_pcput;
  output logic sbr_c_cpunit_npput;
  output logic sbr_c_cpunit_eom;
  output logic [7:0] sbr_c_cpunit_payload;
  output logic sbr_c_cpunit_pccup;
  output logic sbr_c_cpunit_npcup;
  input logic cpunit_sbr_c_pcput;
  input logic cpunit_sbr_c_npput;
  input logic cpunit_sbr_c_eom;
  input logic [7:0] cpunit_sbr_c_payload;

  // Port 7 declarations
  input logic [2:0] legacy_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_legacy_side_ism_fabric;
  input logic legacy_sbr_c_pccup;
  input logic legacy_sbr_c_npcup;
  output logic sbr_c_legacy_pcput;
  output logic sbr_c_legacy_npput;
  output logic sbr_c_legacy_eom;
  output logic [7:0] sbr_c_legacy_payload;
  output logic sbr_c_legacy_pccup;
  output logic sbr_c_legacy_npcup;
  input logic legacy_sbr_c_pcput;
  input logic legacy_sbr_c_npput;
  input logic legacy_sbr_c_eom;
  input logic [7:0] legacy_sbr_c_payload;

  // Port 8 declarations
  input logic [2:0] dfx_lakemore_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_dfx_lakemore_side_ism_fabric;
  input logic dfx_lakemore_sbr_c_pccup;
  input logic dfx_lakemore_sbr_c_npcup;
  output logic sbr_c_dfx_lakemore_pcput;
  output logic sbr_c_dfx_lakemore_npput;
  output logic sbr_c_dfx_lakemore_eom;
  output logic [7:0] sbr_c_dfx_lakemore_payload;
  output logic sbr_c_dfx_lakemore_pccup;
  output logic sbr_c_dfx_lakemore_npcup;
  input logic dfx_lakemore_sbr_c_pcput;
  input logic dfx_lakemore_sbr_c_npput;
  input logic dfx_lakemore_sbr_c_eom;
  input logic [7:0] dfx_lakemore_sbr_c_payload;

  // Port 9 declarations
  input logic [2:0] dfx_omar_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_dfx_omar_side_ism_fabric;
  input logic dfx_omar_sbr_c_pccup;
  input logic dfx_omar_sbr_c_npcup;
  output logic sbr_c_dfx_omar_pcput;
  output logic sbr_c_dfx_omar_npput;
  output logic sbr_c_dfx_omar_eom;
  output logic [7:0] sbr_c_dfx_omar_payload;
  output logic sbr_c_dfx_omar_pccup;
  output logic sbr_c_dfx_omar_npcup;
  input logic dfx_omar_sbr_c_pcput;
  input logic dfx_omar_sbr_c_npput;
  input logic dfx_omar_sbr_c_eom;
  input logic [7:0] dfx_omar_sbr_c_payload;

  // Port 10 declarations
  input logic [2:0] dfx_jtag_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_dfx_jtag_side_ism_fabric;
  input logic dfx_jtag_sbr_c_pccup;
  input logic dfx_jtag_sbr_c_npcup;
  output logic sbr_c_dfx_jtag_pcput;
  output logic sbr_c_dfx_jtag_npput;
  output logic sbr_c_dfx_jtag_eom;
  output logic [7:0] sbr_c_dfx_jtag_payload;
  output logic sbr_c_dfx_jtag_pccup;
  output logic sbr_c_dfx_jtag_npcup;
  input logic dfx_jtag_sbr_c_pcput;
  input logic dfx_jtag_sbr_c_npput;
  input logic dfx_jtag_sbr_c_eom;
  input logic [7:0] dfx_jtag_sbr_c_payload;

  // Port 11 declarations
  input logic [2:0] itunit_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_itunit_side_ism_fabric;
  input logic itunit_sbr_c_pccup;
  input logic itunit_sbr_c_npcup;
  output logic sbr_c_itunit_pcput;
  output logic sbr_c_itunit_npput;
  output logic sbr_c_itunit_eom;
  output logic [7:0] sbr_c_itunit_payload;
  output logic sbr_c_itunit_pccup;
  output logic sbr_c_itunit_npcup;
  input logic itunit_sbr_c_pcput;
  input logic itunit_sbr_c_npput;
  input logic itunit_sbr_c_eom;
  input logic [7:0] itunit_sbr_c_payload;

  // Port 12 declarations
  input logic [2:0] psf_3_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_psf_3_side_ism_fabric;
  input logic psf_3_sbr_c_pccup;
  input logic psf_3_sbr_c_npcup;
  output logic sbr_c_psf_3_pcput;
  output logic sbr_c_psf_3_npput;
  output logic sbr_c_psf_3_eom;
  output logic [7:0] sbr_c_psf_3_payload;
  output logic sbr_c_psf_3_pccup;
  output logic sbr_c_psf_3_npcup;
  input logic psf_3_sbr_c_pcput;
  input logic psf_3_sbr_c_npput;
  input logic psf_3_sbr_c_eom;
  input logic [7:0] psf_3_sbr_c_payload;

  // Port 13 declarations
  input logic [2:0] SAPms_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_SAPms_side_ism_fabric;
  input logic SAPms_sbr_c_pccup;
  input logic SAPms_sbr_c_npcup;
  output logic sbr_c_SAPms_pcput;
  output logic sbr_c_SAPms_npput;
  output logic sbr_c_SAPms_eom;
  output logic [7:0] sbr_c_SAPms_payload;
  output logic sbr_c_SAPms_pccup;
  output logic sbr_c_SAPms_npcup;
  input logic SAPms_sbr_c_pcput;
  input logic SAPms_sbr_c_npput;
  input logic SAPms_sbr_c_eom;
  input logic [7:0] SAPms_sbr_c_payload;

  // Port 14 declarations
  input logic [2:0] itunit2_sbr_c_side_ism_agent;
  output logic [2:0] sbr_c_itunit2_side_ism_fabric;
  input logic itunit2_sbr_c_pccup;
  input logic itunit2_sbr_c_npcup;
  output logic sbr_c_itunit2_pcput;
  output logic sbr_c_itunit2_npput;
  output logic sbr_c_itunit2_eom;
  output logic [7:0] sbr_c_itunit2_payload;
  output logic sbr_c_itunit2_pccup;
  output logic sbr_c_itunit2_npcup;
  input logic itunit2_sbr_c_pcput;
  input logic itunit2_sbr_c_npput;
  input logic itunit2_sbr_c_eom;
  input logic [7:0] itunit2_sbr_c_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_c_sbcportmap;
always_comb sbr_c_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr_c (sbr_c)                                 SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  107 { 17'b0_0000_0000_0000_0000 }},   //   254:148      SBCPORTMAPTABLE
               17'b0_0001_0000_0000_0000,      //   147          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   146          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //   145:144      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   143:140      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   139:136      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   135:132      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   131:128      SBCPORTMAPTABLE
      {   31 { 17'b0_0000_0000_0000_0000 }},   //   127: 97      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    96          SBCPORTMAPTABLE
      {    6 { 17'b0_0000_0000_0000_0000 }},   //    95: 90      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    89: 88      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    87: 86      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0010 }},   //    85: 84      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0000 }},   //    83: 81      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //    80          SBCPORTMAPTABLE
      {   13 { 17'b0_0000_0000_0000_0000 }},   //    79: 67      SBCPORTMAPTABLE
               17'b0_0100_0000_0000_0000,      //    66          SBCPORTMAPTABLE
               17'b0_0010_0000_0000_0000,      //    65          SBCPORTMAPTABLE
               17'b0_0000_1000_0000_0000,      //    64          SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0000 }},   //    63: 59      SBCPORTMAPTABLE
               17'b0_0000_0100_0000_0000,      //    58          SBCPORTMAPTABLE
               17'b0_0000_0010_0000_0000,      //    57          SBCPORTMAPTABLE
               17'b0_0000_0001_0000_0000,      //    56          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0010 }},   //    55: 54      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    53: 52      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //    51: 48      SBCPORTMAPTABLE
      {    9 { 17'b0_0000_0000_0000_0000 }},   //    47: 39      SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_1000_0000 }},   //    38: 32      SBCPORTMAPTABLE
      {   14 { 17'b0_0000_0000_0000_0000 }},   //    31: 18      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    17: 16      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    15: 14      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_1000_0000 }},   //    13: 11      SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //    10          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //     7          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     6:  5      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //     4          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //     3          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //     2          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //     1          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100       //     0          SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      = 14;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p6_pcdstvld;
logic                              p7_pcdstvld;
logic                              p8_pcdstvld;
logic                              p9_pcdstvld;
logic                              p10_pcdstvld;
logic                              p11_pcdstvld;
logic                              p13_pcdstvld;
logic                              p14_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p6_npfence;
logic                              p7_npfence;
logic                              p8_npfence;
logic                              p9_npfence;
logic                              p10_npfence;
logic                              p11_npfence;
logic                              p13_npfence;
logic                              p14_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p6_npdstvld;
logic                              p7_npdstvld;
logic                              p8_npdstvld;
logic                              p9_npdstvld;
logic                              p10_npdstvld;
logic                              p11_npdstvld;
logic                              p13_npdstvld;
logic                              p14_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              p3_ism_idle;
logic                              p3_cg_inprogress;
logic                              p3_credit_reinit;
logic                              p4_ism_idle;
logic                              p4_cg_inprogress;
logic                              p4_credit_reinit;
logic                              p5_ism_idle;
logic                              p5_cg_inprogress;
logic                              p5_credit_reinit;
logic                              p6_ism_idle;
logic                              p6_cg_inprogress;
logic                              p6_credit_reinit;
logic                              p7_ism_idle;
logic                              p7_cg_inprogress;
logic                              p7_credit_reinit;
logic                              p8_ism_idle;
logic                              p8_cg_inprogress;
logic                              p8_credit_reinit;
logic                              p9_ism_idle;
logic                              p9_cg_inprogress;
logic                              p9_credit_reinit;
logic                              p10_ism_idle;
logic                              p10_cg_inprogress;
logic                              p10_credit_reinit;
logic                              p11_ism_idle;
logic                              p11_cg_inprogress;
logic                              p11_credit_reinit;
logic                              p12_ism_idle;
logic                              p12_cg_inprogress;
logic                              p12_credit_reinit;
logic                              p13_ism_idle;
logic                              p13_cg_inprogress;
logic                              p13_credit_reinit;
logic                              p14_ism_idle;
logic                              p14_cg_inprogress;
logic                              p14_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              island0_pok_ff2;
logic                              island2_pok_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = cfg_sbr_c_cgctrl[15];
always_comb cfg_clkgatedef    = cfg_sbr_c_cgctrl[14];
always_comb cfg_idlecnt       = cfg_sbr_c_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = cfg_sbr_c_cgovrd[3];
always_comb jta_force_idle    = cfg_sbr_c_cgovrd[1];
always_comb jta_force_notidle = cfg_sbr_c_cgovrd[0];
always_comb jta_force_creditreq = cfg_sbr_c_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

// Asynchronous port signals
logic                              p2_clkgaten;
logic                              p2_clkgatedef;
logic                              p2_clkgate_ovrd;
logic                              p2_force_idle;
logic                              p2_force_notidle;
logic                              p2_force_creditreq;
logic                              p2_clken;
logic                              p2_gated_clk;
logic                              p2_agent_idle;
logic                              p2_eagent_idle;
logic                              p2_port_idle;
logic                              p2_ififo_idle;
logic                              p2_efifo_idle;
logic                              p2_pctrdy;
logic                              p2_pcirdy;
logic             [INTMAXPLDBIT:0] p2_pcdata;
logic                              p2_pceom;
logic                              p2_nptrdy;
logic                              p2_npirdy;
logic                              p2_npfence;
logic             [INTMAXPLDBIT:0] p2_npdata;
logic                              p2_npeom;
logic                              p2_enpstall;
logic                              p2_epctrdy;
logic                              p2_enptrdy;
logic                              p2_epcirdy;
logic                              p2_enpirdy;
logic                              p2_eom;
logic             [INTMAXPLDBIT:0] p2_data;

logic                              p3_clkgaten;
logic                              p3_clkgatedef;
logic                              p3_clkgate_ovrd;
logic                              p3_force_idle;
logic                              p3_force_notidle;
logic                              p3_force_creditreq;
logic                              p3_clken;
logic                              p3_gated_clk;
logic                              p3_agent_idle;
logic                              p3_eagent_idle;
logic                              p3_port_idle;
logic                              p3_ififo_idle;
logic                              p3_efifo_idle;
logic                              p3_pctrdy;
logic                              p3_pcirdy;
logic             [INTMAXPLDBIT:0] p3_pcdata;
logic                              p3_pceom;
logic                              p3_nptrdy;
logic                              p3_npirdy;
logic                              p3_npfence;
logic             [INTMAXPLDBIT:0] p3_npdata;
logic                              p3_npeom;
logic                              p3_enpstall;
logic                              p3_epctrdy;
logic                              p3_enptrdy;
logic                              p3_epcirdy;
logic                              p3_enpirdy;
logic                              p3_eom;
logic             [INTMAXPLDBIT:0] p3_data;

logic                              p4_clkgaten;
logic                              p4_clkgatedef;
logic                              p4_clkgate_ovrd;
logic                              p4_force_idle;
logic                              p4_force_notidle;
logic                              p4_force_creditreq;
logic                              p4_clken;
logic                              p4_gated_clk;
logic                              p4_agent_idle;
logic                              p4_eagent_idle;
logic                              p4_port_idle;
logic                              p4_ififo_idle;
logic                              p4_efifo_idle;
logic                              p4_pctrdy;
logic                              p4_pcirdy;
logic             [INTMAXPLDBIT:0] p4_pcdata;
logic                              p4_pceom;
logic                              p4_nptrdy;
logic                              p4_npirdy;
logic                              p4_npfence;
logic             [INTMAXPLDBIT:0] p4_npdata;
logic                              p4_npeom;
logic                              p4_enpstall;
logic                              p4_epctrdy;
logic                              p4_enptrdy;
logic                              p4_epcirdy;
logic                              p4_enpirdy;
logic                              p4_eom;
logic             [INTMAXPLDBIT:0] p4_data;

logic                              p5_clkgaten;
logic                              p5_clkgatedef;
logic                              p5_clkgate_ovrd;
logic                              p5_force_idle;
logic                              p5_force_notidle;
logic                              p5_force_creditreq;
logic                              p5_clken;
logic                              p5_gated_clk;
logic                              p5_agent_idle;
logic                              p5_eagent_idle;
logic                              p5_port_idle;
logic                              p5_ififo_idle;
logic                              p5_efifo_idle;
logic                              p5_pctrdy;
logic                              p5_pcirdy;
logic             [INTMAXPLDBIT:0] p5_pcdata;
logic                              p5_pceom;
logic                              p5_nptrdy;
logic                              p5_npirdy;
logic                              p5_npfence;
logic             [INTMAXPLDBIT:0] p5_npdata;
logic                              p5_npeom;
logic                              p5_enpstall;
logic                              p5_epctrdy;
logic                              p5_enptrdy;
logic                              p5_epcirdy;
logic                              p5_enpirdy;
logic                              p5_eom;
logic             [INTMAXPLDBIT:0] p5_data;

logic                              p12_clkgaten;
logic                              p12_clkgatedef;
logic                              p12_clkgate_ovrd;
logic                              p12_force_idle;
logic                              p12_force_notidle;
logic                              p12_force_creditreq;
logic                              p12_clken;
logic                              p12_gated_clk;
logic                              p12_agent_idle;
logic                              p12_eagent_idle;
logic                              p12_port_idle;
logic                              p12_ififo_idle;
logic                              p12_efifo_idle;
logic                              p12_pctrdy;
logic                              p12_pcirdy;
logic             [INTMAXPLDBIT:0] p12_pcdata;
logic                              p12_pceom;
logic                              p12_nptrdy;
logic                              p12_npirdy;
logic                              p12_npfence;
logic             [INTMAXPLDBIT:0] p12_npdata;
logic                              p12_npeom;
logic                              p12_enpstall;
logic                              p12_epctrdy;
logic                              p12_enptrdy;
logic                              p12_epcirdy;
logic                              p12_enpirdy;
logic                              p12_eom;
logic             [INTMAXPLDBIT:0] p12_data;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_c_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_c_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// Async clock reset synchronization
//
//------------------------------------------------------------------------------
logic clk_200_rst_b, clk_200_rst_b_pre;
sbc_doublesync sync_rst_clk_200 (
  .d     ( 1'b1 ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_200 ),
  .q     ( clk_200_rst_b_pre ));

always_comb clk_200_rst_b = fscan_rstbypen ? fscan_byprst_b : clk_200_rst_b_pre;


//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_creditreq               )
);

sbc_doublesync sync_p12_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_force_idle                )
);

sbc_doublesync sync_p12_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_force_notidle             )
);

sbc_doublesync sync_p12_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_force_creditreq           )
);

sbc_doublesync sync_p5_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_force_idle                 )
);

sbc_doublesync sync_p5_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_force_notidle              )
);

sbc_doublesync sync_p5_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_force_creditreq            )
);

sbc_doublesync sync_p4_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_force_idle                 )
);

sbc_doublesync sync_p4_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_force_notidle              )
);

sbc_doublesync sync_p4_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_force_creditreq            )
);

sbc_doublesync sync_p3_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_force_idle                 )
);

sbc_doublesync sync_p3_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_force_notidle              )
);

sbc_doublesync sync_p3_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_force_creditreq            )
);

sbc_doublesync sync_p2_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_force_idle                 )
);

sbc_doublesync sync_p2_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_force_notidle              )
);

sbc_doublesync sync_p2_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_force_creditreq            )
);

//------------------------------------------------------------------------------
//
// Asynchronous port local clock gating
//
//------------------------------------------------------------------------------
// Port 12
sbc_doublesync sync_p12_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_clkgaten                  )
);

sbc_doublesync sync_p12_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_clkgatedef                )
);

sbc_doublesync sync_p12_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p12_clkgate_ovrd              )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p12_clken <= '1;
  else
    p12_clken <= ~p12_clkgate_ovrd &
      (p12_clkgatedef | ~p12_clkgaten | ~p12_cg_inprogress |
       ((psf_3_sbr_c_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_c_psf_3_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (psf_3_sbr_c_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((psf_3_sbr_c_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_c_psf_3_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p12_clkgate  (
  .en                  ( p12_clken                     ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p12_gated_clk                 )
);

// Port 5
sbc_doublesync sync_p5_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_clkgaten                   )
);

sbc_doublesync sync_p5_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_clkgatedef                 )
);

sbc_doublesync sync_p5_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p5_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p5_clken <= '1;
  else
    p5_clken <= ~p5_clkgate_ovrd &
      (p5_clkgatedef | ~p5_clkgaten | ~p5_cg_inprogress |
       ((cunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_c_cunit_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (cunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((cunit_sbr_c_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_c_cunit_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p5_clkgate  (
  .en                  ( p5_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p5_gated_clk                  )
);

// Port 4
sbc_doublesync sync_p4_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_clkgaten                   )
);

sbc_doublesync sync_p4_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_clkgatedef                 )
);

sbc_doublesync sync_p4_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p4_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p4_clken <= '1;
  else
    p4_clken <= ~p4_clkgate_ovrd &
      (p4_clkgatedef | ~p4_clkgaten | ~p4_cg_inprogress |
       ((bunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_c_bunit_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (bunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((bunit_sbr_c_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_c_bunit_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p4_clkgate  (
  .en                  ( p4_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p4_gated_clk                  )
);

// Port 3
sbc_doublesync sync_p3_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_clkgaten                   )
);

sbc_doublesync sync_p3_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_clkgatedef                 )
);

sbc_doublesync sync_p3_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p3_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p3_clken <= '1;
  else
    p3_clken <= ~p3_clkgate_ovrd &
      (p3_clkgatedef | ~p3_clkgaten | ~p3_cg_inprogress |
       ((hunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_c_hunit_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (hunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((hunit_sbr_c_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_c_hunit_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p3_clkgate  (
  .en                  ( p3_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p3_gated_clk                  )
);

// Port 2
sbc_doublesync sync_p2_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_clkgaten                   )
);

sbc_doublesync sync_p2_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_clkgatedef                 )
);

sbc_doublesync sync_p2_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p2_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p2_clken <= '1;
  else
    p2_clken <= ~p2_clkgate_ovrd &
      (p2_clkgatedef | ~p2_clkgaten | ~p2_cg_inprogress |
       ((vtunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_c_vtunit_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (vtunit_sbr_c_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((vtunit_sbr_c_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_c_vtunit_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p2_clkgate  (
  .en                  ( p2_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p2_gated_clk                  )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_island0_pok (
  .d                   ( island0_pok                   ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( island0_pok_ff2               )
);

sbc_doublesync sync_island2_pok (
  .d                   ( island2_pok                   ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( island2_pok_ff2               )
);


always_comb endpoint_pwrgd = { 1'b1,
                          island2_pok_ff2,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          island0_pok_ff2
                        };

logic p13_gated_clk;
sbc_clock_gate p13_pwr_clkgate  (
  .en ( endpoint_pwrgd[13] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p13_gated_clk )
);

logic p0_gated_clk;
sbc_clock_gate p0_pwr_clkgate  (
  .en ( endpoint_pwrgd[0] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p0_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p14_ism_idle | ~endpoint_pwrgd[14])
                  &  (p13_ism_idle | ~endpoint_pwrgd[13])
                  &  p12_efifo_idle
                  &  (p11_ism_idle | ~endpoint_pwrgd[11])
                  &  (p10_ism_idle | ~endpoint_pwrgd[10])
                  &  (p9_ism_idle | ~endpoint_pwrgd[9])
                  &  (p8_ism_idle | ~endpoint_pwrgd[8])
                  &  (p7_ism_idle | ~endpoint_pwrgd[7])
                  &  (p6_ism_idle | ~endpoint_pwrgd[6])
                  &  p5_efifo_idle
                  &  p4_efifo_idle
                  &  p3_efifo_idle
                  &  p2_efifo_idle
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
logic p2_ism_idle_ff2, p2_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p2_ism_idle_pre <= '1;
  else
    p2_ism_idle_pre <= p2_ism_idle;

sbc_doublesync sync_idle_p2 (
  .d ( p2_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p2_ism_idle_ff2 ));

logic p3_ism_idle_ff2, p3_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p3_ism_idle_pre <= '1;
  else
    p3_ism_idle_pre <= p3_ism_idle;

sbc_doublesync sync_idle_p3 (
  .d ( p3_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p3_ism_idle_ff2 ));

logic p4_ism_idle_ff2, p4_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p4_ism_idle_pre <= '1;
  else
    p4_ism_idle_pre <= p4_ism_idle;

sbc_doublesync sync_idle_p4 (
  .d ( p4_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p4_ism_idle_ff2 ));

logic p5_ism_idle_ff2, p5_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p5_ism_idle_pre <= '1;
  else
    p5_ism_idle_pre <= p5_ism_idle;

sbc_doublesync sync_idle_p5 (
  .d ( p5_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p5_ism_idle_ff2 ));

logic p12_ism_idle_ff2, p12_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p12_ism_idle_pre <= '1;
  else
    p12_ism_idle_pre <= p12_ism_idle;

sbc_doublesync sync_idle_p12 (
  .d ( p12_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p12_ism_idle_ff2 ));

// SBR_IDLE signal for PMU
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle &
                  p2_ism_idle_ff2 &
                  p3_ism_idle_ff2 &
                  p4_ism_idle_ff2 &
                  p5_ism_idle_ff2 &
                  p6_ism_idle &
                  p7_ism_idle &
                  p8_ism_idle &
                  p9_ism_idle &
                  p10_ism_idle &
                  p11_ism_idle &
                  p12_ism_idle_ff2 &
                  p13_ism_idle &
                  p14_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p14_npfence,
                 p13_npfence,
                 1'b0,
                 p11_npfence,
                 p10_npfence,
                 p9_npfence,
                 p8_npfence,
                 p7_npfence,
                 p6_npfence,
                 1'b0,
                 1'b0,
                 1'b0,
                 1'b0,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p14_pcdstvld,
                 p13_pcdstvld,
                 pcirdy[12],
                 p11_pcdstvld,
                 p10_pcdstvld,
                 p9_pcdstvld,
                 p8_pcdstvld,
                 p7_pcdstvld,
                 p6_pcdstvld,
                 pcirdy[5],
                 pcirdy[4],
                 pcirdy[3],
                 pcirdy[2],
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p14_npdstvld,
                 p13_npdstvld,
                 npirdy[12],
                 p11_npdstvld,
                 p10_npdstvld,
                 p9_npdstvld,
                 p8_npdstvld,
                 p7_npdstvld,
                 p6_npdstvld,
                 npirdy[5],
                 npirdy[4],
                 npirdy[3],
                 npirdy[2],
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_clk_100 = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk_100                       ),
  .side_rst_b          ( rst_b_100                     ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_clk_100 = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle & agent_idle[0] & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle & p0_side_clk_valid )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_clk_100 = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_clk_100 = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( p0_gated_clk                  ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( sbr_a_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_sbr_a_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_c_sbr_a_pccup             ),
  .tnpcup              ( sbr_c_sbr_a_npcup             ),
  .tpcput              ( sbr_a_sbr_c_pcput             ),
  .tnpput              ( sbr_a_sbr_c_npput             ),
  .teom                ( sbr_a_sbr_c_eom               ),
  .tpayload            ( sbr_a_sbr_c_payload           ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( sbr_a_sbr_c_pccup             ),
  .mnpcup              ( sbr_a_sbr_c_npcup             ),
  .mpcput              ( sbr_c_sbr_a_pcput             ),
  .mnpput              ( sbr_c_sbr_a_npput             ),
  .meom                ( sbr_c_sbr_a_eom               ),
  .mpayload            ( sbr_c_sbr_a_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit & p1_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle & (~agent_idle[1] || ~p1_idle_egress) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle & agent_idle[1] & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle & p1_side_clk_valid )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle )
          p1_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

  always_comb
    begin
      visa_p1_tier1_clk_100 = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_clk_100 = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  1                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( sbr_d_sbr_c_side_ism_fabric   ),
  .side_ism_out        ( sbr_c_sbr_d_side_ism_agent    ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .idle_egress         ( p1_idle_egress                ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_c_sbr_d_pccup             ),
  .tnpcup              ( sbr_c_sbr_d_npcup             ),
  .tpcput              ( sbr_d_sbr_c_pcput             ),
  .tnpput              ( sbr_d_sbr_c_npput             ),
  .teom                ( sbr_d_sbr_c_eom               ),
  .tpayload            ( sbr_d_sbr_c_payload           ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( sbr_d_sbr_c_pccup             ),
  .mnpcup              ( sbr_d_sbr_c_npcup             ),
  .mpcput              ( sbr_c_sbr_d_pcput             ),
  .mnpput              ( sbr_c_sbr_d_npput             ),
  .meom                ( sbr_c_sbr_d_eom               ),
  .mpayload            ( sbr_c_sbr_d_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

// Port 2 (Asynchronous port)
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  logic p2_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit_ff2 & p2_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle_ff2 & (~agent_idle[2] || ~p2_efifo_idle) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle_ff2 & agent_idle[2] & p2_efifo_idle & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle_ff2 & p2_side_clk_valid & ~p2_fab_init_idle_exit )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle_ff2 )
          p2_side_clk_valid <= '1;
      end

logic p2_side_clk_valid_ff2;
sbc_doublesync sync_p2_clk_valid (
  .d     ( p2_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p2_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p2_credit_reinit (
  .d     ( p2_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p2_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

logic [15:0] p2_dbgbus_ing;
logic [15:0] p2_dbgbus_egr;
  always_comb
    begin
      visa_p2_tier1_clk_200 = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_clk_200 = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
      visa_p2_ififo_tier1_clk_100 = { p2_dbgbus_ing[15:14],
                             p2_dbgbus_ing[5:0]};
      visa_p2_ififo_tier2_clk_100 = { p2_dbgbus_ing[13:6] };
      visa_p2_efifo_tier1_clk_100 = { p2_dbgbus_egr[7:0] };
      visa_p2_efifo_tier2_clk_100 = { p2_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p2_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p2_side_clk_valid_ff2         ),
  .side_ism_in         ( vtunit_sbr_c_side_ism_agent   ),
  .side_ism_out        ( sbr_c_vtunit_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( p2_agent_idle                 ),
  .port_idle           ( p2_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_c_vtunit_pccup            ),
  .tnpcup              ( sbr_c_vtunit_npcup            ),
  .tpcput              ( vtunit_sbr_c_pcput            ),
  .tnpput              ( vtunit_sbr_c_npput            ),
  .teom                ( vtunit_sbr_c_eom              ),
  .tpayload            ( vtunit_sbr_c_payload          ),
  .pctrdy              ( p2_pctrdy                     ),
  .pcirdy              ( p2_pcirdy                     ),
  .pcdata              ( p2_pcdata                     ),
  .pceom               ( p2_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p2_nptrdy                     ),
  .npirdy              ( p2_npirdy                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( p2_npdata                     ),
  .npeom               ( p2_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( vtunit_sbr_c_pccup            ),
  .mnpcup              ( vtunit_sbr_c_npcup            ),
  .mpcput              ( sbr_c_vtunit_pcput            ),
  .mnpput              ( sbr_c_vtunit_npput            ),
  .meom                ( sbr_c_vtunit_eom              ),
  .mpayload            ( sbr_c_vtunit_payload          ),
  .enpstall            ( p2_enpstall                   ),
  .epctrdy             ( p2_epctrdy                    ),
  .enptrdy             ( p2_enptrdy                    ),
  .epcirdy             ( p2_epcirdy                    ),
  .enpirdy             ( p2_enpirdy                    ),
  .data                ( p2_data                       ),
  .eom                 ( p2_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p2_clkgaten                   ),
  .force_idle          ( p2_force_idle                 ),
  .force_notidle       ( p2_force_notidle              ),
  .force_creditreq     ( p2_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         ( 10                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress2 (
  .ing_side_clk        ( p2_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p2_port_idle                  ),
  .pcirdy              ( p2_pcirdy                     ),
  .npirdy              ( p2_npirdy                     ),
  .npfence             ( p2_npfence                    ),
  .pceom               ( p2_pceom                      ),
  .pcdata              ( p2_pcdata                     ),
  .npeom               ( p2_npeom                      ),
  .npdata              ( p2_npdata                     ),
  .pctrdy              ( p2_pctrdy                     ),
  .nptrdy              ( p2_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p2_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[2]                     ),
  .enptrdy             ( nptrdy[2]                     ),
  .epcirdy             ( pcirdy[2]                     ),
  .enpirdy             ( npirdy[2]                     ),
  .eom                 ( npeom[2]                      ),
  .data                ( npdata[2]                     ),
  .opceom              ( pceom[2]                      ),
  .opcdata             ( pcdata[2]                     ),
  .agent_idle          ( port_idle[2]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p2_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress2 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[2]                 ),
  .pcirdy              ( epcirdy[2]                    ),
  .npirdy              ( enpirdy[2]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[2]                    ),
  .nptrdy              ( enptrdy[2]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p2_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p2_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p2_enpstall                   ),
  .epctrdy             ( p2_epctrdy                    ),
  .enptrdy             ( p2_enptrdy                    ),
  .epcirdy             ( p2_epcirdy                    ),
  .enpirdy             ( p2_enpirdy                    ),
  .eom                 ( p2_eom                        ),
  .data                ( p2_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p2_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p2_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p2_agent_idle  = p2_eagent_idle & p2_ififo_idle;

// Port 3 (Asynchronous port)
logic p3_side_clk_valid, p3_idle_egress, p3_rst_suppress;
  logic p3_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_rst_suppress <= 1'b1;
    else
      p3_rst_suppress <= p3_credit_reinit_ff2 & p3_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p3_fab_init_idle_exit <= '1;
    else
      if ( ~p3_rst_suppress & (p3_ism_idle_ff2 & (~agent_idle[3] || ~p3_efifo_idle) & ~p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '1;
      else if ( ~p3_rst_suppress & (p3_ism_idle_ff2 & agent_idle[3] & p3_efifo_idle & p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( p3_ism_idle_ff2 & p3_side_clk_valid & ~p3_fab_init_idle_exit )
          p3_side_clk_valid <= '0;
        else if ( (p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack) || ~p3_ism_idle_ff2 )
          p3_side_clk_valid <= '1;
      end

logic p3_side_clk_valid_ff2;
sbc_doublesync sync_p3_clk_valid (
  .d     ( p3_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p3_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p3_credit_reinit (
  .d     ( p3_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p3_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

logic [15:0] p3_dbgbus_ing;
logic [15:0] p3_dbgbus_egr;
  always_comb
    begin
      visa_p3_tier1_clk_200 = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_clk_200 = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
      visa_p3_ififo_tier1_clk_100 = { p3_dbgbus_ing[15:14],
                             p3_dbgbus_ing[5:0]};
      visa_p3_ififo_tier2_clk_100 = { p3_dbgbus_ing[13:6] };
      visa_p3_efifo_tier1_clk_100 = { p3_dbgbus_egr[7:0] };
      visa_p3_efifo_tier2_clk_100 = { p3_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p3_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p3_side_clk_valid_ff2         ),
  .side_ism_in         ( hunit_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_hunit_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( p3_agent_idle                 ),
  .port_idle           ( p3_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p3_ism_idle                   ),
  .credit_reinit       ( p3_credit_reinit              ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_c_hunit_pccup             ),
  .tnpcup              ( sbr_c_hunit_npcup             ),
  .tpcput              ( hunit_sbr_c_pcput             ),
  .tnpput              ( hunit_sbr_c_npput             ),
  .teom                ( hunit_sbr_c_eom               ),
  .tpayload            ( hunit_sbr_c_payload           ),
  .pctrdy              ( p3_pctrdy                     ),
  .pcirdy              ( p3_pcirdy                     ),
  .pcdata              ( p3_pcdata                     ),
  .pceom               ( p3_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p3_nptrdy                     ),
  .npirdy              ( p3_npirdy                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( p3_npdata                     ),
  .npeom               ( p3_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( hunit_sbr_c_pccup             ),
  .mnpcup              ( hunit_sbr_c_npcup             ),
  .mpcput              ( sbr_c_hunit_pcput             ),
  .mnpput              ( sbr_c_hunit_npput             ),
  .meom                ( sbr_c_hunit_eom               ),
  .mpayload            ( sbr_c_hunit_payload           ),
  .enpstall            ( p3_enpstall                   ),
  .epctrdy             ( p3_epctrdy                    ),
  .enptrdy             ( p3_enptrdy                    ),
  .epcirdy             ( p3_epcirdy                    ),
  .enpirdy             ( p3_enpirdy                    ),
  .data                ( p3_data                       ),
  .eom                 ( p3_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p3_clkgaten                   ),
  .force_idle          ( p3_force_idle                 ),
  .force_notidle       ( p3_force_notidle              ),
  .force_creditreq     ( p3_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         ( 10                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress3 (
  .ing_side_clk        ( p3_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p3_port_idle                  ),
  .pcirdy              ( p3_pcirdy                     ),
  .npirdy              ( p3_npirdy                     ),
  .npfence             ( p3_npfence                    ),
  .pceom               ( p3_pceom                      ),
  .pcdata              ( p3_pcdata                     ),
  .npeom               ( p3_npeom                      ),
  .npdata              ( p3_npdata                     ),
  .pctrdy              ( p3_pctrdy                     ),
  .nptrdy              ( p3_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p3_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[3]                     ),
  .enptrdy             ( nptrdy[3]                     ),
  .epcirdy             ( pcirdy[3]                     ),
  .enpirdy             ( npirdy[3]                     ),
  .eom                 ( npeom[3]                      ),
  .data                ( npdata[3]                     ),
  .opceom              ( pceom[3]                      ),
  .opcdata             ( pcdata[3]                     ),
  .agent_idle          ( port_idle[3]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p3_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress3 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[3]                 ),
  .pcirdy              ( epcirdy[3]                    ),
  .npirdy              ( enpirdy[3]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[3]                    ),
  .nptrdy              ( enptrdy[3]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p3_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p3_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p3_enpstall                   ),
  .epctrdy             ( p3_epctrdy                    ),
  .enptrdy             ( p3_enptrdy                    ),
  .epcirdy             ( p3_epcirdy                    ),
  .enpirdy             ( p3_enpirdy                    ),
  .eom                 ( p3_eom                        ),
  .data                ( p3_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p3_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p3_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p3_agent_idle  = p3_eagent_idle & p3_ififo_idle;

// Port 4 (Asynchronous port)
logic p4_side_clk_valid, p4_idle_egress, p4_rst_suppress;
  logic p4_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_rst_suppress <= 1'b1;
    else
      p4_rst_suppress <= p4_credit_reinit_ff2 & p4_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p4_fab_init_idle_exit <= '1;
    else
      if ( ~p4_rst_suppress & (p4_ism_idle_ff2 & (~agent_idle[4] || ~p4_efifo_idle) & ~p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '1;
      else if ( ~p4_rst_suppress & (p4_ism_idle_ff2 & agent_idle[4] & p4_efifo_idle & p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( p4_ism_idle_ff2 & p4_side_clk_valid & ~p4_fab_init_idle_exit )
          p4_side_clk_valid <= '0;
        else if ( (p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack) || ~p4_ism_idle_ff2 )
          p4_side_clk_valid <= '1;
      end

logic p4_side_clk_valid_ff2;
sbc_doublesync sync_p4_clk_valid (
  .d     ( p4_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p4_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p4_credit_reinit (
  .d     ( p4_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p4_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

logic [15:0] p4_dbgbus_ing;
logic [15:0] p4_dbgbus_egr;
  always_comb
    begin
      visa_p4_tier1_clk_200 = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_clk_200 = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
      visa_p4_ififo_tier1_clk_100 = { p4_dbgbus_ing[15:14],
                             p4_dbgbus_ing[5:0]};
      visa_p4_ififo_tier2_clk_100 = { p4_dbgbus_ing[13:6] };
      visa_p4_efifo_tier1_clk_100 = { p4_dbgbus_egr[7:0] };
      visa_p4_efifo_tier2_clk_100 = { p4_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p4_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p4_side_clk_valid_ff2         ),
  .side_ism_in         ( bunit_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_bunit_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( p4_agent_idle                 ),
  .port_idle           ( p4_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p4_ism_idle                   ),
  .credit_reinit       ( p4_credit_reinit              ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_c_bunit_pccup             ),
  .tnpcup              ( sbr_c_bunit_npcup             ),
  .tpcput              ( bunit_sbr_c_pcput             ),
  .tnpput              ( bunit_sbr_c_npput             ),
  .teom                ( bunit_sbr_c_eom               ),
  .tpayload            ( bunit_sbr_c_payload           ),
  .pctrdy              ( p4_pctrdy                     ),
  .pcirdy              ( p4_pcirdy                     ),
  .pcdata              ( p4_pcdata                     ),
  .pceom               ( p4_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p4_nptrdy                     ),
  .npirdy              ( p4_npirdy                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( p4_npdata                     ),
  .npeom               ( p4_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( bunit_sbr_c_pccup             ),
  .mnpcup              ( bunit_sbr_c_npcup             ),
  .mpcput              ( sbr_c_bunit_pcput             ),
  .mnpput              ( sbr_c_bunit_npput             ),
  .meom                ( sbr_c_bunit_eom               ),
  .mpayload            ( sbr_c_bunit_payload           ),
  .enpstall            ( p4_enpstall                   ),
  .epctrdy             ( p4_epctrdy                    ),
  .enptrdy             ( p4_enptrdy                    ),
  .epcirdy             ( p4_epcirdy                    ),
  .enpirdy             ( p4_enpirdy                    ),
  .data                ( p4_data                       ),
  .eom                 ( p4_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p4_clkgaten                   ),
  .force_idle          ( p4_force_idle                 ),
  .force_notidle       ( p4_force_notidle              ),
  .force_creditreq     ( p4_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         ( 10                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress4 (
  .ing_side_clk        ( p4_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p4_port_idle                  ),
  .pcirdy              ( p4_pcirdy                     ),
  .npirdy              ( p4_npirdy                     ),
  .npfence             ( p4_npfence                    ),
  .pceom               ( p4_pceom                      ),
  .pcdata              ( p4_pcdata                     ),
  .npeom               ( p4_npeom                      ),
  .npdata              ( p4_npdata                     ),
  .pctrdy              ( p4_pctrdy                     ),
  .nptrdy              ( p4_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p4_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[4]                     ),
  .enptrdy             ( nptrdy[4]                     ),
  .epcirdy             ( pcirdy[4]                     ),
  .enpirdy             ( npirdy[4]                     ),
  .eom                 ( npeom[4]                      ),
  .data                ( npdata[4]                     ),
  .opceom              ( pceom[4]                      ),
  .opcdata             ( pcdata[4]                     ),
  .agent_idle          ( port_idle[4]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p4_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress4 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[4]                 ),
  .pcirdy              ( epcirdy[4]                    ),
  .npirdy              ( enpirdy[4]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[4]                    ),
  .nptrdy              ( enptrdy[4]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p4_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p4_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p4_enpstall                   ),
  .epctrdy             ( p4_epctrdy                    ),
  .enptrdy             ( p4_enptrdy                    ),
  .epcirdy             ( p4_epcirdy                    ),
  .enpirdy             ( p4_enpirdy                    ),
  .eom                 ( p4_eom                        ),
  .data                ( p4_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p4_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p4_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p4_agent_idle  = p4_eagent_idle & p4_ififo_idle;

// Port 5 (Asynchronous port)
logic p5_side_clk_valid, p5_idle_egress, p5_rst_suppress;
  logic p5_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p5_rst_suppress <= 1'b1;
    else
      p5_rst_suppress <= p5_credit_reinit_ff2 & p5_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p5_fab_init_idle_exit <= '1;
    else
      if ( ~p5_rst_suppress & (p5_ism_idle_ff2 & (~agent_idle[5] || ~p5_efifo_idle) & ~p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '1;
      else if ( ~p5_rst_suppress & (p5_ism_idle_ff2 & agent_idle[5] & p5_efifo_idle & p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p5_side_clk_valid <= 1'b0;
    else
      begin
        if ( p5_ism_idle_ff2 & p5_side_clk_valid & ~p5_fab_init_idle_exit )
          p5_side_clk_valid <= '0;
        else if ( (p5_fab_init_idle_exit & p5_fab_init_idle_exit_ack) || ~p5_ism_idle_ff2 )
          p5_side_clk_valid <= '1;
      end

logic p5_side_clk_valid_ff2;
sbc_doublesync sync_p5_clk_valid (
  .d     ( p5_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p5_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p5_credit_reinit (
  .d     ( p5_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p5_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p5_dbgbus;

logic [15:0] p5_dbgbus_ing;
logic [15:0] p5_dbgbus_egr;
  always_comb
    begin
      visa_p5_tier1_clk_200 = { p5_dbgbus[31],
                            p5_dbgbus[27:24],
                            p5_dbgbus[21:19],
                            p5_dbgbus[15:12],
                            p5_dbgbus[7:4] };
      visa_p5_tier2_clk_200 = { p5_dbgbus[30:28],
                            p5_dbgbus[23:22],
                            p5_dbgbus[18:16],
                            p5_dbgbus[11:8],
                            p5_dbgbus[3:0] };
      visa_p5_ififo_tier1_clk_100 = { p5_dbgbus_ing[15:14],
                             p5_dbgbus_ing[5:0]};
      visa_p5_ififo_tier2_clk_100 = { p5_dbgbus_ing[13:6] };
      visa_p5_efifo_tier1_clk_100 = { p5_dbgbus_egr[7:0] };
      visa_p5_efifo_tier2_clk_100 = { p5_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport5 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p5_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p5_side_clk_valid_ff2         ),
  .side_ism_in         ( cunit_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_cunit_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[5] ),
  .agent_idle          ( p5_agent_idle                 ),
  .port_idle           ( p5_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p5_ism_idle                   ),
  .credit_reinit       ( p5_credit_reinit              ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr_c_cunit_pccup             ),
  .tnpcup              ( sbr_c_cunit_npcup             ),
  .tpcput              ( cunit_sbr_c_pcput             ),
  .tnpput              ( cunit_sbr_c_npput             ),
  .teom                ( cunit_sbr_c_eom               ),
  .tpayload            ( cunit_sbr_c_payload           ),
  .pctrdy              ( p5_pctrdy                     ),
  .pcirdy              ( p5_pcirdy                     ),
  .pcdata              ( p5_pcdata                     ),
  .pceom               ( p5_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p5_nptrdy                     ),
  .npirdy              ( p5_npirdy                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( p5_npdata                     ),
  .npeom               ( p5_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( cunit_sbr_c_pccup             ),
  .mnpcup              ( cunit_sbr_c_npcup             ),
  .mpcput              ( sbr_c_cunit_pcput             ),
  .mnpput              ( sbr_c_cunit_npput             ),
  .meom                ( sbr_c_cunit_eom               ),
  .mpayload            ( sbr_c_cunit_payload           ),
  .enpstall            ( p5_enpstall                   ),
  .epctrdy             ( p5_epctrdy                    ),
  .enptrdy             ( p5_enptrdy                    ),
  .epcirdy             ( p5_epcirdy                    ),
  .enpirdy             ( p5_enpirdy                    ),
  .data                ( p5_data                       ),
  .eom                 ( p5_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p5_clkgaten                   ),
  .force_idle          ( p5_force_idle                 ),
  .force_notidle       ( p5_force_notidle              ),
  .force_creditreq     ( p5_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p5_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         ( 10                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress5 (
  .ing_side_clk        ( p5_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p5_port_idle                  ),
  .pcirdy              ( p5_pcirdy                     ),
  .npirdy              ( p5_npirdy                     ),
  .npfence             ( p5_npfence                    ),
  .pceom               ( p5_pceom                      ),
  .pcdata              ( p5_pcdata                     ),
  .npeom               ( p5_npeom                      ),
  .npdata              ( p5_npdata                     ),
  .pctrdy              ( p5_pctrdy                     ),
  .nptrdy              ( p5_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p5_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[5]                     ),
  .enptrdy             ( nptrdy[5]                     ),
  .epcirdy             ( pcirdy[5]                     ),
  .enpirdy             ( npirdy[5]                     ),
  .eom                 ( npeom[5]                      ),
  .data                ( npdata[5]                     ),
  .opceom              ( pceom[5]                      ),
  .opcdata             ( pcdata[5]                     ),
  .agent_idle          ( port_idle[5]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p5_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress5 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[5]                 ),
  .pcirdy              ( epcirdy[5]                    ),
  .npirdy              ( enpirdy[5]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[5]                    ),
  .nptrdy              ( enptrdy[5]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p5_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p5_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p5_enpstall                   ),
  .epctrdy             ( p5_epctrdy                    ),
  .enptrdy             ( p5_enptrdy                    ),
  .epcirdy             ( p5_epcirdy                    ),
  .enpirdy             ( p5_enpirdy                    ),
  .eom                 ( p5_eom                        ),
  .data                ( p5_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p5_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p5_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p5_agent_idle  = p5_eagent_idle & p5_ififo_idle;

// Port 6
logic p6_side_clk_valid, p6_idle_egress, p6_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p6_rst_suppress <= 1'b1;
    else
      p6_rst_suppress <= p6_credit_reinit & p6_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p6_fab_init_idle_exit <= '1;
    else
      if ( ~p6_rst_suppress & (p6_ism_idle & (~agent_idle[6] || ~p6_idle_egress) & ~p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '1;
      else if ( ~p6_rst_suppress & (p6_ism_idle & agent_idle[6] & p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p6_side_clk_valid <= 1'b0;
    else
      begin
        if ( p6_ism_idle & p6_side_clk_valid )
          p6_side_clk_valid <= '0;
        else if ( (p6_fab_init_idle_exit & p6_fab_init_idle_exit_ack) || ~p6_ism_idle )
          p6_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p6_dbgbus;

  always_comb
    begin
      visa_p6_tier1_clk_100 = { p6_dbgbus[31],
                            p6_dbgbus[27:24],
                            p6_dbgbus[21:19],
                            p6_dbgbus[15:12],
                            p6_dbgbus[7:4] };
      visa_p6_tier2_clk_100 = { p6_dbgbus[30:28],
                            p6_dbgbus[23:22],
                            p6_dbgbus[18:16],
                            p6_dbgbus[11:8],
                            p6_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport6 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p6_side_clk_valid             ),
  .side_ism_in         ( cpunit_sbr_c_side_ism_agent   ),
  .side_ism_out        ( sbr_c_cpunit_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[6] ),
  .agent_idle          ( agent_idle[6]                 ),
  .port_idle           ( port_idle[6]                  ),
  .idle_egress         ( p6_idle_egress                ),
  .ism_idle            ( p6_ism_idle                   ),
  .credit_reinit       ( p6_credit_reinit              ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr_c_cpunit_pccup            ),
  .tnpcup              ( sbr_c_cpunit_npcup            ),
  .tpcput              ( cpunit_sbr_c_pcput            ),
  .tnpput              ( cpunit_sbr_c_npput            ),
  .teom                ( cpunit_sbr_c_eom              ),
  .tpayload            ( cpunit_sbr_c_payload          ),
  .pctrdy              ( pctrdy[6]                     ),
  .pcirdy              ( pcirdy[6]                     ),
  .pcdata              ( pcdata[6]                     ),
  .pceom               ( pceom[6]                      ),
  .pcdstvld            ( p6_pcdstvld                   ),
  .nptrdy              ( nptrdy[6]                     ),
  .npirdy              ( npirdy[6]                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( npdata[6]                     ),
  .npeom               ( npeom[6]                      ),
  .npdstvld            ( p6_npdstvld                   ),
  .mpccup              ( cpunit_sbr_c_pccup            ),
  .mnpcup              ( cpunit_sbr_c_npcup            ),
  .mpcput              ( sbr_c_cpunit_pcput            ),
  .mnpput              ( sbr_c_cpunit_npput            ),
  .meom                ( sbr_c_cpunit_eom              ),
  .mpayload            ( sbr_c_cpunit_payload          ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[6]                    ),
  .enptrdy             ( enptrdy[6]                    ),
  .epcirdy             ( epcirdy[6]                    ),
  .enpirdy             ( enpirdy[6]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p6_dbgbus                     )
);

// Port 7
logic p7_side_clk_valid, p7_idle_egress, p7_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p7_rst_suppress <= 1'b1;
    else
      p7_rst_suppress <= p7_credit_reinit & p7_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p7_fab_init_idle_exit <= '1;
    else
      if ( ~p7_rst_suppress & (p7_ism_idle & (~agent_idle[7] || ~p7_idle_egress) & ~p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '1;
      else if ( ~p7_rst_suppress & (p7_ism_idle & agent_idle[7] & p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p7_side_clk_valid <= 1'b0;
    else
      begin
        if ( p7_ism_idle & p7_side_clk_valid )
          p7_side_clk_valid <= '0;
        else if ( (p7_fab_init_idle_exit & p7_fab_init_idle_exit_ack) || ~p7_ism_idle )
          p7_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p7_dbgbus;

  always_comb
    begin
      visa_p7_tier1_clk_100 = { p7_dbgbus[31],
                            p7_dbgbus[27:24],
                            p7_dbgbus[21:19],
                            p7_dbgbus[15:12],
                            p7_dbgbus[7:4] };
      visa_p7_tier2_clk_100 = { p7_dbgbus[30:28],
                            p7_dbgbus[23:22],
                            p7_dbgbus[18:16],
                            p7_dbgbus[11:8],
                            p7_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport7 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( legacy_sbr_c_side_ism_agent   ),
  .side_ism_out        ( sbr_c_legacy_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[7] ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .idle_egress         ( p7_idle_egress                ),
  .ism_idle            ( p7_ism_idle                   ),
  .credit_reinit       ( p7_credit_reinit              ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr_c_legacy_pccup            ),
  .tnpcup              ( sbr_c_legacy_npcup            ),
  .tpcput              ( legacy_sbr_c_pcput            ),
  .tnpput              ( legacy_sbr_c_npput            ),
  .teom                ( legacy_sbr_c_eom              ),
  .tpayload            ( legacy_sbr_c_payload          ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( legacy_sbr_c_pccup            ),
  .mnpcup              ( legacy_sbr_c_npcup            ),
  .mpcput              ( sbr_c_legacy_pcput            ),
  .mnpput              ( sbr_c_legacy_npput            ),
  .meom                ( sbr_c_legacy_eom              ),
  .mpayload            ( sbr_c_legacy_payload          ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p7_dbgbus                     )
);

// Port 8
logic p8_side_clk_valid, p8_idle_egress, p8_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p8_rst_suppress <= 1'b1;
    else
      p8_rst_suppress <= p8_credit_reinit & p8_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p8_fab_init_idle_exit <= '1;
    else
      if ( ~p8_rst_suppress & (p8_ism_idle & (~agent_idle[8] || ~p8_idle_egress) & ~p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '1;
      else if ( ~p8_rst_suppress & (p8_ism_idle & agent_idle[8] & p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p8_side_clk_valid <= 1'b0;
    else
      begin
        if ( p8_ism_idle & p8_side_clk_valid )
          p8_side_clk_valid <= '0;
        else if ( (p8_fab_init_idle_exit & p8_fab_init_idle_exit_ack) || ~p8_ism_idle )
          p8_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p8_dbgbus;

  always_comb
    begin
      visa_p8_tier1_clk_100 = { p8_dbgbus[31],
                            p8_dbgbus[27:24],
                            p8_dbgbus[21:19],
                            p8_dbgbus[15:12],
                            p8_dbgbus[7:4] };
      visa_p8_tier2_clk_100 = { p8_dbgbus[30:28],
                            p8_dbgbus[23:22],
                            p8_dbgbus[18:16],
                            p8_dbgbus[11:8],
                            p8_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport8 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p8_side_clk_valid             ),
  .side_ism_in         ( dfx_lakemore_sbr_c_side_ism_agent),
  .side_ism_out        ( sbr_c_dfx_lakemore_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[8] ),
  .agent_idle          ( agent_idle[8]                 ),
  .port_idle           ( port_idle[8]                  ),
  .idle_egress         ( p8_idle_egress                ),
  .ism_idle            ( p8_ism_idle                   ),
  .credit_reinit       ( p8_credit_reinit              ),
  .cg_inprogress       ( p8_cg_inprogress              ),
  .tpccup              ( sbr_c_dfx_lakemore_pccup      ),
  .tnpcup              ( sbr_c_dfx_lakemore_npcup      ),
  .tpcput              ( dfx_lakemore_sbr_c_pcput      ),
  .tnpput              ( dfx_lakemore_sbr_c_npput      ),
  .teom                ( dfx_lakemore_sbr_c_eom        ),
  .tpayload            ( dfx_lakemore_sbr_c_payload    ),
  .pctrdy              ( pctrdy[8]                     ),
  .pcirdy              ( pcirdy[8]                     ),
  .pcdata              ( pcdata[8]                     ),
  .pceom               ( pceom[8]                      ),
  .pcdstvld            ( p8_pcdstvld                   ),
  .nptrdy              ( nptrdy[8]                     ),
  .npirdy              ( npirdy[8]                     ),
  .npfence             ( p8_npfence                    ),
  .npdata              ( npdata[8]                     ),
  .npeom               ( npeom[8]                      ),
  .npdstvld            ( p8_npdstvld                   ),
  .mpccup              ( dfx_lakemore_sbr_c_pccup      ),
  .mnpcup              ( dfx_lakemore_sbr_c_npcup      ),
  .mpcput              ( sbr_c_dfx_lakemore_pcput      ),
  .mnpput              ( sbr_c_dfx_lakemore_npput      ),
  .meom                ( sbr_c_dfx_lakemore_eom        ),
  .mpayload            ( sbr_c_dfx_lakemore_payload    ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[8]                    ),
  .enptrdy             ( enptrdy[8]                    ),
  .epcirdy             ( epcirdy[8]                    ),
  .enpirdy             ( enpirdy[8]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p8_dbgbus                     )
);

// Port 9
logic p9_side_clk_valid, p9_idle_egress, p9_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p9_rst_suppress <= 1'b1;
    else
      p9_rst_suppress <= p9_credit_reinit & p9_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p9_fab_init_idle_exit <= '1;
    else
      if ( ~p9_rst_suppress & (p9_ism_idle & (~agent_idle[9] || ~p9_idle_egress) & ~p9_fab_init_idle_exit_ack ))
        p9_fab_init_idle_exit <= '1;
      else if ( ~p9_rst_suppress & (p9_ism_idle & agent_idle[9] & p9_fab_init_idle_exit_ack ))
        p9_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p9_side_clk_valid <= 1'b0;
    else
      begin
        if ( p9_ism_idle & p9_side_clk_valid )
          p9_side_clk_valid <= '0;
        else if ( (p9_fab_init_idle_exit & p9_fab_init_idle_exit_ack) || ~p9_ism_idle )
          p9_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p9_dbgbus;

  always_comb
    begin
      visa_p9_tier1_clk_100 = { p9_dbgbus[31],
                            p9_dbgbus[27:24],
                            p9_dbgbus[21:19],
                            p9_dbgbus[15:12],
                            p9_dbgbus[7:4] };
      visa_p9_tier2_clk_100 = { p9_dbgbus[30:28],
                            p9_dbgbus[23:22],
                            p9_dbgbus[18:16],
                            p9_dbgbus[11:8],
                            p9_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport9 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p9_side_clk_valid             ),
  .side_ism_in         ( dfx_omar_sbr_c_side_ism_agent ),
  .side_ism_out        ( sbr_c_dfx_omar_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[9] ),
  .agent_idle          ( agent_idle[9]                 ),
  .port_idle           ( port_idle[9]                  ),
  .idle_egress         ( p9_idle_egress                ),
  .ism_idle            ( p9_ism_idle                   ),
  .credit_reinit       ( p9_credit_reinit              ),
  .cg_inprogress       ( p9_cg_inprogress              ),
  .tpccup              ( sbr_c_dfx_omar_pccup          ),
  .tnpcup              ( sbr_c_dfx_omar_npcup          ),
  .tpcput              ( dfx_omar_sbr_c_pcput          ),
  .tnpput              ( dfx_omar_sbr_c_npput          ),
  .teom                ( dfx_omar_sbr_c_eom            ),
  .tpayload            ( dfx_omar_sbr_c_payload        ),
  .pctrdy              ( pctrdy[9]                     ),
  .pcirdy              ( pcirdy[9]                     ),
  .pcdata              ( pcdata[9]                     ),
  .pceom               ( pceom[9]                      ),
  .pcdstvld            ( p9_pcdstvld                   ),
  .nptrdy              ( nptrdy[9]                     ),
  .npirdy              ( npirdy[9]                     ),
  .npfence             ( p9_npfence                    ),
  .npdata              ( npdata[9]                     ),
  .npeom               ( npeom[9]                      ),
  .npdstvld            ( p9_npdstvld                   ),
  .mpccup              ( dfx_omar_sbr_c_pccup          ),
  .mnpcup              ( dfx_omar_sbr_c_npcup          ),
  .mpcput              ( sbr_c_dfx_omar_pcput          ),
  .mnpput              ( sbr_c_dfx_omar_npput          ),
  .meom                ( sbr_c_dfx_omar_eom            ),
  .mpayload            ( sbr_c_dfx_omar_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[9]                    ),
  .enptrdy             ( enptrdy[9]                    ),
  .epcirdy             ( epcirdy[9]                    ),
  .enpirdy             ( enpirdy[9]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p9_dbgbus                     )
);

// Port 10
logic p10_side_clk_valid, p10_idle_egress, p10_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p10_rst_suppress <= 1'b1;
    else
      p10_rst_suppress <= p10_credit_reinit & p10_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p10_fab_init_idle_exit <= '1;
    else
      if ( ~p10_rst_suppress & (p10_ism_idle & (~agent_idle[10] || ~p10_idle_egress) & ~p10_fab_init_idle_exit_ack ))
        p10_fab_init_idle_exit <= '1;
      else if ( ~p10_rst_suppress & (p10_ism_idle & agent_idle[10] & p10_fab_init_idle_exit_ack ))
        p10_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p10_side_clk_valid <= 1'b0;
    else
      begin
        if ( p10_ism_idle & p10_side_clk_valid )
          p10_side_clk_valid <= '0;
        else if ( (p10_fab_init_idle_exit & p10_fab_init_idle_exit_ack) || ~p10_ism_idle )
          p10_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p10_dbgbus;

  always_comb
    begin
      visa_p10_tier1_clk_100 = { p10_dbgbus[31],
                            p10_dbgbus[27:24],
                            p10_dbgbus[21:19],
                            p10_dbgbus[15:12],
                            p10_dbgbus[7:4] };
      visa_p10_tier2_clk_100 = { p10_dbgbus[30:28],
                            p10_dbgbus[23:22],
                            p10_dbgbus[18:16],
                            p10_dbgbus[11:8],
                            p10_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport10 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p10_side_clk_valid            ),
  .side_ism_in         ( dfx_jtag_sbr_c_side_ism_agent ),
  .side_ism_out        ( sbr_c_dfx_jtag_side_ism_fabric),
  .int_pok             ( endpoint_pwrgd[10] ),
  .agent_idle          ( agent_idle[10]                ),
  .port_idle           ( port_idle[10]                 ),
  .idle_egress         ( p10_idle_egress               ),
  .ism_idle            ( p10_ism_idle                  ),
  .credit_reinit       ( p10_credit_reinit             ),
  .cg_inprogress       ( p10_cg_inprogress             ),
  .tpccup              ( sbr_c_dfx_jtag_pccup          ),
  .tnpcup              ( sbr_c_dfx_jtag_npcup          ),
  .tpcput              ( dfx_jtag_sbr_c_pcput          ),
  .tnpput              ( dfx_jtag_sbr_c_npput          ),
  .teom                ( dfx_jtag_sbr_c_eom            ),
  .tpayload            ( dfx_jtag_sbr_c_payload        ),
  .pctrdy              ( pctrdy[10]                    ),
  .pcirdy              ( pcirdy[10]                    ),
  .pcdata              ( pcdata[10]                    ),
  .pceom               ( pceom[10]                     ),
  .pcdstvld            ( p10_pcdstvld                  ),
  .nptrdy              ( nptrdy[10]                    ),
  .npirdy              ( npirdy[10]                    ),
  .npfence             ( p10_npfence                   ),
  .npdata              ( npdata[10]                    ),
  .npeom               ( npeom[10]                     ),
  .npdstvld            ( p10_npdstvld                  ),
  .mpccup              ( dfx_jtag_sbr_c_pccup          ),
  .mnpcup              ( dfx_jtag_sbr_c_npcup          ),
  .mpcput              ( sbr_c_dfx_jtag_pcput          ),
  .mnpput              ( sbr_c_dfx_jtag_npput          ),
  .meom                ( sbr_c_dfx_jtag_eom            ),
  .mpayload            ( sbr_c_dfx_jtag_payload        ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[10]                   ),
  .enptrdy             ( enptrdy[10]                   ),
  .epcirdy             ( epcirdy[10]                   ),
  .enpirdy             ( enpirdy[10]                   ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p10_dbgbus                    )
);

// Port 11
logic p11_side_clk_valid, p11_idle_egress, p11_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p11_rst_suppress <= 1'b1;
    else
      p11_rst_suppress <= p11_credit_reinit & p11_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p11_fab_init_idle_exit <= '1;
    else
      if ( ~p11_rst_suppress & (p11_ism_idle & (~agent_idle[11] || ~p11_idle_egress) & ~p11_fab_init_idle_exit_ack ))
        p11_fab_init_idle_exit <= '1;
      else if ( ~p11_rst_suppress & (p11_ism_idle & agent_idle[11] & p11_fab_init_idle_exit_ack ))
        p11_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p11_side_clk_valid <= 1'b0;
    else
      begin
        if ( p11_ism_idle & p11_side_clk_valid )
          p11_side_clk_valid <= '0;
        else if ( (p11_fab_init_idle_exit & p11_fab_init_idle_exit_ack) || ~p11_ism_idle )
          p11_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p11_dbgbus;

  always_comb
    begin
      visa_p11_tier1_clk_100 = { p11_dbgbus[31],
                            p11_dbgbus[27:24],
                            p11_dbgbus[21:19],
                            p11_dbgbus[15:12],
                            p11_dbgbus[7:4] };
      visa_p11_tier2_clk_100 = { p11_dbgbus[30:28],
                            p11_dbgbus[23:22],
                            p11_dbgbus[18:16],
                            p11_dbgbus[11:8],
                            p11_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport11 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p11_side_clk_valid            ),
  .side_ism_in         ( itunit_sbr_c_side_ism_agent   ),
  .side_ism_out        ( sbr_c_itunit_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[11] ),
  .agent_idle          ( agent_idle[11]                ),
  .port_idle           ( port_idle[11]                 ),
  .idle_egress         ( p11_idle_egress               ),
  .ism_idle            ( p11_ism_idle                  ),
  .credit_reinit       ( p11_credit_reinit             ),
  .cg_inprogress       ( p11_cg_inprogress             ),
  .tpccup              ( sbr_c_itunit_pccup            ),
  .tnpcup              ( sbr_c_itunit_npcup            ),
  .tpcput              ( itunit_sbr_c_pcput            ),
  .tnpput              ( itunit_sbr_c_npput            ),
  .teom                ( itunit_sbr_c_eom              ),
  .tpayload            ( itunit_sbr_c_payload          ),
  .pctrdy              ( pctrdy[11]                    ),
  .pcirdy              ( pcirdy[11]                    ),
  .pcdata              ( pcdata[11]                    ),
  .pceom               ( pceom[11]                     ),
  .pcdstvld            ( p11_pcdstvld                  ),
  .nptrdy              ( nptrdy[11]                    ),
  .npirdy              ( npirdy[11]                    ),
  .npfence             ( p11_npfence                   ),
  .npdata              ( npdata[11]                    ),
  .npeom               ( npeom[11]                     ),
  .npdstvld            ( p11_npdstvld                  ),
  .mpccup              ( itunit_sbr_c_pccup            ),
  .mnpcup              ( itunit_sbr_c_npcup            ),
  .mpcput              ( sbr_c_itunit_pcput            ),
  .mnpput              ( sbr_c_itunit_npput            ),
  .meom                ( sbr_c_itunit_eom              ),
  .mpayload            ( sbr_c_itunit_payload          ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[11]                   ),
  .enptrdy             ( enptrdy[11]                   ),
  .epcirdy             ( epcirdy[11]                   ),
  .enpirdy             ( enpirdy[11]                   ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p11_dbgbus                    )
);

// Port 12 (Asynchronous port)
logic p12_side_clk_valid, p12_idle_egress, p12_rst_suppress;
  logic p12_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p12_rst_suppress <= 1'b1;
    else
      p12_rst_suppress <= p12_credit_reinit_ff2 & p12_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p12_fab_init_idle_exit <= '1;
    else
      if ( ~p12_rst_suppress & (p12_ism_idle_ff2 & (~agent_idle[12] || ~p12_efifo_idle) & ~p12_fab_init_idle_exit_ack ))
        p12_fab_init_idle_exit <= '1;
      else if ( ~p12_rst_suppress & (p12_ism_idle_ff2 & agent_idle[12] & p12_efifo_idle & p12_fab_init_idle_exit_ack ))
        p12_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p12_side_clk_valid <= 1'b0;
    else
      begin
        if ( p12_ism_idle_ff2 & p12_side_clk_valid & ~p12_fab_init_idle_exit )
          p12_side_clk_valid <= '0;
        else if ( (p12_fab_init_idle_exit & p12_fab_init_idle_exit_ack) || ~p12_ism_idle_ff2 )
          p12_side_clk_valid <= '1;
      end

logic p12_side_clk_valid_ff2;
sbc_doublesync sync_p12_clk_valid (
  .d     ( p12_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p12_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p12_credit_reinit (
  .d     ( p12_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p12_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p12_dbgbus;

logic [15:0] p12_dbgbus_ing;
logic [15:0] p12_dbgbus_egr;
  always_comb
    begin
      visa_p12_tier1_clk_200 = { p12_dbgbus[31],
                            p12_dbgbus[27:24],
                            p12_dbgbus[21:19],
                            p12_dbgbus[15:12],
                            p12_dbgbus[7:4] };
      visa_p12_tier2_clk_200 = { p12_dbgbus[30:28],
                            p12_dbgbus[23:22],
                            p12_dbgbus[18:16],
                            p12_dbgbus[11:8],
                            p12_dbgbus[3:0] };
      visa_p12_ififo_tier1_clk_100 = { p12_dbgbus_ing[15:14],
                             p12_dbgbus_ing[5:0]};
      visa_p12_ififo_tier2_clk_100 = { p12_dbgbus_ing[13:6] };
      visa_p12_efifo_tier1_clk_100 = { p12_dbgbus_egr[7:0] };
      visa_p12_efifo_tier2_clk_100 = { p12_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport12 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p12_gated_clk                 ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p12_side_clk_valid_ff2        ),
  .side_ism_in         ( psf_3_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_psf_3_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[12] ),
  .agent_idle          ( p12_agent_idle                ),
  .port_idle           ( p12_port_idle                 ),
  .idle_egress         (                               ),
  .ism_idle            ( p12_ism_idle                  ),
  .credit_reinit       ( p12_credit_reinit             ),
  .cg_inprogress       ( p12_cg_inprogress             ),
  .tpccup              ( sbr_c_psf_3_pccup             ),
  .tnpcup              ( sbr_c_psf_3_npcup             ),
  .tpcput              ( psf_3_sbr_c_pcput             ),
  .tnpput              ( psf_3_sbr_c_npput             ),
  .teom                ( psf_3_sbr_c_eom               ),
  .tpayload            ( psf_3_sbr_c_payload           ),
  .pctrdy              ( p12_pctrdy                    ),
  .pcirdy              ( p12_pcirdy                    ),
  .pcdata              ( p12_pcdata                    ),
  .pceom               ( p12_pceom                     ),
  .pcdstvld            (                               ),
  .nptrdy              ( p12_nptrdy                    ),
  .npirdy              ( p12_npirdy                    ),
  .npfence             ( p12_npfence                   ),
  .npdata              ( p12_npdata                    ),
  .npeom               ( p12_npeom                     ),
  .npdstvld            (                               ),
  .mpccup              ( psf_3_sbr_c_pccup             ),
  .mnpcup              ( psf_3_sbr_c_npcup             ),
  .mpcput              ( sbr_c_psf_3_pcput             ),
  .mnpput              ( sbr_c_psf_3_npput             ),
  .meom                ( sbr_c_psf_3_eom               ),
  .mpayload            ( sbr_c_psf_3_payload           ),
  .enpstall            ( p12_enpstall                  ),
  .epctrdy             ( p12_epctrdy                   ),
  .enptrdy             ( p12_enptrdy                   ),
  .epcirdy             ( p12_epcirdy                   ),
  .enpirdy             ( p12_enpirdy                   ),
  .data                ( p12_data                      ),
  .eom                 ( p12_eom                       ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p12_clkgaten                  ),
  .force_idle          ( p12_force_idle                ),
  .force_notidle       ( p12_force_notidle             ),
  .force_creditreq     ( p12_force_creditreq           ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p12_dbgbus                    )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress12 (
  .ing_side_clk        ( p12_gated_clk                 ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p12_port_idle                 ),
  .pcirdy              ( p12_pcirdy                    ),
  .npirdy              ( p12_npirdy                    ),
  .npfence             ( p12_npfence                   ),
  .pceom               ( p12_pceom                     ),
  .pcdata              ( p12_pcdata                    ),
  .npeom               ( p12_npeom                     ),
  .npdata              ( p12_npdata                    ),
  .pctrdy              ( p12_pctrdy                    ),
  .nptrdy              ( p12_nptrdy                    ),
  .npstall             (                               ),
  .fifo_idle           ( p12_ififo_idle                ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[12]                    ),
  .enptrdy             ( nptrdy[12]                    ),
  .epcirdy             ( pcirdy[12]                    ),
  .enpirdy             ( npirdy[12]                    ),
  .eom                 ( npeom[12]                     ),
  .data                ( npdata[12]                    ),
  .opceom              ( pceom[12]                     ),
  .opcdata             ( pcdata[12]                    ),
  .agent_idle          ( port_idle[12]                 ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p12_dbgbus_ing                )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  2                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress12 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[12]                ),
  .pcirdy              ( epcirdy[12]                   ),
  .npirdy              ( enpirdy[12]                   ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[12]                   ),
  .nptrdy              ( enptrdy[12]                   ),
  .npstall             (                               ),
  .fifo_idle           ( p12_efifo_idle                ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p12_gated_clk                 ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p12_enpstall                  ),
  .epctrdy             ( p12_epctrdy                   ),
  .enptrdy             ( p12_enptrdy                   ),
  .epcirdy             ( p12_epcirdy                   ),
  .enpirdy             ( p12_enpirdy                   ),
  .eom                 ( p12_eom                       ),
  .data                ( p12_data                      ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p12_eagent_idle               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p12_dbgbus_egr                ),
  .dbgbus_out          (                               )
);

always_comb p12_agent_idle  = p12_eagent_idle & p12_ififo_idle;

// Port 13
logic p13_side_clk_valid, p13_idle_egress, p13_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p13_rst_suppress <= 1'b1;
    else
      p13_rst_suppress <= p13_credit_reinit & p13_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p13_fab_init_idle_exit <= '1;
    else
      if ( ~p13_rst_suppress & (p13_ism_idle & (~agent_idle[13] || ~p13_idle_egress) & ~p13_fab_init_idle_exit_ack ))
        p13_fab_init_idle_exit <= '1;
      else if ( ~p13_rst_suppress & (p13_ism_idle & agent_idle[13] & p13_fab_init_idle_exit_ack ))
        p13_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p13_side_clk_valid <= 1'b0;
    else
      begin
        if ( p13_ism_idle & p13_side_clk_valid )
          p13_side_clk_valid <= '0;
        else if ( (p13_fab_init_idle_exit & p13_fab_init_idle_exit_ack) || ~p13_ism_idle )
          p13_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p13_dbgbus;

  always_comb
    begin
      visa_p13_tier1_clk_100 = { p13_dbgbus[31],
                            p13_dbgbus[27:24],
                            p13_dbgbus[21:19],
                            p13_dbgbus[15:12],
                            p13_dbgbus[7:4] };
      visa_p13_tier2_clk_100 = { p13_dbgbus[30:28],
                            p13_dbgbus[23:22],
                            p13_dbgbus[18:16],
                            p13_dbgbus[11:8],
                            p13_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport13 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( p13_gated_clk                 ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p13_side_clk_valid            ),
  .side_ism_in         ( SAPms_sbr_c_side_ism_agent    ),
  .side_ism_out        ( sbr_c_SAPms_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[13] ),
  .agent_idle          ( agent_idle[13]                ),
  .port_idle           ( port_idle[13]                 ),
  .idle_egress         ( p13_idle_egress               ),
  .ism_idle            ( p13_ism_idle                  ),
  .credit_reinit       ( p13_credit_reinit             ),
  .cg_inprogress       ( p13_cg_inprogress             ),
  .tpccup              ( sbr_c_SAPms_pccup             ),
  .tnpcup              ( sbr_c_SAPms_npcup             ),
  .tpcput              ( SAPms_sbr_c_pcput             ),
  .tnpput              ( SAPms_sbr_c_npput             ),
  .teom                ( SAPms_sbr_c_eom               ),
  .tpayload            ( SAPms_sbr_c_payload           ),
  .pctrdy              ( pctrdy[13]                    ),
  .pcirdy              ( pcirdy[13]                    ),
  .pcdata              ( pcdata[13]                    ),
  .pceom               ( pceom[13]                     ),
  .pcdstvld            ( p13_pcdstvld                  ),
  .nptrdy              ( nptrdy[13]                    ),
  .npirdy              ( npirdy[13]                    ),
  .npfence             ( p13_npfence                   ),
  .npdata              ( npdata[13]                    ),
  .npeom               ( npeom[13]                     ),
  .npdstvld            ( p13_npdstvld                  ),
  .mpccup              ( SAPms_sbr_c_pccup             ),
  .mnpcup              ( SAPms_sbr_c_npcup             ),
  .mpcput              ( sbr_c_SAPms_pcput             ),
  .mnpput              ( sbr_c_SAPms_npput             ),
  .meom                ( sbr_c_SAPms_eom               ),
  .mpayload            ( sbr_c_SAPms_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[13]                   ),
  .enptrdy             ( enptrdy[13]                   ),
  .epcirdy             ( epcirdy[13]                   ),
  .enpirdy             ( enpirdy[13]                   ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p13_dbgbus                    )
);

// Port 14
logic p14_side_clk_valid, p14_idle_egress, p14_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p14_rst_suppress <= 1'b1;
    else
      p14_rst_suppress <= p14_credit_reinit & p14_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p14_fab_init_idle_exit <= '1;
    else
      if ( ~p14_rst_suppress & (p14_ism_idle & (~agent_idle[14] || ~p14_idle_egress) & ~p14_fab_init_idle_exit_ack ))
        p14_fab_init_idle_exit <= '1;
      else if ( ~p14_rst_suppress & (p14_ism_idle & agent_idle[14] & p14_fab_init_idle_exit_ack ))
        p14_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p14_side_clk_valid <= 1'b0;
    else
      begin
        if ( p14_ism_idle & p14_side_clk_valid )
          p14_side_clk_valid <= '0;
        else if ( (p14_fab_init_idle_exit & p14_fab_init_idle_exit_ack) || ~p14_ism_idle )
          p14_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p14_dbgbus;

  always_comb
    begin
      visa_p14_tier1_clk_100 = { p14_dbgbus[31],
                            p14_dbgbus[27:24],
                            p14_dbgbus[21:19],
                            p14_dbgbus[15:12],
                            p14_dbgbus[7:4] };
      visa_p14_tier2_clk_100 = { p14_dbgbus[30:28],
                            p14_dbgbus[23:22],
                            p14_dbgbus[18:16],
                            p14_dbgbus[11:8],
                            p14_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport14 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p14_side_clk_valid            ),
  .side_ism_in         ( itunit2_sbr_c_side_ism_agent  ),
  .side_ism_out        ( sbr_c_itunit2_side_ism_fabric ),
  .int_pok             ( endpoint_pwrgd[14] ),
  .agent_idle          ( agent_idle[14]                ),
  .port_idle           ( port_idle[14]                 ),
  .idle_egress         ( p14_idle_egress               ),
  .ism_idle            ( p14_ism_idle                  ),
  .credit_reinit       ( p14_credit_reinit             ),
  .cg_inprogress       ( p14_cg_inprogress             ),
  .tpccup              ( sbr_c_itunit2_pccup           ),
  .tnpcup              ( sbr_c_itunit2_npcup           ),
  .tpcput              ( itunit2_sbr_c_pcput           ),
  .tnpput              ( itunit2_sbr_c_npput           ),
  .teom                ( itunit2_sbr_c_eom             ),
  .tpayload            ( itunit2_sbr_c_payload         ),
  .pctrdy              ( pctrdy[14]                    ),
  .pcirdy              ( pcirdy[14]                    ),
  .pcdata              ( pcdata[14]                    ),
  .pceom               ( pceom[14]                     ),
  .pcdstvld            ( p14_pcdstvld                  ),
  .nptrdy              ( nptrdy[14]                    ),
  .npirdy              ( npirdy[14]                    ),
  .npfence             ( p14_npfence                   ),
  .npdata              ( npdata[14]                    ),
  .npeom               ( npeom[14]                     ),
  .npdstvld            ( p14_npdstvld                  ),
  .mpccup              ( itunit2_sbr_c_pccup           ),
  .mnpcup              ( itunit2_sbr_c_npcup           ),
  .mpcput              ( sbr_c_itunit2_pcput           ),
  .mnpput              ( sbr_c_itunit2_npput           ),
  .meom                ( sbr_c_itunit2_eom             ),
  .mpayload            ( sbr_c_itunit2_payload         ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[14]                   ),
  .enptrdy             ( enptrdy[14]                   ),
  .epcirdy             ( epcirdy[14]                   ),
  .enpirdy             ( enpirdy[14]                   ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p14_dbgbus                    )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_c_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_c_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk_100 or negedge rst_b_100)

      if (~rst_b_100) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 1, clk_100, rst_b_100, 0, , 5ns
ClockReset, 0, clk_200, rst_b_200, 0, , 2.5ns
ClockReset, 2, clk_27, rst_b_27, 0, , 18.5ns
Endpoint, SAPms,3, 1, 1, 0, 3, 3, 1, 65, 2, 2, 
Endpoint, adac,0, 1, 1, 0, 3, 3, 1, 129, 2, 2, 
Endpoint, apll,0, 1, 2, 0, 3, 3, 1, 139, 2, 2, 
Endpoint, bunit,2, 1, 0, 0, 3, 3, 1, 03, 2, 2, 
Endpoint, cpunit,2, 1, 1, 0, 3, 3, 1, 10, 2, 2, 
Endpoint, cunit,2, 1, 0, 0, 3, 3, 1, 07, 2, 2, 
Endpoint, ddrio,2, 1, 1, 0, 3, 3, 1, 80, 2, 2, 
Endpoint, dfx_jtag,2, 1, 1, 0, 3, 3, 1, 58, 2, 2, 
Endpoint, dfx_lakemore,2, 1, 1, 0, 3, 3, 1, 56, 2, 2, 
Endpoint, dfx_omar,2, 1, 1, 0, 3, 3, 1, 57, 2, 2, 
Endpoint, dpll,0, 1, 2, 0, 3, 3, 1, 138, 2, 2, 
Endpoint, fpll,0, 1, 2, 0, 3, 3, 1, 136, 2, 2, 
Endpoint, hdmi_rx,0, 1, 1, 0, 3, 3, 1, 131, 2, 2, 
Endpoint, hdmi_tx,0, 1, 1, 0, 3, 3, 1, 130, 2, 2, 
Endpoint, hpll,0, 1, 2, 0, 3, 3, 1, 137, 2, 2, 
Endpoint, hunit,2, 1, 0, 0, 3, 3, 1, 02, 2, 2, 
Endpoint, itunit,2, 1, 1, 0, 3, 3, 1, 64, 2, 2, 
Endpoint, itunit2,2, 1, 1, 0, 3, 3, 1, 66, 2, 2, 
Endpoint, legacy,2, 1, 1, 0, 3, 3, 10, 11,12,13,32,33,34,35,36,37,38, 2, 2, 
Endpoint, mcu,2, 1, 0, 0, 3, 3, 1, 01, 2, 2, 
Endpoint, pcie_afe,4, 1, 1, 0, 3, 3, 1, 17, 2, 2, 
Endpoint, pcie_ctrl,4, 1, 1, 0, 3, 3, 1, 16, 2, 2, 
Endpoint, psf_0_north,4, 1, 0, 0, 3, 3, 1, 50, 2, 2, 
Endpoint, psf_0_south,4, 1, 1, 0, 3, 3, 1, 144, 2, 2, 
Endpoint, psf_1,4, 1, 0, 0, 3, 3, 1, 145, 2, 2, 
Endpoint, psf_3,2, 1, 0, 0, 3, 3, 1, 147, 2, 2, 
Endpoint, punit,1, 1, 2, 0, 3, 3, 1, 04, 2, 2, 
Endpoint, reut_0,2, 1, 1, 0, 3, 3, 1, 84, 2, 2, 
Endpoint, reut_1,2, 1, 1, 0, 3, 3, 1, 85, 2, 2, 
Endpoint, sata_afe,4, 1, 1, 0, 3, 3, 1, 89, 2, 2, 
Endpoint, sata_ctrl,4, 1, 1, 0, 3, 3, 1, 88, 2, 2, 
SyncRouter, sbr_a, sbr_a,1, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 2, 8, sbr_e, sbr_b, sbr_c, dpll, apll, hpll, fpll, punit, , , , , , , , , 
RouterAgentPort, sbr_a, 0
RouterAgentPort, sbr_a, 1
RouterAgentPort, sbr_a, 2
RouterRange, sbr_a, 0, 48,49
SyncRouter, sbr_b, sbr_b,4, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 9, sbr_a, pcie_afe, sata_afe, usb_afe, sata_ctrl, pcie_ctrl, psf_1, psf_0_south, psf_0_north, , , , , , , , 
RouterRange, sbr_b, 0, 51,51
SyncRouter, sbr_c, sbr_c,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 15, sbr_a, sbr_d, vtunit, hunit, bunit, cunit, cpunit, legacy, dfx_lakemore, dfx_omar, dfx_jtag, itunit, psf_3, SAPms, itunit2, , 
RouterAgentPort, sbr_c, 1
RouterRange, sbr_c, 0, 52,52
SyncRouter, sbr_d, sbr_d,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_c, mcu, ddrio, reut_0, reut_1, , , , , , , , , , , , 
RouterRange, sbr_d, 0, 54,55
SyncRouter, sbr_e, sbr_e,5, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_a, vdac, adac, hdmi_tx, hdmi_rx, , , , , , , , , , , , 
Endpoint, usb_afe,4, 1, 1, 0, 3, 3, 1, 96, 2, 2, 
Endpoint, vdac,0, 1, 1, 0, 3, 3, 1, 128, 2, 2, 
Endpoint, vtunit,2, 1, 0, 0, 3, 3, 1, 00, 2, 2, 
AsyncPort, sbr_a, 0, 10, 4, 0, 
AsyncPort, sbr_a, 1, 10, 4, 0, 
AsyncPort, sbr_a, 2, 10, 4, 0, 
AsyncPort, sbr_b, 6, 4, 2, 0, 
AsyncPort, sbr_b, 8, 4, 2, 0, 
AsyncPort, sbr_c, 12, 4, 2, 0, 
AsyncPort, sbr_c, 2, 10, 4, 0, 
AsyncPort, sbr_c, 3, 10, 4, 0, 
AsyncPort, sbr_c, 4, 10, 4, 0, 
AsyncPort, sbr_c, 5, 10, 4, 0, 
AsyncPort, sbr_d, 1, 10, 4, 0, 
PowerWell, 0, 
PowerWell, 1, island0_pok
PowerWell, 2, island1_pok
PowerWell, 3, island2_pok
PowerWell, 4, island3_pok
PowerWell, 5, island8_pok
*/
//------------------------------------------------------------------------------
