
`ifndef INTEL_SVA_OFF

`ifndef HQM_TB_DEFINES
`include "hqm_tb_defines.sv"
`define HQM_TB_DEFINES
`endif

module hqm_assert import hqm_AW_pkg::*, hqm_pkg::*, hqm_core_pkg::*;  ();

  // Insert assertion code here
  // Refer to signals defined in hqm with proper prefix from hqm_tb_defines

`ifdef HQM_MPP
////////////////////////////////////////////////////////////////////////////////////////////////////
//mem_fet_en_b connection ring START
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_0, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_ack_b), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_0 `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_ack_b Not Connected"), SDG_SVA_SOC_SIM) ;
`ifndef HQM_7NM
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_1, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fid_cnt.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_1 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fid_cnt.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_2, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fid_cnt.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_2 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fid_cnt.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_3, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_ap_aqed.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_3 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_ap_aqed.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_4, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_aqed_ap_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_4 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_aqed_ap_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_5, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_aqed_chp_sch.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_5 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_aqed_chp_sch.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_6, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_freelist_return.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_6 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_freelist_return.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_7, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_7 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_lsp_aqed_cmp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_8, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_qed_aqed_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_8 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_qed_aqed_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_9, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_9 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_fifo_qed_aqed_enq_fid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_10, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_10 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_11, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_11 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_12, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_12 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_13, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_13 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_14, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_14 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_15, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_15 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_16, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_16 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_17, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_17 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_cnt_pri3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_18, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_18 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_19, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_19 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_20, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_20 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_21, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_21 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_22, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_22 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_23, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_23 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_24, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_24 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_25, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_25 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_hp_pri3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_26, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_26 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_27, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_27 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_28, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_28 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_29, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_29 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_30, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_30 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_31, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_31 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_32, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_32 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_33, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_33 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_ll_qe_tp_pri3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_34, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_lsp_deq_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_34 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_lsp_deq_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_35, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_35 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_36, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_36 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_37, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b2.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_37 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b2.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_38, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b3.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_38 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid2cqidix.i_rf_b3.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_39, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_39 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_40, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid_fid_limit.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_40 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_aqed_qid_fid_limit.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_41, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_cmp_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_41 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_cmp_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_42, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_fifo_ap_aqed.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_42 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_fifo_ap_aqed.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_43, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_fifo_aqed_ap_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_43 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_atm_fifo_aqed_ap_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_44, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_atm_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_44 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_atm_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_45, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2priov_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_45 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2priov_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_46, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2priov_odd_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_46 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2priov_odd_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_47, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_0_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_47 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_0_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_48, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_0_odd_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_48 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_0_odd_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_49, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_1_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_49 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_1_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_50, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_1_odd_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_50 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq2qid_1_odd_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_51, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_inflight_limit_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_51 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_inflight_limit_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_52, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_inflight_threshold_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_52 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_inflight_threshold_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_53, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_token_depth_select_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_53 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_token_depth_select_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_54, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_54 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_cq_ldb_wu_limit_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_55, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_dir_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_55 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_dir_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_56, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_nalb_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_56 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_nalb_qid_dpth_thrsh_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_57, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_aqed_active_limit_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_57 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_aqed_active_limit_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_58, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_inflight_limit_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_58 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_inflight_limit_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_59, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_59 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_60, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_60 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_61, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_61 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b2.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_62, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_62 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix2_mem.i_rf_b3.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_63, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_63 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_64, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_64 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_65, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_65 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b2.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_66, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_66 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cfg_qid_ldb_qid2cqidix_mem.i_rf_b3.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_67, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_67 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_cmp_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_68, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_68 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_token_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_69, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_atm_pri_arbindex_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_69 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_atm_pri_arbindex_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_70, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_70 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_dir_tot_sch_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_71, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_inflight_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_71 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_inflight_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_72, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_token_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_72 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_token_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_73, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_73 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_tot_sch_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_74, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_wu_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_74 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_ldb_wu_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_75, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_nalb_pri_arbindex_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_75 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_cq_nalb_pri_arbindex_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_76, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_enq_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_76 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_enq_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_77, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_tok_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_77 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_tok_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_78, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_tok_lim_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_78 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dir_tok_lim_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_79, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_79 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_dir_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_80, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_80 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_81, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_enq_nalb_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_81 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_enq_nalb_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_82, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_fid2cqqidix.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_82 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_fid2cqqidix.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_83, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_fid2cqqidix.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_83 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_fid2cqqidix.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_84, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ldb_token_rtn_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_84 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ldb_token_rtn_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_85, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_85 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_86, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_86 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_87, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_87 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_88, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_88 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_89, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_89 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_90, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_90 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_91, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_91 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_92, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_92 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin0_dup3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_93, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_93 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_94, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_94 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_95, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_95 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_96, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_96 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_97, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_97 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_98, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_98 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_99, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_99 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_100, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_100 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin1_dup3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_101, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_101 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_102, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_102 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_103, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_103 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_104, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_104 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_105, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_105 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_106, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_106 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_107, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_107 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_108, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_108 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin2_dup3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_109, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_109 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_110, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_110 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_111, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_111 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_112, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_112 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_113, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_113 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_114, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_114 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_115, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_115 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_116, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_116 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_r_bin3_dup3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_117, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_117 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_118, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_118 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_119, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_119 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_120, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_120 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_121, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_121 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_122, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_122 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_123, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_123 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_124, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_124 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_enq_cnt_s_bin3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_125, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_125 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_126, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_126 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_127, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_127 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_128, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin3.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_128 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hp_bin3.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_129, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_129 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_130, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_130 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_131, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_131 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_132, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_132 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_133, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_133 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_134, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_134 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_135, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_135 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_136, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_136 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_hpnxt_bin3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_137, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_137 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_138, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_138 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_139, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_139 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_140, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin3.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_140 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rdylst_tp_bin3.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_141, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rlst_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_141 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_rlst_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_142, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_142 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_143, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_143 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_144, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_144 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_145, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_145 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_146, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_146 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_147, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_147 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_148, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_148 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_149, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_149 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_sch_cnt_dup3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_150, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_150 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_151, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_151 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_152, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_152 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_153, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin3.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_153 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hp_bin3.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_154, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_154 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_155, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_155 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_156, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_156 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_157, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_157 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_158, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_158 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_159, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_159 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_160, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_160 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_161, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_161 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_hpnxt_bin3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_162, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_162 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_163, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_163 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_164, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_164 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_165, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin3.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_165 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tp_bin3.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_166, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_166 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin0.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_167, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_167 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin0.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_168, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_168 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin1.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_169, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_169 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin1.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_170, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_170 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin2.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_171, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_171 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin2.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_172, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_172 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin3.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_173, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_173 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_schlst_tpprv_bin3.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_174, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_slst_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_174 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_ll_slst_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_175, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_cmp_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_175 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_cmp_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_176, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_176 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_177, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_177 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_178, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_sel_nalb_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_178 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_nalb_sel_nalb_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_179, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qed_lsp_deq_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_179 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qed_lsp_deq_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_180, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_aqed_active_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_180 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_aqed_active_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_181, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atm_active_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_181 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atm_active_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_182, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_182 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atm_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_183, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atq_enqueue_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_183 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_atq_enqueue_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_184, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_max_depth_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_184 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_max_depth_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_185, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_replay_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_185 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_replay_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_186, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_186 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_dir_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_187, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_enqueue_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_187 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_enqueue_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_188, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_inflight_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_188 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_inflight_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_189, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_replay_count_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_189 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_ldb_replay_count_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_190, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_naldb_max_depth_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_190 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_naldb_max_depth_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_191, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_191 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_naldb_tot_enq_cnt_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_192, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_rdylst_clamp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_192 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_qid_rdylst_clamp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_193, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_193 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_rop_lsp_reordercmp_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_194, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_qed_aqed_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_194 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_qed_aqed_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_195, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_195 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_send_atm_to_cq_rx_sync_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_196, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_uno_atm_cmp_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_196 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_rf_pg_cont.i_rf_uno_atm_cmp_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_197, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_197 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_198, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_198 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_199, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed_freelist.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_199 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed_freelist.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_200, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed_ll_qe_hpnxt.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_200 `HQM_LIST_SEL_MEM_PATH.i_hqm_list_sel_mem_hqm_clk_sram_pg_cont.i_sr_aqed_ll_qe_hpnxt.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_201, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_201 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_202, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_202 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_203, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_203 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_atq_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_204, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_204 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_205, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_205 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_206, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_206 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_207, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_207 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_208, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_208 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_replay_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_209, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_209 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_210, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_210 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_211, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_211 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_rofrag_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_212, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_212 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dir_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_213, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_dqed.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_213 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_dqed.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_214, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_dir.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_214 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_dir.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_215, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_215 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_dp_lsp_enq_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_216, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_dp_sch_dir.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_216 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_dp_sch_dir.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_217, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_dp_sch_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_217 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_dp_sch_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_218, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_atq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_218 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_atq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_219, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_219 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_220, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_unoord.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_220 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_lsp_nalb_sch_unoord.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_221, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_221 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_222, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_222 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_223, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_223 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_224, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_unoord.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_224 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_lsp_enq_unoord.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_225, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_qed.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_225 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_qed.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_226, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_226 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_227, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_227 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_228, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_228 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_replay_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_229, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_cnt.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_229 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_cnt.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_230, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_hp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_230 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_hp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_231, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_231 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_rofrag_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_232, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_tp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_232 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_nalb_tp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_233, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_data.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_233 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_data.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_234, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_dp_enq_dir.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_234 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_dp_enq_dir.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_235, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_dp_enq_ro.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_235 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_dp_enq_ro.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_236, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_nalb_enq_ro.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_236 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_nalb_enq_ro.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_237, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_nalb_enq_unoord.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_237 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rop_nalb_enq_unoord.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_238, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_dp_dqed_data.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_238 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_dp_dqed_data.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_239, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_239 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_dp_sch_dir.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_240, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_240 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_dp_sch_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_241, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_241 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_atq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_242, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_242 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_rorply.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_243, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_243 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_lsp_nalb_sch_unoord.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_244, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_nalb_qed_data.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_244 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_nalb_qed_data.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_245, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_dp_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_245 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_dp_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_246, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_nalb_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_246 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_nalb_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_247, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_247 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_rf_pg_cont.i_rf_rx_sync_rop_qed_dqed_enq.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_248, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_248 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_249, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_249 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_250, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b2.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_250 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b2.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_251, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b3.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_251 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_dir_nxthp.i_sram_b3.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_252, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_252 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_253, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_253 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_254, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b2.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_254 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b2.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_255, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b3.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_255 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_nalb_nxthp.i_sram_b3.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_256, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_0.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_256 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_0.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_257, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_0.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_257 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_0.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_258, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_1.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_258 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_1.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_259, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_1.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_259 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_1.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_260, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_2.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_260 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_2.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_261, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_2.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_261 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_2.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_262, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_3.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_262 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_3.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_263, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_3.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_263 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_3.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_264, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_4.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_264 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_4.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_265, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_4.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_265 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_4.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_266, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_5.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_266 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_5.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_267, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_5.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_267 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_5.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_268, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_6.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_268 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_6.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_269, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_6.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_269 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_6.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_270, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_7.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_270 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_7.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_271, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_7.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_271 `HQM_QED_MEM_PATH.i_hqm_qed_mem_hqm_clk_sram_pg_cont.i_sr_qed_7.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_272, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_272 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_273, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_273 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_274, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_274 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_alarm_vf_synd2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_275, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_aqed_chp_sch_rx_sync_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_275 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_aqed_chp_sch_rx_sync_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_276, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_chp_rop_hcw_fifo_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_276 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_chp_rop_hcw_fifo_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_277, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_chp_rop_hcw_fifo_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_277 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_chp_rop_hcw_fifo_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_278, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_278 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_ap_cmp_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_279, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_tok_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_279 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_lsp_tok_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_280, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_280 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_sys_tx_fifo_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_281, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_281 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_chp_sys_tx_fifo_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_282, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_cmp_id_chk_enbl_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_282 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_cmp_id_chk_enbl_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_283, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_count_rmw_pipe_dir_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_283 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_count_rmw_pipe_dir_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_284, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_count_rmw_pipe_ldb_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_284 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_count_rmw_pipe_ldb_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_285, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_depth.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_285 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_depth.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_286, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_intr_thresh.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_286 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_intr_thresh.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_287, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_token_depth_select.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_287 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_token_depth_select.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_288, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_wptr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_288 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_cq_wptr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_289, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_rply_req_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_289 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_rply_req_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_290, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_290 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_291, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_291 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_292, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_292 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_dir_wb2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_293, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hcw_enq_w_rx_sync_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_293 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hcw_enq_w_rx_sync_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_294, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_a_minmax.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_294 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_a_minmax.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_295, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_a_ptr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_295 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_a_ptr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_296, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_minmax.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_296 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_minmax.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_297, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_ptr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_297 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_hist_list_ptr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_298, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_depth.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_298 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_depth.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_299, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_intr_thresh.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_299 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_intr_thresh.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_300, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_on_off_threshold.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_300 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_on_off_threshold.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_301, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_token_depth_select.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_301 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_token_depth_select.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_302, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_wptr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_302 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_cq_wptr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_303, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_rply_req_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_303 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_rply_req_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_304, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_304 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_305, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_305 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_306, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_306 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ldb_wb2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_307, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lsp_reordercmp_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_307 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lsp_reordercmp_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_308, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq2vf_pf_ro.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_308 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq2vf_pf_ro.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_309, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_addr_l.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_309 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_addr_l.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_310, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_addr_u.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_310 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_addr_u.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_311, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_addr_l.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_311 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_addr_l.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_312, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_addr_u.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_312 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_addr_u.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_313, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_data.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_313 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_ai_data.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_314, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_isr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_314 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_isr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_315, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_pasid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_315 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_cq_pasid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_316, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_pp2vas.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_316 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_pp2vas.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_317, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_pp_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_317 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_pp_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_318, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_vasqid_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_318 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_dir_vasqid_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_319, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq2vf_pf_ro.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_319 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq2vf_pf_ro.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_320, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_addr_l.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_320 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_addr_l.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_321, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_addr_u.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_321 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_addr_u.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_322, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_addr_l.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_322 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_addr_l.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_323, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_addr_u.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_323 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_addr_u.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_324, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_data.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_324 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_ai_data.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_325, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_isr.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_325 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_isr.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_326, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_pasid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_326 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_cq_pasid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_327, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_pp2vas.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_327 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_pp2vas.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_328, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_qid2vqid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_328 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_qid2vqid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_329, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_vasqid_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_329 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_ldb_vasqid_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_330, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vpp2pp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_330 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vpp2pp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_331, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vpp_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_331 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vpp_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_332, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vqid2qid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_332 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vqid2qid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_333, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vqid_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_333 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_dir_vqid_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_334, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vpp2pp.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_334 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vpp2pp.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_335, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vpp_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_335 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vpp_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_336, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vqid2qid.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_336 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vqid2qid.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_337, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vqid_v.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_337 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_lut_vf_ldb_vqid_v.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_338, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word0.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_338 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word0.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_339, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word1.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_339 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word1.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_340, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word2.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_340 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_msix_tbl_word2.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_341, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ord_qid_sn.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_341 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ord_qid_sn.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_342, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ord_qid_sn_map.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_342 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_ord_qid_sn_map.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_343, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_outbound_hcw_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_343 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_outbound_hcw_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_344, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_344 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_flid_ret_rx_sync_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_345, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_rx_sync_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_345 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_chp_sch_rx_sync_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_346, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_to_cq_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_346 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_qed_to_cq_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_347, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_cnt_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_347 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_cnt_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_348, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_cnt_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_348 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_cnt_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_349, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirhp_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_349 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirhp_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_350, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirhp_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_350 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirhp_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_351, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirtp_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_351 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirtp_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_352, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirtp_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_352 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_dirtp_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_353, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbhp_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_353 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbhp_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_354, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbhp_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_354 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbhp_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_355, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbtp_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_355 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbtp_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_356, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbtp_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_356 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_lbtp_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_357, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_st_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_357 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_st_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_358, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_st_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_358 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_reord_st_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_359, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_rop_chp_rop_hcw_fifo_mem.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_359 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_rop_chp_rop_hcw_fifo_mem.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_360, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_rop_chp_rop_hcw_fifo_mem.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_360 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_rop_chp_rop_hcw_fifo_mem.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_361, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sch_out_fifo.i_rf_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_361 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sch_out_fifo.i_rf_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_362, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sch_out_fifo.i_rf_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_362 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sch_out_fifo.i_rf_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_363, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn0_order_shft_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_363 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn0_order_shft_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_364, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn1_order_shft_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_364 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn1_order_shft_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_365, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn_complete_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_365 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn_complete_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_366, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn_ordered_fifo_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_366 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_sn_ordered_fifo_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_367, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_threshold_r_pipe_dir_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_367 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_threshold_r_pipe_dir_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_368, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_threshold_r_pipe_ldb_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_368 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_rf_pg_cont.i_rf_threshold_r_pipe_ldb_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_369, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_0.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_369 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_0.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_370, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_1.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_370 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_1.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_371, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_2.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_371 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_2.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_372, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_3.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_372 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_3.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_373, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_4.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_373 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_4.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_374, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_5.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_374 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_5.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_375, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_6.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_375 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_6.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_376, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_7.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_376 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_freelist_7.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_377, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_hist_list.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_377 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_hist_list.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_378, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_hist_list_a.i_sram.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_378 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_hist_list_a.i_sram.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_379, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_rob_mem.i_sram_b0.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_379 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_rob_mem.i_sram_b0.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_380, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_rob_mem.i_sram_b1.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_380 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_hqm_clk_sram_pg_cont.i_sr_rob_mem.i_sram_b1.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_381, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_pgcb_clk_rf_pg_cont.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_381 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_pgcb_clk_rf_pg_cont.i_rf_count_rmw_pipe_wd_dir_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_382, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_pgcb_clk_rf_pg_cont.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_382 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_pgcb_clk_rf_pg_cont.i_rf_count_rmw_pipe_wd_ldb_mem.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`HQM_SDG_ASSERTS_FORBIDDEN( PGCB_MEM_FET_EN_383, (`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_pm_unit.pgcb_fet_en_b != `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_prim_clk_rf_dc_pg_cont.i_rf_hcw_enq_fifo.i_rf.PWR_MGMT_OUT), `HQM_SIF_PATH.prim_freerun_clk, `HQM_SIF_PATH.prim_gated_rst_b, `HQM_SVA_ERR_MSG("PGCB_MEM_FET_EN_383 `HQM_SYSTEM_MEM_PATH.i_hqm_system_mem_prim_clk_rf_dc_pg_cont.i_rf_hcw_enq_fifo.i_rf.PWR_MGMT_OUT Not Connected"), SDG_SVA_SOC_SIM) ;
`endif
//mem_fet_en_b connection ring END
`endif



////////////////////////////////////////////////////////////////////////////////////////////////////
//CFG access & not pipedile

logic chp_collision_mask ;

assign chp_collision_mask = 1'b0 ; 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_chp
                      , (   ( `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.cfg_unit_idle_reg_f.pipe_idle === 1'b0 )
                          & ( `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                          & ~ chp_collision_mask
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_chp: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_rop
                      , (   ( `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_reorder_pipe_func.cfg_unit_idle_f.pipe_idle === 1'b0 )
                          & ( `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_rop: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_ap
                      , (   ( `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.cfg_unit_idle_f.pipe_idle === 1'b0 )
                          & ( `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_ap: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_aqed
                      , (   ( `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.cfg_unit_idle_f.pipe_idle === 1'b0 )
                          & ( `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_aqed: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_qed
                      , (   ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.cfg_unit_idle_reg_f.pipe_idle === 1'b0 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_qed: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_nalb
                      , (   ( ~`HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_nalb_pipe_core.cfg_unit_idle_f.pipe_idle === 1'b0 )
                          & ( ~`HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_nalb_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_nalb_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_nalb_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~`HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_nalb: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_collision_dp
                      , (   ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_dir_pipe_core.cfg_unit_idle_f.pipe_idle === 1'b0 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_dir_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.err === 1'b0 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_dir_pipe_core.i_hqm_AW_cfg_sc.ctrl_f.idlepipe === 1'b1 )
                          & ( `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.i_hqm_dir_pipe_core.i_hqm_AW_cfg_sc.assert_working_nc === 1'b1 )
                        )
                      , posedge `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_clk
                      , ~ `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.i_hqm_cfg_master_sys2cfg.prim_gated_rst_b_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_collision_dp: cfg request issued when pipe is active" )
                      , SDG_SVA_SOC_SIM) 


////////////////////////////////////////////////////////////////////////////////////////////////////
// Check that hqm_gated_rst_b width is wide enough to be synchronized to slower pgcb_clk domain
`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_hqm_gated_rst_b_sync_pgcb_clk
                      , ( 
                          ( $rose(`HQM_MASTER_PATH.hqm_gated_rst_b) & `HQM_CHP_HQM_GATED_RST_PGCB_SYNC_N_PATH.rst_n_sync)
                        )
                      , posedge `HQM_SIF_PATH.pgcb_clk
                      , ~`HQM_MASTER_HQM_CLK_RPTR_RST_SYNC_N_PATH.rst_n_sync
                      , `HQM_SVA_ERR_MSG( "Error: par_hqm_system.sv  assert_forbidden_hqm_gated_rst_b_sync_pgcb_clk: hqm_gated_rst_b pulse width not sufficient for synchronization to pgcb_clk " )
                      , SDG_SVA_SOC_SIM)
////////////////////////////////////////////////////////////////////////////////////////////////////
`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_hqm_cdc_clk_isolation_on_with_rcb_and_lcb_set
                      , (
                          ( ~`HQM_MASTER_PATH.pgcb_isol_en_b  & `HQM_MASTER_HQM_CLK_RPTR_RST_SYNC_N_PATH.rst_n_sync & `HQM_MASTER_HQM_CDC_CLK_ENABLE_RPTR_PATH.data_q)
                        )
                      , posedge `HQM_MASTER_PATH.hqm_fullrate_clk
                      , ~`HQM_MASTER_HQM_CLK_RPTR_RST_SYNC_N_PATH.rst_n_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_hqm_cdc_clk_isolation_on_with_rcb_or_lcb_set: clock_enable while isolation active " )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_hqm_freerun_clk_isolation_on_with_rcb_set
                      , (
                          ( ~`HQM_MASTER_PATH.pgcb_isol_en_b  & `HQM_MASTER_HQM_FREERUN_CLK_ENABLE_RPTR_PATH.data_q )
                        )
                      , posedge `HQM_MASTER_PATH.hqm_fullrate_clk
                      , ~`HQM_MASTER_HQM_CLK_RPTR_RST_SYNC_N_PATH.rst_n_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_hqm_freerun_clk_isolation_on_with_lcb_or_lcb_set: clock_enable while isolation active " )
                      , SDG_SVA_SOC_SIM) 

`HQM_SDG_ASSERTS_FORBIDDEN    ( assert_forbidden_hqm_inp_gated_clk_isolation_on_with_rcb_set
                      , (
                          ( ~`HQM_MASTER_PATH.pgcb_isol_en_b  & `HQM_MASTER_HQM_INP_GATED_CLK_ENABLE_RPTR_PATH.data_q)
                        )
                      , negedge `HQM_MASTER_PATH.hqm_fullrate_clk
                      , ~`HQM_MASTER_HQM_CLK_RPTR_RST_SYNC_N_PATH.rst_n_sync
                      , `HQM_SVA_ERR_MSG( "Error: hqm_pkg.sv  assert_forbidden_hqm_inp_gated_clk_isolation_on_with_lcb_or_lcb_set: clock_enable while isolation active " )
                      , SDG_SVA_SOC_SIM) 

////////////////////////////////////////////////////////////////////////////////////////////////////
// For any core non-FUNC_PF, non-FUNC_VF CSR access, verify this is actually a CSR bar access

`HQM_SDG_ASSERTS_FORBIDDEN(
                       assert_forbidden_non_csr_bar_csr_access
                      ,~( ((`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.iosfsb[0]) ?
                           (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.bar == 3'h2)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.fid == 8'h00)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:32]   == 32'h00000000)
                           ) :
                           (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:32] ==
                            `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.csr_pf_bar[63:32]
                           )
                          )
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[31:28] >= 4'h1)
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[31:28] <= 4'h9)
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_decode_val[0]
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr_mmio
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.mem_req_good
                        )
                      ,negedge `HQM_SYSTEM_PATH.hqm_gated_clk
                      ,~(      `HQM_SYSTEM_PATH.hqm_gated_rst_b_sys
                         &     `HQM_SYSTEM_PATH.hqm_inp_gated_rst_b
                         & |{  `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.unit_cfg_req_write
                            ,  `HQM_AQED_PIPE_PATH.i_hqm_aqed_pipe_core.unit_cfg_req_read
                            ,  `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.unit_cfg_req_write
                            ,  `HQM_ATM_PIPE_PATH.i_hqm_list_sel_pipe_core.i_hqm_lsp_atm_pipe.unit_cfg_req_read
                            ,  `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.unit_cfg_req_write
                            ,  `HQM_CREDIT_HIST_PIPE_PATH.i_hqm_credit_hist_pipe_core.unit_cfg_req_read
                            ,  `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.unit_cfg_req_write
                            ,  `HQM_DIR_PIPE_PATH.i_hqm_dir_pipe_core.unit_cfg_req_read
                            ,  `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.unit_cfg_req_write
                            ,  `HQM_LIST_SEL_PIPE_PATH.i_hqm_list_sel_pipe_core.unit_cfg_req_read
                            ,  `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.unit_cfg_req_write
                            ,  `HQM_NALB_PIPE_PATH.i_hqm_nalb_pipe_core.unit_cfg_req_read
                            ,  `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.unit_cfg_req_write
                            ,  `HQM_QED_PIPE_PATH.i_hqm_qed_pipe_core.unit_cfg_req_read
                            ,  `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.unit_cfg_req_write
                            ,  `HQM_REORDER_PIPE_PATH.i_hqm_reorder_pipe_core.unit_cfg_req_read
                            ,  `HQM_SYSTEM_PATH.i_hqm_system_core.hqm_system_csr_req.valid
                            }
                        )
                      ,`HQM_SVA_ERR_MSG("Error: hqm_core CSR accessed by non-CSR transaction")
                      ,SDG_SVA_SOC_SIM
)

`HQM_SDG_ASSERTS_FORBIDDEN(
                       assert_forbidden_non_csr_bar_csr_access_prim
                      ,~( ((`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.iosfsb[0]) ?
                           (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.bar == 3'h2)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.fid == 8'h00)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:32]   == 32'h00000000)
                           ) :
                           (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:32] ==
                            `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.csr_pf_bar[63:32]
                           )
                          )
                         & (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[31:28] == 4'h0)
                            | (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[31:28] == 4'ha)
                           )
                         & `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_decode_val[0]
                         & `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr_mmio
                         & `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.mem_req_good
                        )
                      ,negedge `HQM_SIF_PATH.i_hqm_sif_core.prim_nonflr_clk
                      ,~(      `HQM_SIF_PATH.i_hqm_sif_core.prim_gated_rst_b
                         & |{  `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.cfg_req_internal_write
                            ,  `HQM_MASTER_PATH.i_hqm_master_core.i_hqm_cfg_master.cfg_req_internal_read
                            ,  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_sif_csr_wrap.hqm_csr_int_mmio_req.valid
                            }
                        )
                      ,`HQM_SVA_ERR_MSG("Error: hqm_sif or hqm_master CSR accessed by non-CSR transaction")
                      ,SDG_SVA_SOC_SIM
)

////////////////////////////////////////////////////////////////////////////////////////////////////
// For any MSI-X table access, verify this is actually a valid FUNC_PF MMIO access to the MSI-X table

`HQM_SDG_ASSERTS_FORBIDDEN(
                       assert_forbidden_non_func_pf_msix_table_access
                      ,~( ((   `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.iosfsb[0]) ?
                           (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.bar == 3'h0)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.fid == 8'h00)
                            & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:26]   == 38'h0000000000)
                           ) :
                           (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:26] ==
                            `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.func_pf_bar[63:26]
                           )
                          )
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_decode_val[0]
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr_mmio
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.mem_req_good
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[25:11] == 15'h2000)
                         // Only 16B table entries 0-64 are valid
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[10: 4] <=  7'h40)
                        )
                      ,negedge `HQM_SYSTEM_PATH.hqm_gated_clk
                      ,~(      `HQM_SYSTEM_PATH.hqm_gated_rst_b_sys
                         &     `HQM_SYSTEM_PATH.hqm_inp_gated_rst_b
                         & (   `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_re_v.msg_addr_l
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_we_v.msg_addr_l
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_re_v.msg_addr_u
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_we_v.msg_addr_u
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_re_v.msg_data
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_we_v.msg_data
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_re_v.vector_ctrl
                            |  `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_alarm.cfg_we_v.vector_ctrl
                           )
                        )
                      ,`HQM_SVA_ERR_MSG("Error: MSI-X table accessed by non-FUNC_PF transaction")
                      ,SDG_SVA_SOC_SIM
)

////////////////////////////////////////////////////////////////////////////////////////////////////
// For any MSIX PBA access, verify this is actually a valid FUNC_PF MMIO access to the PBA 

`HQM_SDG_ASSERTS_FORBIDDEN(
                       assert_forbidden_non_func_pf_msix_pba_access
                      ,~(  ((   `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.iosfsb[0]) ?
                            (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.bar == 3'h0)
                             & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.sb_cds_msg.fid == 8'h00)
                             & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:26]   == 38'h0000000000)
                            ) :
                            (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:26] ==
                             `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.func_pf_bar[63:26]
                            )
                           )
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_decode_val[0]
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr_mmio
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.mem_req_good
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[25: 4] == 22'h100100)
                         // Only 3 PBA entries are valid
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[ 3: 2] <=  2'd2)
                        )
                      ,negedge `HQM_SYSTEM_PATH.hqm_gated_clk
                      ,~(      `HQM_SYSTEM_PATH.hqm_gated_rst_b_sys
                         &     `HQM_SYSTEM_PATH.hqm_inp_gated_rst_b
                         &     `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_msix_mem_wrap.i_hqm_msix_mem.req.valid
                         & (   `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_msix_mem_wrap.i_hqm_msix_mem.req.addr.mem.offset[47: 4] == 44'h0000_0100_100)
                         & (   `HQM_SYSTEM_PATH.i_hqm_system_core.i_hqm_system_msix_mem_wrap.i_hqm_msix_mem.req.addr.mem.offset[ 3: 2] >= 2'd2)
                        )
                      ,`HQM_SVA_ERR_MSG("Error: MSI-X PBA accessed by non-FUNC_PF transaction")
                      ,SDG_SVA_SOC_SIM
)

////////////////////////////////////////////////////////////////////////////////////////////////////
// For any PF HCW enqueue, verify this is actually a valid FUNC_PF MMIO HCW region access

`HQM_SDG_ASSERTS_FORBIDDEN(
                       assert_forbidden_non_func_pf_hcw_access
                      ,~(// No GPSB access
                         ~`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.iosfsb[0]
                         // Must be a write
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.posted
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_decode_val[0]
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr_mmio
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.mem_req_good
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[63:26] ==
                            `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.func_pf_bar[63:26]
                           )
                         &  `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[25]
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[24:22] == 3'd0)
                         // [21] is non-maskable
                         & ((`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[20]) ? // LDB/DIR PPs
                            (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[19:12] <  8'd64) :
                            (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[19:12] <  8'd128)
                           )
                         // Cannot access more than first 16 64B cache lines (1024B) within each PP's 4KB range
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[11:10] == 2'd0)
                         // [9:6] allows any of first 16 64B cache lines
                         // [5:0] is offset within 64B cache line.  Access must be modulo-16B aligned and within 64B cache line
                         & (  (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[5:2] == 4'hc)
                               & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length    == 10'd4)
                              )
                            | (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[5:2] == 4'h8)
                               & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length    <= 10'd8)
                              )
                            | (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[5:2] == 4'h4)
                               & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length    <= 10'd12)
                              )
                            | (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.addr[5:2] == 4'h0)
                               & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length    <= 10'd16)
                              )
                           )
                         // Length must be 4, 8, 12, or 16 DW
                         & (  (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length == 10'd4)
                            | (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length == 10'd8)
                            | (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length == 10'd12)
                            | (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.length == 10'd16)
                           )
                         // All byte enables must be on
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.endbe   == 4'hf)
                         & (`HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.cbd_hdr.startbe == 4'hf)
                        )
                      ,negedge `HQM_SIF_PATH.i_hqm_sif_core.prim_nonflr_clk
                      ,~(  `HQM_SIF_PATH.i_hqm_sif_core.prim_gated_rst_b
                         & `HQM_SIF_PATH.i_hqm_sif_core.i_hqm_ri.i_ri_cds.hcw_wr_wp
                        )
                      ,`HQM_SVA_ERR_MSG("Error: PF HCW enqueued by non-FUNC_PF transaction")
                      ,SDG_SVA_SOC_SIM
)

////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule

bind hqm_sip hqm_assert i_hqm_assert();

`endif
