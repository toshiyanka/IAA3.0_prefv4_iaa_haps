package rcfwl_picker_pkg;

import ovm_pkg::*;
import ConfigDB::*;
import systeminit::*;
import base_picker_pkg::*;

`include "rcfwl_picker.sv" 

// Reusable constraints
`include "default_rcfwl_constraints.sv"

endpackage: rcfwl_picker_pkg
