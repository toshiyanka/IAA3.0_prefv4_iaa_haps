
agent_compliance #
(.MAXPCMSTR(MAXPCMSTR),
 .MAXNPMSTR(MAXNPMSTR),
 .MAXPCTRGT(MAXPCTRGT),
 .MAXNPTRGT(MAXNPTRGT),
 .MAXTRGTADDR(MAXTRGTADDR),
 .MAXTRGTDATA(MAXTRGTDATA),
 .MAXMSTRADDR(MAXMSTRADDR),
 .MAXMSTRDATA(MAXMSTRDATA),
 .NUM_TX_EXT_HEADERS(NUM_TX_EXT_HEADERS),
 .NUM_RX_EXT_HEADERS(NUM_RX_EXT_HEADERS),
 .TX_EXT_HEADER_SUPPORT(TX_EXT_HEADER_SUPPORT),
 .RX_EXT_HEADER_SUPPORT(RX_EXT_HEADER_SUPPORT))
