/*
================================================================================
  Copyright (c) 2011 Intel Corporation, all rights reserved.

  THIS PROGRAM IS AN UNPUBLISHED WORK FULLY PROTECTED BY COPYRIGHT LAWS AND IS 
  CONSIDERED A TRADE SECRET BELONGING TO THE INTEL CORPORATION.
================================================================================

  Author          : 
  Email           : 
  Phone           : 
  Date            : 

================================================================================
  Description     : One line description of this class
  
Write your wordy description here.
================================================================================
*/

//Minimum Subset an Agent should contain
`include "CCAgentTypes.svh"
`include "CCAgentDriver.svh"
//col change
`include "CCAgentDriver_Col.svh"
//END col change
`include "CCAgentSeqItem.svh"
`include "CCAgentSequencer.svh"
`include "CCAgentResponder.svh"
`include "CCAgentSIPResponder.svh"
`include "CCAgentSeqLib.svh"
`include "CCAgent.svh"
`include "CCAgentResponseSeqItem.svh"
`include "CCAgentArbiter.svh"
`include "CCAgentSIPFSM.svh"
`include "CCAgentFabricFSM.svh"
//col change
`include "CCAgentSIPFSM_Col.svh"
`include "CCAgentFabricFSM_Col.svh"
//END col change


