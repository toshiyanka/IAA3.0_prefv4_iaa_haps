`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

(* inserted_by="VISA IT" *) logic [29:0] visaPrbsFrom_hqm_master_visa_block;



`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
