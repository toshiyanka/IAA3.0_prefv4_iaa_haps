VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf054b256e1r1w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf054b256e1r1w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 43.2 BY 25.92 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 13.8 19.028 15 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 11.88 22.072 13.08 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 13.8 19.928 15 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 13.8 20.016 15 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 13.8 20.272 15 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 13.8 20.528 15 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 13.8 20.616 15 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 13.8 20.828 15 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 13.8 20.916 15 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 13.8 21.172 15 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 13.8 19.116 15 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 13.8 19.372 15 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 13.8 19.628 15 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 13.8 19.716 15 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.184 11.88 23.228 13.08 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.272 11.88 23.316 13.08 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.484 11.88 23.528 13.08 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.572 11.88 23.616 13.08 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 23.828 11.88 23.872 13.08 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 11.88 18.472 13.08 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.88 18.728 13.08 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 11.88 18.816 13.08 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 11.88 22.328 13.08 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 11.88 22.416 13.08 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 0.24 18.472 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 3.84 22.716 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 3.84 22.972 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 4.56 19.116 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 4.56 19.372 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 5.28 20.272 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 5.28 20.528 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 6 20.916 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 6 21.172 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 6.72 21.728 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 6.72 21.816 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 0.24 18.728 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 7.44 22.416 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 7.44 22.628 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 8.16 18.472 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 8.16 18.728 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 8.88 19.928 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 8.88 20.016 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 9.6 20.616 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 9.6 20.828 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 10.32 21.428 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 10.32 21.516 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 0.96 19.928 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 15.84 18.472 17.04 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 15.84 18.728 17.04 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 16.56 19.716 17.76 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 16.56 19.928 17.76 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 17.28 20.616 18.48 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 17.28 20.828 18.48 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 18 21.428 19.2 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 18 21.516 19.2 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 18.72 22.072 19.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 18.72 22.328 19.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 0.96 20.016 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 19.44 22.716 20.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 19.44 22.972 20.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 20.16 19.116 21.36 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.328 20.16 19.372 21.36 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 20.88 20.272 22.08 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 20.88 20.528 22.08 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 21.6 20.916 22.8 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 21.6 21.172 22.8 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 22.32 21.728 23.52 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 22.32 21.816 23.52 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.68 20.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 23.04 22.416 24.24 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 23.04 22.628 24.24 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 23.76 18.472 24.96 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 23.76 18.728 24.96 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.884 24.48 19.928 25.68 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 24.48 20.016 25.68 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 1.68 20.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 2.4 21.428 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 2.4 21.516 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 3.12 22.072 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 3.12 22.328 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 11.88 22.716 13.08 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 11.88 22.972 13.08 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 11.88 22.628 13.08 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 3.84 18.472 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 3.84 18.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 4.56 19.628 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 4.56 19.716 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 5.28 20.616 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 5.28 20.828 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 6 21.428 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 6 21.516 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 6.72 22.072 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 6.72 22.328 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 7.44 22.716 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 7.44 22.972 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.16 18.816 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.16 19.028 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 8.88 20.272 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 8.88 20.528 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 9.6 20.916 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 9.6 21.172 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 10.32 21.728 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 10.32 21.816 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 0.96 20.272 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 15.84 18.816 17.04 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 15.84 21.428 17.04 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 16.56 20.016 17.76 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 16.56 20.272 17.76 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 17.28 20.916 18.48 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 17.28 21.172 18.48 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 18 21.728 19.2 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 18 21.816 19.2 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 18.72 22.416 19.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 18.72 22.628 19.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 0.96 20.528 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 19.44 18.472 20.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 19.44 18.728 20.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 20.16 19.628 21.36 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 20.16 19.716 21.36 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 20.88 20.616 22.08 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 20.88 20.828 22.08 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 21.6 21.428 22.8 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 21.6 21.516 22.8 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.028 22.32 22.072 23.52 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.284 22.32 22.328 23.52 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 1.68 20.916 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.672 23.04 22.716 24.24 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.928 23.04 22.972 24.24 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 23.76 18.816 24.96 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 23.76 19.028 24.96 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 24.48 20.272 25.68 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 24.48 20.528 25.68 ;
    END
  END rddatap0[55]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 1.68 21.172 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 2.4 21.728 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.4 21.816 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.372 3.12 22.416 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 22.584 3.12 22.628 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 25.86 ;
        RECT 2.662 0.06 2.738 25.86 ;
        RECT 4.462 0.06 4.538 25.86 ;
        RECT 6.262 0.06 6.338 25.86 ;
        RECT 8.062 0.06 8.138 25.86 ;
        RECT 9.862 0.06 9.938 25.86 ;
        RECT 11.662 0.06 11.738 25.86 ;
        RECT 13.462 0.06 13.538 25.86 ;
        RECT 15.262 0.06 15.338 25.86 ;
        RECT 17.062 0.06 17.138 25.86 ;
        RECT 18.862 0.06 18.938 25.86 ;
        RECT 20.662 0.06 20.738 25.86 ;
        RECT 22.462 0.06 22.538 25.86 ;
        RECT 24.262 0.06 24.338 25.86 ;
        RECT 26.062 0.06 26.138 25.86 ;
        RECT 27.862 0.06 27.938 25.86 ;
        RECT 29.662 0.06 29.738 25.86 ;
        RECT 31.462 0.06 31.538 25.86 ;
        RECT 33.262 0.06 33.338 25.86 ;
        RECT 35.062 0.06 35.138 25.86 ;
        RECT 36.862 0.06 36.938 25.86 ;
        RECT 38.662 0.06 38.738 25.86 ;
        RECT 40.462 0.06 40.538 25.86 ;
        RECT 42.262 0.06 42.338 25.86 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 25.86 ;
        RECT 3.562 0.06 3.638 25.86 ;
        RECT 5.362 0.06 5.438 25.86 ;
        RECT 7.162 0.06 7.238 25.86 ;
        RECT 8.962 0.06 9.038 25.86 ;
        RECT 10.762 0.06 10.838 25.86 ;
        RECT 12.562 0.06 12.638 25.86 ;
        RECT 14.362 0.06 14.438 25.86 ;
        RECT 16.162 0.06 16.238 25.86 ;
        RECT 17.962 0.06 18.038 25.86 ;
        RECT 19.762 0.06 19.838 25.86 ;
        RECT 21.562 0.06 21.638 25.86 ;
        RECT 23.362 0.06 23.438 25.86 ;
        RECT 25.162 0.06 25.238 25.86 ;
        RECT 26.962 0.06 27.038 25.86 ;
        RECT 28.762 0.06 28.838 25.86 ;
        RECT 30.562 0.06 30.638 25.86 ;
        RECT 32.362 0.06 32.438 25.86 ;
        RECT 34.162 0.06 34.238 25.86 ;
        RECT 35.962 0.06 36.038 25.86 ;
        RECT 37.762 0.06 37.838 25.86 ;
        RECT 39.562 0.06 39.638 25.86 ;
        RECT 41.362 0.06 41.438 25.86 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 43.216 25.934 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 43.22 25.94 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 43.2705 25.958 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 43.235 25.99 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 43.27 25.958 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 43.259 26.01 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 43.29 25.982 ;
    LAYER m7 SPACING 0 ;
      RECT 42.338 25.98 43.24 26.04 ;
      RECT 42.338 -0.06 43.292 25.98 ;
      RECT 42.338 -0.12 43.24 -0.06 ;
      RECT 41.438 -0.12 42.262 26.04 ;
      RECT 40.538 -0.12 41.362 26.04 ;
      RECT 39.638 -0.12 40.462 26.04 ;
      RECT 38.738 -0.12 39.562 26.04 ;
      RECT 37.838 -0.12 38.662 26.04 ;
      RECT 36.938 -0.12 37.762 26.04 ;
      RECT 36.038 -0.12 36.862 26.04 ;
      RECT 35.138 -0.12 35.962 26.04 ;
      RECT 34.238 -0.12 35.062 26.04 ;
      RECT 33.338 -0.12 34.162 26.04 ;
      RECT 32.438 -0.12 33.262 26.04 ;
      RECT 31.538 -0.12 32.362 26.04 ;
      RECT 30.638 -0.12 31.462 26.04 ;
      RECT 29.738 -0.12 30.562 26.04 ;
      RECT 28.838 -0.12 29.662 26.04 ;
      RECT 27.938 -0.12 28.762 26.04 ;
      RECT 27.038 -0.12 27.862 26.04 ;
      RECT 26.138 -0.12 26.962 26.04 ;
      RECT 25.238 -0.12 26.062 26.04 ;
      RECT 24.338 -0.12 25.162 26.04 ;
      RECT 23.438 13.08 24.262 26.04 ;
      RECT 23.438 11.88 23.484 13.08 ;
      RECT 23.528 11.88 23.572 13.08 ;
      RECT 23.616 11.88 23.828 13.08 ;
      RECT 23.872 11.88 24.262 13.08 ;
      RECT 23.438 -0.12 24.262 11.88 ;
      RECT 22.538 24.24 23.362 26.04 ;
      RECT 22.538 23.04 22.584 24.24 ;
      RECT 22.628 23.04 22.672 24.24 ;
      RECT 22.716 23.04 22.928 24.24 ;
      RECT 22.972 23.04 23.362 24.24 ;
      RECT 22.538 20.64 23.362 23.04 ;
      RECT 22.538 19.92 22.672 20.64 ;
      RECT 22.716 19.44 22.928 20.64 ;
      RECT 22.972 19.44 23.362 20.64 ;
      RECT 22.628 19.44 22.672 19.92 ;
      RECT 22.538 18.72 22.584 19.92 ;
      RECT 22.628 18.72 23.362 19.44 ;
      RECT 22.538 13.08 23.362 18.72 ;
      RECT 22.538 11.88 22.584 13.08 ;
      RECT 22.628 11.88 22.672 13.08 ;
      RECT 22.716 11.88 22.928 13.08 ;
      RECT 22.972 11.88 23.184 13.08 ;
      RECT 23.228 11.88 23.272 13.08 ;
      RECT 23.316 11.88 23.362 13.08 ;
      RECT 22.538 8.64 23.362 11.88 ;
      RECT 22.538 7.44 22.584 8.64 ;
      RECT 22.628 7.44 22.672 8.64 ;
      RECT 22.716 7.44 22.928 8.64 ;
      RECT 22.972 7.44 23.362 8.64 ;
      RECT 22.538 5.04 23.362 7.44 ;
      RECT 22.538 4.32 22.672 5.04 ;
      RECT 22.716 3.84 22.928 5.04 ;
      RECT 22.972 3.84 23.362 5.04 ;
      RECT 22.628 3.84 22.672 4.32 ;
      RECT 22.538 3.12 22.584 4.32 ;
      RECT 22.628 3.12 23.362 3.84 ;
      RECT 22.538 -0.12 23.362 3.12 ;
      RECT 21.638 24.24 22.462 26.04 ;
      RECT 21.638 23.52 22.372 24.24 ;
      RECT 22.416 23.04 22.462 24.24 ;
      RECT 22.328 23.04 22.372 23.52 ;
      RECT 21.638 22.32 21.684 23.52 ;
      RECT 21.728 22.32 21.772 23.52 ;
      RECT 21.816 22.32 22.028 23.52 ;
      RECT 22.072 22.32 22.284 23.52 ;
      RECT 22.328 22.32 22.462 23.04 ;
      RECT 21.638 19.92 22.462 22.32 ;
      RECT 21.638 19.2 22.028 19.92 ;
      RECT 22.072 18.72 22.284 19.92 ;
      RECT 22.328 18.72 22.372 19.92 ;
      RECT 22.416 18.72 22.462 19.92 ;
      RECT 21.816 18.72 22.028 19.2 ;
      RECT 21.638 18 21.684 19.2 ;
      RECT 21.728 18 21.772 19.2 ;
      RECT 21.816 18 22.462 18.72 ;
      RECT 21.638 13.08 22.462 18 ;
      RECT 21.638 11.88 22.028 13.08 ;
      RECT 22.072 11.88 22.284 13.08 ;
      RECT 22.328 11.88 22.372 13.08 ;
      RECT 22.416 11.88 22.462 13.08 ;
      RECT 21.638 11.52 22.462 11.88 ;
      RECT 21.638 10.32 21.684 11.52 ;
      RECT 21.728 10.32 21.772 11.52 ;
      RECT 21.816 10.32 22.462 11.52 ;
      RECT 21.638 8.64 22.462 10.32 ;
      RECT 21.638 7.92 22.372 8.64 ;
      RECT 22.416 7.44 22.462 8.64 ;
      RECT 22.328 7.44 22.372 7.92 ;
      RECT 21.638 6.72 21.684 7.92 ;
      RECT 21.728 6.72 21.772 7.92 ;
      RECT 21.816 6.72 22.028 7.92 ;
      RECT 22.072 6.72 22.284 7.92 ;
      RECT 22.328 6.72 22.462 7.44 ;
      RECT 21.638 4.32 22.462 6.72 ;
      RECT 21.638 3.6 22.028 4.32 ;
      RECT 22.072 3.12 22.284 4.32 ;
      RECT 22.328 3.12 22.372 4.32 ;
      RECT 22.416 3.12 22.462 4.32 ;
      RECT 21.816 3.12 22.028 3.6 ;
      RECT 21.638 2.4 21.684 3.6 ;
      RECT 21.728 2.4 21.772 3.6 ;
      RECT 21.816 2.4 22.462 3.12 ;
      RECT 21.638 -0.12 22.462 2.4 ;
      RECT 20.738 22.8 21.562 26.04 ;
      RECT 20.738 22.08 20.872 22.8 ;
      RECT 20.916 21.6 21.128 22.8 ;
      RECT 21.172 21.6 21.384 22.8 ;
      RECT 21.428 21.6 21.472 22.8 ;
      RECT 21.516 21.6 21.562 22.8 ;
      RECT 20.828 21.6 20.872 22.08 ;
      RECT 20.738 20.88 20.784 22.08 ;
      RECT 20.828 20.88 21.562 21.6 ;
      RECT 20.738 19.2 21.562 20.88 ;
      RECT 20.738 18.48 21.384 19.2 ;
      RECT 21.428 18 21.472 19.2 ;
      RECT 21.516 18 21.562 19.2 ;
      RECT 21.172 18 21.384 18.48 ;
      RECT 20.738 17.28 20.784 18.48 ;
      RECT 20.828 17.28 20.872 18.48 ;
      RECT 20.916 17.28 21.128 18.48 ;
      RECT 21.172 17.28 21.562 18 ;
      RECT 20.738 17.04 21.562 17.28 ;
      RECT 20.738 15.84 21.384 17.04 ;
      RECT 21.428 15.84 21.562 17.04 ;
      RECT 20.738 15 21.562 15.84 ;
      RECT 20.738 13.8 20.784 15 ;
      RECT 20.828 13.8 20.872 15 ;
      RECT 20.916 13.8 21.128 15 ;
      RECT 21.172 13.8 21.562 15 ;
      RECT 20.738 11.52 21.562 13.8 ;
      RECT 20.738 10.8 21.384 11.52 ;
      RECT 21.428 10.32 21.472 11.52 ;
      RECT 21.516 10.32 21.562 11.52 ;
      RECT 21.172 10.32 21.384 10.8 ;
      RECT 20.738 9.6 20.784 10.8 ;
      RECT 20.828 9.6 20.872 10.8 ;
      RECT 20.916 9.6 21.128 10.8 ;
      RECT 21.172 9.6 21.562 10.32 ;
      RECT 20.738 7.2 21.562 9.6 ;
      RECT 20.738 6.48 20.872 7.2 ;
      RECT 20.916 6 21.128 7.2 ;
      RECT 21.172 6 21.384 7.2 ;
      RECT 21.428 6 21.472 7.2 ;
      RECT 21.516 6 21.562 7.2 ;
      RECT 20.828 6 20.872 6.48 ;
      RECT 20.738 5.28 20.784 6.48 ;
      RECT 20.828 5.28 21.562 6 ;
      RECT 20.738 3.6 21.562 5.28 ;
      RECT 20.738 2.88 21.384 3.6 ;
      RECT 21.428 2.4 21.472 3.6 ;
      RECT 21.516 2.4 21.562 3.6 ;
      RECT 21.172 2.4 21.384 2.88 ;
      RECT 20.738 1.68 20.784 2.88 ;
      RECT 20.828 1.68 20.872 2.88 ;
      RECT 20.916 1.68 21.128 2.88 ;
      RECT 21.172 1.68 21.562 2.4 ;
      RECT 20.738 -0.12 21.562 1.68 ;
      RECT 19.838 25.68 20.662 26.04 ;
      RECT 19.838 24.48 19.884 25.68 ;
      RECT 19.928 24.48 19.972 25.68 ;
      RECT 20.016 24.48 20.228 25.68 ;
      RECT 20.272 24.48 20.484 25.68 ;
      RECT 20.528 24.48 20.662 25.68 ;
      RECT 19.838 22.08 20.662 24.48 ;
      RECT 19.838 20.88 20.228 22.08 ;
      RECT 20.272 20.88 20.484 22.08 ;
      RECT 20.528 20.88 20.572 22.08 ;
      RECT 20.616 20.88 20.662 22.08 ;
      RECT 19.838 18.48 20.662 20.88 ;
      RECT 19.838 17.76 20.572 18.48 ;
      RECT 20.616 17.28 20.662 18.48 ;
      RECT 20.272 17.28 20.572 17.76 ;
      RECT 19.838 16.56 19.884 17.76 ;
      RECT 19.928 16.56 19.972 17.76 ;
      RECT 20.016 16.56 20.228 17.76 ;
      RECT 20.272 16.56 20.662 17.28 ;
      RECT 19.838 15 20.662 16.56 ;
      RECT 19.838 13.8 19.884 15 ;
      RECT 19.928 13.8 19.972 15 ;
      RECT 20.016 13.8 20.228 15 ;
      RECT 20.272 13.8 20.484 15 ;
      RECT 20.528 13.8 20.572 15 ;
      RECT 20.616 13.8 20.662 15 ;
      RECT 19.838 10.8 20.662 13.8 ;
      RECT 19.838 10.08 20.572 10.8 ;
      RECT 20.616 9.6 20.662 10.8 ;
      RECT 20.528 9.6 20.572 10.08 ;
      RECT 19.838 8.88 19.884 10.08 ;
      RECT 19.928 8.88 19.972 10.08 ;
      RECT 20.016 8.88 20.228 10.08 ;
      RECT 20.272 8.88 20.484 10.08 ;
      RECT 20.528 8.88 20.662 9.6 ;
      RECT 19.838 6.48 20.662 8.88 ;
      RECT 19.838 5.28 20.228 6.48 ;
      RECT 20.272 5.28 20.484 6.48 ;
      RECT 20.528 5.28 20.572 6.48 ;
      RECT 20.616 5.28 20.662 6.48 ;
      RECT 19.838 2.88 20.662 5.28 ;
      RECT 19.838 2.16 20.572 2.88 ;
      RECT 20.616 1.68 20.662 2.88 ;
      RECT 20.528 1.68 20.572 2.16 ;
      RECT 19.838 0.96 19.884 2.16 ;
      RECT 19.928 0.96 19.972 2.16 ;
      RECT 20.016 0.96 20.228 2.16 ;
      RECT 20.272 0.96 20.484 2.16 ;
      RECT 20.528 0.96 20.662 1.68 ;
      RECT 19.838 -0.12 20.662 0.96 ;
      RECT 18.938 24.96 19.762 26.04 ;
      RECT 18.938 23.76 18.984 24.96 ;
      RECT 19.028 23.76 19.762 24.96 ;
      RECT 18.938 21.36 19.762 23.76 ;
      RECT 18.938 20.16 19.072 21.36 ;
      RECT 19.116 20.16 19.328 21.36 ;
      RECT 19.372 20.16 19.584 21.36 ;
      RECT 19.628 20.16 19.672 21.36 ;
      RECT 19.716 20.16 19.762 21.36 ;
      RECT 18.938 17.76 19.762 20.16 ;
      RECT 18.938 16.56 19.672 17.76 ;
      RECT 19.716 16.56 19.762 17.76 ;
      RECT 18.938 15 19.762 16.56 ;
      RECT 18.938 13.8 18.984 15 ;
      RECT 19.028 13.8 19.072 15 ;
      RECT 19.116 13.8 19.328 15 ;
      RECT 19.372 13.8 19.584 15 ;
      RECT 19.628 13.8 19.672 15 ;
      RECT 19.716 13.8 19.762 15 ;
      RECT 18.938 9.36 19.762 13.8 ;
      RECT 18.938 8.16 18.984 9.36 ;
      RECT 19.028 8.16 19.762 9.36 ;
      RECT 18.938 5.76 19.762 8.16 ;
      RECT 18.938 4.56 19.072 5.76 ;
      RECT 19.116 4.56 19.328 5.76 ;
      RECT 19.372 4.56 19.584 5.76 ;
      RECT 19.628 4.56 19.672 5.76 ;
      RECT 19.716 4.56 19.762 5.76 ;
      RECT 18.938 1.44 19.762 4.56 ;
      RECT 18.938 0.24 18.984 1.44 ;
      RECT 19.028 0.24 19.762 1.44 ;
      RECT 18.938 -0.12 19.762 0.24 ;
      RECT 18.038 24.96 18.862 26.04 ;
      RECT 18.038 23.76 18.428 24.96 ;
      RECT 18.472 23.76 18.684 24.96 ;
      RECT 18.728 23.76 18.772 24.96 ;
      RECT 18.816 23.76 18.862 24.96 ;
      RECT 18.038 20.64 18.862 23.76 ;
      RECT 18.038 19.44 18.428 20.64 ;
      RECT 18.472 19.44 18.684 20.64 ;
      RECT 18.728 19.44 18.862 20.64 ;
      RECT 18.038 17.04 18.862 19.44 ;
      RECT 18.038 15.84 18.428 17.04 ;
      RECT 18.472 15.84 18.684 17.04 ;
      RECT 18.728 15.84 18.772 17.04 ;
      RECT 18.816 15.84 18.862 17.04 ;
      RECT 18.038 13.08 18.862 15.84 ;
      RECT 18.038 11.88 18.428 13.08 ;
      RECT 18.472 11.88 18.684 13.08 ;
      RECT 18.728 11.88 18.772 13.08 ;
      RECT 18.816 11.88 18.862 13.08 ;
      RECT 18.038 9.36 18.862 11.88 ;
      RECT 18.038 8.16 18.428 9.36 ;
      RECT 18.472 8.16 18.684 9.36 ;
      RECT 18.728 8.16 18.772 9.36 ;
      RECT 18.816 8.16 18.862 9.36 ;
      RECT 18.038 5.04 18.862 8.16 ;
      RECT 18.038 3.84 18.428 5.04 ;
      RECT 18.472 3.84 18.684 5.04 ;
      RECT 18.728 3.84 18.862 5.04 ;
      RECT 18.038 1.44 18.862 3.84 ;
      RECT 18.038 0.24 18.428 1.44 ;
      RECT 18.472 0.24 18.684 1.44 ;
      RECT 18.728 0.24 18.772 1.44 ;
      RECT 18.816 0.24 18.862 1.44 ;
      RECT 18.038 -0.12 18.862 0.24 ;
      RECT 17.138 -0.12 17.962 26.04 ;
      RECT 16.238 -0.12 17.062 26.04 ;
      RECT 15.338 -0.12 16.162 26.04 ;
      RECT 14.438 -0.12 15.262 26.04 ;
      RECT 13.538 -0.12 14.362 26.04 ;
      RECT 12.638 -0.12 13.462 26.04 ;
      RECT 11.738 -0.12 12.562 26.04 ;
      RECT 10.838 -0.12 11.662 26.04 ;
      RECT 9.938 -0.12 10.762 26.04 ;
      RECT 9.038 -0.12 9.862 26.04 ;
      RECT 8.138 -0.12 8.962 26.04 ;
      RECT 7.238 -0.12 8.062 26.04 ;
      RECT 6.338 -0.12 7.162 26.04 ;
      RECT 5.438 -0.12 6.262 26.04 ;
      RECT 4.538 -0.12 5.362 26.04 ;
      RECT 3.638 -0.12 4.462 26.04 ;
      RECT 2.738 -0.12 3.562 26.04 ;
      RECT 1.838 -0.12 2.662 26.04 ;
      RECT 0.938 -0.12 1.762 26.04 ;
      RECT -0.04 25.98 0.862 26.04 ;
      RECT -0.092 -0.06 0.862 25.98 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 42.458 0 43.12 25.92 ;
      RECT 41.558 0 42.142 25.92 ;
      RECT 40.658 0 41.242 25.92 ;
      RECT 39.758 0 40.342 25.92 ;
      RECT 38.858 0 39.442 25.92 ;
      RECT 37.958 0 38.542 25.92 ;
      RECT 37.058 0 37.642 25.92 ;
      RECT 36.158 0 36.742 25.92 ;
      RECT 35.258 0 35.842 25.92 ;
      RECT 34.358 0 34.942 25.92 ;
      RECT 33.458 0 34.042 25.92 ;
      RECT 32.558 0 33.142 25.92 ;
      RECT 31.658 0 32.242 25.92 ;
      RECT 30.758 0 31.342 25.92 ;
      RECT 29.858 0 30.442 25.92 ;
      RECT 28.958 0 29.542 25.92 ;
      RECT 28.058 0 28.642 25.92 ;
      RECT 27.158 0 27.742 25.92 ;
      RECT 26.258 0 26.842 25.92 ;
      RECT 25.358 0 25.942 25.92 ;
      RECT 24.458 0 25.042 25.92 ;
      RECT 23.558 13.2 24.142 25.92 ;
      RECT 23.992 11.76 24.142 13.2 ;
      RECT 23.558 0 24.142 11.76 ;
      RECT 22.658 24.36 23.242 25.92 ;
      RECT 23.092 22.92 23.242 24.36 ;
      RECT 22.658 20.76 23.242 22.92 ;
      RECT 23.092 19.32 23.242 20.76 ;
      RECT 22.748 18.6 23.242 19.32 ;
      RECT 22.658 13.2 23.242 18.6 ;
      RECT 21.758 24.36 22.342 25.92 ;
      RECT 21.758 23.64 22.252 24.36 ;
      RECT 20.858 22.92 21.442 25.92 ;
      RECT 19.958 25.8 20.542 25.92 ;
      RECT 19.058 25.08 19.642 25.92 ;
      RECT 19.148 23.64 19.642 25.08 ;
      RECT 19.058 21.48 19.642 23.64 ;
      RECT 18.158 25.08 18.742 25.92 ;
      RECT 18.158 23.64 18.308 25.08 ;
      RECT 18.158 20.76 18.742 23.64 ;
      RECT 18.158 19.32 18.308 20.76 ;
      RECT 18.158 17.16 18.742 19.32 ;
      RECT 18.158 15.72 18.308 17.16 ;
      RECT 18.158 13.2 18.742 15.72 ;
      RECT 18.158 11.76 18.308 13.2 ;
      RECT 18.158 9.48 18.742 11.76 ;
      RECT 18.158 8.04 18.308 9.48 ;
      RECT 18.158 5.16 18.742 8.04 ;
      RECT 18.158 3.72 18.308 5.16 ;
      RECT 18.158 1.56 18.742 3.72 ;
      RECT 18.158 0.12 18.308 1.56 ;
      RECT 18.158 0 18.742 0.12 ;
      RECT 17.258 0 17.842 25.92 ;
      RECT 16.358 0 16.942 25.92 ;
      RECT 15.458 0 16.042 25.92 ;
      RECT 14.558 0 15.142 25.92 ;
      RECT 13.658 0 14.242 25.92 ;
      RECT 12.758 0 13.342 25.92 ;
      RECT 11.858 0 12.442 25.92 ;
      RECT 10.958 0 11.542 25.92 ;
      RECT 10.058 0 10.642 25.92 ;
      RECT 9.158 0 9.742 25.92 ;
      RECT 8.258 0 8.842 25.92 ;
      RECT 7.358 0 7.942 25.92 ;
      RECT 6.458 0 7.042 25.92 ;
      RECT 5.558 0 6.142 25.92 ;
      RECT 4.658 0 5.242 25.92 ;
      RECT 3.758 0 4.342 25.92 ;
      RECT 2.858 0 3.442 25.92 ;
      RECT 1.958 0 2.542 25.92 ;
      RECT 1.058 0 1.642 25.92 ;
      RECT 0.08 0 0.742 25.92 ;
      RECT 19.958 22.2 20.542 24.36 ;
      RECT 19.958 20.76 20.108 22.2 ;
      RECT 19.958 18.6 20.542 20.76 ;
      RECT 19.958 17.88 20.452 18.6 ;
      RECT 20.392 17.16 20.452 17.88 ;
      RECT 20.392 16.44 20.542 17.16 ;
      RECT 19.958 15.12 20.542 16.44 ;
      RECT 21.758 20.04 22.342 22.2 ;
      RECT 21.758 19.32 21.908 20.04 ;
      RECT 20.948 20.76 21.442 21.48 ;
      RECT 20.858 19.32 21.442 20.76 ;
      RECT 20.858 18.6 21.264 19.32 ;
      RECT 19.058 17.88 19.642 20.04 ;
      RECT 19.058 16.44 19.552 17.88 ;
      RECT 19.058 15.12 19.642 16.44 ;
      RECT 21.936 17.88 22.342 18.6 ;
      RECT 21.758 13.2 22.342 17.88 ;
      RECT 21.758 11.76 21.908 13.2 ;
      RECT 21.758 11.64 22.342 11.76 ;
      RECT 21.936 10.2 22.342 11.64 ;
      RECT 21.758 8.76 22.342 10.2 ;
      RECT 21.758 8.04 22.252 8.76 ;
      RECT 21.292 17.16 21.442 17.88 ;
      RECT 20.858 15.72 21.264 17.16 ;
      RECT 20.858 15.12 21.442 15.72 ;
      RECT 21.292 13.68 21.442 15.12 ;
      RECT 20.858 11.64 21.442 13.68 ;
      RECT 20.858 10.92 21.264 11.64 ;
      RECT 19.958 10.92 20.542 13.68 ;
      RECT 19.958 10.2 20.452 10.92 ;
      RECT 19.058 9.48 19.642 13.68 ;
      RECT 19.148 8.04 19.642 9.48 ;
      RECT 19.058 5.88 19.642 8.04 ;
      RECT 22.658 8.76 23.242 11.76 ;
      RECT 23.092 7.32 23.242 8.76 ;
      RECT 22.658 5.16 23.242 7.32 ;
      RECT 23.092 3.72 23.242 5.16 ;
      RECT 22.748 3 23.242 3.72 ;
      RECT 22.658 0 23.242 3 ;
      RECT 21.292 9.48 21.442 10.2 ;
      RECT 20.858 7.32 21.442 9.48 ;
      RECT 19.958 6.6 20.542 8.76 ;
      RECT 19.958 5.16 20.108 6.6 ;
      RECT 19.958 3 20.542 5.16 ;
      RECT 19.958 2.28 20.452 3 ;
      RECT 21.758 4.44 22.342 6.6 ;
      RECT 21.758 3.72 21.908 4.44 ;
      RECT 20.948 5.16 21.442 5.88 ;
      RECT 20.858 3.72 21.442 5.16 ;
      RECT 20.858 3 21.264 3.72 ;
      RECT 19.058 1.56 19.642 4.44 ;
      RECT 19.148 0.12 19.642 1.56 ;
      RECT 19.058 0 19.642 0.12 ;
      RECT 21.936 2.28 22.342 3 ;
      RECT 21.758 0 22.342 2.28 ;
      RECT 21.292 1.56 21.442 2.28 ;
      RECT 20.858 0 21.442 1.56 ;
      RECT 19.958 0 20.542 0.84 ;
    LAYER m0 ;
      RECT 0 0.002 43.2 25.918 ;
    LAYER m1 ;
      RECT 0 0 43.2 25.92 ;
    LAYER m2 ;
      RECT 0 0.015 43.2 25.905 ;
    LAYER m3 ;
      RECT 0.015 0 43.185 25.92 ;
    LAYER m4 ;
      RECT 0 0.02 43.2 25.9 ;
    LAYER m5 ;
      RECT 0.012 0 43.188 25.92 ;
    LAYER m6 ;
      RECT 0 0.012 43.2 25.908 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf054b256e1r1w0cbbeheaa4acw

END LIBRARY
