//Place any new sequences in the SeqLib directory & `include them here. This file `included in your main include file.
`include "SeqLib/PGCBAgentBaseSequence.svh"
`include "SeqLib/PGCBAgentDefaultSequence.svh"
//`include "SeqLib/PGCBAgentBaseResponseVSeq.svh"
