//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// hqm_list_sel_pipe
//
// The list select pipe consists of 5 essentially independent pipelines:
// - LBARB      : Load-balanced arbitration/scheduling, including CQ selection, for Unordered, Ordered
//                and ATM requests.  ATM scheduling splits off earlier in the pipe for performance,
//                and works off sched/ready list status provided by AP rather than seeing enqueues directly.
// - ATQ        : ATQ -> ATM requests
// - DIRENQ     : Directed scheduling based on Directed enqueue requests
// - LBRPL      : Load-balanced reorder -> replay requests
// - DIRRPL     : Directed reorder -> replay requests
//
// 
// The overall flow is:
//                                       +----------+
//                               +-+     |          |
// chp_lsp_cmp         --------->|A|---->|          |
// rop_lsp_reordercmp  --------->|R|     |          |
//                               |B|     |          |-------------------------------> lsp_nalb_sch_unoord
//                               +-+     |  LBARB   |
// chp_lsp_token       --+-------------->|          |
//                       |               |          |
// +----+                |       +-+     |          |
// |    |  rlst_*      --|------>|A|---->|          |
// | AP |  slst_*      --|------>|R|     +--+-------+                      +----+
// +----+                |       |B|        |                              |    |
// nalb_lsp_enq_lb     --|---+-->| |        +-------------- lsp_ap_atm --> | AP |
//                       |   |   +-+                                       +----+
//                       |   |           +----------+
//                       |   +---------->| ATQ      |-------------------------------> lsp_nalb_sch_atq
// aqed_lsp_sch        --|-------------->|          |
//                       |               +----------+
//                       |        
//                       |               +----------+
// nalb_lsp_enq_rorply --|-------------->| LBRPL    |-------------------------------> lsp_nalb_sch_rorply
//                       |               +----------+
//                       |
//                       |               +----------+
//                       +-------------->| DIRENQ   |-------------------------------> lsp_dp_sch_dir
// dp_lsp_enq_dir      ----------------->|          |
//                                       +----------+
//                                
//                                       +----------+
// dp_lsp_enq_rorply   ----------------->| DIRRPL   |-------------------------------> lsp_dp_sch_rorply
//                                       +----------+
//
// rtl organization is:
//   LBARB
//   ATQ
//   DIRENQ
//   LBRPL
//   DIRRPL
//-----------------------------------------------------------------------------------------------------

module hqm_list_sel_pipe_core
import hqm_AW_pkg::*, hqm_pkg::*, hqm_core_pkg::*;
(

  input  logic hqm_gated_clk
, input  logic hqm_inp_gated_clk
, output logic hqm_proc_clk_en_lsp
, input  logic hqm_rst_prep_lsp
, input  logic hqm_gated_rst_b_lsp
, input  logic hqm_inp_gated_rst_b_lsp

, input  logic hqm_rst_prep_atm
, input  logic hqm_gated_rst_b_atm
, input  logic hqm_inp_gated_rst_b_atm

, input  logic hqm_gated_rst_b_start_lsp
, input  logic hqm_gated_rst_b_active_lsp
, output logic hqm_gated_rst_b_done_lsp

, input  logic hqm_gated_rst_b_start_atm
, input  logic hqm_gated_rst_b_active_atm
, output logic hqm_gated_rst_b_done_atm

, input logic aqed_clk_idle
, input logic aqed_unit_idle
, output logic aqed_clk_enable

, output logic                  lsp_unit_idle
, output logic                  lsp_unit_pipeidle
, output logic                  lsp_reset_done

, output logic                  ap_unit_idle
, output logic                  ap_unit_pipeidle
, output logic                  ap_reset_done

// CFG interface
, input  logic                  lsp_cfg_req_up_read
, input  logic                  lsp_cfg_req_up_write
, input  cfg_req_t              lsp_cfg_req_up
, input  logic                  lsp_cfg_rsp_up_ack
, input  cfg_rsp_t              lsp_cfg_rsp_up
, output logic                  lsp_cfg_req_down_read
, output logic                  lsp_cfg_req_down_write
, output cfg_req_t              lsp_cfg_req_down
, output logic                  lsp_cfg_rsp_down_ack
, output cfg_rsp_t              lsp_cfg_rsp_down

, input  logic                  ap_cfg_req_up_read
, input  logic                  ap_cfg_req_up_write
, input  cfg_req_t              ap_cfg_req_up
, input  logic                  ap_cfg_rsp_up_ack
, input  cfg_rsp_t              ap_cfg_rsp_up
, output logic                  ap_cfg_req_down_read
, output logic                  ap_cfg_req_down_write
, output cfg_req_t              ap_cfg_req_down
, output logic                  ap_cfg_rsp_down_ack
, output cfg_rsp_t              ap_cfg_rsp_down

// interrupt interface
, input  logic                  lsp_alarm_up_v
, output logic                  lsp_alarm_up_ready
, input  aw_alarm_t             lsp_alarm_up_data

, output logic                  lsp_alarm_down_v
, input  logic                  lsp_alarm_down_ready
, output aw_alarm_t             lsp_alarm_down_data

, input  logic                  ap_alarm_up_v
, output logic                  ap_alarm_up_ready
, input  aw_alarm_t             ap_alarm_up_data

, output logic                  ap_alarm_down_v
, input  logic                  ap_alarm_down_ready
, output aw_alarm_t             ap_alarm_down_data


, output logic                           lsp_aqed_cmp_v
, input  logic                           lsp_aqed_cmp_ready
, output lsp_aqed_cmp_t                  lsp_aqed_cmp_data

, input  logic                           aqed_lsp_dec_fid_cnt_v

// chp lsp PALB (Power Aware Load Balancing) interface
, input  logic [ HQM_NUM_LB_CQ - 1 : 0 ] chp_lsp_ldb_cq_off

// chp_lsp_cmp interface
, input  logic                  chp_lsp_cmp_v
, output logic                  chp_lsp_cmp_ready
, input  chp_lsp_cmp_t          chp_lsp_cmp_data

// qed_lsp_deq interface
, input  logic                  qed_lsp_deq_v
, input  qed_lsp_deq_t          qed_lsp_deq_data

// aqed_lsp_deq interface
, input  logic                  aqed_lsp_deq_v
, input  aqed_lsp_deq_t         aqed_lsp_deq_data

// chp_lsp_token interface
, input  logic                  chp_lsp_token_v
, output logic                  chp_lsp_token_ready
, input  chp_lsp_token_t        chp_lsp_token_data

// lsp_nalb_sch_unoord interface
, output logic                  lsp_nalb_sch_unoord_v
, input  logic                  lsp_nalb_sch_unoord_ready
, output lsp_nalb_sch_unoord_t  lsp_nalb_sch_unoord_data

// lsp_dp_sch_dir interface
, output logic                  lsp_dp_sch_dir_v
, input  logic                  lsp_dp_sch_dir_ready
, output lsp_dp_sch_dir_t       lsp_dp_sch_dir_data

// lsp_nalb_sch_rorply interface
, output logic                  lsp_nalb_sch_rorply_v
, input  logic                  lsp_nalb_sch_rorply_ready
, output lsp_nalb_sch_rorply_t  lsp_nalb_sch_rorply_data

// lsp_dp_sch_rorply interface
, output logic                  lsp_dp_sch_rorply_v
, input  logic                  lsp_dp_sch_rorply_ready
, output lsp_dp_sch_rorply_t    lsp_dp_sch_rorply_data

// lsp_nalb_sch_atq interface
, output logic                  lsp_nalb_sch_atq_v
, input  logic                  lsp_nalb_sch_atq_ready
, output lsp_nalb_sch_atq_t     lsp_nalb_sch_atq_data

// nalb_lsp_enq_lb interface
, input  logic                  nalb_lsp_enq_lb_v
, output logic                  nalb_lsp_enq_lb_ready
, input  nalb_lsp_enq_lb_t      nalb_lsp_enq_lb_data

// nalb_lsp_enq_rorpl interface
, input  logic                  nalb_lsp_enq_rorply_v
, output logic                  nalb_lsp_enq_rorply_ready
, input  nalb_lsp_enq_rorply_t  nalb_lsp_enq_rorply_data

// dp_lsp_enq_dir interface
, input  logic                  dp_lsp_enq_dir_v
, output logic                  dp_lsp_enq_dir_ready
, input  dp_lsp_enq_dir_t       dp_lsp_enq_dir_data

// dp_lsp_enq_rorply interface
, input  logic                  dp_lsp_enq_rorply_v
, output logic                  dp_lsp_enq_rorply_ready
, input  dp_lsp_enq_rorply_t    dp_lsp_enq_rorply_data

// rop_lsp_reordercmp interface
, input  logic                  rop_lsp_reordercmp_v
, output logic                  rop_lsp_reordercmp_ready
, input  rop_lsp_reordercmp_t   rop_lsp_reordercmp_data

// aqed_lsp_sch interface
, input  logic                  aqed_lsp_sch_v
, output logic                  aqed_lsp_sch_ready
, input  aqed_lsp_sch_t         aqed_lsp_sch_data

// ap_aqed interface
, output logic                  ap_aqed_v
, input  logic                  ap_aqed_ready
, output ap_aqed_t              ap_aqed_data

// aqed_ap_enq interface
, input  logic                  aqed_ap_enq_v
, output logic                  aqed_ap_enq_ready
, input  aqed_ap_enq_t          aqed_ap_enq_data

// aqed_lsp_fid_cnt_upd interface
, input logic                   aqed_lsp_fid_cnt_upd_v
, input logic                   aqed_lsp_fid_cnt_upd_val
, input logic [6:0]             aqed_lsp_fid_cnt_upd_qid
, input logic                   aqed_lsp_stop_atqatm

// Spares

, input  logic [1:0]            spare_qed_lsp
, input  logic [1:0]            spare_sys_lsp

, output logic [1:0]            spare_lsp_qed
, output logic [1:0]            spare_lsp_sys

// BEGIN HQM_MEMPORT_DECL hqm_list_sel_pipe_core
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_re
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_rclk
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_aqed_lsp_deq_fifo_mem_raddr
    ,output logic [(       5)-1:0] rf_aqed_lsp_deq_fifo_mem_waddr
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_we
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_wclk
    ,output logic                  rf_aqed_lsp_deq_fifo_mem_wclk_rst_n
    ,output logic [(       9)-1:0] rf_aqed_lsp_deq_fifo_mem_wdata
    ,input  logic [(       9)-1:0] rf_aqed_lsp_deq_fifo_mem_rdata

    ,output logic                  rf_atm_cmp_fifo_mem_re
    ,output logic                  rf_atm_cmp_fifo_mem_rclk
    ,output logic                  rf_atm_cmp_fifo_mem_rclk_rst_n
    ,output logic [(       3)-1:0] rf_atm_cmp_fifo_mem_raddr
    ,output logic [(       3)-1:0] rf_atm_cmp_fifo_mem_waddr
    ,output logic                  rf_atm_cmp_fifo_mem_we
    ,output logic                  rf_atm_cmp_fifo_mem_wclk
    ,output logic                  rf_atm_cmp_fifo_mem_wclk_rst_n
    ,output logic [(      55)-1:0] rf_atm_cmp_fifo_mem_wdata
    ,input  logic [(      55)-1:0] rf_atm_cmp_fifo_mem_rdata

    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_re
    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_rclk
    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_atm_qid_dpth_thrsh_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_atm_qid_dpth_thrsh_mem_waddr
    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_we
    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_wclk
    ,output logic                  rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n
    ,output logic [(      16)-1:0] rf_cfg_atm_qid_dpth_thrsh_mem_wdata
    ,input  logic [(      16)-1:0] rf_cfg_atm_qid_dpth_thrsh_mem_rdata

    ,output logic                  rf_cfg_cq2priov_mem_re
    ,output logic                  rf_cfg_cq2priov_mem_rclk
    ,output logic                  rf_cfg_cq2priov_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2priov_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2priov_mem_waddr
    ,output logic                  rf_cfg_cq2priov_mem_we
    ,output logic                  rf_cfg_cq2priov_mem_wclk
    ,output logic                  rf_cfg_cq2priov_mem_wclk_rst_n
    ,output logic [(      33)-1:0] rf_cfg_cq2priov_mem_wdata
    ,input  logic [(      33)-1:0] rf_cfg_cq2priov_mem_rdata

    ,output logic                  rf_cfg_cq2priov_odd_mem_re
    ,output logic                  rf_cfg_cq2priov_odd_mem_rclk
    ,output logic                  rf_cfg_cq2priov_odd_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2priov_odd_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2priov_odd_mem_waddr
    ,output logic                  rf_cfg_cq2priov_odd_mem_we
    ,output logic                  rf_cfg_cq2priov_odd_mem_wclk
    ,output logic                  rf_cfg_cq2priov_odd_mem_wclk_rst_n
    ,output logic [(      33)-1:0] rf_cfg_cq2priov_odd_mem_wdata
    ,input  logic [(      33)-1:0] rf_cfg_cq2priov_odd_mem_rdata

    ,output logic                  rf_cfg_cq2qid_0_mem_re
    ,output logic                  rf_cfg_cq2qid_0_mem_rclk
    ,output logic                  rf_cfg_cq2qid_0_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_0_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_0_mem_waddr
    ,output logic                  rf_cfg_cq2qid_0_mem_we
    ,output logic                  rf_cfg_cq2qid_0_mem_wclk
    ,output logic                  rf_cfg_cq2qid_0_mem_wclk_rst_n
    ,output logic [(      29)-1:0] rf_cfg_cq2qid_0_mem_wdata
    ,input  logic [(      29)-1:0] rf_cfg_cq2qid_0_mem_rdata

    ,output logic                  rf_cfg_cq2qid_0_odd_mem_re
    ,output logic                  rf_cfg_cq2qid_0_odd_mem_rclk
    ,output logic                  rf_cfg_cq2qid_0_odd_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_0_odd_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_0_odd_mem_waddr
    ,output logic                  rf_cfg_cq2qid_0_odd_mem_we
    ,output logic                  rf_cfg_cq2qid_0_odd_mem_wclk
    ,output logic                  rf_cfg_cq2qid_0_odd_mem_wclk_rst_n
    ,output logic [(      29)-1:0] rf_cfg_cq2qid_0_odd_mem_wdata
    ,input  logic [(      29)-1:0] rf_cfg_cq2qid_0_odd_mem_rdata

    ,output logic                  rf_cfg_cq2qid_1_mem_re
    ,output logic                  rf_cfg_cq2qid_1_mem_rclk
    ,output logic                  rf_cfg_cq2qid_1_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_1_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_1_mem_waddr
    ,output logic                  rf_cfg_cq2qid_1_mem_we
    ,output logic                  rf_cfg_cq2qid_1_mem_wclk
    ,output logic                  rf_cfg_cq2qid_1_mem_wclk_rst_n
    ,output logic [(      29)-1:0] rf_cfg_cq2qid_1_mem_wdata
    ,input  logic [(      29)-1:0] rf_cfg_cq2qid_1_mem_rdata

    ,output logic                  rf_cfg_cq2qid_1_odd_mem_re
    ,output logic                  rf_cfg_cq2qid_1_odd_mem_rclk
    ,output logic                  rf_cfg_cq2qid_1_odd_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_1_odd_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_cq2qid_1_odd_mem_waddr
    ,output logic                  rf_cfg_cq2qid_1_odd_mem_we
    ,output logic                  rf_cfg_cq2qid_1_odd_mem_wclk
    ,output logic                  rf_cfg_cq2qid_1_odd_mem_wclk_rst_n
    ,output logic [(      29)-1:0] rf_cfg_cq2qid_1_odd_mem_wdata
    ,input  logic [(      29)-1:0] rf_cfg_cq2qid_1_odd_mem_rdata

    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_re
    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_rclk
    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_inflight_limit_mem_raddr
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_inflight_limit_mem_waddr
    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_we
    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_wclk
    ,output logic                  rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n
    ,output logic [(      14)-1:0] rf_cfg_cq_ldb_inflight_limit_mem_wdata
    ,input  logic [(      14)-1:0] rf_cfg_cq_ldb_inflight_limit_mem_rdata

    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_re
    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_rclk
    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_inflight_threshold_mem_raddr
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_inflight_threshold_mem_waddr
    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_we
    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_wclk
    ,output logic                  rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n
    ,output logic [(      14)-1:0] rf_cfg_cq_ldb_inflight_threshold_mem_wdata
    ,input  logic [(      14)-1:0] rf_cfg_cq_ldb_inflight_threshold_mem_rdata

    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_re
    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_rclk
    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_token_depth_select_mem_raddr
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_token_depth_select_mem_waddr
    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_we
    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_wclk
    ,output logic                  rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_cq_ldb_token_depth_select_mem_wdata
    ,input  logic [(       5)-1:0] rf_cfg_cq_ldb_token_depth_select_mem_rdata

    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_re
    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_rclk
    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_wu_limit_mem_raddr
    ,output logic [(       6)-1:0] rf_cfg_cq_ldb_wu_limit_mem_waddr
    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_we
    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_wclk
    ,output logic                  rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_cfg_cq_ldb_wu_limit_mem_wdata
    ,input  logic [(      17)-1:0] rf_cfg_cq_ldb_wu_limit_mem_rdata

    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_re
    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_rclk
    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cfg_dir_qid_dpth_thrsh_mem_raddr
    ,output logic [(       6)-1:0] rf_cfg_dir_qid_dpth_thrsh_mem_waddr
    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_we
    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_wclk
    ,output logic                  rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n
    ,output logic [(      16)-1:0] rf_cfg_dir_qid_dpth_thrsh_mem_wdata
    ,input  logic [(      16)-1:0] rf_cfg_dir_qid_dpth_thrsh_mem_rdata

    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_re
    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_rclk
    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_nalb_qid_dpth_thrsh_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_nalb_qid_dpth_thrsh_mem_waddr
    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_we
    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_wclk
    ,output logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n
    ,output logic [(      16)-1:0] rf_cfg_nalb_qid_dpth_thrsh_mem_wdata
    ,input  logic [(      16)-1:0] rf_cfg_nalb_qid_dpth_thrsh_mem_rdata

    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_re
    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_rclk
    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_qid_aqed_active_limit_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_qid_aqed_active_limit_mem_waddr
    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_we
    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_wclk
    ,output logic                  rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n
    ,output logic [(      13)-1:0] rf_cfg_qid_aqed_active_limit_mem_wdata
    ,input  logic [(      13)-1:0] rf_cfg_qid_aqed_active_limit_mem_rdata

    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_re
    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_rclk
    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_inflight_limit_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_inflight_limit_mem_waddr
    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_we
    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_wclk
    ,output logic                  rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n
    ,output logic [(      13)-1:0] rf_cfg_qid_ldb_inflight_limit_mem_wdata
    ,input  logic [(      13)-1:0] rf_cfg_qid_ldb_inflight_limit_mem_rdata

    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_re
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_rclk
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_qid2cqidix2_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_qid2cqidix2_mem_waddr
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_we
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_wclk
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n
    ,output logic [(     528)-1:0] rf_cfg_qid_ldb_qid2cqidix2_mem_wdata
    ,input  logic [(     528)-1:0] rf_cfg_qid_ldb_qid2cqidix2_mem_rdata

    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_re
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_rclk
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_qid2cqidix_mem_raddr
    ,output logic [(       5)-1:0] rf_cfg_qid_ldb_qid2cqidix_mem_waddr
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_we
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_wclk
    ,output logic                  rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n
    ,output logic [(     528)-1:0] rf_cfg_qid_ldb_qid2cqidix_mem_wdata
    ,input  logic [(     528)-1:0] rf_cfg_qid_ldb_qid2cqidix_mem_rdata

    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_re
    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk
    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr
    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_we
    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk
    ,output logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      73)-1:0] rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata
    ,input  logic [(      73)-1:0] rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata

    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_re
    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_rclk
    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_chp_lsp_token_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_chp_lsp_token_rx_sync_fifo_mem_waddr
    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_we
    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_wclk
    ,output logic                  rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      25)-1:0] rf_chp_lsp_token_rx_sync_fifo_mem_wdata
    ,input  logic [(      25)-1:0] rf_chp_lsp_token_rx_sync_fifo_mem_rdata

    ,output logic                  rf_cq_atm_pri_arbindex_mem_re
    ,output logic                  rf_cq_atm_pri_arbindex_mem_rclk
    ,output logic                  rf_cq_atm_pri_arbindex_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cq_atm_pri_arbindex_mem_raddr
    ,output logic [(       5)-1:0] rf_cq_atm_pri_arbindex_mem_waddr
    ,output logic                  rf_cq_atm_pri_arbindex_mem_we
    ,output logic                  rf_cq_atm_pri_arbindex_mem_wclk
    ,output logic                  rf_cq_atm_pri_arbindex_mem_wclk_rst_n
    ,output logic [(      96)-1:0] rf_cq_atm_pri_arbindex_mem_wdata
    ,input  logic [(      96)-1:0] rf_cq_atm_pri_arbindex_mem_rdata

    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_re
    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_rclk
    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cq_dir_tot_sch_cnt_mem_raddr
    ,output logic [(       6)-1:0] rf_cq_dir_tot_sch_cnt_mem_waddr
    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_we
    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_wclk
    ,output logic                  rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n
    ,output logic [(      66)-1:0] rf_cq_dir_tot_sch_cnt_mem_wdata
    ,input  logic [(      66)-1:0] rf_cq_dir_tot_sch_cnt_mem_rdata

    ,output logic                  rf_cq_ldb_inflight_count_mem_re
    ,output logic                  rf_cq_ldb_inflight_count_mem_rclk
    ,output logic                  rf_cq_ldb_inflight_count_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cq_ldb_inflight_count_mem_raddr
    ,output logic [(       6)-1:0] rf_cq_ldb_inflight_count_mem_waddr
    ,output logic                  rf_cq_ldb_inflight_count_mem_we
    ,output logic                  rf_cq_ldb_inflight_count_mem_wclk
    ,output logic                  rf_cq_ldb_inflight_count_mem_wclk_rst_n
    ,output logic [(      15)-1:0] rf_cq_ldb_inflight_count_mem_wdata
    ,input  logic [(      15)-1:0] rf_cq_ldb_inflight_count_mem_rdata

    ,output logic                  rf_cq_ldb_token_count_mem_re
    ,output logic                  rf_cq_ldb_token_count_mem_rclk
    ,output logic                  rf_cq_ldb_token_count_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cq_ldb_token_count_mem_raddr
    ,output logic [(       6)-1:0] rf_cq_ldb_token_count_mem_waddr
    ,output logic                  rf_cq_ldb_token_count_mem_we
    ,output logic                  rf_cq_ldb_token_count_mem_wclk
    ,output logic                  rf_cq_ldb_token_count_mem_wclk_rst_n
    ,output logic [(      13)-1:0] rf_cq_ldb_token_count_mem_wdata
    ,input  logic [(      13)-1:0] rf_cq_ldb_token_count_mem_rdata

    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_re
    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_rclk
    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cq_ldb_tot_sch_cnt_mem_raddr
    ,output logic [(       6)-1:0] rf_cq_ldb_tot_sch_cnt_mem_waddr
    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_we
    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_wclk
    ,output logic                  rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n
    ,output logic [(      66)-1:0] rf_cq_ldb_tot_sch_cnt_mem_wdata
    ,input  logic [(      66)-1:0] rf_cq_ldb_tot_sch_cnt_mem_rdata

    ,output logic                  rf_cq_ldb_wu_count_mem_re
    ,output logic                  rf_cq_ldb_wu_count_mem_rclk
    ,output logic                  rf_cq_ldb_wu_count_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_cq_ldb_wu_count_mem_raddr
    ,output logic [(       6)-1:0] rf_cq_ldb_wu_count_mem_waddr
    ,output logic                  rf_cq_ldb_wu_count_mem_we
    ,output logic                  rf_cq_ldb_wu_count_mem_wclk
    ,output logic                  rf_cq_ldb_wu_count_mem_wclk_rst_n
    ,output logic [(      19)-1:0] rf_cq_ldb_wu_count_mem_wdata
    ,input  logic [(      19)-1:0] rf_cq_ldb_wu_count_mem_rdata

    ,output logic                  rf_cq_nalb_pri_arbindex_mem_re
    ,output logic                  rf_cq_nalb_pri_arbindex_mem_rclk
    ,output logic                  rf_cq_nalb_pri_arbindex_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_cq_nalb_pri_arbindex_mem_raddr
    ,output logic [(       5)-1:0] rf_cq_nalb_pri_arbindex_mem_waddr
    ,output logic                  rf_cq_nalb_pri_arbindex_mem_we
    ,output logic                  rf_cq_nalb_pri_arbindex_mem_wclk
    ,output logic                  rf_cq_nalb_pri_arbindex_mem_wclk_rst_n
    ,output logic [(      96)-1:0] rf_cq_nalb_pri_arbindex_mem_wdata
    ,input  logic [(      96)-1:0] rf_cq_nalb_pri_arbindex_mem_rdata

    ,output logic                  rf_dir_enq_cnt_mem_re
    ,output logic                  rf_dir_enq_cnt_mem_rclk
    ,output logic                  rf_dir_enq_cnt_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_dir_enq_cnt_mem_raddr
    ,output logic [(       6)-1:0] rf_dir_enq_cnt_mem_waddr
    ,output logic                  rf_dir_enq_cnt_mem_we
    ,output logic                  rf_dir_enq_cnt_mem_wclk
    ,output logic                  rf_dir_enq_cnt_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_dir_enq_cnt_mem_wdata
    ,input  logic [(      17)-1:0] rf_dir_enq_cnt_mem_rdata

    ,output logic                  rf_dir_tok_cnt_mem_re
    ,output logic                  rf_dir_tok_cnt_mem_rclk
    ,output logic                  rf_dir_tok_cnt_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_dir_tok_cnt_mem_raddr
    ,output logic [(       6)-1:0] rf_dir_tok_cnt_mem_waddr
    ,output logic                  rf_dir_tok_cnt_mem_we
    ,output logic                  rf_dir_tok_cnt_mem_wclk
    ,output logic                  rf_dir_tok_cnt_mem_wclk_rst_n
    ,output logic [(      13)-1:0] rf_dir_tok_cnt_mem_wdata
    ,input  logic [(      13)-1:0] rf_dir_tok_cnt_mem_rdata

    ,output logic                  rf_dir_tok_lim_mem_re
    ,output logic                  rf_dir_tok_lim_mem_rclk
    ,output logic                  rf_dir_tok_lim_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_dir_tok_lim_mem_raddr
    ,output logic [(       6)-1:0] rf_dir_tok_lim_mem_waddr
    ,output logic                  rf_dir_tok_lim_mem_we
    ,output logic                  rf_dir_tok_lim_mem_wclk
    ,output logic                  rf_dir_tok_lim_mem_wclk_rst_n
    ,output logic [(       8)-1:0] rf_dir_tok_lim_mem_wdata
    ,input  logic [(       8)-1:0] rf_dir_tok_lim_mem_rdata

    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re
    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk
    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr
    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we
    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk
    ,output logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(       8)-1:0] rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata
    ,input  logic [(       8)-1:0] rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata

    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re
    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk
    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr
    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we
    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk
    ,output logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      23)-1:0] rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata
    ,input  logic [(      23)-1:0] rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata

    ,output logic                  rf_enq_nalb_fifo_mem_re
    ,output logic                  rf_enq_nalb_fifo_mem_rclk
    ,output logic                  rf_enq_nalb_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_enq_nalb_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_enq_nalb_fifo_mem_waddr
    ,output logic                  rf_enq_nalb_fifo_mem_we
    ,output logic                  rf_enq_nalb_fifo_mem_wclk
    ,output logic                  rf_enq_nalb_fifo_mem_wclk_rst_n
    ,output logic [(      10)-1:0] rf_enq_nalb_fifo_mem_wdata
    ,input  logic [(      10)-1:0] rf_enq_nalb_fifo_mem_rdata

    ,output logic                  rf_ldb_token_rtn_fifo_mem_re
    ,output logic                  rf_ldb_token_rtn_fifo_mem_rclk
    ,output logic                  rf_ldb_token_rtn_fifo_mem_rclk_rst_n
    ,output logic [(       3)-1:0] rf_ldb_token_rtn_fifo_mem_raddr
    ,output logic [(       3)-1:0] rf_ldb_token_rtn_fifo_mem_waddr
    ,output logic                  rf_ldb_token_rtn_fifo_mem_we
    ,output logic                  rf_ldb_token_rtn_fifo_mem_wclk
    ,output logic                  rf_ldb_token_rtn_fifo_mem_wclk_rst_n
    ,output logic [(      25)-1:0] rf_ldb_token_rtn_fifo_mem_wdata
    ,input  logic [(      25)-1:0] rf_ldb_token_rtn_fifo_mem_rdata

    ,output logic                  rf_nalb_cmp_fifo_mem_re
    ,output logic                  rf_nalb_cmp_fifo_mem_rclk
    ,output logic                  rf_nalb_cmp_fifo_mem_rclk_rst_n
    ,output logic [(       3)-1:0] rf_nalb_cmp_fifo_mem_raddr
    ,output logic [(       3)-1:0] rf_nalb_cmp_fifo_mem_waddr
    ,output logic                  rf_nalb_cmp_fifo_mem_we
    ,output logic                  rf_nalb_cmp_fifo_mem_wclk
    ,output logic                  rf_nalb_cmp_fifo_mem_wclk_rst_n
    ,output logic [(      18)-1:0] rf_nalb_cmp_fifo_mem_wdata
    ,input  logic [(      18)-1:0] rf_nalb_cmp_fifo_mem_rdata

    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re
    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk
    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr
    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we
    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk
    ,output logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      10)-1:0] rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata
    ,input  logic [(      10)-1:0] rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata

    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re
    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk
    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr
    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we
    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk
    ,output logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      27)-1:0] rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata
    ,input  logic [(      27)-1:0] rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata

    ,output logic                  rf_nalb_sel_nalb_fifo_mem_re
    ,output logic                  rf_nalb_sel_nalb_fifo_mem_rclk
    ,output logic                  rf_nalb_sel_nalb_fifo_mem_rclk_rst_n
    ,output logic [(       4)-1:0] rf_nalb_sel_nalb_fifo_mem_raddr
    ,output logic [(       4)-1:0] rf_nalb_sel_nalb_fifo_mem_waddr
    ,output logic                  rf_nalb_sel_nalb_fifo_mem_we
    ,output logic                  rf_nalb_sel_nalb_fifo_mem_wclk
    ,output logic                  rf_nalb_sel_nalb_fifo_mem_wclk_rst_n
    ,output logic [(      27)-1:0] rf_nalb_sel_nalb_fifo_mem_wdata
    ,input  logic [(      27)-1:0] rf_nalb_sel_nalb_fifo_mem_rdata

    ,output logic                  rf_qed_lsp_deq_fifo_mem_re
    ,output logic                  rf_qed_lsp_deq_fifo_mem_rclk
    ,output logic                  rf_qed_lsp_deq_fifo_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qed_lsp_deq_fifo_mem_raddr
    ,output logic [(       5)-1:0] rf_qed_lsp_deq_fifo_mem_waddr
    ,output logic                  rf_qed_lsp_deq_fifo_mem_we
    ,output logic                  rf_qed_lsp_deq_fifo_mem_wclk
    ,output logic                  rf_qed_lsp_deq_fifo_mem_wclk_rst_n
    ,output logic [(       9)-1:0] rf_qed_lsp_deq_fifo_mem_wdata
    ,input  logic [(       9)-1:0] rf_qed_lsp_deq_fifo_mem_rdata

    ,output logic                  rf_qid_aqed_active_count_mem_re
    ,output logic                  rf_qid_aqed_active_count_mem_rclk
    ,output logic                  rf_qid_aqed_active_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_aqed_active_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_aqed_active_count_mem_waddr
    ,output logic                  rf_qid_aqed_active_count_mem_we
    ,output logic                  rf_qid_aqed_active_count_mem_wclk
    ,output logic                  rf_qid_aqed_active_count_mem_wclk_rst_n
    ,output logic [(      14)-1:0] rf_qid_aqed_active_count_mem_wdata
    ,input  logic [(      14)-1:0] rf_qid_aqed_active_count_mem_rdata

    ,output logic                  rf_qid_atm_active_mem_re
    ,output logic                  rf_qid_atm_active_mem_rclk
    ,output logic                  rf_qid_atm_active_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_atm_active_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_atm_active_mem_waddr
    ,output logic                  rf_qid_atm_active_mem_we
    ,output logic                  rf_qid_atm_active_mem_wclk
    ,output logic                  rf_qid_atm_active_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_qid_atm_active_mem_wdata
    ,input  logic [(      17)-1:0] rf_qid_atm_active_mem_rdata

    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_re
    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_rclk
    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_atm_tot_enq_cnt_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_atm_tot_enq_cnt_mem_waddr
    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_we
    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_wclk
    ,output logic                  rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n
    ,output logic [(      66)-1:0] rf_qid_atm_tot_enq_cnt_mem_wdata
    ,input  logic [(      66)-1:0] rf_qid_atm_tot_enq_cnt_mem_rdata

    ,output logic                  rf_qid_atq_enqueue_count_mem_re
    ,output logic                  rf_qid_atq_enqueue_count_mem_rclk
    ,output logic                  rf_qid_atq_enqueue_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_atq_enqueue_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_atq_enqueue_count_mem_waddr
    ,output logic                  rf_qid_atq_enqueue_count_mem_we
    ,output logic                  rf_qid_atq_enqueue_count_mem_wclk
    ,output logic                  rf_qid_atq_enqueue_count_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_qid_atq_enqueue_count_mem_wdata
    ,input  logic [(      17)-1:0] rf_qid_atq_enqueue_count_mem_rdata

    ,output logic                  rf_qid_dir_max_depth_mem_re
    ,output logic                  rf_qid_dir_max_depth_mem_rclk
    ,output logic                  rf_qid_dir_max_depth_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_qid_dir_max_depth_mem_raddr
    ,output logic [(       6)-1:0] rf_qid_dir_max_depth_mem_waddr
    ,output logic                  rf_qid_dir_max_depth_mem_we
    ,output logic                  rf_qid_dir_max_depth_mem_wclk
    ,output logic                  rf_qid_dir_max_depth_mem_wclk_rst_n
    ,output logic [(      15)-1:0] rf_qid_dir_max_depth_mem_wdata
    ,input  logic [(      15)-1:0] rf_qid_dir_max_depth_mem_rdata

    ,output logic                  rf_qid_dir_replay_count_mem_re
    ,output logic                  rf_qid_dir_replay_count_mem_rclk
    ,output logic                  rf_qid_dir_replay_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_dir_replay_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_dir_replay_count_mem_waddr
    ,output logic                  rf_qid_dir_replay_count_mem_we
    ,output logic                  rf_qid_dir_replay_count_mem_wclk
    ,output logic                  rf_qid_dir_replay_count_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_qid_dir_replay_count_mem_wdata
    ,input  logic [(      17)-1:0] rf_qid_dir_replay_count_mem_rdata

    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_re
    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_rclk
    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n
    ,output logic [(       6)-1:0] rf_qid_dir_tot_enq_cnt_mem_raddr
    ,output logic [(       6)-1:0] rf_qid_dir_tot_enq_cnt_mem_waddr
    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_we
    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_wclk
    ,output logic                  rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n
    ,output logic [(      66)-1:0] rf_qid_dir_tot_enq_cnt_mem_wdata
    ,input  logic [(      66)-1:0] rf_qid_dir_tot_enq_cnt_mem_rdata

    ,output logic                  rf_qid_ldb_enqueue_count_mem_re
    ,output logic                  rf_qid_ldb_enqueue_count_mem_rclk
    ,output logic                  rf_qid_ldb_enqueue_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_ldb_enqueue_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_ldb_enqueue_count_mem_waddr
    ,output logic                  rf_qid_ldb_enqueue_count_mem_we
    ,output logic                  rf_qid_ldb_enqueue_count_mem_wclk
    ,output logic                  rf_qid_ldb_enqueue_count_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_qid_ldb_enqueue_count_mem_wdata
    ,input  logic [(      17)-1:0] rf_qid_ldb_enqueue_count_mem_rdata

    ,output logic                  rf_qid_ldb_inflight_count_mem_re
    ,output logic                  rf_qid_ldb_inflight_count_mem_rclk
    ,output logic                  rf_qid_ldb_inflight_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_ldb_inflight_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_ldb_inflight_count_mem_waddr
    ,output logic                  rf_qid_ldb_inflight_count_mem_we
    ,output logic                  rf_qid_ldb_inflight_count_mem_wclk
    ,output logic                  rf_qid_ldb_inflight_count_mem_wclk_rst_n
    ,output logic [(      14)-1:0] rf_qid_ldb_inflight_count_mem_wdata
    ,input  logic [(      14)-1:0] rf_qid_ldb_inflight_count_mem_rdata

    ,output logic                  rf_qid_ldb_replay_count_mem_re
    ,output logic                  rf_qid_ldb_replay_count_mem_rclk
    ,output logic                  rf_qid_ldb_replay_count_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_ldb_replay_count_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_ldb_replay_count_mem_waddr
    ,output logic                  rf_qid_ldb_replay_count_mem_we
    ,output logic                  rf_qid_ldb_replay_count_mem_wclk
    ,output logic                  rf_qid_ldb_replay_count_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_qid_ldb_replay_count_mem_wdata
    ,input  logic [(      17)-1:0] rf_qid_ldb_replay_count_mem_rdata

    ,output logic                  rf_qid_naldb_max_depth_mem_re
    ,output logic                  rf_qid_naldb_max_depth_mem_rclk
    ,output logic                  rf_qid_naldb_max_depth_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_naldb_max_depth_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_naldb_max_depth_mem_waddr
    ,output logic                  rf_qid_naldb_max_depth_mem_we
    ,output logic                  rf_qid_naldb_max_depth_mem_wclk
    ,output logic                  rf_qid_naldb_max_depth_mem_wclk_rst_n
    ,output logic [(      15)-1:0] rf_qid_naldb_max_depth_mem_wdata
    ,input  logic [(      15)-1:0] rf_qid_naldb_max_depth_mem_rdata

    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_re
    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_rclk
    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_naldb_tot_enq_cnt_mem_raddr
    ,output logic [(       5)-1:0] rf_qid_naldb_tot_enq_cnt_mem_waddr
    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_we
    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_wclk
    ,output logic                  rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n
    ,output logic [(      66)-1:0] rf_qid_naldb_tot_enq_cnt_mem_wdata
    ,input  logic [(      66)-1:0] rf_qid_naldb_tot_enq_cnt_mem_rdata

    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re
    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk
    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       3)-1:0] rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr
    ,output logic [(       3)-1:0] rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr
    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we
    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk
    ,output logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      17)-1:0] rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata
    ,input  logic [(      17)-1:0] rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata

    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_re
    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_rclk
    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n
    ,output logic [(       2)-1:0] rf_send_atm_to_cq_rx_sync_fifo_mem_raddr
    ,output logic [(       2)-1:0] rf_send_atm_to_cq_rx_sync_fifo_mem_waddr
    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_we
    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_wclk
    ,output logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n
    ,output logic [(      35)-1:0] rf_send_atm_to_cq_rx_sync_fifo_mem_wdata
    ,input  logic [(      35)-1:0] rf_send_atm_to_cq_rx_sync_fifo_mem_rdata

    ,output logic                  rf_uno_atm_cmp_fifo_mem_re
    ,output logic                  rf_uno_atm_cmp_fifo_mem_rclk
    ,output logic                  rf_uno_atm_cmp_fifo_mem_rclk_rst_n
    ,output logic [(       3)-1:0] rf_uno_atm_cmp_fifo_mem_raddr
    ,output logic [(       3)-1:0] rf_uno_atm_cmp_fifo_mem_waddr
    ,output logic                  rf_uno_atm_cmp_fifo_mem_we
    ,output logic                  rf_uno_atm_cmp_fifo_mem_wclk
    ,output logic                  rf_uno_atm_cmp_fifo_mem_wclk_rst_n
    ,output logic [(      20)-1:0] rf_uno_atm_cmp_fifo_mem_wdata
    ,input  logic [(      20)-1:0] rf_uno_atm_cmp_fifo_mem_rdata

// END HQM_MEMPORT_DECL hqm_list_sel_pipe_core
// BEGIN HQM_MEMPORT_DECL hqm_lsp_atm_pipe
    ,output logic                  rf_aqed_qid2cqidix_re
    ,output logic                  rf_aqed_qid2cqidix_rclk
    ,output logic                  rf_aqed_qid2cqidix_rclk_rst_n
    ,output logic [(       5)-1:0] rf_aqed_qid2cqidix_raddr
    ,output logic [(       5)-1:0] rf_aqed_qid2cqidix_waddr
    ,output logic                  rf_aqed_qid2cqidix_we
    ,output logic                  rf_aqed_qid2cqidix_wclk
    ,output logic                  rf_aqed_qid2cqidix_wclk_rst_n
    ,output logic [(     528)-1:0] rf_aqed_qid2cqidix_wdata
    ,input  logic [(     528)-1:0] rf_aqed_qid2cqidix_rdata

    ,output logic                  rf_atm_fifo_ap_aqed_re
    ,output logic                  rf_atm_fifo_ap_aqed_rclk
    ,output logic                  rf_atm_fifo_ap_aqed_rclk_rst_n
    ,output logic [(       4)-1:0] rf_atm_fifo_ap_aqed_raddr
    ,output logic [(       4)-1:0] rf_atm_fifo_ap_aqed_waddr
    ,output logic                  rf_atm_fifo_ap_aqed_we
    ,output logic                  rf_atm_fifo_ap_aqed_wclk
    ,output logic                  rf_atm_fifo_ap_aqed_wclk_rst_n
    ,output logic [(      45)-1:0] rf_atm_fifo_ap_aqed_wdata
    ,input  logic [(      45)-1:0] rf_atm_fifo_ap_aqed_rdata

    ,output logic                  rf_atm_fifo_aqed_ap_enq_re
    ,output logic                  rf_atm_fifo_aqed_ap_enq_rclk
    ,output logic                  rf_atm_fifo_aqed_ap_enq_rclk_rst_n
    ,output logic [(       5)-1:0] rf_atm_fifo_aqed_ap_enq_raddr
    ,output logic [(       5)-1:0] rf_atm_fifo_aqed_ap_enq_waddr
    ,output logic                  rf_atm_fifo_aqed_ap_enq_we
    ,output logic                  rf_atm_fifo_aqed_ap_enq_wclk
    ,output logic                  rf_atm_fifo_aqed_ap_enq_wclk_rst_n
    ,output logic [(      24)-1:0] rf_atm_fifo_aqed_ap_enq_wdata
    ,input  logic [(      24)-1:0] rf_atm_fifo_aqed_ap_enq_rdata

    ,output logic                  rf_fid2cqqidix_re
    ,output logic                  rf_fid2cqqidix_rclk
    ,output logic                  rf_fid2cqqidix_rclk_rst_n
    ,output logic [(      11)-1:0] rf_fid2cqqidix_raddr
    ,output logic [(      11)-1:0] rf_fid2cqqidix_waddr
    ,output logic                  rf_fid2cqqidix_we
    ,output logic                  rf_fid2cqqidix_wclk
    ,output logic                  rf_fid2cqqidix_wclk_rst_n
    ,output logic [(      12)-1:0] rf_fid2cqqidix_wdata
    ,input  logic [(      12)-1:0] rf_fid2cqqidix_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_re
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup0_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup0_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_we
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup0_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup0_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_re
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup1_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup1_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_we
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup1_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup1_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_re
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup2_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup2_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_we
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup2_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup2_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_re
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup3_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin0_dup3_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_we
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup3_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin0_dup3_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_re
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup0_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup0_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_we
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup0_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup0_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_re
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup1_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup1_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_we
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup1_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup1_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_re
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup2_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup2_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_we
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup2_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup2_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_re
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup3_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin1_dup3_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_we
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup3_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin1_dup3_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_re
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup0_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup0_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_we
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup0_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup0_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_re
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup1_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup1_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_we
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup1_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup1_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_re
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup2_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup2_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_we
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup2_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup2_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_re
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup3_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin2_dup3_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_we
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup3_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin2_dup3_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_re
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup0_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup0_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_we
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup0_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup0_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_re
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup1_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup1_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_we
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup1_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup1_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_re
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup2_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup2_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_we
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup2_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup2_rdata

    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_re
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_rclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup3_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_r_bin3_dup3_waddr
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_we
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_wclk
    ,output logic                  rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup3_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_r_bin3_dup3_rdata

    ,output logic                  rf_ll_enq_cnt_s_bin0_re
    ,output logic                  rf_ll_enq_cnt_s_bin0_rclk
    ,output logic                  rf_ll_enq_cnt_s_bin0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin0_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin0_waddr
    ,output logic                  rf_ll_enq_cnt_s_bin0_we
    ,output logic                  rf_ll_enq_cnt_s_bin0_wclk
    ,output logic                  rf_ll_enq_cnt_s_bin0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_s_bin0_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_s_bin0_rdata

    ,output logic                  rf_ll_enq_cnt_s_bin1_re
    ,output logic                  rf_ll_enq_cnt_s_bin1_rclk
    ,output logic                  rf_ll_enq_cnt_s_bin1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin1_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin1_waddr
    ,output logic                  rf_ll_enq_cnt_s_bin1_we
    ,output logic                  rf_ll_enq_cnt_s_bin1_wclk
    ,output logic                  rf_ll_enq_cnt_s_bin1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_s_bin1_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_s_bin1_rdata

    ,output logic                  rf_ll_enq_cnt_s_bin2_re
    ,output logic                  rf_ll_enq_cnt_s_bin2_rclk
    ,output logic                  rf_ll_enq_cnt_s_bin2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin2_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin2_waddr
    ,output logic                  rf_ll_enq_cnt_s_bin2_we
    ,output logic                  rf_ll_enq_cnt_s_bin2_wclk
    ,output logic                  rf_ll_enq_cnt_s_bin2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_s_bin2_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_s_bin2_rdata

    ,output logic                  rf_ll_enq_cnt_s_bin3_re
    ,output logic                  rf_ll_enq_cnt_s_bin3_rclk
    ,output logic                  rf_ll_enq_cnt_s_bin3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin3_raddr
    ,output logic [(      11)-1:0] rf_ll_enq_cnt_s_bin3_waddr
    ,output logic                  rf_ll_enq_cnt_s_bin3_we
    ,output logic                  rf_ll_enq_cnt_s_bin3_wclk
    ,output logic                  rf_ll_enq_cnt_s_bin3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_enq_cnt_s_bin3_wdata
    ,input  logic [(      16)-1:0] rf_ll_enq_cnt_s_bin3_rdata

    ,output logic                  rf_ll_rdylst_hp_bin0_re
    ,output logic                  rf_ll_rdylst_hp_bin0_rclk
    ,output logic                  rf_ll_rdylst_hp_bin0_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin0_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin0_waddr
    ,output logic                  rf_ll_rdylst_hp_bin0_we
    ,output logic                  rf_ll_rdylst_hp_bin0_wclk
    ,output logic                  rf_ll_rdylst_hp_bin0_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_hp_bin0_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_hp_bin0_rdata

    ,output logic                  rf_ll_rdylst_hp_bin1_re
    ,output logic                  rf_ll_rdylst_hp_bin1_rclk
    ,output logic                  rf_ll_rdylst_hp_bin1_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin1_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin1_waddr
    ,output logic                  rf_ll_rdylst_hp_bin1_we
    ,output logic                  rf_ll_rdylst_hp_bin1_wclk
    ,output logic                  rf_ll_rdylst_hp_bin1_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_hp_bin1_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_hp_bin1_rdata

    ,output logic                  rf_ll_rdylst_hp_bin2_re
    ,output logic                  rf_ll_rdylst_hp_bin2_rclk
    ,output logic                  rf_ll_rdylst_hp_bin2_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin2_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin2_waddr
    ,output logic                  rf_ll_rdylst_hp_bin2_we
    ,output logic                  rf_ll_rdylst_hp_bin2_wclk
    ,output logic                  rf_ll_rdylst_hp_bin2_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_hp_bin2_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_hp_bin2_rdata

    ,output logic                  rf_ll_rdylst_hp_bin3_re
    ,output logic                  rf_ll_rdylst_hp_bin3_rclk
    ,output logic                  rf_ll_rdylst_hp_bin3_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin3_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_hp_bin3_waddr
    ,output logic                  rf_ll_rdylst_hp_bin3_we
    ,output logic                  rf_ll_rdylst_hp_bin3_wclk
    ,output logic                  rf_ll_rdylst_hp_bin3_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_hp_bin3_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_hp_bin3_rdata

    ,output logic                  rf_ll_rdylst_hpnxt_bin0_re
    ,output logic                  rf_ll_rdylst_hpnxt_bin0_rclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin0_raddr
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin0_waddr
    ,output logic                  rf_ll_rdylst_hpnxt_bin0_we
    ,output logic                  rf_ll_rdylst_hpnxt_bin0_wclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin0_wdata
    ,input  logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin0_rdata

    ,output logic                  rf_ll_rdylst_hpnxt_bin1_re
    ,output logic                  rf_ll_rdylst_hpnxt_bin1_rclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin1_raddr
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin1_waddr
    ,output logic                  rf_ll_rdylst_hpnxt_bin1_we
    ,output logic                  rf_ll_rdylst_hpnxt_bin1_wclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin1_wdata
    ,input  logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin1_rdata

    ,output logic                  rf_ll_rdylst_hpnxt_bin2_re
    ,output logic                  rf_ll_rdylst_hpnxt_bin2_rclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin2_raddr
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin2_waddr
    ,output logic                  rf_ll_rdylst_hpnxt_bin2_we
    ,output logic                  rf_ll_rdylst_hpnxt_bin2_wclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin2_wdata
    ,input  logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin2_rdata

    ,output logic                  rf_ll_rdylst_hpnxt_bin3_re
    ,output logic                  rf_ll_rdylst_hpnxt_bin3_rclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin3_raddr
    ,output logic [(      11)-1:0] rf_ll_rdylst_hpnxt_bin3_waddr
    ,output logic                  rf_ll_rdylst_hpnxt_bin3_we
    ,output logic                  rf_ll_rdylst_hpnxt_bin3_wclk
    ,output logic                  rf_ll_rdylst_hpnxt_bin3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin3_wdata
    ,input  logic [(      16)-1:0] rf_ll_rdylst_hpnxt_bin3_rdata

    ,output logic                  rf_ll_rdylst_tp_bin0_re
    ,output logic                  rf_ll_rdylst_tp_bin0_rclk
    ,output logic                  rf_ll_rdylst_tp_bin0_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin0_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin0_waddr
    ,output logic                  rf_ll_rdylst_tp_bin0_we
    ,output logic                  rf_ll_rdylst_tp_bin0_wclk
    ,output logic                  rf_ll_rdylst_tp_bin0_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_tp_bin0_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_tp_bin0_rdata

    ,output logic                  rf_ll_rdylst_tp_bin1_re
    ,output logic                  rf_ll_rdylst_tp_bin1_rclk
    ,output logic                  rf_ll_rdylst_tp_bin1_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin1_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin1_waddr
    ,output logic                  rf_ll_rdylst_tp_bin1_we
    ,output logic                  rf_ll_rdylst_tp_bin1_wclk
    ,output logic                  rf_ll_rdylst_tp_bin1_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_tp_bin1_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_tp_bin1_rdata

    ,output logic                  rf_ll_rdylst_tp_bin2_re
    ,output logic                  rf_ll_rdylst_tp_bin2_rclk
    ,output logic                  rf_ll_rdylst_tp_bin2_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin2_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin2_waddr
    ,output logic                  rf_ll_rdylst_tp_bin2_we
    ,output logic                  rf_ll_rdylst_tp_bin2_wclk
    ,output logic                  rf_ll_rdylst_tp_bin2_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_tp_bin2_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_tp_bin2_rdata

    ,output logic                  rf_ll_rdylst_tp_bin3_re
    ,output logic                  rf_ll_rdylst_tp_bin3_rclk
    ,output logic                  rf_ll_rdylst_tp_bin3_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin3_raddr
    ,output logic [(       5)-1:0] rf_ll_rdylst_tp_bin3_waddr
    ,output logic                  rf_ll_rdylst_tp_bin3_we
    ,output logic                  rf_ll_rdylst_tp_bin3_wclk
    ,output logic                  rf_ll_rdylst_tp_bin3_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_rdylst_tp_bin3_wdata
    ,input  logic [(      14)-1:0] rf_ll_rdylst_tp_bin3_rdata

    ,output logic                  rf_ll_rlst_cnt_re
    ,output logic                  rf_ll_rlst_cnt_rclk
    ,output logic                  rf_ll_rlst_cnt_rclk_rst_n
    ,output logic [(       5)-1:0] rf_ll_rlst_cnt_raddr
    ,output logic [(       5)-1:0] rf_ll_rlst_cnt_waddr
    ,output logic                  rf_ll_rlst_cnt_we
    ,output logic                  rf_ll_rlst_cnt_wclk
    ,output logic                  rf_ll_rlst_cnt_wclk_rst_n
    ,output logic [(      56)-1:0] rf_ll_rlst_cnt_wdata
    ,input  logic [(      56)-1:0] rf_ll_rlst_cnt_rdata

    ,output logic                  rf_ll_sch_cnt_dup0_re
    ,output logic                  rf_ll_sch_cnt_dup0_rclk
    ,output logic                  rf_ll_sch_cnt_dup0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup0_raddr
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup0_waddr
    ,output logic                  rf_ll_sch_cnt_dup0_we
    ,output logic                  rf_ll_sch_cnt_dup0_wclk
    ,output logic                  rf_ll_sch_cnt_dup0_wclk_rst_n
    ,output logic [(      17)-1:0] rf_ll_sch_cnt_dup0_wdata
    ,input  logic [(      17)-1:0] rf_ll_sch_cnt_dup0_rdata

    ,output logic                  rf_ll_sch_cnt_dup1_re
    ,output logic                  rf_ll_sch_cnt_dup1_rclk
    ,output logic                  rf_ll_sch_cnt_dup1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup1_raddr
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup1_waddr
    ,output logic                  rf_ll_sch_cnt_dup1_we
    ,output logic                  rf_ll_sch_cnt_dup1_wclk
    ,output logic                  rf_ll_sch_cnt_dup1_wclk_rst_n
    ,output logic [(      17)-1:0] rf_ll_sch_cnt_dup1_wdata
    ,input  logic [(      17)-1:0] rf_ll_sch_cnt_dup1_rdata

    ,output logic                  rf_ll_sch_cnt_dup2_re
    ,output logic                  rf_ll_sch_cnt_dup2_rclk
    ,output logic                  rf_ll_sch_cnt_dup2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup2_raddr
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup2_waddr
    ,output logic                  rf_ll_sch_cnt_dup2_we
    ,output logic                  rf_ll_sch_cnt_dup2_wclk
    ,output logic                  rf_ll_sch_cnt_dup2_wclk_rst_n
    ,output logic [(      17)-1:0] rf_ll_sch_cnt_dup2_wdata
    ,input  logic [(      17)-1:0] rf_ll_sch_cnt_dup2_rdata

    ,output logic                  rf_ll_sch_cnt_dup3_re
    ,output logic                  rf_ll_sch_cnt_dup3_rclk
    ,output logic                  rf_ll_sch_cnt_dup3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup3_raddr
    ,output logic [(      11)-1:0] rf_ll_sch_cnt_dup3_waddr
    ,output logic                  rf_ll_sch_cnt_dup3_we
    ,output logic                  rf_ll_sch_cnt_dup3_wclk
    ,output logic                  rf_ll_sch_cnt_dup3_wclk_rst_n
    ,output logic [(      17)-1:0] rf_ll_sch_cnt_dup3_wdata
    ,input  logic [(      17)-1:0] rf_ll_sch_cnt_dup3_rdata

    ,output logic                  rf_ll_schlst_hp_bin0_re
    ,output logic                  rf_ll_schlst_hp_bin0_rclk
    ,output logic                  rf_ll_schlst_hp_bin0_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin0_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin0_waddr
    ,output logic                  rf_ll_schlst_hp_bin0_we
    ,output logic                  rf_ll_schlst_hp_bin0_wclk
    ,output logic                  rf_ll_schlst_hp_bin0_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_hp_bin0_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_hp_bin0_rdata

    ,output logic                  rf_ll_schlst_hp_bin1_re
    ,output logic                  rf_ll_schlst_hp_bin1_rclk
    ,output logic                  rf_ll_schlst_hp_bin1_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin1_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin1_waddr
    ,output logic                  rf_ll_schlst_hp_bin1_we
    ,output logic                  rf_ll_schlst_hp_bin1_wclk
    ,output logic                  rf_ll_schlst_hp_bin1_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_hp_bin1_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_hp_bin1_rdata

    ,output logic                  rf_ll_schlst_hp_bin2_re
    ,output logic                  rf_ll_schlst_hp_bin2_rclk
    ,output logic                  rf_ll_schlst_hp_bin2_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin2_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin2_waddr
    ,output logic                  rf_ll_schlst_hp_bin2_we
    ,output logic                  rf_ll_schlst_hp_bin2_wclk
    ,output logic                  rf_ll_schlst_hp_bin2_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_hp_bin2_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_hp_bin2_rdata

    ,output logic                  rf_ll_schlst_hp_bin3_re
    ,output logic                  rf_ll_schlst_hp_bin3_rclk
    ,output logic                  rf_ll_schlst_hp_bin3_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin3_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_hp_bin3_waddr
    ,output logic                  rf_ll_schlst_hp_bin3_we
    ,output logic                  rf_ll_schlst_hp_bin3_wclk
    ,output logic                  rf_ll_schlst_hp_bin3_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_hp_bin3_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_hp_bin3_rdata

    ,output logic                  rf_ll_schlst_hpnxt_bin0_re
    ,output logic                  rf_ll_schlst_hpnxt_bin0_rclk
    ,output logic                  rf_ll_schlst_hpnxt_bin0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin0_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin0_waddr
    ,output logic                  rf_ll_schlst_hpnxt_bin0_we
    ,output logic                  rf_ll_schlst_hpnxt_bin0_wclk
    ,output logic                  rf_ll_schlst_hpnxt_bin0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin0_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin0_rdata

    ,output logic                  rf_ll_schlst_hpnxt_bin1_re
    ,output logic                  rf_ll_schlst_hpnxt_bin1_rclk
    ,output logic                  rf_ll_schlst_hpnxt_bin1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin1_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin1_waddr
    ,output logic                  rf_ll_schlst_hpnxt_bin1_we
    ,output logic                  rf_ll_schlst_hpnxt_bin1_wclk
    ,output logic                  rf_ll_schlst_hpnxt_bin1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin1_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin1_rdata

    ,output logic                  rf_ll_schlst_hpnxt_bin2_re
    ,output logic                  rf_ll_schlst_hpnxt_bin2_rclk
    ,output logic                  rf_ll_schlst_hpnxt_bin2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin2_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin2_waddr
    ,output logic                  rf_ll_schlst_hpnxt_bin2_we
    ,output logic                  rf_ll_schlst_hpnxt_bin2_wclk
    ,output logic                  rf_ll_schlst_hpnxt_bin2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin2_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin2_rdata

    ,output logic                  rf_ll_schlst_hpnxt_bin3_re
    ,output logic                  rf_ll_schlst_hpnxt_bin3_rclk
    ,output logic                  rf_ll_schlst_hpnxt_bin3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin3_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_hpnxt_bin3_waddr
    ,output logic                  rf_ll_schlst_hpnxt_bin3_we
    ,output logic                  rf_ll_schlst_hpnxt_bin3_wclk
    ,output logic                  rf_ll_schlst_hpnxt_bin3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin3_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_hpnxt_bin3_rdata

    ,output logic                  rf_ll_schlst_tp_bin0_re
    ,output logic                  rf_ll_schlst_tp_bin0_rclk
    ,output logic                  rf_ll_schlst_tp_bin0_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin0_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin0_waddr
    ,output logic                  rf_ll_schlst_tp_bin0_we
    ,output logic                  rf_ll_schlst_tp_bin0_wclk
    ,output logic                  rf_ll_schlst_tp_bin0_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_tp_bin0_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_tp_bin0_rdata

    ,output logic                  rf_ll_schlst_tp_bin1_re
    ,output logic                  rf_ll_schlst_tp_bin1_rclk
    ,output logic                  rf_ll_schlst_tp_bin1_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin1_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin1_waddr
    ,output logic                  rf_ll_schlst_tp_bin1_we
    ,output logic                  rf_ll_schlst_tp_bin1_wclk
    ,output logic                  rf_ll_schlst_tp_bin1_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_tp_bin1_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_tp_bin1_rdata

    ,output logic                  rf_ll_schlst_tp_bin2_re
    ,output logic                  rf_ll_schlst_tp_bin2_rclk
    ,output logic                  rf_ll_schlst_tp_bin2_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin2_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin2_waddr
    ,output logic                  rf_ll_schlst_tp_bin2_we
    ,output logic                  rf_ll_schlst_tp_bin2_wclk
    ,output logic                  rf_ll_schlst_tp_bin2_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_tp_bin2_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_tp_bin2_rdata

    ,output logic                  rf_ll_schlst_tp_bin3_re
    ,output logic                  rf_ll_schlst_tp_bin3_rclk
    ,output logic                  rf_ll_schlst_tp_bin3_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin3_raddr
    ,output logic [(       9)-1:0] rf_ll_schlst_tp_bin3_waddr
    ,output logic                  rf_ll_schlst_tp_bin3_we
    ,output logic                  rf_ll_schlst_tp_bin3_wclk
    ,output logic                  rf_ll_schlst_tp_bin3_wclk_rst_n
    ,output logic [(      14)-1:0] rf_ll_schlst_tp_bin3_wdata
    ,input  logic [(      14)-1:0] rf_ll_schlst_tp_bin3_rdata

    ,output logic                  rf_ll_schlst_tpprv_bin0_re
    ,output logic                  rf_ll_schlst_tpprv_bin0_rclk
    ,output logic                  rf_ll_schlst_tpprv_bin0_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin0_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin0_waddr
    ,output logic                  rf_ll_schlst_tpprv_bin0_we
    ,output logic                  rf_ll_schlst_tpprv_bin0_wclk
    ,output logic                  rf_ll_schlst_tpprv_bin0_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_tpprv_bin0_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_tpprv_bin0_rdata

    ,output logic                  rf_ll_schlst_tpprv_bin1_re
    ,output logic                  rf_ll_schlst_tpprv_bin1_rclk
    ,output logic                  rf_ll_schlst_tpprv_bin1_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin1_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin1_waddr
    ,output logic                  rf_ll_schlst_tpprv_bin1_we
    ,output logic                  rf_ll_schlst_tpprv_bin1_wclk
    ,output logic                  rf_ll_schlst_tpprv_bin1_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_tpprv_bin1_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_tpprv_bin1_rdata

    ,output logic                  rf_ll_schlst_tpprv_bin2_re
    ,output logic                  rf_ll_schlst_tpprv_bin2_rclk
    ,output logic                  rf_ll_schlst_tpprv_bin2_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin2_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin2_waddr
    ,output logic                  rf_ll_schlst_tpprv_bin2_we
    ,output logic                  rf_ll_schlst_tpprv_bin2_wclk
    ,output logic                  rf_ll_schlst_tpprv_bin2_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_tpprv_bin2_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_tpprv_bin2_rdata

    ,output logic                  rf_ll_schlst_tpprv_bin3_re
    ,output logic                  rf_ll_schlst_tpprv_bin3_rclk
    ,output logic                  rf_ll_schlst_tpprv_bin3_rclk_rst_n
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin3_raddr
    ,output logic [(      11)-1:0] rf_ll_schlst_tpprv_bin3_waddr
    ,output logic                  rf_ll_schlst_tpprv_bin3_we
    ,output logic                  rf_ll_schlst_tpprv_bin3_wclk
    ,output logic                  rf_ll_schlst_tpprv_bin3_wclk_rst_n
    ,output logic [(      16)-1:0] rf_ll_schlst_tpprv_bin3_wdata
    ,input  logic [(      16)-1:0] rf_ll_schlst_tpprv_bin3_rdata

    ,output logic                  rf_ll_slst_cnt_re
    ,output logic                  rf_ll_slst_cnt_rclk
    ,output logic                  rf_ll_slst_cnt_rclk_rst_n
    ,output logic [(       9)-1:0] rf_ll_slst_cnt_raddr
    ,output logic [(       9)-1:0] rf_ll_slst_cnt_waddr
    ,output logic                  rf_ll_slst_cnt_we
    ,output logic                  rf_ll_slst_cnt_wclk
    ,output logic                  rf_ll_slst_cnt_wclk_rst_n
    ,output logic [(      60)-1:0] rf_ll_slst_cnt_wdata
    ,input  logic [(      60)-1:0] rf_ll_slst_cnt_rdata

    ,output logic                  rf_qid_rdylst_clamp_re
    ,output logic                  rf_qid_rdylst_clamp_rclk
    ,output logic                  rf_qid_rdylst_clamp_rclk_rst_n
    ,output logic [(       5)-1:0] rf_qid_rdylst_clamp_raddr
    ,output logic [(       5)-1:0] rf_qid_rdylst_clamp_waddr
    ,output logic                  rf_qid_rdylst_clamp_we
    ,output logic                  rf_qid_rdylst_clamp_wclk
    ,output logic                  rf_qid_rdylst_clamp_wclk_rst_n
    ,output logic [(       6)-1:0] rf_qid_rdylst_clamp_wdata
    ,input  logic [(       6)-1:0] rf_qid_rdylst_clamp_rdata

// END HQM_MEMPORT_DECL hqm_lsp_atm_pipe
) ;


typedef struct packed {
  logic                                         qid_p ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]         qid ;
} lsp_lb_qid_t ;

typedef struct packed {
  logic                                         qid_p ;
  logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]        qid ;
} lsp_dir_qid_t ;

localparam      HQM_LSP_ARCH_CNT_MEM_WIDTH              = $bits( lsp_arch_cnt_t ) ;

localparam      HQM_LSP_CFG_DIAG_0_SLIST_V              = 0 ;
localparam      HQM_LSP_CFG_DIAG_0_SLIST_BLAST          = 1 ;
localparam      HQM_LSP_CFG_DIAG_0_RLIST_V              = 2 ;
localparam      HQM_LSP_CFG_DIAG_0_RLIST_BLAST          = 3 ;
localparam      HQM_LSP_CFG_DIAG_0_NALB_V               = 4 ;
localparam      HQM_LSP_CFG_DIAG_0_NALB_BLAST           = 5 ;
localparam      HQM_LSP_CFG_DIAG_0_CMPBLAST_CHKV        = 6 ;
localparam      HQM_LSP_CFG_DIAG_0_CMPBLAST             = 7 ;
localparam      HQM_LSP_CFG_DIAG_0_ATQ_QID_DIS          = 8 ;
localparam      HQM_LSP_CFG_DIAG_0_CQ_BUSY              = 9 ;
localparam      HQM_LSP_CFG_DIAG_0_CQ_NO_SPACE          = 10 ;
localparam      HQM_LSP_CFG_DIAG_0_DIR_TOK_V            = 11 ;
localparam      HQM_LSP_CFG_DIAG_0_ATQ_ACT_V            = 12 ;
localparam      HQM_LSP_CFG_DIAG_0_ATM_HASWORK_V        = 13 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_TOK_V             = 14 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_CMP_V             = 15 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT0       = 16 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT1       = 17 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT2       = 18 ;
localparam      HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT3       = 19 ;

localparam      HQM_LSP_CFG_DIAG_0_QED_CRED_AFULL       = 20 ;
localparam      HQM_LSP_CFG_DIAG_0_AQED_CRED_AFULL      = 21 ;
localparam      HQM_LSP_CFG_DIAG_0_LBA_OW_ANY           = 22 ;
localparam      HQM_LSP_CFG_DIAG_0_STOP_ATQATM          = 23 ;
localparam      HQM_LSP_CFG_DIAG_0_NSN_FCERR_RPTD       = 24 ;
localparam      HQM_LSP_CFG_DIAG_0_AQED_EMPTY           = 25 ;
localparam      HQM_LSP_CFG_DIAG_0_ATM_IF_V             = 26 ;
localparam      HQM_LSP_CFG_DIAG_0_TOT_IF_V             = 27 ;
localparam      HQM_LSP_CFG_DIAG_0_LBWU_P1_V            = 28 ;
localparam      HQM_LSP_CFG_DIAG_0_LBWU_P2_V            = 29 ;
localparam      HQM_LSP_CFG_DIAG_0_LBWU_P3_V            = 30 ;
localparam      HQM_LSP_CFG_DIAG_0_LBWU_P4_V            = 31 ;

localparam      HQM_LSP_VF_RESET_CMD_INIT_RESET         = 12'h001 ;     // Should never go here from other state, only (hw) reset
localparam      HQM_LSP_VF_RESET_CMD_START              = 12'h001 ;
localparam      HQM_LSP_VF_RESET_CMD_DIR_CQ_WRITE       = 12'h002 ;
localparam      HQM_LSP_VF_RESET_CMD_DIR_QID_WRITE      = 12'h004 ;
localparam      HQM_LSP_VF_RESET_CMD_LDB_CQ_READ        = 12'h008 ;
localparam      HQM_LSP_VF_RESET_CMD_LDB_QID_READ       = 12'h010 ;
localparam      HQM_LSP_VF_RESET_CMD_LDB_CQ_WRITE       = 12'h020 ;
localparam      HQM_LSP_VF_RESET_CMD_LDB_QID_WRITE      = 12'h040 ;
localparam      HQM_LSP_VF_RESET_CMD_DONE               = 12'h080 ;
localparam      HQM_LSP_VF_RESET_CMD_UNSUPPORTED        = 12'h100 ;

localparam      HQM_LSP_SMON0_WIDTH                     = 24 ;

localparam      HQM_QID_PER_CQ_2X			= ( HQM_QID_PER_CQ << 1 ) ;
localparam      HQM_LSP_NUM_LB_CQQIDIX_2X               = ( HQM_LSP_NUM_LB_CQQIDIX << 1 ) ;

//------------------------------------------------------------------------------------------------
// LBARB pipe structs, enums, params
typedef enum logic [2:0] {
    HQM_LSP_LBA_ARB_STATE_WAIT_FOR_WORK         = 3'b001
  , HQM_LSP_LBA_ARB_STATE_SCHED                 = 3'b010
  , HQM_LSP_LBA_ARB_STATE_WAIT_FOR_BLAST        = 3'b100
} lba_arb_state_t;

typedef struct packed {
  logic                                 sch_v ;
  logic                                 sch_nalb_v ;
  logic                                 sch_atm_v ;
  logic                                 sch_atm_rlist ;
  logic [15:0]                          sch_rlist_qidixv ;                      //JTC
  logic [15:0]                          sch_slist_qidixv ;                      //JTC
  logic [15:0]                          sch_nalb_qidixv ;                       //JTC
  logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]  sch_cq ;
  logic                                 sch_cq_p ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] sch_qid ;
  logic                                 sch_qidix_msb ;
  logic [2:0]                           sch_qidix ;
  logic [15:0]                          sch_cmpblast_qidixv ;                   //JTC
  logic                                 enq_v ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] enq_qid ;
  logic                                 enq_qid_p ;
  logic                                 tok_v ;
  logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]  tok_cq ;
  logic                                 tok_cq_p ;
  logic [10:0]                          tok_cnt ;
  logic [1:0]                           tok_cnt_res ;
  logic                                 cq_cmp_v ;
  logic                                 qid_cmp_v ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] cmp_qid ;
  logic                                 cmp_qid_p ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] cmp_qid_atm ;           // In case atm cmp paired with uno/rop "qid" completion (for different qid)
  logic                                 cmp_qid_atm_p ;
  logic                                 cmp_qid_no_dec ;
  logic                                 cmp_cq_no_dec ;
  logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]  cmp_cq ;
  logic                                 cmp_cq_p ;
  logic                                 cmp_qidix_msb ;
  logic [2:0]                           cmp_qidix ;
  logic [2:0]                           cmp_qpri ;
  logic                                 cmp_p ;
  logic [HQM_LSP_ARCH_NUM_FIDB2-1:0]    cmp_fid ;
  logic                                 cmp_fid_p ;
  logic [15:0]                          cmp_hid ;
  logic                                 cmp_hid_p ;
  logic                                 cmp_atm ;
  logic                                 qid_if_dec_v ;
} lba_ctrl_pipe_t ;

typedef struct packed {
  logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]  cq ;
  logic                                 slot_msb ;
  logic [2:0]                           slot ;
  logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] qid ;  
  logic                                 parity ;                // cq / total parity
  logic [1:0]                           cm_code ;
} lba_sch_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_cfg_cq2priov_t                            data_priov ;
  lsp_cfg_cq2qid_t                              data_qid_ms ;
  lsp_cfg_cq2qid_t                              data_qid_ls ;
} lba_cq2qid_rw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]     pcq ;           // paired cq
  lsp_cfg_cq2priov_t                            data_priov_odd ;
  lsp_cfg_cq2priov_t                            data_priov_even ;
  lsp_cfg_cq2qid_t                              data_qid_ms_odd ;
  lsp_cfg_cq2qid_t                              data_qid_ms_even ;
  lsp_cfg_cq2qid_t                              data_qid_ls_odd ;
  lsp_cfg_cq2qid_t                              data_qid_ls_even ;
} lba_cq2qid2x_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_lb_qid_enq_cnt_t                          data ;
} lba_qid_enq_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_lb_qid_dpth_thrsh_t                       data ;
} lba_qid_dpth_thrsh_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_lb_qid_if_cnt_t                           data ;
} lba_qid_if_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_lb_qid_if_lim_t                           data ;
} lba_qid_if_lim_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_lb_cq_tok_cnt_t                           data ;
} lba_cq_tok_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_lb_cq_tok_lim_t                           data ;
} lba_cq_tok_lim_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_lb_cq_if_cnt_t                            data ;
} lba_cq_if_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_lb_cq_if_lim_t                            data ;
} lba_cq_if_lim_rw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_lb_cq_if_thr_t                            data ;
} lba_cq_if_thr_rw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_cfg_qid2cqidix_t                          data ;
} lba_qid2cqidix_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_arch_cnt_t                                data ;
} lba_tot_enq_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]         cq ;
  lsp_arch_cnt_t                                data ;
} lba_tot_sch_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]      data ;
} lba_max_enq_depth_rmw_pipe_t ;

localparam      HQM_LSP_PRI_BIN_FACTOR                  = 0 ;   // Number of priority bits ignored
localparam      HQM_LSP_NUM_PRI_BINS                    = ( HQM_NUM_PRI >> HQM_LSP_PRI_BIN_FACTOR ) ;
localparam      HQM_LSP_NUM_PRI_BINSB2                  = AW_logb2 ( HQM_LSP_NUM_PRI_BINS - 1 ) + 1 ;

localparam      HQM_LSP_NUM_LDB_WRR_COUNT               = 8 ;
localparam      HQM_LSP_NUM_LDB_WRR_COUNTB2             = AW_logb2 ( HQM_LSP_NUM_LDB_WRR_COUNT - 1 ) + 1 ;

typedef struct packed {
  logic  [(HQM_QID_PER_CQ*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]     counts ;
  logic  [(HQM_LSP_NUM_PRI_BINS*HQM_QIDIX)-1:0]                 indexes ;
} lba_ldb_arb_index_t ;

typedef struct packed {
  logic  [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]     counts ;
  logic  [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]                  indexes ;
} lba_ldb_arb_index_pcm_t ;

typedef struct packed {
  logic  [(HQM_QID_PER_CQ*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]     counts_odd ;
  logic  [(HQM_LSP_NUM_PRI_BINS*HQM_QIDIX)-1:0]                 indexes_odd ;
  logic  [(HQM_QID_PER_CQ*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]     counts_even ;
  logic  [(HQM_LSP_NUM_PRI_BINS*HQM_QIDIX)-1:0]                 indexes_even ;
} lba_ldb_arb_index2x_t ;


localparam      HQM_LSP_AP_LSP_CMD_CMP                  = 2'h0 ;
localparam      HQM_LSP_AP_LSP_CMD_SCH_RLIST            = 2'h1 ;
localparam      HQM_LSP_AP_LSP_CMD_SCH_SLIST            = 2'h2 ;

localparam      HQM_LSP_LB_QID_ENQ_CNT_MEM_WIDTH        = $bits( lsp_lb_qid_enq_cnt_t ) ;
localparam      HQM_LSP_LB_QID_DPTH_THRSH_MEM_WIDTH     = $bits( lsp_lb_qid_dpth_thrsh_t ) ;
localparam      HQM_LSP_LB_QID_IF_CNT_MEM_WIDTH         = $bits( lsp_lb_qid_if_cnt_t ) ;
localparam      HQM_LSP_LB_QID_IF_LIM_MEM_WIDTH         = $bits( lsp_lb_qid_if_lim_t ) ;
localparam      HQM_LSP_LB_CQ_TOK_CNT_MEM_WIDTH         = $bits( lsp_lb_cq_tok_cnt_t ) ;
localparam      HQM_LSP_LB_CQ_TOK_LIM_SEL_MEM_WIDTH     = $bits( lsp_lb_cq_tok_lim_t ) ;
localparam      HQM_LSP_LB_CQ_IF_CNT_MEM_WIDTH          = $bits( lsp_lb_cq_if_cnt_t ) ;
localparam      HQM_LSP_LB_CQ_IF_LIM_MEM_WIDTH          = $bits( lsp_lb_cq_if_lim_t ) ;
localparam      HQM_LSP_LB_CQ_IF_THR_MEM_WIDTH          = $bits( lsp_lb_cq_if_thr_t ) ;
localparam      HQM_LSP_LB_CQ2PRIOV_MEM_WIDTH           = $bits( lsp_cfg_cq2priov_t ) ;
localparam      HQM_LSP_LB_CQ2QID_MEM_WIDTH             = $bits( lsp_cfg_cq2qid_t ) ;
localparam      HQM_LSP_LB_QID2CQIDIX_MEM_WIDTH         = $bits( lsp_cfg_qid2cqidix_t ) ;
localparam      HQM_LSP_LB_ARBINDEX_MEM_WIDTH           = $bits( lba_ldb_arb_index2x_t ) ;

localparam      HQM_LSP_LBA_CQ_ARB_ATM                  = 1'b0 ;
localparam      HQM_LSP_LBA_CQ_ARB_NALB                 = 1'b1 ;
localparam      HQM_LSP_LBA_QID_ARB_ORD                 = 1'b0 ;
localparam      HQM_LSP_LBA_QID_ARB_UNO_ATM             = 1'b1 ;
localparam      HQM_LSP_LBA_EC_ARB_CMP                  = 1'b0 ;
localparam      HQM_LSP_LBA_EC_ARB_ENQ                  = 1'b1 ;

localparam      HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR         = 6 ;

//------------------------------------------------------------------------------------------------
// ATQ pipe structs, enums, params

typedef struct packed {
  logic                                 sch_v ;
  logic                                 sch_qid_p ;
  logic                                 enq_v ;
  logic                                 enq_qid_p ;
  logic                                 cmp_v ;
  logic                                 cmp_qid_p ;
  logic                                 blast_enq ;
  logic                                 blast_cmp ;
} atq_ctrl_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_atq_enq_cnt_t                             data ;
} atq_enq_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_atq_atm_active_t                          data ;
} atq_atm_active_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_atq_qid_dpth_thrsh_t                      data ;
} atq_qid_dpth_thrsh_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_atq_aqed_act_cnt_t                        data ;
} atq_aqed_act_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_atq_aqed_act_lim_t                        data ;
} atq_aqed_act_lim_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_arch_cnt_t                                data ;
} atq_tot_enq_cnt_rmw_pipe_t ;

localparam      HQM_LSP_ATQ_ENQ_CNT_MEM_WIDTH           = $bits( lsp_atq_enq_cnt_t ) ;
localparam      HQM_LSP_ATQ_ATM_ACTIVE_MEM_WIDTH        = $bits( lsp_atq_atm_active_t ) ;
localparam      HQM_LSP_ATQ_QID_DPTH_THRSH_MEM_WIDTH    = $bits( lsp_atq_qid_dpth_thrsh_t ) ;
localparam      HQM_LSP_ATQ_AQED_ACT_CNT_MEM_WIDTH      = $bits( lsp_atq_aqed_act_cnt_t ) ;
localparam      HQM_LSP_ATQ_AQED_ACT_LIM_MEM_WIDTH      = $bits( lsp_atq_aqed_act_lim_t ) ;

//------------------------------------------------------------------------------------------------
// DIRENQ pipe structs, enums, params

localparam      HQM_LSP_DIR_TOK_DELTA_WIDTH = 11 ;      // struct has ms unused bits

// Same as lsp_dp_sch_dir_t, with additional fields for num_beats/wbo on-the-fly calculation
typedef struct packed {
  logic [7:0]           cq ;                    // Same as lsp_dp_sch_dir
  logic [6:0]           qid ;                   // Same as lsp_dp_sch_dir
  logic [2:0]           qidix ;                 // Same as lsp_dp_sch_dir
  logic                 parity ;                // Same as lsp_dp_sch_dir
  hqm_core_flags_t      hqm_core_flags ;        // Same as lsp_dp_sch_dir
  logic                 fill_in_progress ;
  logic [2:0]           qid_v ;
  logic [2:0]           cq_avail ;
  logic [1:0]           wp ;
  logic                 disab_opt ;
} direnq_lsp_dp_sch_dir_t;

typedef struct packed {
  logic  [1:0]  cnt_res ;
  logic  [HQM_LSP_DIR_TOK_DELTA_WIDTH-1:0] cnt ;
} direnq_tok_delta_t ;

typedef struct packed {
  logic                                 sch_v ;
  logic                                 sch_qid_p ;
  logic [2:0]                           sch_beats ;
  logic                                 enq_v ;
  logic                                 enq_qid_p ;
  logic                                 tok_v ;
  logic                                 tok_cq_p ;
  direnq_tok_delta_t                    tok_delta ;
  logic                                 blast_enq ;
  logic                                 blast_tok ;
} direnq_ctrl_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]       qid ;
  lsp_direnq_enq_cnt_t                          data ;
} direnq_enq_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]       qid ;
  lsp_direnq_dpth_thrsh_t                       data ;
} direnq_dpth_thrsh_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]        cq ;
  lsp_direnq_tok_cnt_t                          data ; } direnq_tok_cnt_rmw_pipe_t ; 
typedef struct packed {
  aw_rwpipe_cmd_t                               rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]        cq ;
  lsp_direnq_tok_lim_t                          data ;
} direnq_tok_lim_rw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]       qid ;
  lsp_arch_cnt_t                                data ;
} direnq_tot_enq_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]        cq ;
  lsp_arch_cnt_t                                data ;
} direnq_tot_sch_cnt_rmw_pipe_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]        qid ;
  logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]      data ;
} direnq_max_enq_depth_rmw_pipe_t ;

typedef struct packed {
  logic [2:0]   cq_avail ;              // 0, 1, 2, 3 or >= 4
  logic [2:0]   qid_v ;                 // 0, 1, 2, 3 or >= 4
} direnq_arb_stat_t ;

localparam      HQM_LSP_DIRENQ_ENQ_CNT_MEM_WIDTH        = $bits( lsp_direnq_enq_cnt_t ) ;
localparam      HQM_LSP_DIRENQ_DPTH_THRSH_MEM_WIDTH     = $bits( lsp_direnq_dpth_thrsh_t ) ;
localparam      HQM_LSP_DIRENQ_TOK_CNT_MEM_WIDTH        = $bits( lsp_direnq_tok_cnt_t ) ;
localparam      HQM_LSP_DIRENQ_TOK_LIM_MEM_WIDTH        = $bits( lsp_direnq_tok_lim_t ) ;

localparam      HQM_LSP_CFG_RST_PFMAX                   = 256 ;         // Deepest RAM no deeper than this
localparam      HQM_LSP_CFG_RST_PFMAXB2                 = ( AW_logb2(HQM_LSP_CFG_RST_PFMAX-1)+1);

//------------------------------------------------------------------------------------------------
// LBRPL pipe structs, enums, params

typedef struct packed {
  logic                                 enq_v ;
  logic                                 qid_p ;
  logic [1:0]                           frag_cnt_res ;
  logic [12:0]                          frag_cnt ;      // Max count = 4K
  logic                                 sch_v ;
  logic                                 blast_enq ;
} dirrpl_ctrl_pipe_t ;

typedef struct packed {
  logic                                 enq_v ;
  logic                                 qid_p ;
  logic [1:0]                           frag_cnt_res ;
  logic [14:0]                          frag_cnt ;      // Max count = 16K
  logic                                 sch_v ;
  logic                                 blast_enq ;
} lbrpl_ctrl_pipe_t ;

typedef struct packed {
  logic         qid_v ;
} rpl_arb_stat_t ;

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_lbrpl_enq_cnt_t                           data ;
} lbrpl_enq_cnt_rmw_pipe_t ;

localparam      HQM_LSP_LBRPL_ENQ_CNT_MEM_WIDTH = $bits( lsp_lbrpl_enq_cnt_t ) ;


//------------------------------------------------------------------------------------------------
// DIRRPL pipe structs, enums, params

typedef struct packed {
  aw_rmwpipe_cmd_t                              rw_cmd ;
  logic  [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]        qid ;
  lsp_dirrpl_enq_cnt_t                          data ;
} dirrpl_enq_cnt_rmw_pipe_t ;

localparam      HQM_LSP_DIRRPL_ENQ_CNT_MEM_WIDTH        = $bits( lsp_dirrpl_enq_cnt_t ) ;

//------------------------------------------------------------------------------------------------
// PALB (Power Aware Load Balancing) Interface declarations 

logic [ HQM_NUM_LB_CQ - 1 : 0 ] core_chp_lsp_ldb_cq_off_f ;

//------------------------------------------------------------------------------------------------
// Interface declarations

logic                  disable_smon ;
assign disable_smon = 1'b0 ;

// chp_lsp_cmp
logic                           core_chp_lsp_cmp_v ;
logic                           core_chp_lsp_cmp_ready ;
chp_lsp_cmp_t                   core_chp_lsp_cmp_data ;
aw_fifo_status_t                chp_lsp_cmp_fifo_status_pnc ;

// qed_lsp_deq and aqed_lsp_deq are inside hqm_lsp_wu_pipe

// chp_lsp_token
logic                           core_chp_lsp_token_v ;
logic                           core_chp_lsp_token_ready ;
chp_lsp_token_t                 core_chp_lsp_token_data ;
aw_fifo_status_t                chp_lsp_token_fifo_status_pnc ;

// nalb_lsp_enq_lb
logic                           core_nalb_lsp_enq_lb_v ;
logic                           core_nalb_lsp_enq_lb_ready ;
nalb_lsp_enq_lb_t               core_nalb_lsp_enq_lb_data ;
aw_fifo_status_t                nalb_lsp_enq_lb_fifo_status_pnc ;

// nalb_lsp_enq_rorply
logic                           core_nalb_lsp_enq_rorply_v ;
logic                           core_nalb_lsp_enq_rorply_ready ;
nalb_lsp_enq_rorply_t           core_nalb_lsp_enq_rorply_data ;
aw_fifo_status_t                nalb_lsp_enq_rorply_fifo_status_pnc ;

// dp_lsp_enq_dir
logic                           core_dp_lsp_enq_dir_v ;
logic                           core_dp_lsp_enq_dir_ready ;
dp_lsp_enq_dir_t                core_dp_lsp_enq_dir_data ;
aw_fifo_status_t                dp_lsp_enq_dir_fifo_status_pnc ;

// dp_lsp_enq_rorply
logic                           core_dp_lsp_enq_rorply_v ;
logic                           core_dp_lsp_enq_rorply_ready ;
dp_lsp_enq_rorply_t             core_dp_lsp_enq_rorply_data ;
aw_fifo_status_t                dp_lsp_enq_rorply_fifo_status_pnc ;

// rop_lsp_reordercmp
logic                           core_rop_lsp_reordercmp_v ;
logic                           core_rop_lsp_reordercmp_ready ;
rop_lsp_reordercmp_t            core_rop_lsp_reordercmp_data ;
aw_fifo_status_t                rop_lsp_reordercmp_fifo_status_pnc ;

// aqed_lsp_sch
logic                           send_atm_to_cq_v ;
logic                           send_atm_to_cq_ready ;
aqed_lsp_sch_t                  send_atm_to_cq_data ;
aw_fifo_status_t                send_atm_to_cq_fifo_status_pnc ;

//------------------------------------------------------------------------------------------------
// Input buffering declarations
logic                                           dir_tokrtn_fifo_push ;
logic                                           dir_tokrtn_fifo_pop ;
chp_lsp_token_t                                 dir_tokrtn_fifo_push_data ;
chp_lsp_token_t                                 dir_tokrtn_fifo_pop_data ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]           dir_tokrtn_fifo_pop_data_cq ;
logic                                           dir_tokrtn_fifo_pop_data_v ;
logic                                           dir_tokrtn_fifo_pop_data_vreq ;
logic [1:0]                                     dir_tokrtn_fifo_pop_data_count_ms_nc ;
logic                                           dir_tokrtn_fifo_afull ;
logic                                           dir_tokrtn_fifo_empty ;
logic                                           dir_tokrtn_fifo_pop_data_cq_p ;
//                      Actually a DB
logic [6:0]                                     dir_tokrtn_db_status_pnc ;
logic                                           dir_tokrtn_db_in_ready ;
logic                                           dir_tokrtn_db_out_valid ;

//------------------------------------------------------------------------------------------------
logic                                           ldb_token_rtn_fifo_push ;
logic                                           ldb_token_rtn_fifo_pop ;
lsp_ldb_token_rtn_t                             ldb_token_rtn_fifo_push_data ;
lsp_ldb_token_rtn_t                             ldb_token_rtn_fifo_pop_data ;
logic                                           ldb_token_rtn_fifo_pop_data_v ;
logic                                           ldb_token_rtn_fifo_pop_data_vreq ;
logic [1:0]                                     ldb_token_rtn_fifo_pop_data_nc ;
logic                                           ldb_token_rtn_fifo_afull ;
logic                                           ldb_token_rtn_fifo_full_nc ;
logic                                           ldb_token_rtn_fifo_empty ;
logic                                           ldb_token_rtn_fifo_of ;
logic                                           ldb_token_rtn_fifo_uf ;
logic [HQM_LSP_LDB_TOKEN_RTN_FIFO_WMWIDTH-1:0]  ldb_token_rtn_fifo_hwm ;
logic [31:0]                                    ldb_token_rtn_fifo_status_pnc ;

//------------------------------------------------------------------------------------------------
logic                                           uno_atm_cmp_fifo_push ;
logic                                           uno_atm_cmp_fifo_pop ;
lsp_uno_atm_cmp_t                               uno_atm_cmp_fifo_push_data ;
lsp_uno_atm_cmp_t                               uno_atm_cmp_fifo_pop_data ;
logic                                           uno_atm_cmp_fifo_pop_data_v ;
logic                                           uno_atm_cmp_fifo_pop_data_vreq ;
logic                                           uno_atm_cmp_fifo_pop_data_qid_p ;
logic [1:0]                                     uno_atm_cmp_fifo_pop_data_nc ;
logic                                           uno_atm_cmp_fifo_afull ;
logic                                           uno_atm_cmp_fifo_full_nc ;
logic                                           uno_atm_cmp_fifo_empty ;
logic                                           uno_atm_cmp_fifo_of ;
logic                                           uno_atm_cmp_fifo_uf ;
logic [HQM_LSP_UNO_ATM_CMP_FIFO_WMWIDTH-1:0]    uno_atm_cmp_fifo_hwm ;
logic [31:0]                                    uno_atm_cmp_fifo_status_pnc ;
logic                                           core_chp_lsp_cmp_atm_v ;
logic                                           core_chp_lsp_cmp_uno_v ;
logic                                           core_chp_lsp_cmp_nalb_v ;
logic                                           core_chp_lsp_cmp_rel_v ;
logic                                           uno_atm_cmp_fifo_ready ;
logic                                           atm_cmp_fifo_ready ;
logic                                           nalb_cmp_fifo_ready ;

//------------------------------------------------------------------------------------------------
logic                                           nalb_cmp_fifo_push ;
logic                                           nalb_cmp_fifo_pop ;
lsp_nalb_cmp_t                                  nalb_cmp_fifo_push_data ;
lsp_nalb_cmp_t                                  nalb_cmp_fifo_pop_data ;
logic                                           nalb_cmp_fifo_pop_data_v ;
logic                                           nalb_cmp_fifo_pop_data_vreq ;
logic                                           nalb_cmp_fifo_pop_data_cq_p ;
logic                                           nalb_cmp_fifo_pop_data_cq_wt_p ;
logic [1:0]                                     nalb_cmp_fifo_pop_data_cq_ms_nc ;
logic                                           nalb_cmp_fifo_afull ;
logic                                           nalb_cmp_fifo_full_nc ;
logic                                           nalb_cmp_fifo_empty ;
logic                                           nalb_cmp_fifo_of ;
logic                                           nalb_cmp_fifo_uf ;
logic [HQM_LSP_NALB_CMP_FIFO_WMWIDTH-1:0]       nalb_cmp_fifo_hwm ;
logic [31:0]                                    nalb_cmp_fifo_status_pnc ;

//------------------------------------------------------------------------------------------------
logic                                           core_chp_lsp_cmp_data_ap_p ;
logic                                           core_chp_lsp_cmp_data_cmp_p ;
logic                                           core_chp_lsp_cmp_data_fid_p ;
logic                                           core_chp_lsp_cmp_data_cq_qid_p ;

logic                                           atm_cmp_fifo_push ;
logic                                           atm_cmp_fifo_pop ;
lsp_atm_cmp_t                                   atm_cmp_fifo_push_data ;
lsp_atm_cmp_t                                   atm_cmp_fifo_pop_data ;
logic                                           atm_cmp_fifo_pop_data_v ;
logic                                           atm_cmp_fifo_pop_data_vreq ;
logic                                           atm_cmp_fifo_afull ;
logic                                           atm_cmp_fifo_full_nc ;
logic                                           atm_cmp_fifo_empty ;
logic                                           atm_cmp_fifo_of ;
logic                                           atm_cmp_fifo_uf ;
logic [HQM_LSP_ATM_CMP_FIFO_WMWIDTH-1:0]        atm_cmp_fifo_hwm ;
logic [31:0]                                    atm_cmp_fifo_status_pnc ;

logic                                           atm_cmp_fifo_pop_data_cq_p ;
logic                                           atm_cmp_fifo_pop_data_qid_p ;
logic                                           atm_cmp_fifo_pop_data_cq_wt_p ;

logic                                           atm_cmp_fifo_single_op_hold ;
logic                                           atm_cmp_wait_for_ap_cmp_nxt ;
logic                                           atm_cmp_wait_for_ap_cmp_f ;

//------------------------------------------------------------------------------------------------
logic                                           rop_lsp_reordercmp_fifo_pop ;
rop_lsp_reordercmp_t                            rop_lsp_reordercmp_fifo_pop_data ;
logic                                           rop_lsp_reordercmp_fifo_pop_data_vreq ;
logic                                           rop_lsp_reordercmp_fifo_pop_data_qid_p ;

//------------------------------------------------------------------------------------------------
logic                                           enq_nalb_fifo_push ;
logic                                           enq_nalb_fifo_pop ;
nalb_lsp_enq_lb_t                               enq_nalb_fifo_push_data ;
nalb_lsp_enq_lb_t                               enq_nalb_fifo_pop_data ;
logic                                           enq_nalb_fifo_pop_data_v ;
logic                                           enq_nalb_fifo_pop_data_vreq ;
logic                                           enq_nalb_fifo_afull ;
logic                                           enq_nalb_fifo_full_nc ;
logic                                           enq_nalb_fifo_empty ;
logic                                           enq_nalb_fifo_of ;
logic                                           enq_nalb_fifo_uf ;
logic [HQM_LSP_ENQ_NALB_FIFO_WMWIDTH-1:0]       enq_nalb_fifo_hwm ;
logic [31:0]                                    enq_nalb_fifo_status_pnc ;

//------------------------------------------------------------------------------------------------
logic                                           nalbrpl_fifo_pop ;
logic                                           nalbrpl_fifo_pop_data_v ;
logic                                           nalbrpl_fifo_pop_data_vreq ;
nalb_lsp_enq_rorply_t                           nalbrpl_fifo_pop_data  ;
//------------------------------------------------------------------------------------------------
logic                                           dp_lsp_enq_dir_fifo_pop ;
dp_lsp_enq_dir_t                                dp_lsp_enq_dir_fifo_pop_data ;
logic                                           dp_lsp_enq_dir_fifo_pop_data_v ;
logic                                           dp_lsp_enq_dir_fifo_pop_data_vreq ;

//------------------------------------------------------------------------------------------------
logic                                           dirrpl_fifo_pop ;
logic                                           dirrpl_fifo_pop_data_v ;
logic                                           dirrpl_fifo_pop_data_vreq ;
dp_lsp_enq_rorply_t                             dirrpl_fifo_pop_data  ;
//------------------------------------------------------------------------------------------------
logic                                           send_atm_to_cq_fifo_pop ;
logic                                           send_atm_to_cq_fifo_pop_data_v ;
logic                                           send_atm_to_cq_fifo_pop_data_vreq ;
aqed_lsp_sch_t                                  send_atm_to_cq_fifo_pop_data  ;
logic                                           send_atm_to_cq_fifo_pop_data_qid_p  ;
logic [15:0]                                    send_atm_to_cq_fifo_pop_data_flid_nc ;

//------------------------------------------------------------------------------------------------
// Internal buffering declarations
logic [6:0]                                     enq_atq_db_status_pnc ;
logic                                           enq_atq_db_in_ready ;
logic                                           enq_atq_db_in_valid ;
nalb_lsp_enq_lb_t                               enq_atq_db_in_data ;
logic                                           enq_atq_db_out_ready ;
logic                                           enq_atq_db_out_valid ;
nalb_lsp_enq_lb_t                               enq_atq_db_out_data ;

logic                                           enq_atq_fifo_pop_data_v ;
logic                                           enq_atq_fifo_pop_data_vreq ;
logic                                           enq_atq_fifo_pop ;
nalb_lsp_enq_lb_t                               enq_atq_fifo_pop_data ;
logic                                           enq_atq_fifo_pop_data_qid_p ;

//------------------------------------------------------------------------------------------------
// Output buffering declarations
logic                                           dir_sel_dp_fifo_push ;
direnq_lsp_dp_sch_dir_t                         dir_sel_dp_fifo_push_data ;
logic                                           dir_sel_dp_fifo_afull ;
logic                                           dir_sel_dp_fifo_empty ;
logic                                           dir_sel_dp_fifo_hold ;


direnq_lsp_dp_sch_dir_t                         lsp_dp_sch_dir_pre_data ;
logic [1:0]                                     lsp_dp_sch_dir_data_write_buffer_optimization ;

logic                                           dir_sel_dp_db_in_valid ;
direnq_lsp_dp_sch_dir_t                         dir_sel_dp_db_in_data ;
logic                                           dir_sel_dp_db_in_ready ;
logic [6:0]                                     dir_sel_dp_db_status_nc ;

//------------------------------------------------------------------------------------------------
// Config / Alarm /sidecar declarations


logic                                           cfg_idle ;

logic   [ ( $bits(lsp_alarm_down_data.unit) -1 ) : 0]   lsp_uid ;

logic   [ ( HQM_LSP_ALARM_NUM_INF ) -1 : 0]             int_inf_v ;
aw_alarm_syn_t [ ( HQM_LSP_ALARM_NUM_INF ) -1 : 0]      int_inf_data ;
logic   [ ( HQM_LSP_ALARM_NUM_COR) -1 : 0]              int_cor_v ;
aw_alarm_syn_t [ ( HQM_LSP_ALARM_NUM_COR) -1 : 0]       int_cor_data ;
logic   [ ( HQM_LSP_ALARM_NUM_UNC ) -1 : 0]             int_unc_v ;
aw_alarm_syn_t [ ( HQM_LSP_ALARM_NUM_UNC ) -1 : 0]      int_unc_data ;
logic   [ ( 32 ) -1 : 0]                                int_serializer_status_pnc ;
logic [2:0]                                             int_serializer_status_up ;
logic [2:0]                                             int_serializer_status_down ;
logic                                                   int_idle ;
logic [30:0]                                            err_hw_class_01 ;
logic                                                   err_hw_class_01_v ;
logic [30:0]                                            err_hw_class_02 ;
logic                                                   err_hw_class_02_v ;
logic [30:0]                                            err_hw_class_03 ;
logic                                                   err_hw_class_03_v ;
logic [30:0]                                            err_hw_class_04 ;
logic                                                   err_hw_class_04_v ;
logic [30:0]                                            err_hw_class_05 ;
logic                                                   err_hw_class_05_v ;


// Note: Since the LB and DIR pipes share the token return FIFO, there is nothing to be gained by trying
// to keep the dir pipe alive while doing a LB config access, etc.  The only truly-independent pipes are
// the two replay pipes, and it is not worth the complexity/risk to try to optimize just them.
// cause_pipe_idle needs to prevent new upstream requests from being processed, and needs to prevent
// LSP from generating any new traffic (schedules).
logic                                                   cause_pipe_idle ;

logic [31:0]                                            cfg_control_general_0_nxt ;
logic [31:0]                                            cfg_control_general_0_f ;
logic                                                   cfg_control_disable_atq_empty_arb ;
logic                                                   cfg_control_include_tok_unit_idle ;
logic                                                   cfg_control_disable_rlist_pri ;
logic                                                   cfg_control_include_cmp_unit_idle ;
logic                                                   cfg_control_enable_inflight_thresh ;
logic                                                   cfg_control_single_op_direnq ;
logic                                                   cfg_control_half_bw_direnq ;
logic                                                   cfg_control_single_out_direnq ;
logic                                                   cfg_control_disable_multi_op_direnq ;
logic                                                   cfg_control_single_op_atq ;
logic                                                   cfg_control_half_bw_atq ;
logic                                                   cfg_control_single_out_atq ;
logic                                                   cfg_control_disable_multi_op_atq ;
logic                                                   cfg_control_single_op_dirrpl ;
logic                                                   cfg_control_half_bw_dirrpl ;
logic                                                   cfg_control_single_out_dirrpl ;
logic                                                   cfg_control_single_op_lbrpl ;
logic                                                   cfg_control_half_bw_lbrpl ;
logic                                                   cfg_control_single_out_lbrpl ;
logic                                                   cfg_control_single_op_lba ;
logic                                                   cfg_control_half_bw_lba ;
logic                                                   cfg_control_disable_multi_op_lba ;
logic                                                   cfg_control_single_op_atm_sched ;
logic                                                   cfg_control_single_op_atm_cmp ;
logic                                                   cfg_control_ldb_ce_tog_arb ;
logic [1:0]                                             cfg_smon0_v_sel ;
logic                                                   cfg_smon0_value_sel ;
logic [1:0]                                             cfg_smon0_comp_sel ;

logic [31:0]                                            cfg_control_general_1_nxt ;
logic [31:0]                                            cfg_control_general_1_f ;
logic [1:0]                                             cfg_control_qe_wt_frc_val ;
logic                                                   cfg_control_qe_wt_frc_v ;
logic                                                   cfg_control_qe_wt_blk ;
logic [4:0]                                             cfg_control_qed_lsp_deq_high_pri_wm ;
logic [4:0]                                             cfg_control_aqed_lsp_deq_high_pri_wm ;
logic                                                   cfg_control_disable_wu_res_chk ;

logic                                                   direnq_upipe_idle_nxt ;
logic                                                   direnq_upipe_idle_f ;
logic                                                   atq_upipe_idle_nxt ;
logic                                                   atq_upipe_idle_f ;
logic                                                   dirrpl_upipe_idle_nxt ;
logic                                                   dirrpl_upipe_idle_f ;
logic                                                   lbrpl_upipe_idle_nxt ;
logic                                                   lbrpl_upipe_idle_f ;
logic                                                   lba_pipe_idle_nxt ;
logic                                                   lba_pipe_idle_f ;


logic [31:0]                                            cfg_control_pipeline_credits_nxt ;
logic [31:0]                                            cfg_control_pipeline_credits_f ;
logic [7:0]                                             cfg_lba_pipeline_credit_limit ;
logic [7:0]                                             cfg_atm_pipeline_credit_limit ;
logic [7:0]                                             cfg_qed_deq_pipeline_credit_limit_pnc ;
logic [7:0]                                             cfg_aqed_deq_pipeline_credit_limit_pnc ;

logic [HQM_NUM_LB_CQ-1:0]                               cfg_cq_ldb_disable_f ;
logic [HQM_NUM_LB_CQ-1:0]                               cfg_cq_ldb_enable_pcm_f ;

logic                                                   p2_lba_inp_tok_cq_disable ;
logic                                                   p3_lba_cq2qid_cq_disable ;
logic                                                   p3_lba_cq2qid_cq_disable_odd ;
logic                                                   p3_lba_cq2qid_cq_disable_even ;
logic                                                   p3_lba_cq2qid_cq_disable_x ;
logic                                                   p7_lba_if_cnt_cq_disable ;
logic                                                   p7_lba_tok_cnt_cq_disable ;

logic [HQM_NUM_DIR_CQ-1:0]                              cfg_cq_dir_disable_nxt ;
logic [HQM_NUM_DIR_CQ-1:0]                              cfg_cq_dir_disable_f ;

logic                                                   p0_direnq_inp_tok_cq_disable ;
logic                                                   p2_direnq_enq_cnt_cq_disable ;
logic                                                   p2_direnq_tok_cnt_cq_disable ;

logic [31:0]                                            cfg_lsp_csr_control_nxt ;
logic [31:0]                                            cfg_lsp_csr_control_f ;
logic                                                   cfg_control_disable_tok_uflow_interrupt ;
logic                                                   cfg_control_disable_tok_uflow_synd_load ;
logic                                                   cfg_control_disable_cq_if_uflow_interrupt ;
logic                                                   cfg_control_disable_cq_if_uflow_synd_load ;
logic                                                   cfg_control_disable_hwerr_interrupt ;
logic                                                   cfg_control_disable_hwerr_synd_load ;
logic                                                   cfg_control_disable_qid_if_uflow_interrupt ;
logic                                                   cfg_control_disable_qid_if_uflow_synd_load ;
logic                                                   cfg_control_disable_non_mc_interrupt ;
logic                                                   cfg_control_disable_non_mc_synd_load ;
logic [HQM_LSP_NUM_LDB_WRR_COUNTB2-1:0]                 cfg_control_ldb_wrr_count_base ;
logic                                                   cfg_control_atm_cq_qid_priority_prot ;

logic [31:0]                                            cfg_ldb_sched_control_nxt ;
logic [31:0]                                            cfg_ldb_sched_control_f_pnc ;
logic [5:0]                                             cfg_ldb_sched_control_cq ;
logic [2:0]                                             cfg_ldb_sched_control_qidix ;
logic                                                   cfg_ldb_sched_control_value ;
logic                                                   cfg_ldb_sched_control_nalb_haswork_v ;
logic                                                   cfg_ldb_sched_control_rlist_haswork_v ;
logic                                                   cfg_ldb_sched_control_slist_haswork_v ;
logic                                                   cfg_ldb_sched_control_inflight_ok_v ;
logic                                                   cfg_ldb_sched_control_aqed_nfull_v ;
logic [8:0]                                             cfg_ldb_sched_control_cq_qidix ;
logic [6:0]                                             cfg_ldb_sched_control_qid ;

logic [31:0]                                            cfg_arb_weight_ldb_qid_0_nxt ;
logic [31:0]                                            cfg_arb_weight_ldb_qid_0_f ;
logic [31:0]                                            cfg_arb_weight_ldb_qid_1_nxt ;
logic [31:0]                                            cfg_arb_weight_ldb_qid_1_f ;

logic [31:0]                                            cfg_arb_weight_atm_nalb_qid_0_nxt ;
logic [31:0]                                            cfg_arb_weight_atm_nalb_qid_0_f ;
logic [31:0]                                            cfg_arb_weight_atm_nalb_qid_1_nxt ;
logic [31:0]                                            cfg_arb_weight_atm_nalb_qid_1_f ;

logic [31:0]                                            cfg_arb_weight_ldb_issue_0_nxt ;
logic [31:0]                                            cfg_arb_weight_ldb_issue_0_f ;

logic                                                   cfg_qid_atq_sch_v_nxt ;
logic                                                   cfg_qid_dir_replay_v_nxt ;
logic                                                   cfg_qid_ldb_replay_v_nxt ;
logic                                                   cfg_qid_atq_sch_v_f ;
logic                                                   cfg_qid_dir_replay_v_f ;
logic                                                   cfg_qid_ldb_replay_v_f ;

logic [31:0]                                            cfg_detect_feature_0_set ;
logic [31:0]                                            cfg_detect_feature_0_nxt ;
logic [31:0]                                            cfg_detect_feature_0_f ;
logic [31:0]                                            cfg_detect_feature_1_set ;
logic [31:0]                                            cfg_detect_feature_1_nxt ;
logic [31:0]                                            cfg_detect_feature_1_f ;


logic [31:0]                                            cfg_agitate_control_nxt ;
logic [31:0]                                            cfg_agitate_control_f ;
logic [31:0]                                            cfg_agitate_select_nxt ;
logic [31:0]                                            cfg_agitate_select_f ;

logic                                                   cfg_lbwu_pipe_idle ;

idle_status_t                                           cfg_unit_idle_nxt ;
idle_status_t                                           cfg_unit_idle_f ;

logic                                                   cfg_lba_cq_arb_reqs_nxt ;
logic                                                   cfg_lba_cq_arb_reqs_f ;
logic                                                   cfg_direnq_arb_reqs_nxt ;
logic                                                   cfg_direnq_arb_reqs_f ;
logic                                                   cfg_atq_arb_winner_v_nxt ;
logic                                                   cfg_atq_arb_winner_v_f ;

// Replicated to reduce fanout
idle_status_t                                           cfg_unit_idle_1_f_pnc ;         // Selected bits used to decrease transitive fanout
idle_status_t                                           cfg_unit_idle_2_f_pnc ;         // Selected bits used to decrease transitive fanout

logic [31:0]                                            cfg_error_inject_nxt ;
logic [31:0]                                            cfg_error_inject_f ;

logic                                                   cfg_ldb_sched_perf_cq_disabled ;
logic                                                   cfg_ldb_sched_perf_no_work ;
logic                                                   cfg_ldb_sched_perf_no_space ;
logic                                                   cfg_ldb_sched_perf_sched ;
logic                                                   cfg_ldb_sched_perf_pipe_frict_not_wait_work ;
logic                                                   cfg_ldb_sched_perf_pipe_frict_wait_work_hold ;
logic                                                   cfg_ldb_sched_perf_wait_blast ;
logic                                                   cfg_ldb_sched_perf_pipe_frict_cause_pipe_idle ;
logic                                                   cfg_ldb_sched_perf_3_inc ;
logic                                                   cfg_ldb_sched_perf_wait_tot_inflight ;
logic                                                   cfg_ldb_sched_perf_wait_cq_busy ;
logic                                                   cfg_ldb_sched_perf_wait_atq_fid_unavail ;
logic                                                   cfg_ldb_sched_perf_overworked ;

logic [31:0]                            cfg_pipe_health_hold_0_nxt ;
logic [31:0]                            cfg_pipe_health_hold_1_nxt ;

logic [31:0]                            cfg_pipe_health_valid_0_nxt ;
logic [31:0]                            cfg_pipe_health_valid_1_nxt ;

logic                                   cfg_syndrome0_capture_v ;
logic [30:0]                            cfg_syndrome0_capture_data ;
logic                                   cfg_syndrome1_capture_v ;
logic [30:0]                            cfg_syndrome1_capture_data ;

logic [31:0]                            cfg_diag_status_0_nxt ;
logic [31:0]                            cfg_diag_status_0_f ;

logic                                   cfg_lba_rlist_v ;
logic                                   cfg_lba_rlist_blast ;
logic                                   cfg_lba_slist_v ;
logic                                   cfg_lba_slist_blast ;
logic                                   cfg_lba_nalb_v ;
logic                                   cfg_lba_nalb_blast ;
logic                                   cfg_lba_cmpblast_chkv ;
logic                                   cfg_lba_cmpblast ;
logic                                   cfg_atq_qid_dis ;
logic                                   cfg_lba_cq_busy ;
logic                                   cfg_lba_cq_no_space ;
logic                                   cfg_direnq_tok_cnt_v ;
logic                                   cfg_atq_aqed_act_v ;
logic                                   cfg_lba_atm_haswork ;
logic                                   cfg_lba_cq_tok_cnt_v ;
logic                                   cfg_lba_cq_if_cnt_v ;
logic                                   cfg_lba_atm_if_v ;
logic                                   cfg_lba_ow_any ;

logic [31:0]                            cfg_diag_status_2_nxt ;
logic [31:0]                            cfg_diag_status_2_f ;                                   // For non-synth checking code only
logic                                   cfg_diag_status_2_allow_load ;

logic [31:0]                            cfg_diag_status_4_nxt ;
logic [31:0]                            cfg_diag_status_4_f_nc ;                                // For non-synth checking code only

logic                                   p0_lba_cmpblast_ap_val_nxt ;
logic                                   p0_lba_cmpblast_ap_val_f ;
logic                                   p0_lba_cmpblast_ap_rst_v_nxt ;
logic                                   p0_lba_cmpblast_ap_rst_v_f ;
logic                                   p0_lba_cmpblast_lsp_set_v_nxt ;
logic                                   p0_lba_cmpblast_lsp_set_v_f ;
logic                                   p0_lba_cmpblast_lsp_val_nxt ;
logic                                   p0_lba_cmpblast_lsp_val_f ;
logic                                   p0_lba_cmpblast_ap_rst_err ;
logic                                   p0_lba_cmpblast_lsp_set_err ;

logic [HQM_NUM_DIR_QID-1:0]             p3_qid_dir_sch_v_status ;
logic [HQM_NUM_DIR_CQ-1:0]              p3_cq_dir_tok_v_status ;

logic [511:0]                           cfg_qid_ldb_if_v_status ;
logic [511:0]                           cfg_qid_ldb_sch_v_status ;

logic [HQM_NUM_LB_CQ-1:0]               cfg_cq_ldb_if_v_status ;
logic [HQM_NUM_LB_CQ-1:0]               cfg_cq_ldb_thr_v_status ;
logic [HQM_NUM_LB_CQ-1:0]               cfg_cq_ldb_tok_v_status ;

logic [HQM_NUM_LB_QID-1:0]              cfg_qid_atq_sch_v_status ;
logic [HQM_NUM_LB_QID-1:0]              cfg_qid_atq_aqed_avail_status ;
logic                                   cfg_qid_atq_aqed_empty ;

logic [HQM_NUM_LB_QID-1:0]              cfg_qid_dir_replay_v_status ;
logic [HQM_NUM_LB_QID-1:0]              cfg_qid_ldb_replay_v_status ;

//------------------------------------------------------------------------------------------------
// LBARB pipe declarations

logic [HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR-1:0]     p0_lba_pop_cq ;
logic                                           p1_lba_issue_sched_cond ;
logic                                           p1_lba_issue_sched ;
lba_arb_state_t                                 p0_lba_sch_state_nxt ;
lba_arb_state_t                                 p0_lba_sch_state_f ;
logic                                           p0_lba_sch_state_ready_for_work ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_slist_cq_v ;
logic [511:0]                           p0_lba_slist_v_nxt ;
logic [511:0]                           p0_lba_slist_v_f ;
logic [511:0]                           p0_lba_slist_blast_nxt ;
logic [511:0]                           p0_lba_slist_blast_f ;
logic [511:0]                           p0_lba_slist_v_blasted ;
logic [511:0]                           p1_lba_sch_slist_v_nxt ;
logic [511:0]                           p1_lba_sch_slist_v_f ;
logic [7:0]                             p1_lba_sch_slist_v_ar [HQM_NUM_LB_CQ-1:0] ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_has_space_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_has_space_f ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_busy_sch_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_busy_sch_f ;

logic [511:0]                           p0_lba_atm_if_v_nxt ;
logic [511:0]                           p0_lba_atm_if_v_f ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_rlist_cq_v ;
logic [511:0]                           p0_lba_rlist_v_nxt ;
logic [511:0]                           p0_lba_rlist_v_f ;
logic [511:0]                           p0_lba_rlist_blast_nxt ;
logic [511:0]                           p0_lba_rlist_blast_f ;
logic [511:0]                           p0_lba_rlist_v_blasted ;
logic [511:0]                           p1_lba_sch_rlist_v_nxt ;
logic [511:0]                           p1_lba_sch_rlist_v_f ;
logic [7:0]                             p1_lba_sch_rlist_v_ar [HQM_NUM_LB_CQ-1:0] ;

logic [511:0]                           p0_lba_cmpblast_nxt ;
logic [511:0]                           p0_lba_cmpblast_f ;
logic [511:0]                           p0_lba_cmpblast_chkv_nxt ;
logic [511:0]                           p0_lba_cmpblast_chkv_f ;

logic [511:0]                           p0_lba_nalb_v_nxt ;
logic [511:0]                           p0_lba_nalb_v_f ;
logic [511:0]                           p0_lba_nalb_blast_nxt ;
logic [511:0]                           p0_lba_nalb_blast_f ;
logic [511:0]                           p0_lba_nalb_v_blasted ;
logic [511:0]                           p1_lba_sch_nalb_v_nxt ;
logic [511:0]                           p1_lba_sch_nalb_v_f ;
logic [7:0]                             p1_lba_sch_nalb_v_ar [HQM_NUM_LB_CQ-1:0] ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_arb_slist_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_arb_rlist_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_arb_nalb_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_arb_any_has_work ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_arb_reqs ;
logic                                   p0_lba_cq_arb_update ;
logic [HQM_NUM_LB_CQB2-1:0]             p0_lba_cq_arb_winner ;
logic [HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR-1:0]     p0_lba_cq_arb_winner_pre_v ;
logic [HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR-1:0]     p0_lba_cq_arb_winner_v ;

//--------
// V2 cq_cos arbiter declarations
logic [31:0]                                    cfg_range_cos0_reg_nxt ;
logic [31:0]                                    cfg_range_cos0_reg_f ;
logic [31:0]                                    cfg_range_cos1_reg_nxt ;
logic [31:0]                                    cfg_range_cos1_reg_f ;
logic [31:0]                                    cfg_range_cos2_reg_nxt ;
logic [31:0]                                    cfg_range_cos2_reg_f ;
logic [31:0]                                    cfg_range_cos3_reg_nxt ;
logic [31:0]                                    cfg_range_cos3_reg_f ;
logic [8:0]                                     cfg_range_cos0_f ;
logic [8:0]                                     cfg_range_cos1_f ;
logic [8:0]                                     cfg_range_cos2_f ;
logic [8:0]                                     cfg_range_cos3_f ;
logic [15:0]                                    cfg_credit_sat_cos0_f ;
logic [15:0]                                    cfg_credit_sat_cos1_f ;
logic [15:0]                                    cfg_credit_sat_cos2_f ;
logic [15:0]                                    cfg_credit_sat_cos3_f ;
logic [15:0]                                    cfg_credit_cnt_cos0 ;
logic [15:0]                                    cfg_credit_cnt_cos1 ;
logic [15:0]                                    cfg_credit_cnt_cos2 ;
logic [15:0]                                    cfg_credit_cnt_cos3 ;
logic                                           cfg_no_extra_credit0_f ;
logic                                           cfg_no_extra_credit1_f ;
logic                                           cfg_no_extra_credit2_f ;
logic                                           cfg_no_extra_credit3_f ;
logic [10:0]                                    cfg_starv_avoid_cnt_cos0 ;
logic [10:0]                                    cfg_starv_avoid_cnt_cos1 ;
logic [10:0]                                    cfg_starv_avoid_cnt_cos2 ;
logic [10:0]                                    cfg_starv_avoid_cnt_cos3 ;
logic                                           cfg_starv_avoid_enable_f ;
logic [9:0]                                     cfg_starv_avoid_thresh_min_f ;
logic [9:0]                                     cfg_starv_avoid_thresh_max_f ;
logic                                           cfg_shdw_ctrl_load ;
logic [30:0]                                    cfg_shdw_ctrl_load_spare_nc ;
logic [3:0]                                     cfg_schd_cos ;
logic [3:0]                                     cfg_rdy_cos ;
logic [3:0]                                     cfg_rnd_loss_cos ;
logic [3:0]                                     cfg_cnt_win_cos ;
logic [63:0]                                    hqm_lsp_target_cfg_sch_rdy_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_schd_cos0_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_schd_cos1_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_schd_cos2_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_schd_cos3_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rdy_cos0_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rdy_cos1_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rdy_cos2_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rdy_cos3_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rnd_loss_cos0_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rnd_loss_cos1_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rnd_loss_cos2_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_rnd_loss_cos3_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_cnt_win_cos0_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_cnt_win_cos1_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_cnt_win_cos2_count_nc ;
logic [63:0]                                    hqm_lsp_target_cfg_cnt_win_cos3_count_nc ;
logic [31:0]                                    hqm_lsp_target_cfg_credit_cnt_cos0_nc ;
logic [31:0]                                    hqm_lsp_target_cfg_credit_cnt_cos1_nc ;
logic [31:0]                                    hqm_lsp_target_cfg_credit_cnt_cos2_nc ;
logic [31:0]                                    hqm_lsp_target_cfg_credit_cnt_cos3_nc ;
//--------

logic [511:0]                           p0_nxt_lba_slist_v_blasted_nc ;
logic [511:0]                           p0_nxt_lba_rlist_v_blasted_nc ;
logic [511:0]                           p0_nxt_lba_nalb_v_blasted_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_nxt_lba_cq_arb_slist_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_nxt_lba_cq_arb_rlist_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_nxt_lba_cq_arb_nalb_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_nxt_lba_cq_arb_any_has_work_nc ;
logic [HQM_NUM_LB_CQ-1:0]               p0_nxt_lba_cq_arb_reqs ;

logic                                   p0_lba_cq_arb_error_f ;
logic [3:0]                             p0_lba_cq_arb_status ;

logic                                   p0_lba_cq_gp ;
logic [15:0]                            p1_lba_sch_cmpblast_qidixv_nxt ;
logic [15:0]                            p1_lba_sch_cmpblast_qidixv_f ;

logic                                   p0_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p1_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p2_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p3_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p4_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p5_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p6_lba_ctrl_pipe_cmpblast_cond ;
logic                                   p7_lba_ctrl_pipe_cmpblast_cond ;

logic [15:0]                            p0_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p1_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p2_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p3_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p4_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p5_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p6_lba_sch_cmpblast_qidixv_blasted ;
logic [15:0]                            p7_lba_sch_cmpblast_qidixv_blasted ;

logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   lbi_inp_enq_qid ;
logic                                   lbi_inp_enq_qid_p ;
logic                                   lbi_enq_req_taken ;

logic [HQM_NUM_LB_CQB2-1:0]             lbi_inp_tok_cq ;
logic                                   lbi_inp_tok_cq_p ;
logic                                   lbi_inp_tok_cnt_uflow_cond ;
logic [10:0]                            lbi_inp_tok_cnt ;
logic [1:0]                             lbi_inp_tok_cnt_res ;

logic                                   lbi_tok_req_taken ;

logic                                   lbi_inp_cq_cmp_no_dec ;
logic [HQM_NUM_LB_CQB2-1:0]             lbi_inp_cq_cmp_cq ;
logic [1:0]                             lbi_inp_cq_cmp_qe_wt ;
logic                                   lbi_inp_cq_cmp_cq_wt_p ;
logic                                   lbi_inp_cq_cmp_cq_p ;
logic                                   lbi_cq_cmp_arb_atm_v ;
logic [1:0]                             lbi_cq_cmp_arb_reqs ;
logic                                   lbi_cq_cmp_arb_winner ;
logic                                   lbi_cq_cmp_arb_winner_v ;
logic                                   lbi_cq_cmp_req_taken ;
logic                                   p0_lba_supress_cq_cmp ;
logic [7:0]                             cfg_lbi_cq_cmp_arb_weight_atm ;
logic [7:0]                             cfg_lbi_cq_cmp_arb_weight_nalb ;


logic                                   lbi_inp_cmp_qidix_msb ;
logic [2:0]                             lbi_inp_cmp_qidix ;
logic [2:0]                             lbi_inp_cmp_qpri ;
logic [HQM_LSP_ARCH_NUM_FIDB2-1:0]      lbi_inp_cmp_fid ;
logic                                   lbi_inp_cmp_fid_p ;
logic [15:0]                            lbi_inp_cmp_hid ;
logic                                   lbi_inp_cmp_hid_p ;
logic                                   lbi_inp_cmp_p ;

logic                                   lbi_inp_qid_cmp_no_dec ;
logic                                   lbi_inp_qid_cmp_dec_only ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   lbi_inp_qid_cmp_qid ;
logic                                   lbi_inp_qid_cmp_qid_p ;
logic [1:0]                             lbi_qid_cmp_arb_reqs ;
logic                                   lbi_qid_cmp_arb_winner ;
logic                                   lbi_qid_cmp_arb_winner_v ;
logic                                   lbi_qid_cmp_req_taken ;
logic [7:0]                             cfg_lbi_qid_cmp_arb_weight_ord ;
logic [7:0]                             cfg_lbi_qid_cmp_arb_weight_uno_atm ;

logic [1:0]                             lbi_ec_arb_reqs ;
logic                                   lbi_ec_arb_strict_winner ;
logic                                   lbi_ec_arb_strict_winner_v ;
logic                                   lbi_ec_arb_tog_winner ;
logic                                   lbi_ec_arb_tog_winner_v ;
logic                                   lbi_ec_arb_winner ;
logic                                   lbi_ec_arb_winner_v ;
logic                                   lbi_ec_arb_enq_v ;
logic                                   lbi_ec_arb_cmp_v;       // include RELEASE
logic                                   lbi_ec_arb_update ;
logic                                   lbi_ec_arb_tie ;
logic                                   lbi_ec_arb_tie_broken ;
logic                                   lbi_ec_arb_tog_nxt ;
logic                                   lbi_ec_arb_tog_f ;

logic                                   p0_lba_atm_credit_count_inc ;
logic [4:0]                             p0_lba_atm_credit_count_nxt ;
logic [4:0]                             p0_lba_atm_credit_count_f ;
logic [4:0]                             p0_lba_atm_credit_count_px ;
logic [2:0]                             p0_lba_atm_credit_count_dec_amt ;
logic                                   p0_lba_atm_credit_count_eq_0 ;
logic                                   p4_lba_atm_credit_count_dec_miss ;

logic                                   p0_lba_nalb_credit_count_inc ;
logic                                   p0_lba_nalb_credit_count_dec_hit ;
logic [4:0]                             p0_lba_nalb_credit_count_nxt ;
logic [4:0]                             p0_lba_nalb_credit_count_f ;
logic [4:0]                             p0_lba_nalb_credit_count_p1 ;
logic [4:0]                             p0_lba_nalb_credit_count_m1 ;
logic [4:0]                             p0_lba_nalb_credit_count_m2 ;
logic                                   p0_lba_nalb_credit_count_eq_0 ;
logic                                   p4_lba_nalb_credit_count_dec_miss ;

logic                                   p0_lba_nalb_credit_hold_cond ;
logic                                   p0_lba_atm_credit_hold_cond ;
logic                                   p0_lba_ctrl_pipe_sch_hold_cond ;
logic                                   p0_lba_restrict_bw_hold_cond ;

logic                                   p0_lba_arb_winner_pre_v ;
logic                                   p0_lba_arb_winner_v ;

logic                                   p0_lba_arb_sch_v ;
logic                                   p0_lba_arb_pre_enq_v_cond ;
logic                                   p0_lba_arb_pre_enq_v ;
logic                                   p0_lba_arb_enq_v ;
logic                                   p0_lba_arb_pre_tok_v_cond ;
logic                                   p0_lba_arb_pre_tok_v ;
logic                                   p0_lba_arb_tok_v ;
logic                                   p0_lba_arb_pre_cq_cmp_v_cond ;
logic                                   p0_lba_arb_pre_cq_cmp_v ;
logic                                   p0_lba_arb_cq_cmp_v ;
logic                                   p0_lba_arb_pre_qid_cmp_v_cond ; // includes RELEASE
logic                                   p0_lba_arb_pre_qid_cmp_v ;      // includes RELEASE
logic                                   p0_lba_arb_qid_cmp_v ;          // includes RELEASE
logic                                   p0_lba_arb_cmp_atm_v ;
logic [3:0]                             p0_lba_mop_arb_reqs ;
logic                                   p0_lba_mop_arb_update ;
logic [1:0]                             p0_lba_mop_arb_winner ;
logic                                   p0_lba_mop_arb_winner_pre_v ;
logic                                   p0_lba_mop_arb_winner_v ;


lsp_pipe_ctrl_t                         p0_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p1_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p2_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p3_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p4_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p5_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p6_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p7_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p8_lba_ctrl_pipe ;
lsp_pipe_ctrl_t                         p9_lba_ctrl_pipe ;


logic                                   p1_lba_ctrl_pipe_v_nxt ;
logic                                   p1_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p1_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p1_lba_ctrl_pipe_f ;


logic                                   p2_lba_ctrl_pipe_v_nxt ;
logic                                   p2_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p2_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p2_lba_ctrl_pipe_f ;

logic                                   p3_lba_ctrl_pipe_v_nxt ;
logic                                   p3_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p3_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p3_lba_ctrl_pipe_f ;

logic                                   p4_lba_ctrl_pipe_v_nxt ;
logic                                   p4_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p4_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p4_lba_ctrl_pipe_f ;
logic                                   p4_from_p5_hold ;
logic                                   p4_lba_atm_sch_hold ;
logic                                   p4_lba_ctrl_pipe_cmp_p ;

logic                                   p5_lba_ctrl_pipe_v_nxt ;
logic                                   p5_lba_ctrl_pipe_v_nxt_gated ;
logic                                   p5_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p5_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p5_lba_ctrl_pipe_f ;

logic                                   p6_lba_ctrl_pipe_v_f ;
lba_ctrl_pipe_t                         p6_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p6_lba_ctrl_pipe_f ;
lba_sch_pipe_t                          p8_lba_sch_pipe_nxt ;
lba_sch_pipe_t                          p8_lba_sch_pipe_f ;
logic                                   p8_lba_sch_pipe_gp ;

logic                                   p7_lba_ctrl_pipe_v_f ;
logic                                   p7_lba_ctrl_pipe_v_1_f ;                // Replicated for drive
lba_ctrl_pipe_t                         p7_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p7_lba_ctrl_pipe_f ;

logic                                   p8_lba_ctrl_pipe_v_f ;

// Replicated for drive
logic                                   p8_lba_ctrl_pipe_v_1_f_nnc ;
lba_ctrl_pipe_t                         p8_lba_ctrl_pipe_nxt ;
lba_ctrl_pipe_t                         p8_lba_ctrl_pipe_f ;


logic                                   lba_cq2qid_rw_pipe_status ;
logic                                   p1_lba_ctrl_pipe_v_nxt_gated ;

lba_cq2qid2x_rw_pipe_t                  p1_lba_cq2qid_rw_pipe_nxt ;
lba_cq2qid2x_rw_pipe_t                  p3_lba_cq2qid_rw_pipe_f_pnc ;
logic [55:0]                            p3_lba_cq2qid_rw_pipe_qid_8_odd ;
logic [55:0]                            p3_lba_cq2qid_rw_pipe_qid_8_even ;
logic [55:0]                            p3_lba_cq2qid_rw_pipe_qid_8_x ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   p3_lba_cq2qid_qid_8_upper_ar [7:0] ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   p3_lba_cq2qid_qid_8_ar [7:0] ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]      p3_lba_cq2qid_rw_pipe_pri_scaled [HQM_QID_PER_CQ-1:0] ;
lba_cq2qid2x_rw_pipe_t                  p4_lba_cq2qid_rw_pipe_f_nc ;

aw_rwpipe_cmd_t                         p3_lba_cq2qid_rw_pipe_rw_cmd_f_nc ;

logic                                   p1_lba_cq2qid_rw_pipe_v_f_nc ;
logic                                   p2_lba_cq2qid_rw_pipe_v_f_nc ;
logic                                   p3_lba_cq2qid_rw_pipe_v_f_nc ;
logic                                   p4_lba_cq2qid_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p1_lba_cq2qid_rw_pipe_rw_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p1_lba_cq2qid_rw_pipe_addr_f_nc ;
logic [181:0]                           p1_lba_cq2qid_rw_pipe_data_f_nc ;
aw_rwpipe_cmd_t                         p2_lba_cq2qid_rw_pipe_rw_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p2_lba_cq2qid_rw_pipe_addr_f_nc ;
logic [181:0]                           p2_lba_cq2qid_rw_pipe_data_f_nc ;

logic                                   p7_lba_inp_enq_qid_par_chk_en ;
logic                                   p7_lba_inp_cmp_qid_par_chk_en ;
logic                                   p7_lba_inp_enq_qid_par_err_cond ;
logic                                   p7_lba_inp_cmp_qid_par_err_cond ;
logic                                   p7_lba_inp_qid_par_err_cond ;
logic                                   p7_lba_inp_tok_cq_par_chk_en ;
logic                                   p7_lba_inp_cmp_cq_par_chk_en ;
logic                                   p7_lba_inp_tok_cq_par_err_cond ;
logic                                   p7_lba_inp_cmp_cq_par_err_cond ;
logic                                   p7_lba_inp_cq_par_err_cond ;
logic                                   p8_lba_inp_qid_par_err_nxt ;
logic                                   p8_lba_inp_cq_par_err_nxt ;
logic                                   p3_lba_inp_tok_cnt_res_err_nxt ;
logic                                   p8_lba_inp_qid_par_err_f ;
logic                                   p8_lba_inp_cq_par_err_f ;
logic                                   p3_lba_inp_tok_cnt_res_err_f ;

logic                                   p3_lba_cq2qid_priov_par_err_cond ;
logic                                   p3_lba_cq2qid_qid0_par_err_cond ;
logic                                   p3_lba_cq2qid_qid1_par_err_cond ;
logic                                   p3_lba_cq2qid_v_err_cond ;
logic                                   p3_lba_cq2qid_v_err ;
logic                                   p4_lba_cq2qid_priov_par_err_nxt ;
logic                                   p4_lba_cq2qid_qid0_par_err_nxt ;
logic                                   p4_lba_cq2qid_qid1_par_err_nxt ;
logic                                   p4_lba_cq2qid_priov_par_err_f ;
logic                                   p4_lba_cq2qid_qid0_par_err_f ;
logic                                   p4_lba_cq2qid_qid1_par_err_f ;

lba_qid_enq_cnt_rmw_pipe_t              p5_lba_qid_enq_cnt_rmw_pipe_nxt ;
lba_qid_enq_cnt_rmw_pipe_t              p7_lba_qid_enq_cnt_rmw_pipe_f ;
logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]        p7_lba_qid_enq_cnt_p1 ;
logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]        p7_lba_qid_enq_cnt_m1 ;
lsp_lb_qid_enq_cnt_t                    p7_lba_qid_enq_cnt_upd ;
logic                                   p7_lba_qid_enq_cnt_upd_v ;
logic                                   p7_lba_qid_enq_cnt_upd_gt0 ;
logic [1:0]                             p7_lba_qid_enq_cnt_res_p1 ;
logic [1:0]                             p7_lba_qid_enq_cnt_res_m1 ;
logic                                   p7_lba_qid_enq_cnt_p1_carry ;
logic                                   p7_lba_qid_enq_cnt_m1_borrow ;
logic                                   p7_lba_qid_enq_cnt_oflow_cond ;
logic                                   p7_lba_qid_enq_cnt_uflow_cond ;
logic                                   p7_lba_qid_enq_cnt_res_chk_en ;
logic                                   p7_lba_qid_enq_cnt_res_err_cond ;

logic                                   lba_qid_enq_cnt_rmw_pipe_status_nc ;
logic                                   p5_lba_qid_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p5_lba_qid_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_qid_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_ENQ_CNT_WIDTH+2)-1:0]    p5_lba_qid_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                   p6_lba_qid_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p6_lba_qid_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_qid_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_ENQ_CNT_WIDTH+2)-1:0]    p6_lba_qid_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                   p7_lba_qid_enq_cnt_rmw_pipe_v_f_nc ;
logic                                   p8_lba_qid_enq_cnt_rmw_pipe_v_f_nc ;

lba_qid_enq_cnt_rmw_pipe_t              p8_lba_qid_enq_cnt_rmw_pipe_f_nc ;
logic                                   p8_lba_qid_enq_cnt_uflow_err_nxt ;
logic                                   p8_lba_qid_enq_cnt_oflow_err_nxt ;
logic                                   p8_lba_qid_enq_cnt_uflow_err_f ;
logic                                   p8_lba_qid_enq_cnt_oflow_err_f ;
logic                                   p8_lba_qid_enq_cnt_res_err_nxt ;
logic                                   p8_lba_qid_enq_cnt_res_err_f ;

lba_qid_dpth_thrsh_rw_pipe_t                    p5_lba_qid_dpth_thrsh_rw_pipe_nxt ;
lba_qid_dpth_thrsh_rw_pipe_t                    p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc ;
logic                                           p7_lba_qid_dpth_thrsh_par_chk_en ;
logic                                           p7_lba_qid_dpth_thrsh_par_err_cond ;
logic                                           p8_lba_qid_dpth_thrsh_par_err_nxt ;
logic                                           p8_lba_qid_dpth_thrsh_par_err_f ;
logic [1:0]                                     p7_lba_qid_dpth_thrsh_cm_code ;

logic                                           lba_qid_dpth_thrsh_rw_pipe_status_nc ;
logic                                           p5_lba_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p5_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p5_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_DPTH_THRSH_WIDTH+1)-1:0] p5_lba_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity
logic                                           p6_lba_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p6_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p6_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_DPTH_THRSH_WIDTH+1)-1:0] p6_lba_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity
logic                                           p7_lba_qid_dpth_thrsh_rw_pipe_v_f_nc ;
logic                                           p8_lba_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p8_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p8_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_DPTH_THRSH_WIDTH+1)-1:0] p8_lba_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity


lba_qid_if_cnt_rmw_pipe_t               p5_lba_qid_if_cnt_rmw_pipe_nxt ;
lba_qid_if_cnt_rmw_pipe_t               p7_lba_qid_if_cnt_rmw_pipe_f ;
logic [HQM_LSP_LB_QID_IF_CNT_WIDTH-1:0]        p7_lba_qid_if_cnt_p1 ;
logic [HQM_LSP_LB_QID_IF_CNT_WIDTH-1:0]        p7_lba_qid_if_cnt_m1 ;
lsp_lb_qid_if_cnt_t                     p7_lba_qid_if_cnt_upd ;
logic                                   p7_lba_qid_if_cnt_upd_v ;
logic                                   p7_lba_qid_if_cnt_upd_lt_lim ;
logic [1:0]                             p7_lba_qid_if_cnt_res_p1 ;
logic [1:0]                             p7_lba_qid_if_cnt_res_m1  ;
logic                                   p7_lba_qid_if_cnt_p1_carry ;
logic                                   p7_lba_qid_if_cnt_m1_borrow ;
logic                                   p7_lba_qid_if_cnt_oflow_cond ;
logic                                   p7_lba_qid_if_cnt_uflow_cond ;
logic                                   p7_lba_qid_if_cnt_res_chk_en ;
logic                                   p7_lba_qid_if_cnt_res_err_cond ;

logic                                   lba_qid_if_cnt_rmw_pipe_status_nc ;
logic                                   p5_lba_qid_if_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p5_lba_qid_if_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_qid_if_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_IF_CNT_WIDTH+2)-1:0]     p5_lba_qid_if_cnt_rmw_pipe_data_f_nc ;          // +2 for residue
logic                                   p6_lba_qid_if_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p6_lba_qid_if_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_qid_if_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_IF_CNT_WIDTH+2)-1:0]     p6_lba_qid_if_cnt_rmw_pipe_data_f_nc ;          // +2 for residue
logic                                   p7_lba_qid_if_cnt_rmw_pipe_v_f_nc ;
logic                                   p8_lba_qid_if_cnt_rmw_pipe_v_f_nc ;

lba_qid_if_cnt_rmw_pipe_t               p8_lba_qid_if_cnt_rmw_pipe_f_pnc ;
logic                                   p8_lba_qid_if_cnt_uflow_err_nxt ;
logic                                   p8_lba_qid_if_cnt_oflow_err_nxt ;
logic                                   p8_lba_qid_if_cnt_uflow_err_f ;
logic [7:0]                             p8_lba_qid_if_cnt_uflow_err_rid ;
logic                                   p8_lba_qid_if_cnt_oflow_err_f ;
logic                                   p8_lba_qid_if_cnt_res_err_nxt ;
logic                                   p8_lba_qid_if_cnt_res_err_f ;

lba_qid_if_lim_rw_pipe_t                p5_lba_qid_if_lim_rw_pipe_nxt ;
lba_qid_if_lim_rw_pipe_t                p7_lba_qid_if_lim_rw_pipe_f_pnc ;
logic                                   p7_lba_qid_if_lim_par_chk_en ;
logic                                   p7_lba_qid_if_lim_par_err_cond ;
logic                                   p8_lba_qid_if_lim_par_err_nxt ;
logic                                   p8_lba_qid_if_lim_par_err_f ;

logic                                   lba_qid_if_lim_rw_pipe_status_nc ;
logic                                   p5_lba_qid_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p5_lba_qid_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_qid_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_IF_LIM_WIDTH+1)-1:0]     p5_lba_qid_if_lim_rw_pipe_data_f_nc ;           // +1 for parity
logic                                   p6_lba_qid_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_qid_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_qid_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_IF_LIM_WIDTH+1)-1:0]     p6_lba_qid_if_lim_rw_pipe_data_f_nc ;           // +1 for parity
logic                                   p7_lba_qid_if_lim_rw_pipe_v_f_nc ;
logic                                   p8_lba_qid_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p8_lba_qid_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p8_lba_qid_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_QID_IF_LIM_WIDTH+1)-1:0]     p8_lba_qid_if_lim_rw_pipe_data_f_nc ;           // +1 for parity

logic                                   p2_lba_inp_tok_cnt_res_chk_en ;
logic                                   p2_lba_inp_tok_cnt_res_err_cond ;
logic                                   lba_cq_tok_cnt_rmw_pipe_status ;
lba_cq_tok_cnt_rmw_pipe_t               p5_lba_cq_tok_cnt_rmw_pipe_nxt ;
lba_cq_tok_cnt_rmw_pipe_t               p7_lba_cq_tok_cnt_rmw_pipe_f ;
logic [HQM_LSP_LB_CQ_TOK_CNT_WIDTH-1:0] p7_lba_cq_tok_cnt_p1 ;
logic [HQM_LSP_LB_CQ_TOK_CNT_WIDTH-1:0] p7_lba_cq_tok_cnt_mn ;
lsp_lb_cq_tok_cnt_t                     p7_lba_cq_tok_cnt_upd_cnt ;
logic                                   p7_lba_cq_tok_cnt_upd_v ;
logic                                   p7_lba_cq_tok_cnt_upd_lt_lim_next ;
logic                                   p7_lba_cq_tok_cnt_upd_gt_0 ;
logic [1:0]                             p7_lba_cq_tok_cnt_res_p1 ;
logic [1:0]                             p7_lba_cq_tok_cnt_res_mn ;
logic                                   p7_lba_cq_tok_cnt_p1_carry ;
logic                                   p7_lba_cq_tok_cnt_mn_borrow ;
logic                                   p7_lba_cq_tok_cnt_oflow_cond ;
logic                                   p7_lba_cq_tok_cnt_uflow_cond ;
logic                                   p7_lba_cq_tok_cnt_res_chk_en ;
logic                                   p7_lba_cq_tok_cnt_res_err_cond ;

aw_rmwpipe_cmd_t                        p5_lba_cq_tok_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_cq_tok_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_TOK_CNT_WIDTH+2)-1:0]     p5_lba_cq_tok_cnt_rmw_pipe_data_f_nc ;          // +2 for residue
aw_rmwpipe_cmd_t                        p6_lba_cq_tok_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_cq_tok_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_TOK_CNT_WIDTH+2)-1:0]     p6_lba_cq_tok_cnt_rmw_pipe_data_f_nc ;          // +2 for residue

lba_cq_tok_cnt_rmw_pipe_t               p8_lba_cq_tok_cnt_rmw_pipe_f_pnc ;
logic                                   p8_lba_cq_tok_cnt_oflow_err_nxt ;
logic                                   p8_lba_cq_tok_cnt_uflow_err_nxt ;
logic                                   p8_lba_cq_tok_cnt_oflow_err_f ;
logic                                   p8_lba_cq_tok_cnt_uflow_err_f ;
logic [7:0]                             p8_lba_cq_tok_cnt_uflow_err_rid  ;
logic                                   p8_lba_cq_tok_cnt_res_err_nxt ;
logic                                   p8_lba_cq_tok_cnt_res_err_f ;

lba_cq_tok_lim_rw_pipe_t                p5_lba_cq_tok_lim_rw_pipe_nxt ;
lba_cq_tok_lim_rw_pipe_t                p7_lba_cq_tok_lim_rw_pipe_f_pnc ;
logic [HQM_LSP_LB_CQ_TOK_CNT_WIDTH-1:0] p7_lba_cq_tok_limit ;
logic                                   p7_lba_cq_tok_lim_par_chk_en ;
logic                                   p7_lba_cq_tok_lim_par_err_cond ;

logic                                   p8_lba_cq_tok_lim_par_err_nxt ;
logic                                   p8_lba_cq_tok_lim_par_err_f ;
logic                                   lba_cq_tok_lim_rw_pipe_status_nc ;
logic                                   p5_lba_cq_tok_lim_rw_pipe_v_f_nc ;

aw_rwpipe_cmd_t                         p5_lba_cq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_cq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_TOK_LIM_SEL_WIDTH+1)-1:0] p5_lba_cq_tok_lim_rw_pipe_data_f_nc ;           // +1 for parity
logic                                   p6_lba_cq_tok_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_cq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_cq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_TOK_LIM_SEL_WIDTH+1)-1:0] p6_lba_cq_tok_lim_rw_pipe_data_f_nc ;           // +1 for parity
aw_rwpipe_cmd_t                         p8_lba_cq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p8_lba_cq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_TOK_LIM_SEL_WIDTH+1)-1:0] p8_lba_cq_tok_lim_rw_pipe_data_f_nc ;           // +1 for parity

lba_cq_if_cnt_rmw_pipe_t                p5_lba_cq_if_cnt_rmw_pipe_nxt ;
lba_cq_if_cnt_rmw_pipe_t                p7_lba_cq_if_cnt_rmw_pipe_f ;
logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  p7_lba_cq_if_cnt_p1 ;
logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  p7_lba_cq_if_cnt_m1 ;
lsp_lb_cq_if_cnt_t                      p7_lba_cq_if_cnt_upd_cnt ;
logic                                   p7_lba_cq_if_cnt_upd_v ;
logic                                   p7_lba_cq_if_cnt_upd_lt_lim ;
logic                                   p7_lba_cq_if_cnt_upd_le_thr ;
logic                                   p7_lba_cq_if_cnt_upd_gt_0 ;
logic [1:0]                             p7_lba_cq_if_cnt_res_p1 ;
logic [1:0]                             p7_lba_cq_if_cnt_res_m1 ;
logic                                   p7_lba_cq_if_cnt_p1_carry ;
logic                                   p7_lba_cq_if_cnt_m1_borrow ;
logic                                   p7_lba_cq_if_cnt_oflow_cond ;
logic                                   p7_lba_cq_if_cnt_uflow_cond ;
logic                                   p7_lba_cq_if_cnt_res_chk_en ;
logic                                   p7_lba_cq_if_cnt_res_err_cond ;

logic                                   lba_cq_if_cnt_rmw_pipe_status_nc ;
logic                                   p5_lba_cq_if_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p5_lba_cq_if_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_cq_if_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_CNT_WIDTH+2)-1:0]      p5_lba_cq_if_cnt_rmw_pipe_data_f_nc ;           // +2 for residue
logic                                   p6_lba_cq_if_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p6_lba_cq_if_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_cq_if_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_CNT_WIDTH+2)-1:0]      p6_lba_cq_if_cnt_rmw_pipe_data_f_nc ;           // +2 for residue
logic                                   p7_lba_cq_if_cnt_rmw_pipe_v_f_nc ;
logic                                   p8_lba_cq_if_cnt_rmw_pipe_v_f_nc ;

lba_cq_if_cnt_rmw_pipe_t                p8_lba_cq_if_cnt_rmw_pipe_f_pnc ;
logic                                   p8_lba_cq_if_cnt_uflow_err_nxt ;
logic                                   p8_lba_cq_if_cnt_oflow_err_nxt ;
logic                                   p8_lba_cq_if_cnt_uflow_err_f ;
logic [7:0]                             p8_lba_cq_if_cnt_uflow_err_rid ;
logic                                   p8_lba_cq_if_cnt_oflow_err_f ;
logic                                   p8_lba_cq_if_cnt_res_err_nxt ;
logic                                   p8_lba_cq_if_cnt_res_err_f ;

logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  p7_lba_tot_if_cnt_p1 ;
logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  p7_lba_tot_if_cnt_m1 ;
lsp_lb_cq_if_cnt_t                      p7_lba_tot_if_cnt_upd_cnt ;
logic                                   p7_lba_tot_if_cnt_upd_lt_lim ;
logic [1:0]                             p7_lba_tot_if_cnt_res_p1 ;
logic [1:0]                             p7_lba_tot_if_cnt_res_m1 ;
logic                                   p7_lba_tot_if_cnt_p1_carry ;
logic                                   p7_lba_tot_if_cnt_m1_borrow ;
logic                                   p7_lba_tot_if_cnt_oflow_cond ;
logic                                   p7_lba_tot_if_cnt_uflow_cond ;
lsp_lb_cq_if_cnt_t                      cfg_cq_ldb_tot_inflight_count_nxt ;
lsp_lb_cq_if_cnt_t                      cfg_cq_ldb_tot_inflight_count_f ;
logic [(32-HQM_LSP_LB_CQ_IF_CNT_WIDTH)-1:0]     cfg_cq_ldb_tot_inflight_count_f_nc ;
logic [1:0]                             cfg_cq_ldb_tot_inflight_count_res_nxt ;
logic [1:0]                             cfg_cq_ldb_tot_inflight_count_res_f ;
lsp_lb_cq_if_cnt_t                      p7_lba_tot_if_cnt_f ;
logic                                   p7_lba_tot_if_cnt_res_err_cond ;
logic                                   p8_lba_tot_if_cnt_res_err_nxt ;
logic                                   p8_lba_tot_if_cnt_res_err_f ;

logic                                   p8_lba_tot_if_cnt_uflow_err_nxt ;
logic                                   p8_lba_tot_if_cnt_oflow_err_nxt ;
logic                                   p8_lba_tot_if_cnt_uflow_err_f ;
logic                                   p8_lba_tot_if_cnt_oflow_err_f ;
logic [7:0]                             p8_lba_tot_if_cnt_uflow_err_rid ;

logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  cfg_cq_ldb_tot_inflight_limit_nxt ;
logic [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]  cfg_cq_ldb_tot_inflight_limit_f ;
logic [(32-HQM_LSP_LB_CQ_IF_CNT_WIDTH)-1:0]     cfg_cq_ldb_tot_inflight_limit_f_nc ;

lba_cq_if_lim_rw_pipe_t                 p5_lba_cq_if_lim_rw_pipe_nxt ;
lba_cq_if_lim_rw_pipe_t                 p7_lba_cq_if_lim_rw_pipe_f_pnc ;
logic                                   p7_lba_cq_if_lim_par_chk_en ;
logic                                   p7_lba_cq_if_lim_par_err_cond ;
logic                                   p8_lba_cq_if_lim_par_err_nxt ;
logic                                   p8_lba_cq_if_lim_par_err_f ;

logic                                   lba_cq_if_lim_rw_pipe_status_nc ;
logic                                   p5_lba_cq_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p5_lba_cq_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_cq_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_LIM_WIDTH+1)-1:0]      p5_lba_cq_if_lim_rw_pipe_data_f_nc ;            // +1 for parity
logic                                   p6_lba_cq_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_cq_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_cq_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_LIM_WIDTH+1)-1:0]      p6_lba_cq_if_lim_rw_pipe_data_f_nc ;            // +1 for parity
logic                                   p7_lba_cq_if_lim_rw_pipe_v_f_nc ;
logic                                   p8_lba_cq_if_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p8_lba_cq_if_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p8_lba_cq_if_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_LIM_WIDTH+1)-1:0]      p8_lba_cq_if_lim_rw_pipe_data_f_nc ;            // +1 for parity

lba_cq_if_thr_rw_pipe_t                 p5_lba_cq_if_thr_rw_pipe_nxt ;
lba_cq_if_thr_rw_pipe_t                 p7_lba_cq_if_thr_rw_pipe_f_pnc ;
logic                                   p7_lba_cq_if_thr_par_chk_en ;
logic                                   p7_lba_cq_if_thr_par_err_cond ;

logic                                   lba_cq_if_thr_rw_pipe_status_nc ;
logic                                   p5_lba_cq_if_thr_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p5_lba_cq_if_thr_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_cq_if_thr_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_THR_WIDTH+1)-1:0]      p5_lba_cq_if_thr_rw_pipe_data_f_nc ;            // +1 for parity
logic                                   p6_lba_cq_if_thr_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_cq_if_thr_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_cq_if_thr_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_THR_WIDTH+1)-1:0]      p6_lba_cq_if_thr_rw_pipe_data_f_nc ;            // +1 for parity
logic                                   p7_lba_cq_if_thr_rw_pipe_v_f_nc ;
logic                                   p8_lba_cq_if_thr_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p8_lba_cq_if_thr_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p8_lba_cq_if_thr_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_LB_CQ_IF_THR_WIDTH+1)-1:0]      p8_lba_cq_if_thr_rw_pipe_data_f_nc ;            // +1 for parity

logic [8:0]                             p7_lba_qid2cqidix_ix ;
logic [7:0]                             p7_lba_qid2cqidix_v_qidix ;
logic                                   p7_lba_qid2cqidix_sch_v_err_cond ;
logic                                   p7_lba_qid2cqidix_sch_v_err ;
logic                                   p7_lba_qid2cqidix_enq_v_err_cond ;
logic                                   p7_lba_qid2cqidix_enq_v_err ;

logic [HQM_QID_PER_CQ-1:0]                              p3_lba_sch_atm_req_upper ;
logic [HQM_QID_PER_CQ-1:0]                              p3_lba_sch_atm_req ;
logic [HQM_LSP_NUM_PRI_BINS-1:0]                        p3_lba_sch_atm_arb_pri_reqs_upper [HQM_QID_PER_CQ-1:0] ;
logic [HQM_LSP_NUM_PRI_BINS-1:0]                        p3_lba_sch_atm_arb_pri_reqs [HQM_QID_PER_CQ-1:0] ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_PRI_BINS)-1:0]       p3_lba_sch_atm_arb_reqs ;
logic                                                   p3_lba_sch_atm_arb_winner_v ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]                      p3_lba_sch_atm_arb_winner_pri ;
logic                                                   p3_lba_sch_atm_arb_winner_msb ;
logic [HQM_QIDIX-1:0]                                   p3_lba_sch_atm_arb_winner ;
logic                                                   p3_lba_sch_atm_arb_winner_in_seq ;
logic                                                   p3_lba_sch_atm_arb_winner_boosted ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]                p3_lba_sch_atm_index_upd_pcm ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]   p3_lba_sch_atm_count_upd_pcm ;

logic [HQM_QID_PER_CQ-1:0]                              p3_lba_sch_nalb_req_upper ;
logic [HQM_QID_PER_CQ-1:0]                              p3_lba_sch_nalb_req ;
logic [HQM_LSP_NUM_PRI_BINS-1:0]                        p3_lba_sch_nalb_arb_pri_reqs_upper [HQM_QID_PER_CQ-1:0] ;
logic [HQM_LSP_NUM_PRI_BINS-1:0]                        p3_lba_sch_nalb_arb_pri_reqs [HQM_QID_PER_CQ-1:0] ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_PRI_BINS)-1:0]       p3_lba_sch_nalb_arb_reqs ;
logic                                                   p3_lba_sch_nalb_arb_winner_v ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]                      p3_lba_sch_nalb_arb_winner_pri ;
logic                                                   p3_lba_sch_nalb_arb_winner_msb ;
logic [HQM_QIDIX-1:0]                                   p3_lba_sch_nalb_arb_winner ;
logic                                                   p3_lba_sch_nalb_arb_winner_in_seq ;
logic                                                   p3_lba_sch_nalb_arb_winner_boosted ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]                p3_lba_sch_nalb_index_upd_pcm ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]   p3_lba_sch_nalb_count_upd_pcm ;

logic                                   p3_lba_sch_atm_rlist_v ;
logic                                   p3_lba_sch_atm_slist_v ;
logic                                   p3_lba_sch_atm_rlist_slist_collide ;
logic [HQM_QID_PER_CQ_2X-1:0]           p2_lba_cq_rpri ;
logic [HQM_QID_PER_CQ_2X-1:0]           p3_lba_cq_rpri_nxt ;
logic [HQM_QID_PER_CQ_2X-1:0]           p3_lba_cq_rpri_f ;
logic                                   p3_lba_cq_qidix_rpri ;
logic                                   p3_lba_rpri_set_cond ;
logic                                   p3_lba_rpri_reset_cond ;
logic                                   p4_lba_rpri_set_nxt ;
logic                                   p4_lba_rpri_set_f ;
logic                                   p4_lba_rpri_reset_nxt ;
logic                                   p4_lba_rpri_reset_f ;
logic                                   p5_lba_rpri_set_nxt ;
logic                                   p5_lba_rpri_set_f ;
logic                                   p5_lba_rpri_reset_nxt ;
logic                                   p5_lba_rpri_reset_f ;
logic [HQM_LSP_NUM_LB_CQQIDIXB2-1:0]    p5_lba_ctrl_pipe_sch_cq_qidix ;
logic [HQM_LSP_NUM_LB_CQQIDIX-1:0]      p6_lba_rpri_nxt ;
logic [HQM_LSP_NUM_LB_CQQIDIX-1:0]      p6_lba_rpri_f ;
logic [HQM_LSP_NUM_LB_CQQIDIXB2-1:0]    p7_lba_ctrl_pipe_sch_cq_qidix ;


logic                                   p4_lba_sch_arb_winner_v ;

logic                                   p4_lba_sch_arb_atm_nalb_collide_cond_nc ;       // Used by coverage

logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   p4_lba_sch_arb_winner_qid ;
logic                                   p4_lba_sch_arb_winner_qidix_msb ;
logic [HQM_QIDIX-1:0]                   p4_lba_sch_arb_winner_qidix ;
logic [1:0]                             p4_lba_sch_arb_winner_cm_code ;

logic                                   p4_lba_nalb_sch_arb_update ;
logic                                   p4_lba_atm_sch_arb_update ;

logic                                   p4_lba_sch_arb_atm_cond ;
logic                                   p4_lba_sch_arb_atm ;
logic                                   p4_lba_sch_arb_nalb ;


logic                                                           p4_lba_sch_arb_tog_nxt ;
logic                                                           p4_lba_sch_arb_tog_f ;

logic                                           p4_lba_sch_atm_v_nxt ;
logic                                           p4_lba_sch_atm_v_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p4_lba_sch_atm_qid_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p4_lba_sch_atm_qid_f ;
logic                                           p4_lba_sch_atm_qidix_msb_nxt ;
logic                                           p4_lba_sch_atm_qidix_msb_f ;
logic [HQM_QIDIX-1:0]                           p4_lba_sch_atm_qidix_nxt ;
logic [HQM_QIDIX-1:0]                           p4_lba_sch_atm_qidix_f ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]              p4_lba_sch_atm_pri_nxt ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]              p4_lba_sch_atm_pri_f ;
logic [HQM_NUM_PRIB2-1:0]                       p4_lba_sch_atm_pri_scaled_pnc ;
logic                                           p4_lba_sch_atm_in_seq_nxt ;
logic                                           p4_lba_sch_atm_in_seq_f ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]    p4_lba_sch_atm_index_upd_pcm_nxt ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]    p4_lba_sch_atm_index_upd_pcm_f ;
logic [(HQM_LSP_NUM_PRI_BINS*HQM_QIDIX)-1:0]    p4_lba_sch_atm_index_upd ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_atm_count_upd_pcm_nxt ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_atm_count_upd_pcm_f ;
logic [(HQM_QID_PER_CQ*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_atm_count_upd ;
logic                                           p4_lba_sch_atm_rlist_nxt ;
logic                                           p4_lba_sch_atm_rlist_f ;
logic                                           p4_lba_sch_atm_in_seq ;
logic [(1+HQM_LSP_NUM_PRI_BINSB2+1)-1:0]        p4_lba_sch_atm_sel_pri ;

logic                                           p4_lba_sch_nalb_v_nxt ;
logic                                           p4_lba_sch_nalb_v_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p4_lba_sch_nalb_qid_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p4_lba_sch_nalb_qid_f ;
logic                                           p4_lba_sch_nalb_qidix_msb_nxt ;
logic                                           p4_lba_sch_nalb_qidix_msb_f ;
logic [HQM_QIDIX-1:0]                           p4_lba_sch_nalb_qidix_nxt ;
logic [HQM_QIDIX-1:0]                           p4_lba_sch_nalb_qidix_f ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]              p4_lba_sch_nalb_pri_nxt ;
logic [HQM_LSP_NUM_PRI_BINSB2-1:0]              p4_lba_sch_nalb_pri_f ;
logic                                           p4_lba_sch_nalb_in_seq_nxt ;
logic                                           p4_lba_sch_nalb_in_seq_f ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]    p4_lba_sch_nalb_index_upd_pcm_nxt ;
logic [(HQM_LSP_NUM_PRI_BINS*(HQM_QIDIX+1))-1:0]    p4_lba_sch_nalb_index_upd_pcm_f ;
logic [(HQM_LSP_NUM_PRI_BINS*HQM_QIDIX)-1:0]    p4_lba_sch_nalb_index_upd ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_nalb_count_upd_pcm_f ;
logic [(HQM_QID_PER_CQ_2X*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_nalb_count_upd_pcm_nxt ;
logic [(HQM_QID_PER_CQ*HQM_LSP_NUM_LDB_WRR_COUNTB2)-1:0]        p4_lba_sch_nalb_count_upd ;
logic                                           p4_lba_sch_nalb_in_seq ;
logic [(1+HQM_LSP_NUM_PRI_BINSB2+1)-1:0]        p4_lba_sch_nalb_sel_pri ;


logic                                   p3_lba_cq2qid0_par_chk_en_odd ;
logic                                   p3_lba_cq2qid1_par_chk_en_odd ;
logic                                   p3_lba_cq2qid0_par_chk_en_even ;
logic                                   p3_lba_cq2qid1_par_chk_en_even ;
logic                                   p3_lba_cq2qid0_par_chk_en_x ;
logic                                   p3_lba_cq2qid1_par_chk_en_x ;
logic                                   p3_lba_cq2qid_par_chk_en ;
logic [15:0]                            p3_lba_cq2qid_rw_pipe_data_priov_v_16 ;
lsp_cfg_cq2priov_t                      p3_lba_cq2qid_rw_pipe_data_priov_x ;
lsp_cfg_cq2qid_t                        p3_lba_cq2qid_rw_pipe_data_qid_ls_x ;
lsp_cfg_cq2qid_t                        p3_lba_cq2qid_rw_pipe_data_qid_ms_x ;

logic                                   lba_qid2cqidix_rw_pipe_status;
lba_qid2cqidix_rw_pipe_t                p5_lba_qid2cqidix_rw_pipe_nxt ;
lba_qid2cqidix_rw_pipe_t                p7_lba_qid2cqidix_rw_pipe_f ;
lba_qid2cqidix_rw_pipe_t                p8_lba_qid2cqidix_rw_pipe_f_nc ;

logic                                   p5_lba_qid2cqidix_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p5_lba_qid2cqidix_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_qid2cqidix_rw_pipe_addr_f_nc ;
logic [(512+16)-1:0]                    p5_lba_qid2cqidix_rw_pipe_data_f_nc ;
logic                                   p6_lba_qid2cqidix_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_qid2cqidix_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_qid2cqidix_rw_pipe_addr_f_nc ;
logic [(512+16)-1:0]                    p6_lba_qid2cqidix_rw_pipe_data_f_nc ;
logic                                   p7_lba_qid2cqidix_rw_pipe_v_f_nc ;
logic                                   p8_lba_qid2cqidix_rw_pipe_v_f_nc ;

logic                                   p7_lba_qid2cqidix_par_chk_en ;
logic [15:0]                            p7_lba_qid2cqidix_par_err_cond ;

logic [15:0]                            p8_lba_qid2cqidix_par_err_nxt ;
logic [15:0]                            p8_lba_qid2cqidix_par_err_f ;
logic                                   p8_lba_qid2cqidix_par_err_any ;

lba_qid2cqidix_rw_pipe_t                p5_lba_blast_qid2cqidix_rw_pipe_nxt ;
lba_qid2cqidix_rw_pipe_t                p7_lba_blast_qid2cqidix_rw_pipe_f_pnc ;
lba_qid2cqidix_rw_pipe_t                p8_lba_blast_qid2cqidix_rw_pipe_f_nc ;

logic                                   lba_blast_qid2cqidix_rmw_pipe_status_nc ;
logic                                   p5_lba_blast_qid2cqidix_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p5_lba_blast_qid2cqidix_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_blast_qid2cqidix_rw_pipe_addr_f_nc ;
logic [(512+16)-1:0]                    p5_lba_blast_qid2cqidix_rw_pipe_data_f_nc ;             // +16 for parity bits
logic                                   p6_lba_blast_qid2cqidix_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                         p6_lba_blast_qid2cqidix_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_blast_qid2cqidix_rw_pipe_addr_f_nc ;
logic [(512+16)-1:0]                    p6_lba_blast_qid2cqidix_rw_pipe_data_f_nc ;             // +16 for parity bits
logic                                   p7_lba_blast_qid2cqidix_rw_pipe_v_f_nc ;
logic                                   p8_lba_blast_qid2cqidix_rw_pipe_v_f_nc ;

logic                                   p7_lba_blast_qid2cqidix_par_chk_en ;
logic [15:0]                            p7_lba_blast_qid2cqidix_par_err_cond ;

logic [15:0]                            p8_lba_blast_qid2cqidix_par_err_nxt ;
logic [15:0]                            p8_lba_blast_qid2cqidix_par_err_f ;
logic                                   p8_lba_blast_qid2cqidix_par_err_any ;

logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_has_space ;

logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_tok_v_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_tok_v_f ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_if_v_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_if_v_f ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_thr_v_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_thr_v_f ;
logic                                   p8_lba_tot_if_v_nxt ;
logic                                   p8_lba_tot_if_v_f ;

logic                                   p7_lba_cq_tok_v_upd ;
logic                                   p8_lba_cq_tok_v_upd_nxt ;
logic                                   p8_lba_cq_tok_v_upd_f ;
logic                                   p7_lba_cq_if_v_upd ;
logic                                   p8_lba_cq_if_v_upd_nxt ;
logic                                   p8_lba_cq_if_v_upd_f ;

logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_tok_cnt_v_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_tok_cnt_v_f ;

logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_if_cnt_v_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p8_lba_cq_if_cnt_v_f ;

logic [511:0]                           p7_lba_qid2cqidix_v ;
logic [15:0]                            p7_lba_qid2cqidix_p ;

logic [511:0]                           p8_lba_qidix_if_v_nxt ;
logic [511:0]                           p8_lba_qidix_if_v_f ;
logic                                   p7_lba_qidix_if_v_upd ;
logic                                   p8_lba_qidix_if_v_upd_nxt ;
logic                                   p8_lba_qidix_if_v_upd_f ;

logic [511:0]                           p8_lba_qidix_sch_v_nxt ;
logic [511:0]                           p8_lba_qidix_sch_v_f ;
logic                                   p7_lba_qidix_sch_v_upd ;
logic                                   p8_lba_qidix_sch_v_upd_nxt ;
logic                                   p8_lba_qidix_sch_v_upd_f ;

logic [511:0]                           p8_lba_qidix_has_work ;

logic                                   p7_lba_blast_slist ;
logic                                   p7_lba_blast_rlist ;
logic                                   p7_lba_blast_nalb ;
logic                                   p7_lba_set_cmpblast ;
logic [511:0]                           p7_lba_blast_qid2cqidix_v ;
logic [15:0]                            p7_lba_blast_qid2cqidix_p ;
logic                                   p7_lba_sched ;

logic [511:0]                           p8_lba_blast_qid2cqidix_v_nxt ;
logic [511:0]                           p8_lba_blast_qid2cqidix_v_f ;

logic                                   nalb_sel_nalb_fifo_credit_err_cond ;
logic                                   nalb_sel_nalb_fifo_cerr_reported_nxt ;
logic                                   nalb_sel_nalb_fifo_cerr_reported_f ;
logic                                   p9_lba_nalb_sch_err_nxt ;
logic                                   p9_lba_nalb_sch_err_f ;

logic [6:0]                             lsp_nalb_sch_unoord_status_pnc ;
logic                                   lsp_nalb_sch_unoord_in_ready ;

logic                                   p7_lba_tot_enq_cnt_upd_v ;
lsp_arch_cnt_t                          p7_lba_tot_enq_cnt_upd ;
logic [HQM_LSP_ARCH_CNT_WIDTH-1:0]      p7_lba_tot_enq_cnt_p1 ;
logic [1:0]                             p7_lba_tot_enq_cnt_res_p1 ;
lba_tot_enq_cnt_rmw_pipe_t              p5_lba_tot_enq_cnt_rmw_pipe_nxt ;
lba_tot_enq_cnt_rmw_pipe_t              p7_lba_tot_enq_cnt_rmw_pipe_f_pnc ;

lba_tot_enq_cnt_rmw_pipe_t              p8_lba_tot_enq_cnt_rmw_pipe_f_pnc ;
logic                                   p8_lba_tot_enq_cnt_res_chk_en ;
logic                                   p9_lba_tot_enq_cnt_res_err_nxt ;
logic                                   p9_lba_tot_enq_cnt_res_err_f ;

logic                                   lba_tot_enq_cnt_rmw_pipe_status_nc ;
logic                                   p5_lba_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p5_lba_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p5_lba_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]  p5_lba_tot_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                   p6_lba_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p6_lba_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]            p6_lba_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]  p6_lba_tot_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                   p7_lba_tot_enq_cnt_rmw_pipe_v_f_nc ;
logic                                   p8_lba_tot_enq_cnt_rmw_pipe_v_f_nc ;

logic                                   p7_lba_tot_sch_cnt_upd_v ;
lsp_arch_cnt_t                          p7_lba_tot_sch_cnt_upd ;
logic [HQM_LSP_ARCH_CNT_WIDTH-1:0]      p7_lba_tot_sch_cnt_p1 ;
logic [1:0]                             p7_lba_tot_sch_cnt_res_p1 ;
lba_tot_sch_cnt_rmw_pipe_t              p5_lba_tot_sch_cnt_rmw_pipe_nxt ;
lba_tot_sch_cnt_rmw_pipe_t              p7_lba_tot_sch_cnt_rmw_pipe_f_pnc ;

lba_tot_sch_cnt_rmw_pipe_t              p8_lba_tot_sch_cnt_rmw_pipe_f_pnc ;
logic                                   p8_lba_tot_sch_cnt_res_chk_en ;
logic                                   p9_lba_tot_sch_cnt_res_err_nxt ;
logic                                   p9_lba_tot_sch_cnt_res_err_f ;

logic                                   lba_tot_sch_cnt_rmw_pipe_status_nc ;
logic                                   p5_lba_tot_sch_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p5_lba_tot_sch_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p5_lba_tot_sch_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]  p5_lba_tot_sch_cnt_rmw_pipe_datav_f_nc ;        // +2 for residue
logic                                   p6_lba_tot_sch_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                        p6_lba_tot_sch_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]             p6_lba_tot_sch_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]  p6_lba_tot_sch_cnt_rmw_pipe_datav_f_nc ;        // +2 for residue
logic                                   p7_lba_tot_sch_cnt_rmw_pipe_v_f_nc ;
logic                                   p8_lba_tot_sch_cnt_rmw_pipe_v_f_nc ;

logic                                   p7_lba_perf_sch_count_upd_v ;

logic                                           p7_lba_enq_cnt_gt_max_depth ;
logic                                           p7_lba_max_enq_depth_upd_v ;
logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]        p7_lba_max_enq_depth_upd ;
lba_max_enq_depth_rmw_pipe_t                    p5_lba_max_enq_depth_rmw_pipe_nxt ;
lba_max_enq_depth_rmw_pipe_t                    p7_lba_max_enq_depth_rmw_pipe_f ;
lba_max_enq_depth_rmw_pipe_t                    p8_lba_max_enq_depth_rmw_pipe_f_nc ;

logic                                           lba_max_enq_depth_rmw_pipe_status_nc ;
logic                                           p5_lba_max_enq_depth_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p5_lba_max_enq_depth_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p5_lba_max_enq_depth_rmw_pipe_addr_f_nc ;
logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]        p5_lba_max_enq_depth_rmw_pipe_data_f_nc ;
logic                                           p6_lba_max_enq_depth_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p6_lba_max_enq_depth_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p6_lba_max_enq_depth_rmw_pipe_addr_f_nc ;
logic [HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0]        p6_lba_max_enq_depth_rmw_pipe_data_f_nc ;
logic                                           p7_lba_max_enq_depth_rmw_pipe_v_f_nc ;
logic                                           p8_lba_max_enq_depth_rmw_pipe_v_f_nc ;


logic                                           p1_lba_ctrl_pipe_f_pcm_nxt ;		// piared CQ Mode
logic                                           p1_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p2_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p3_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p4_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p5_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p6_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p7_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic                                           p8_lba_ctrl_pipe_f_pcm ;		// piared CQ Mode
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p1_lba_ctrl_pipe_nxt_sch_pcq ;          // paired CQ, 1 less bit
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p1_lba_ctrl_pipe_f_sch_pcq ;            // paired CQ, 1 less bit
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p4_lba_ctrl_pipe_f_sch_pcq ;            // paired CQ, 1 less bit

logic                                           p1_lba_nalb_index_v_f_nc ;
logic                                           p2_lba_nalb_index_v_f_nc ;
logic                                           p3_lba_nalb_index_v_f_nc ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       p3_lba_nalb_index_rw_pipe_data_f ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       p3_lba_nalb_index_rw_pipe_data_nobyp_f_nc ;
lba_ldb_arb_index2x_t                           p3_lba_nalb_index_rw_pipe_data_struct ;
lba_ldb_arb_index_t                             p3_lba_nalb_index_rw_pipe_data_odd ;
lba_ldb_arb_index_t                             p3_lba_nalb_index_rw_pipe_data_even ;
lba_ldb_arb_index_t                             p3_lba_nalb_index_rw_pipe_data_x ;
lba_ldb_arb_index_pcm_t                         p3_lba_nalb_index_rw_pipe_data_pcm ;
lba_ldb_arb_index_t                             p3_lba_nalb_index_rw_pipe_data_unch ;
lba_ldb_arb_index_t                             p4_lba_nalb_index_rw_pipe_data_unch_nxt ;
lba_ldb_arb_index_t                             p4_lba_nalb_index_rw_pipe_data_unch_f ;
lba_ldb_arb_index2x_t                           p4_lba_nalb_index_rw_pipe_data_struct ;

logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p1_lba_nalb_index_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p2_lba_nalb_index_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p3_lba_nalb_index_rw_pipe_addr_f_nc ;

logic                                           pw_lba_nalb_index_v_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        pw_lba_nalb_index_rw_pipe_addr_f_nc ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       pw_lba_nalb_index_rw_pipe_data_f_nc ;

logic                                           lba_nalb_pri_arbindex_pipe_status ;

logic                                           p1_lba_atm_index_v_f_nc ;
logic                                           p2_lba_atm_index_v_f_nc ;
logic                                           p3_lba_atm_index_v_f_nc ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       p3_lba_atm_index_rw_pipe_data_f ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       p3_lba_atm_index_rw_pipe_data_nobyp_f_nc ;
lba_ldb_arb_index2x_t                           p3_lba_atm_index_rw_pipe_data_struct ;
lba_ldb_arb_index_t                             p3_lba_atm_index_rw_pipe_data_odd ;
lba_ldb_arb_index_t                             p3_lba_atm_index_rw_pipe_data_even ;
lba_ldb_arb_index_t                             p3_lba_atm_index_rw_pipe_data_x ;
lba_ldb_arb_index_pcm_t                         p3_lba_atm_index_rw_pipe_data_pcm ;
lba_ldb_arb_index_t                             p3_lba_atm_index_rw_pipe_data_unch ;
lba_ldb_arb_index_t                             p4_lba_atm_index_rw_pipe_data_unch_nxt ;
lba_ldb_arb_index_t                             p4_lba_atm_index_rw_pipe_data_unch_f ;
lba_ldb_arb_index2x_t                           p4_lba_atm_index_rw_pipe_data_struct ;

logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p1_lba_atm_index_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p2_lba_atm_index_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        p3_lba_atm_index_rw_pipe_addr_f_nc ;

logic                                           pw_lba_atm_index_v_f_nc ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        pw_lba_atm_index_rw_pipe_addr_f_nc ;
logic [HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0]       pw_lba_atm_index_rw_pipe_data_f_nc ;

logic                                           lba_atm_pri_arbindex_pipe_status ;

logic                                   qed_deq_credit_error ;
logic                                   qed_deq_credit_empty ;
logic                                   qed_deq_credit_afull ;

logic                                   aqed_deq_credit_error ;
logic                                   aqed_deq_credit_empty ;
logic                                   aqed_deq_credit_afull ;

logic                                   p1_lbwu_ctrl_pipe_v_f ;
logic                                   p2_lbwu_ctrl_pipe_v_f ;
logic                                   p3_lbwu_ctrl_pipe_v_f ;
logic                                   p4_lbwu_ctrl_pipe_v_f ;

logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_ow_nxt ;
logic [HQM_NUM_LB_CQ-1:0]               p0_lba_cq_ow_f ;

logic                                   lbwu_cq_wu_cnt_rmw_pipe_status ;
logic                                   p3_lbwu_cq_wu_cnt_upd_v_func ;
logic                                   p4_lbwu_cq_wu_cnt_upd_v_f ;
logic [HQM_NUM_LB_CQB2-1:0]             p4_lbwu_cq_wu_cnt_upd_cq_f ;
logic                                   p4_lbwu_cq_wu_cnt_upd_gt_lim_f ;

logic                                   p3_lbwu_cq_wu_cnt_res_err_cond ;
logic                                   p4_lbwu_cq_wu_cnt_res_err_nxt ;
logic                                   p4_lbwu_cq_wu_cnt_res_err_f ;

logic                                   p3_lbwu_cq_wu_lim_par_err_cond ;
logic                                   p4_lbwu_cq_wu_lim_par_err_nxt ;
logic                                   p4_lbwu_cq_wu_lim_par_err_f ;

logic                                   p3_lbwu_inp_par_err_cond ;
logic                                   p4_lbwu_inp_par_err_nxt ;
logic                                   p4_lbwu_inp_par_err_f ;

logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count_nc ;

logic                   cfg_sched_slot_count_en ;
logic                   cfg_sched_slot_count_clr ;
logic [7:0]             cfg_sched_slot_count_cq ;
logic                   cfg_sched_slot_count_trigger ;

logic [7:0]             cfg_sched_slot_count_inc_nxt ;
logic [7:0]             cfg_sched_slot_count_inc_f ;
logic                   cfg_sched_slot_count_prev_slot_v_nxt ;
logic                   cfg_sched_slot_count_prev_slot_v_f ;
logic [2:0]             cfg_sched_slot_count_prev_slot_nxt ;
logic [2:0]             cfg_sched_slot_count_prev_slot_f ;

//------------------------------------------------------------------------------------------------
// ATQ pipe declarations
logic                                           atq_input_arb_new_both ;
logic                                           atq_input_arb_new_either ;
logic [1:0]                                     atq_input_arb_reqs ;
logic                                           atq_input_arb_update ;
logic                                           atq_input_arb_winner_pre_v ;
logic                                           atq_input_arb_winner_v ;
logic                                           atq_input_arb_winner ;
logic                                           atq_input_arb_sch ;
logic                                           atq_input_arb_pre_enq ;
logic                                           atq_input_arb_enq ;
logic                                           atq_input_arb_pre_cmp ;
logic                                           atq_input_arb_cmp ;
lsp_lb_qid_t                                    atq_input_arb_sch_qid ;
logic                                           atq_input_arb_tog_nxt ;
logic                                           atq_input_arb_tog_f ;


lsp_pipe_ctrl_t                                 p0_atq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p1_atq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p2_atq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p3_atq_ctrl_pipe ;
logic                                           p4_atq_ctrl_pipe_en ;

logic                                           p0_atq_ctrl_pipe_v_nxt ;
logic                                           p0_atq_ctrl_pipe_v_nxt_gated ;
logic                                           p0_atq_ctrl_pipe_v_f ;
atq_ctrl_pipe_t                                 p0_atq_ctrl_pipe_nxt ;
atq_ctrl_pipe_t                                 p0_atq_ctrl_pipe_f ;

logic                                           p1_atq_ctrl_pipe_v_f ;
atq_ctrl_pipe_t                                 p1_atq_ctrl_pipe_nxt ;
atq_ctrl_pipe_t                                 p1_atq_ctrl_pipe_f ;

logic                                           p2_atq_ctrl_pipe_v_f ;
atq_ctrl_pipe_t                                 p2_atq_ctrl_pipe_nxt ;
atq_ctrl_pipe_t                                 p2_atq_ctrl_pipe_f ;

logic                                           p3_atq_ctrl_pipe_v_f ;

logic                                           atq_input_req_v ;

logic                                           p2_atq_inp_enq_qid_p ;
logic                                           p2_atq_inp_cmp_qid_p ;
logic                                           p2_atq_inp_enq_qid_par_chk_en ;
logic                                           p2_atq_inp_cmp_qid_par_chk_en ;
logic                                           p2_atq_inp_enq_qid_par_err_cond ;
logic                                           p2_atq_inp_cmp_qid_par_err_cond ;
logic                                           p2_atq_inp_qid_par_err_cond ;
logic                                           p3_atq_inp_qid_par_err_nxt ;
logic                                           p3_atq_inp_qid_par_err_f ;

logic                                           p2_atq_enq_cnt_upd_v ;
lsp_atq_enq_cnt_t                               p2_atq_enq_cnt_upd ;
logic [HQM_LSP_ATQ_ENQ_CNT_WIDTH-1:0]           p2_atq_enq_cnt_p1 ;
logic [HQM_LSP_ATQ_ENQ_CNT_WIDTH-1:0]           p2_atq_enq_cnt_m1 ;
logic                                           p2_atq_enq_cnt_upd_gt0 ;
logic [1:0]                                     p2_atq_enq_cnt_res_p1 ;
logic [1:0]                                     p2_atq_enq_cnt_res_m1 ;
logic                                           p2_atq_enq_cnt_p1_carry ;
logic                                           p2_atq_enq_cnt_m1_borrow ;
logic                                           p2_atq_enq_cnt_oflow_cond ;
logic                                           p2_atq_enq_cnt_uflow_cond ;
logic                                           atq_enq_cnt_rmw_pipe_status ;
atq_enq_cnt_rmw_pipe_t                          p0_atq_enq_cnt_rmw_pipe_nxt ;
atq_enq_cnt_rmw_pipe_t                          p0_atq_enq_cnt_rmw_pipe_f_pnc ;
atq_enq_cnt_rmw_pipe_t                          p1_atq_enq_cnt_rmw_pipe_f_pnc ;
atq_enq_cnt_rmw_pipe_t                          p2_atq_enq_cnt_rmw_pipe_f ;
atq_enq_cnt_rmw_pipe_t                          p3_atq_enq_cnt_rmw_pipe_f_nc ;
logic                                           p2_atq_enq_cnt_res_chk_en ;
logic                                           p2_atq_enq_cnt_res_err_cond ;
logic                                           p3_atq_enq_cnt_uflow_err_nxt ;
logic                                           p3_atq_enq_cnt_oflow_err_nxt ;
logic                                           p3_atq_enq_cnt_uflow_err_f ;
logic                                           p3_atq_enq_cnt_oflow_err_f ;
logic                                           p3_atq_enq_cnt_res_err_nxt ;
logic                                           p3_atq_enq_cnt_res_err_f ;

lsp_atq_atm_active_t                            p2_atq_atm_active_curr ;
logic                                           p3_atq_atm_active_bypdata_sel_nxt ;
lsp_atq_atm_active_t                            p3_atq_atm_active_bypdata_nxt ;
logic                                           p3_atq_atm_active_bypaddr_sel_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p3_atq_atm_active_bypaddr_nxt ;
atq_atm_active_rmw_pipe_t                       p0_atq_atm_active_rmw_pipe_nxt ;
aw_rmwpipe_cmd_t                                p0_atq_atm_active_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p0_atq_atm_active_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_ATM_ACTIVE_WIDTH+2)-1:0]    p0_atq_atm_active_rmw_pipe_data_f_nc ;          // +2 for residue
aw_rmwpipe_cmd_t                                p1_atq_atm_active_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p1_atq_atm_active_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_ATM_ACTIVE_WIDTH+2)-1:0]    p1_atq_atm_active_rmw_pipe_data_f_nc ;          // +2 for residue
atq_atm_active_rmw_pipe_t                       p2_atq_atm_active_rmw_pipe_f_pnc ;
atq_atm_active_rmw_pipe_t                       p3_atq_atm_active_rmw_pipe_f_nc ;
logic                                           atq_atm_active_rmw_pipe_status_nc ;
logic                                           p0_atq_atm_active_rmw_pipe_v_f_nc ;
logic                                           p1_atq_atm_active_rmw_pipe_v_f_nc ;
logic                                           p2_atq_atm_active_rmw_pipe_v_f_nc ;
logic                                           p3_atq_atm_active_rmw_pipe_v_f_nc ;

atq_qid_dpth_thrsh_rw_pipe_t                            p0_atq_qid_dpth_thrsh_rw_pipe_nxt ;
atq_qid_dpth_thrsh_rw_pipe_t                            p2_atq_qid_dpth_thrsh_rw_pipe_f_pnc ;

logic                                                   atq_qid_dpth_thrsh_rw_pipe_status_nc ;
logic                                                   p0_atq_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                         p0_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                   p0_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH+1)-1:0]        p0_atq_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity
logic                                                   p1_atq_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                         p1_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                   p1_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH+1)-1:0]        p1_atq_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity
logic                                                   p2_atq_qid_dpth_thrsh_rw_pipe_v_f_nc ;
logic                                                   p3_atq_qid_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                         p3_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                   p3_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH+1)-1:0]        p3_atq_qid_dpth_thrsh_rw_pipe_data_f_nc ;       // +1 for parity

logic                                           p2_atq_atm_active_sum_v ;
lsp_atq_aqed_act_cnt_t                          p3_atq_aqed_act_cnt_upd_nxt ;
lsp_atq_aqed_act_cnt_t                          p3_atq_aqed_act_cnt_upd_f ;
lsp_atq_atm_active_t                            p3_atq_atm_active_curr_nxt ;
lsp_atq_atm_active_t                            p3_atq_atm_active_curr_f ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_aqed_act_cnt_qid_nxt ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_aqed_act_cnt_qid_f ;
lsp_atq_qid_dpth_thrsh_t                        p3_atq_qid_dpth_thrsh_nxt ;
lsp_atq_qid_dpth_thrsh_t                        p3_atq_qid_dpth_thrsh_f ;
logic                                           p3_atq_atm_active_sum_v_nxt ;
logic                                           p3_atq_atm_active_sum_v_f ;
lsp_atq_atm_active_t                            p3_atq_atm_active_sum ;
logic                                           p3_atq_atm_active_sum_carry ;
lsp_atq_atm_active_t                            p3_atq_atm_active_tot ;
logic [1:0]                                     p3_atq_qid_dpth_thrsh_cm_code ;
logic                                           p3_atq_atm_active_oflow_cond ;
logic                                           p4_atq_atm_active_oflow_err_nxt ;
logic                                           p4_atq_atm_active_oflow_err_f ;
logic                                           p3_atq_atm_active_res_chk_en ;
logic                                           p3_atq_atm_active_res_err_cond ;
logic                                           p4_atq_atm_active_res_err_nxt ;
logic                                           p4_atq_atm_active_res_err_f ;
logic                                           p3_atq_qid_dpth_thrsh_par_chk_en ;
logic                                           p3_atq_qid_dpth_thrsh_par_err_cond ;
logic                                           p4_atq_qid_dpth_thrsh_par_err_nxt ;
logic                                           p4_atq_qid_dpth_thrsh_par_err_f ;

logic                                           p2_atq_aqed_act_cnt_upd_v ;
lsp_atq_aqed_act_cnt_t                          p2_atq_aqed_act_cnt_upd ;
logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      p2_atq_aqed_act_cnt_p1 ;
logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      p2_atq_aqed_act_cnt_m1 ;
logic                                           p2_atq_aqed_act_cnt_upd_lt_lim ;
logic                                           p2_atq_aqed_act_cnt_upd_gt_0 ;
logic                                           p2_atq_aqed_act_cnt_upd_eq_0 ;
logic [1:0]                                     p2_atq_aqed_act_cnt_res_p1 ;
logic [1:0]                                     p2_atq_aqed_act_cnt_res_m1 ;
logic                                           p2_atq_aqed_act_cnt_p1_carry ;
logic                                           p2_atq_aqed_act_cnt_m1_borrow ;
logic                                           p2_atq_aqed_act_cnt_oflow_cond ;
logic                                           p2_atq_aqed_act_cnt_uflow_cond ;
atq_aqed_act_cnt_rmw_pipe_t                     p0_atq_aqed_act_cnt_rmw_pipe_nxt ;
atq_aqed_act_cnt_rmw_pipe_t                     p0_atq_aqed_act_cnt_rmw_pipe_f_pnc ;
atq_aqed_act_cnt_rmw_pipe_t                     p1_atq_aqed_act_cnt_rmw_pipe_f_pnc ;
atq_aqed_act_cnt_rmw_pipe_t                     p2_atq_aqed_act_cnt_rmw_pipe_f ;
atq_aqed_act_cnt_rmw_pipe_t                     p3_atq_aqed_act_cnt_rmw_pipe_f_nc ;
logic                                           p2_atq_aqed_act_cnt_res_chk_en ;
logic                                           p2_atq_aqed_act_cnt_res_err_cond ;
logic                                           p3_atq_aqed_act_cnt_uflow_err_nxt ;
logic                                           p3_atq_aqed_act_cnt_oflow_err_nxt ;
logic                                           p3_atq_aqed_act_cnt_uflow_err_f ;
logic                                           p3_atq_aqed_act_cnt_oflow_err_f ;
logic                                           p3_atq_aqed_act_cnt_res_err_nxt ;
logic                                           p3_atq_aqed_act_cnt_res_err_f ;

logic                                           aqed_lsp_dec_fid_cnt_v_f ;
logic                                           aqed_lsp_dec_fid_cnt_v_last_nxt ;
logic                                           aqed_lsp_dec_fid_cnt_v_last_f ;
logic                                           p3_atq_fid_inflight_cnt_upd_inc ;
logic                                           p3_atq_fid_inflight_cnt_upd_dec ;
logic                                           p3_atq_fid_inflight_cnt_upd_v ;

logic [11:0]                                    p3_atq_fid_inflight_cnt_m1 ;
logic [11:0]                                    p3_atq_fid_inflight_cnt_p1 ;
logic [1:0]                                     p3_atq_fid_inflight_cnt_res_m1 ;
logic [1:0]                                     p3_atq_fid_inflight_cnt_res_p1 ;
logic                                           p3_atq_fid_inflight_cnt_p1_carry ;
logic                                           p3_atq_fid_inflight_cnt_m1_borrow ;
lsp_atq_fid_if_cnt_t                            p3_atq_fid_inflight_cnt_upd ;
logic                                           p3_atq_fid_inflight_cnt_oflow_cond ;
logic                                           p3_atq_fid_inflight_cnt_uflow_cond ;

logic                                           p3_atq_fid_inflight_cnt_lt_lim ;
logic                                           p3_atq_fid_inflight_cnt_eq_lim ;
logic                                           p3_atq_fid_inflight_cnt_gt_lim ;

logic                                           p4_atq_fid_inflight_cnt_oflow_err_nxt ;
logic                                           p4_atq_fid_inflight_cnt_oflow_err_f ;
logic                                           p4_atq_fid_inflight_cnt_uflow_err_nxt ;
logic                                           p4_atq_fid_inflight_cnt_uflow_err_f ;
logic                                           p3_atq_fid_inflight_cnt_res_err_cond ;
logic                                           p4_atq_fid_inflight_cnt_res_err_nxt ;
logic                                           p4_atq_fid_inflight_cnt_res_err_f ;

logic                                           atq_aqed_act_cnt_rmw_pipe_status_nc ;
logic                                           p0_atq_aqed_act_cnt_rmw_pipe_v_f_nc ;
logic                                           p1_atq_aqed_act_cnt_rmw_pipe_v_f_nc ;
logic                                           p2_atq_aqed_act_cnt_rmw_pipe_v_f_nc ;
logic                                           p3_atq_aqed_act_cnt_rmw_pipe_v_f_nc ;

lsp_atq_aqed_act_cnt_t                          cfg_aqed_tot_enqueue_count_nxt ;
lsp_atq_aqed_act_cnt_t                          cfg_aqed_tot_enqueue_count_f ;
logic [(32-HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH)-1:0]         cfg_aqed_tot_enqueue_count_f_nc ;
logic [1:0]                                     cfg_aqed_tot_enqueue_count_res_nxt ;
logic [1:0]                                     cfg_aqed_tot_enqueue_count_res_f ;

lsp_atq_aqed_act_cnt_t                          p3_atq_tot_act_cnt_f ;
lsp_atq_aqed_act_cnt_t                          p3_atq_tot_act_cnt_upd ;
logic [1:0]                                     p3_atq_tot_act_cnt_res_p1 ;
logic [1:0]                                     p3_atq_tot_act_cnt_res_m1 ;
logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      p3_atq_tot_act_cnt_p1 ;
logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      p3_atq_tot_act_cnt_m1 ;
logic                                           p3_atq_tot_act_cnt_p1_carry ;
logic                                           p3_atq_tot_act_cnt_m1_borrow ;
logic                                           p3_atq_tot_act_cnt_oflow_cond ;
logic                                           p3_atq_tot_act_cnt_uflow_cond ;
logic                                           p3_atq_tot_act_cnt_upd_inc ;
logic                                           p3_atq_tot_act_cnt_upd_dec ;
logic                                           p3_atq_tot_act_cnt_upd_v ;

logic                                           p3_atq_tot_act_cnt_lt_lim ;
logic                                           p3_atq_tot_act_cnt_eq_lim ;
logic                                           p3_atq_tot_act_cnt_gt_lim ;

logic                                           p4_atq_tot_act_cnt_oflow_err_nxt ;
logic                                           p4_atq_tot_act_cnt_uflow_err_nxt ;
logic                                           p4_atq_tot_act_cnt_oflow_err_f ;
logic                                           p4_atq_tot_act_cnt_uflow_err_f ;
logic                                           p3_atq_aqed_tot_enq_cnt_res_err_cond ;
logic                                           p4_atq_aqed_tot_enq_cnt_res_err_nxt ;
logic                                           p4_atq_aqed_tot_enq_cnt_res_err_f ;

lsp_atq_fid_if_cnt_t                            cfg_fid_inflight_count_nxt ;
lsp_atq_fid_if_cnt_t                            cfg_fid_inflight_count_f ;
logic [(32-HQM_LSP_ATQ_FID_IF_CNT_WIDTH)-1:0]            cfg_fid_inflight_count_f_nc ;
logic [1:0]                                     cfg_fid_inflight_count_res_nxt ;
logic [1:0]                                     cfg_fid_inflight_count_res_f ;
logic [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0]        cfg_fid_inflight_limit_nxt ;
logic [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0]        cfg_fid_inflight_limit_f ;
logic [(32-HQM_LSP_ATQ_FID_IF_CNT_WIDTH)-1:0]   cfg_fid_inflight_limit_f_nc ;

logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      cfg_aqed_tot_enqueue_limit_nxt ;
logic [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]      cfg_aqed_tot_enqueue_limit_f ;
logic [(32-HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH)-1:0] cfg_aqed_tot_enqueue_limit_f_nc ;

atq_aqed_act_lim_rw_pipe_t                      p0_atq_aqed_act_lim_rw_pipe_nxt ;
atq_aqed_act_lim_rw_pipe_t                      p2_atq_aqed_act_lim_rw_pipe_f_pnc ;
logic                                           p2_atq_aqed_act_lim_par_chk_en ;
logic                                           p2_atq_aqed_act_lim_par_err_cond ;
logic                                           p3_atq_aqed_act_lim_par_err_nxt ;
logic                                           p3_atq_aqed_act_lim_par_err_f ;

logic                                           atq_aqed_act_lim_rw_pipe_status_nc ;
logic                                           p0_atq_aqed_act_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p0_atq_aqed_act_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p0_atq_aqed_act_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH+1)-1:0]  p0_atq_aqed_act_lim_rw_pipe_data_f_nc ;                 // +1 for parity
logic                                           p1_atq_aqed_act_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p1_atq_aqed_act_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p1_atq_aqed_act_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH+1)-1:0]  p1_atq_aqed_act_lim_rw_pipe_data_f_nc ;                 // +1 for parity
logic                                           p2_atq_aqed_act_lim_rw_pipe_v_f_nc ;
logic                                           p3_atq_aqed_act_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p3_atq_aqed_act_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p3_atq_aqed_act_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH+1)-1:0]  p3_atq_aqed_act_lim_rw_pipe_data_f_nc ;                 // +1 for parity

logic [HQM_NUM_LB_QID-1:0]                      p3_atq_sch_hit ;

logic [HQM_NUM_LB_QID-1:0]                      p3_atq_p2_enq_hit ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_p2_cmp_hit ;

logic [HQM_NUM_LB_QID-1:0]                      p3_atq_qid_v_nxt ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_qid_v_f ;
logic                                           p3_atq_qid_v_any ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_nfull_nxt ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_nfull_f ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_empty_nxt ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_empty_f ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_act_v_nxt ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_aqed_act_v_f ;

logic [1:0]                                     p4_atq_cm_code_nxt [HQM_NUM_LB_QID-1:0] ;
logic [1:0]                                     p4_atq_cm_code_f [HQM_NUM_LB_QID-1:0] ;

logic [HQM_NUM_LB_QID-1:0]                      p3_atq_qid_avail ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_index_0_nxt ;        // Duplicated for drive, goes to 2 arbiters
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_index_0_f ;          // Duplicated for drive, goes to 2 arbiters
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_index_1_nxt ;        // Duplicated for drive, goes to 2 arbiters
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_index_1_f ;          // Duplicated for drive, goes to 2 arbiters
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_nfull_arb_reqs ;
logic                                           p3_atq_nfull_arb_winner_v ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_nfull_arb_winner ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_empty_arb_reqs ;
logic                                           p3_atq_empty_arb_winner_pre_v ;
logic                                           p3_atq_empty_arb_winner_v ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_empty_arb_winner ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_winner_p1 ;          // wrap ok


logic                                           p3_atq_arb_update ;
logic                                           p3_atq_arb_winner_pre_v ;
logic                                           p3_atq_arb_winner_v ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_atq_arb_winner ;
logic                                           p3_atq_arb_winner_gp ;
logic                                           p3_atq_sch_req ;
lsp_lb_qid_t                                    p3_atq_sch_req_qid ;
logic                                           p3_atq_sch_stall_smon ;
logic                                           p3_atq_sch_start ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p3_atq_sch_start_qid ;
logic                                           p4_atq_sch_v_nxt ;
logic                                           p4_atq_sch_v_f ;
lsp_lb_qid_t                                    p4_atq_sch_qid_nxt ;
lsp_lb_qid_t                                    p4_atq_sch_qid_f ;
logic                                           p4_atq_sch_hold ;

logic [6:0]                                     atq_sel_ap_db_status_pnc ;
logic                                           atq_sel_ap_db_in_ready ;
logic                                           atq_sel_ap_db_in_valid ;
lsp_nalb_sch_atq_t                              atq_sel_ap_db_in_data ;

lsp_nalb_sch_atq_t                              atq_sel_ap_fifo_push_data ;
logic                                           atq_sel_ap_fifo_push ;
logic                                           atq_sel_ap_fifo_afull ;
logic                                           atq_sel_ap_fifo_empty ;
logic                                           atq_sel_ap_fifo_hold ;

logic                                           p2_atq_tot_enq_cnt_upd_v ;
lsp_arch_cnt_t                                  p2_atq_tot_enq_cnt_upd ;
logic [HQM_LSP_ARCH_CNT_WIDTH-1:0]              p2_atq_tot_enq_cnt_p1 ;
logic [1:0]                                     p2_atq_tot_enq_cnt_res_p1 ;
atq_tot_enq_cnt_rmw_pipe_t                      p0_atq_tot_enq_cnt_rmw_pipe_nxt ;
atq_tot_enq_cnt_rmw_pipe_t                      p2_atq_tot_enq_cnt_rmw_pipe_f_pnc ;

atq_tot_enq_cnt_rmw_pipe_t                      p3_atq_tot_enq_cnt_rmw_pipe_f_pnc ;
logic                                           p3_atq_tot_enq_cnt_res_chk_en ;
logic                                           p4_atq_tot_enq_cnt_res_err_nxt ;
logic                                           p4_atq_tot_enq_cnt_res_err_f ;

logic                                           atq_tot_enq_cnt_rmw_pipe_status_nc ;
logic                                           p0_atq_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p0_atq_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p0_atq_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p0_atq_tot_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                           p1_atq_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p1_atq_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]                    p1_atq_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p1_atq_tot_enq_cnt_rmw_pipe_data_f_nc ;         // +2 for residue
logic                                           p2_atq_tot_enq_cnt_rmw_pipe_v_f_nc ;
logic                                           p3_atq_tot_enq_cnt_rmw_pipe_v_f_nc ;

logic                                           atq_fid_cnt_upd_v_nxt ;
logic                                           atq_fid_cnt_upd_v_f ;
logic                                           atq_fid_cnt_upd_last_v_nxt ;
logic                                           atq_fid_cnt_upd_last_v_f ;
logic                                           atq_fid_cnt_upd_val_nxt ;
logic                                           atq_fid_cnt_upd_val_f ;
logic [6:0]                                     atq_fid_cnt_upd_qid_nxt ;
logic [6:0]                                     atq_fid_cnt_upd_qid_f ;

logic                                           atq_stop_atqatm_nxt ;
logic                                           atq_stop_atqatm_f ;
logic                                           atq_stop_atqatm_last_nxt ;
logic                                           atq_stop_atqatm_last_f ;
logic                                           atq_stop_atqatm_change ;

logic [HQM_NUM_LB_QID-1:0]                      p3_atq_qid_en_nxt ;
logic [HQM_NUM_LB_QID-1:0]                      p3_atq_qid_en_f ;

//------------------------------------------------------------------------------------------------
// DIRENQ pipe declarations

logic                                           direnq_input_arb_new_both ;
logic                                           direnq_input_arb_new_either ;
logic [1:0]                                     direnq_input_arb_reqs ;
logic                                           direnq_input_arb_update ;
logic                                           direnq_input_arb_winner_pre_v ;
logic                                           direnq_input_arb_winner_v ;
logic                                           direnq_input_arb_winner ;
logic                                           direnq_input_arb_sch ;
logic                                           direnq_input_arb_pre_enq ;
logic                                           direnq_input_arb_enq ;
logic                                           direnq_input_arb_pre_tok ;
logic                                           direnq_input_arb_tok ;
lsp_dir_qid_t                                   direnq_input_arb_sch_qid ;
logic [2:0]                                     direnq_input_arb_sch_beats ;            // 1..4
logic                                           direnq_input_req_v ;
logic                                           direnq_input_arb_tog_nxt ;
logic                                           direnq_input_arb_tog_f ;

logic                                           p3_direnq_inp_qid_cq_par_err_nxt ;
logic                                           p3_direnq_inp_qid_cq_par_err_f ;

direnq_enq_cnt_rmw_pipe_t                       p0_direnq_enq_cnt_rmw_pipe_nxt ;
direnq_enq_cnt_rmw_pipe_t                       p0_direnq_enq_cnt_rmw_pipe_f_pnc ;
direnq_enq_cnt_rmw_pipe_t                       p1_direnq_enq_cnt_rmw_pipe_f_pnc ;
direnq_enq_cnt_rmw_pipe_t                       p2_direnq_enq_cnt_rmw_pipe_f ;
logic                                           direnq_enq_cnt_rmw_pipe_status ;
lsp_direnq_enq_cnt_t                            p2_direnq_enq_cnt_upd ;
logic                                           p2_direnq_enq_cnt_upd_v ;
direnq_enq_cnt_rmw_pipe_t                       p3_direnq_enq_cnt_rmw_pipe_f_nc ;
logic                                           p3_direnq_enq_cnt_uflow_err_nxt ;
logic                                           p3_direnq_enq_cnt_oflow_err_nxt ;
logic                                           p3_direnq_enq_cnt_uflow_err_f ;
logic                                           p3_direnq_enq_cnt_oflow_err_f ;
logic                                           p3_direnq_enq_cnt_res_err_nxt ;
logic                                           p3_direnq_enq_cnt_res_err_f ;

direnq_dpth_thrsh_rw_pipe_t                     p0_direnq_dpth_thrsh_rw_pipe_nxt ;
direnq_dpth_thrsh_rw_pipe_t                     p2_direnq_dpth_thrsh_rw_pipe_f_pnc ;
logic                                           p2_direnq_dpth_thrsh_par_chk_en ;
logic                                           p2_direnq_dpth_thrsh_par_err_cond ;
logic                                           p3_direnq_dpth_thrsh_par_err_nxt ;
logic                                           p3_direnq_dpth_thrsh_par_err_f ;
logic [1:0]                                     p2_direnq_dpth_thrsh_cm_code ;

logic                                           direnq_dpth_thrsh_rw_pipe_status_nc ;
logic                                           p0_direnq_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p0_direnq_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          p0_direnq_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH+1)-1:0] p0_direnq_dpth_thrsh_rw_pipe_data_f_nc ;        // +1 for parity
logic                                           p1_direnq_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p1_direnq_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          p1_direnq_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH+1)-1:0] p1_direnq_dpth_thrsh_rw_pipe_data_f_nc ;        // +1 for parity
logic                                           p2_direnq_dpth_thrsh_rw_pipe_v_f_nc ;
logic                                           p3_direnq_dpth_thrsh_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p3_direnq_dpth_thrsh_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          p3_direnq_dpth_thrsh_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH+1)-1:0] p3_direnq_dpth_thrsh_rw_pipe_data_f_nc ;        // +1 for parity

lsp_pipe_ctrl_t                                 p0_direnq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p1_direnq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p2_direnq_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p3_direnq_ctrl_pipe ;
logic                                           p4_direnq_ctrl_pipe_en ;

logic                                           p0_direnq_ctrl_pipe_v_nxt ;
logic                                           p0_direnq_ctrl_pipe_v_nxt_gated ;
logic                                           p0_direnq_ctrl_pipe_v_f ;
direnq_ctrl_pipe_t                              p0_direnq_ctrl_pipe_nxt ;
direnq_ctrl_pipe_t                              p0_direnq_ctrl_pipe_f ;

logic                                           p1_direnq_ctrl_pipe_v_f ;
direnq_ctrl_pipe_t                              p1_direnq_ctrl_pipe_nxt ;
direnq_ctrl_pipe_t                              p1_direnq_ctrl_pipe_f ;

logic                                           p2_direnq_ctrl_pipe_v_f ;
direnq_ctrl_pipe_t                              p2_direnq_ctrl_pipe_nxt ;
direnq_ctrl_pipe_t                              p2_direnq_ctrl_pipe_f ;

logic                                           p3_direnq_ctrl_pipe_v_f ;

logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p2_direnq_ctrl_pipe_enq_delta ;
logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]        p2_direnq_ctrl_pipe_sch_delta ;
logic [1:0]                                     p2_direnq_ctrl_pipe_sch_delta_res ;

logic                                           p2_direnq_enq_cnt_upd_ge4 ;

logic [1:0]                                     p2_direnq_enq_cnt_res_p1 ;
logic [1:0]                                     p2_direnq_enq_cnt_res_mn ;
logic                                           p2_direnq_enq_cnt_oflow_cond ;
logic                                           p2_direnq_enq_cnt_uflow_cond ;
logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p2_direnq_enq_cnt_p1 ;
logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p2_direnq_enq_cnt_mn ;
logic                                           p2_direnq_enq_cnt_p1_carry ;
logic                                           p2_direnq_enq_cnt_mn_borrow ;
logic                                           p2_direnq_enq_cnt_res_chk_en ;
logic                                           p2_direnq_enq_cnt_res_err_cond ;

logic                                           p0_direnq_inp_tok_cnt_res_chk_en ;
logic                                           p0_direnq_inp_tok_cnt_res_err_cond ;
logic                                           p1_direnq_inp_tok_cnt_res_err_nxt ;
logic                                           p1_direnq_inp_tok_cnt_res_err_f ;

direnq_tok_cnt_rmw_pipe_t                       p0_direnq_tok_cnt_rmw_pipe_nxt ;
direnq_tok_cnt_rmw_pipe_t                       p0_direnq_tok_cnt_rmw_pipe_f_pnc ;
direnq_tok_cnt_rmw_pipe_t                       p1_direnq_tok_cnt_rmw_pipe_f_pnc ;
direnq_tok_cnt_rmw_pipe_t                       p2_direnq_tok_cnt_rmw_pipe_f ;
lsp_direnq_tok_cnt_t                            p2_direnq_tok_cnt_upd ;
logic                                           p2_direnq_tok_cnt_upd_v ;
direnq_tok_cnt_rmw_pipe_t                       p3_direnq_tok_cnt_rmw_pipe_f_pnc ;
logic                                           p2_direnq_tok_cnt_res_chk_en ;
logic                                           p2_direnq_tok_cnt_res_err_cond ;
logic                                           p3_direnq_tok_cnt_uflow_err_nxt ;
logic                                           p3_direnq_tok_cnt_oflow_err_nxt ;
logic                                           p3_direnq_tok_cnt_uflow_err_f ;
logic [7:0]                                     p3_direnq_tok_cnt_uflow_err_rid ;
logic                                           p3_direnq_tok_cnt_oflow_err_f ;
logic                                           p3_direnq_tok_cnt_res_err_nxt ;
logic                                           p3_direnq_tok_cnt_res_err_f ;

logic                                           direnq_tok_cnt_rmw_pipe_status_nc ;
logic                                           p0_direnq_tok_cnt_rmw_pipe_v_f_nc ;
logic                                           p1_direnq_tok_cnt_rmw_pipe_v_f_nc ;
logic                                           p2_direnq_tok_cnt_rmw_pipe_v_f_nc ;
logic                                           p3_direnq_tok_cnt_rmw_pipe_v_f_nc ;

logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]        p2_direnq_tok_limit ;
logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH:0]          p2_direnq_tok_cnt_upd_space_sub ;               // extra bit for borrow
logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]        p2_direnq_tok_cnt_upd_space ;
logic                                           p2_direnq_tok_cnt_upd_space_ge4 ;
logic                                           p2_direnq_tok_cnt_upd_gt_0 ;
logic                                           p2_direnq_tok_lim_par_chk_en ;
logic                                           p2_direnq_tok_lim_par_err_cond ;

direnq_tok_lim_rw_pipe_t                        p0_direnq_tok_lim_rw_pipe_nxt ;
direnq_tok_lim_rw_pipe_t                        p2_direnq_tok_lim_rw_pipe_f_pnc ;
logic                                           p3_direnq_tok_lim_par_err_nxt ;
logic                                           p3_direnq_tok_lim_par_err_f ;

logic                                           direnq_tok_lim_rw_pipe_status_nc ;
logic                                           p0_direnq_tok_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p0_direnq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]                    p0_direnq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_TOK_LIM_SEL_WIDTH+4)-1:0]        p0_direnq_tok_lim_rw_pipe_data_f_nc ;   // +4 for 2 control, 1 spare, 1 parity
logic                                           p1_direnq_tok_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p1_direnq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]                    p1_direnq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_TOK_LIM_SEL_WIDTH+4)-1:0]        p1_direnq_tok_lim_rw_pipe_data_f_nc ;   // +4 for 2 control, 1 spare, 1 parity
logic                                           p2_direnq_tok_lim_rw_pipe_v_f_nc ;
logic                                           p3_direnq_tok_lim_rw_pipe_v_f_nc ;
aw_rwpipe_cmd_t                                 p3_direnq_tok_lim_rw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]                    p3_direnq_tok_lim_rw_pipe_addr_f_nc ;
logic [(HQM_LSP_DIRENQ_TOK_LIM_SEL_WIDTH+4)-1:0]        p3_direnq_tok_lim_rw_pipe_data_f_nc ;   // +4 for 2 control, 1 spare, 1 parity

logic [1:0]                                     p2_direnq_tok_cnt_res_pn ;
logic [1:0]                                     p2_direnq_tok_cnt_res_mn ;
logic                                           p2_direnq_tok_cnt_oflow_cond ;
logic                                           p2_direnq_tok_cnt_uflow_cond ;
logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]        p2_direnq_tok_cnt_pn ;
logic [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]        p2_direnq_tok_cnt_mn ;
logic                                           p2_direnq_tok_cnt_pn_carry ;
logic                                           p2_direnq_tok_cnt_mn_borrow ;

logic [1:0]                                     p3_direnq_cm_code_nxt [HQM_NUM_DIR_QID-1:0] ;
logic [1:0]                                     p3_direnq_cm_code_f [HQM_NUM_DIR_QID-1:0] ;
logic [HQM_NUM_DIR_CQ-1:0]                      p3_direnq_wp_en ;
logic [1:0]                                     p3_direnq_wp_nxt [HQM_NUM_DIR_CQ-1:0] ;
logic [1:0]                                     p3_direnq_wp_f [HQM_NUM_DIR_CQ-1:0] ;
logic [HQM_NUM_DIR_CQ-1:0]                      cfg_dir_tok_lim_disab_opt_nxt ;
logic [HQM_NUM_DIR_CQ-1:0]                      cfg_dir_tok_lim_disab_opt_f ;           // Need copy of RAM in reg - can't do RAM read on sch

logic   [HQM_NUM_DIR_CQ-1:0]                    p3_direnq_sch_hit ;
logic   [HQM_NUM_DIR_CQ-1:0]                    p3_direnq_p2_enq_hit ;
logic   [HQM_NUM_DIR_CQ-1:0]                    p3_direnq_p2_tok_hit ;
direnq_arb_stat_t                               p3_direnq_arb_stat_nxt [HQM_NUM_DIR_QID-1:0] ;
direnq_arb_stat_t                               p3_direnq_arb_stat_f [HQM_NUM_DIR_QID-1:0] ;

logic                                           p3_direnq_fill_in_progress ;

logic   [HQM_NUM_DIR_CQ-1:0]                    p3_direnq_tok_cnt_v_nxt ;
logic   [HQM_NUM_DIR_CQ-1:0]                    p3_direnq_tok_cnt_v_f ;

logic   [HQM_NUM_DIR_QID-1:0]                   p3_direnq_arb_reqs ;
logic                                           p3_direnq_arb_update ;
logic                                           p3_direnq_arb_winner_pre_v ;
logic                                           p3_direnq_arb_winner_v ;
logic   [HQM_NUM_DIR_QIDB2-1:0]                 p3_direnq_arb_winner ;

lsp_dir_qid_t                                   p3_direnq_arb_winner_qid ;

logic [2:0]                                     p3_direnq_arb_winner_qid_v ;
logic [2:0]                                     p3_direnq_arb_winner_cq_avail ;
logic [1:0]                                     p3_direnq_arb_winner_cm_code ;
logic [1:0]                                     p3_direnq_arb_winner_wp ;
logic                                           p3_direnq_arb_winner_disab_opt ;

logic [1:0]                                     p3_direnq_rem_beats ;                   // Remaining beats, after this clock
logic [1:0]                                     p3_direnq_rem_beats_m1 ;

logic [1:0]                                     p4_direnq_sch_rem_beats_nxt ;
logic [2:0]                                     p4_direnq_sch_qid_v_nxt ;
logic [2:0]                                     p4_direnq_sch_cq_avail_nxt ;
logic [1:0]                                     p4_direnq_sch_wp_nxt ;
lsp_dir_qid_t                                   p4_direnq_sch_qid_nxt ;
logic [1:0]                                     p4_direnq_sch_cm_code_nxt ;
logic                                           p4_direnq_sch_disab_opt_nxt ;
logic                                           p4_direnq_sch_first_beat_nxt ;
logic                                           p4_direnq_sch_first_clock_nxt ;

logic [1:0]                                     p4_direnq_sch_rem_beats_f ;
logic [2:0]                                     p4_direnq_sch_qid_v_f ;
logic [2:0]                                     p4_direnq_sch_cq_avail_f ;
logic [1:0]                                     p4_direnq_sch_wp_f ;
lsp_dir_qid_t                                   p4_direnq_sch_qid_f ;
logic [1:0]                                     p4_direnq_sch_cm_code_f ;
logic                                           p4_direnq_sch_disab_opt_f ;
logic                                           p4_direnq_sch_first_beat_f ;
logic                                           p4_direnq_sch_first_clock_f ;

logic [1:0]                                     p4_direnq_calc_rem_beats_enab ;
logic [1:0]                                     p4_direnq_calc_rem_beats ;
logic [1:0]                                     p4_direnq_sch_rem_beats_m1 ;

logic                                           p3_direnq_sch_req ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          p3_direnq_sch_req_qid ;
logic                                           p3_direnq_sch_start ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          p3_direnq_sch_start_qid ;
logic                                           p3_direnq_sch_out ;
logic [HQM_NUM_DIR_QIDB2-1:0]                   p3_direnq_sch_out_qid ;
logic [1:0]                                     p3_direnq_sch_out_cm_code ;
logic                                           p4_direnq_sch_v_nxt ;
logic                                           p4_direnq_sch_v_f ;

logic                                           p4_direnq_sch_hold ;

logic                                           p2_direnq_inp_enq_qid_p ;
logic                                           p2_direnq_inp_tok_cq_p ;
logic                                           p2_direnq_inp_enq_qid_par_chk_en ;
logic                                           p2_direnq_inp_tok_cq_par_chk_en ;
logic                                           p2_direnq_inp_enq_qid_par_err_cond ;
logic                                           p2_direnq_inp_tok_cq_par_err_cond ;
logic                                           p2_direnq_inp_qid_cq_par_err_cond ;

logic                                           p2_direnq_tot_enq_cnt_upd_v ;
lsp_arch_cnt_t                                  p2_direnq_tot_enq_cnt_upd ;
logic [HQM_LSP_ARCH_CNT_WIDTH-1:0]              p2_direnq_tot_enq_cnt_p1 ;
logic [1:0]                                     p2_direnq_tot_enq_cnt_res_p1 ;
direnq_tot_enq_cnt_rmw_pipe_t                   p0_direnq_tot_enq_cnt_rmw_pipe_nxt ;
direnq_tot_enq_cnt_rmw_pipe_t                   p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc ;

direnq_tot_enq_cnt_rmw_pipe_t                   p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc ;
logic                                           p3_direnq_tot_enq_cnt_res_chk_en ;
logic                                           p4_direnq_tot_enq_cnt_res_err_nxt ;
logic                                           p4_direnq_tot_enq_cnt_res_err_f ;

logic                                           direnq_tot_enq_cnt_rmw_pipe_status_nc ;
logic                                           p0_direnq_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p0_direnq_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]                   p0_direnq_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p0_direnq_tot_enq_cnt_rmw_pipe_data_f_nc ;              // +2 for residue
logic                                           p1_direnq_tot_enq_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p1_direnq_tot_enq_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]                   p1_direnq_tot_enq_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p1_direnq_tot_enq_cnt_rmw_pipe_data_f_nc ;              // +2 for residue
logic                                           p2_direnq_tot_enq_cnt_rmw_pipe_v_f_nc ;
logic                                           p3_direnq_tot_enq_cnt_rmw_pipe_v_f_nc ;

logic                                           p2_direnq_tot_sch_cnt_upd_v ;
lsp_arch_cnt_t                                  p2_direnq_tot_sch_cnt_upd ;
logic [HQM_LSP_ARCH_CNT_WIDTH-1:0]              p2_direnq_tot_sch_cnt_pn ;
logic [1:0]                                     p2_direnq_tot_sch_cnt_res_pn ;
direnq_tot_sch_cnt_rmw_pipe_t                   p0_direnq_tot_sch_cnt_rmw_pipe_nxt ;
direnq_tot_sch_cnt_rmw_pipe_t                   p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc ;

direnq_tot_sch_cnt_rmw_pipe_t                   p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc ;
logic                                           p3_direnq_tot_sch_cnt_res_chk_en ;
logic                                           p4_direnq_tot_sch_cnt_res_err_nxt ;
logic                                           p4_direnq_tot_sch_cnt_res_err_f ;

logic                                           direnq_tot_sch_cnt_rmw_pipe_status_nc ;
logic                                           p0_direnq_tot_sch_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p0_direnq_tot_sch_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]                    p0_direnq_tot_sch_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p0_direnq_tot_sch_cnt_rmw_pipe_data_f_nc ;              // +2 for residue
logic                                           p1_direnq_tot_sch_cnt_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p1_direnq_tot_sch_cnt_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]                    p1_direnq_tot_sch_cnt_rmw_pipe_addr_f_nc ;
logic [(HQM_LSP_ARCH_CNT_WIDTH+2)-1:0]          p1_direnq_tot_sch_cnt_rmw_pipe_data_f_nc ;              // +2 for residue
logic                                           p2_direnq_tot_sch_cnt_rmw_pipe_v_f_nc ;
logic                                           p3_direnq_tot_sch_cnt_rmw_pipe_v_f_nc ;

logic                                           p2_direnq_enq_cnt_gt_max_depth ;
logic                                           p2_direnq_max_enq_depth_upd_v ;
logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p2_direnq_max_enq_depth_upd ;
direnq_max_enq_depth_rmw_pipe_t                 p0_direnq_max_enq_depth_rmw_pipe_nxt ;
direnq_max_enq_depth_rmw_pipe_t                 p2_direnq_max_enq_depth_rmw_pipe_f ;
direnq_max_enq_depth_rmw_pipe_t                 p3_direnq_max_enq_depth_rmw_pipe_f_nc ;

logic                                           direnq_max_enq_depth_rmw_pipe_status_nc ;
logic                                           p0_direnq_max_enq_depth_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p0_direnq_max_enq_depth_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]                   p0_direnq_max_enq_depth_rmw_pipe_addr_f_nc ;
logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p0_direnq_max_enq_depth_rmw_pipe_data_f_nc ;
logic                                           p1_direnq_max_enq_depth_rmw_pipe_v_f_nc ;
aw_rmwpipe_cmd_t                                p1_direnq_max_enq_depth_rmw_pipe_rw_f_nc ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]                   p1_direnq_max_enq_depth_rmw_pipe_addr_f_nc ;
logic [HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0]        p1_direnq_max_enq_depth_rmw_pipe_data_f_nc ;
logic                                           p2_direnq_max_enq_depth_rmw_pipe_v_f_nc ;
logic                                           p3_direnq_max_enq_depth_rmw_pipe_v_f_nc ;

//------------------------------------------------------------------------------------------------
// LBRPL pipe declarations
logic [1:0]                                     lbrpl_input_arb_reqs ;
logic                                           lbrpl_input_arb_winner_pre_v ;
logic                                           lbrpl_input_arb_winner_v ;
logic                                           lbrpl_input_arb_winner ;
logic                                           lbrpl_input_arb_sch ;
lsp_lb_qid_t                                    lbrpl_input_arb_sch_qid ;
logic                                           lbrpl_input_arb_enq ;

lsp_pipe_ctrl_t                                 p0_lbrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p1_lbrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p2_lbrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p3_lbrpl_ctrl_pipe ;

logic                                           p0_lbrpl_ctrl_pipe_v_nxt ;
logic                                           p0_lbrpl_ctrl_pipe_v_nxt_gated ;
logic                                           p0_lbrpl_ctrl_pipe_v_f ;
lbrpl_ctrl_pipe_t                               p0_lbrpl_ctrl_pipe_nxt ;
lbrpl_ctrl_pipe_t                               p0_lbrpl_ctrl_pipe_f ;

logic                                           p1_lbrpl_ctrl_pipe_v_f ;
lbrpl_ctrl_pipe_t                               p1_lbrpl_ctrl_pipe_nxt ;
lbrpl_ctrl_pipe_t                               p1_lbrpl_ctrl_pipe_f ;

logic                                           p2_lbrpl_ctrl_pipe_v_f ;
lbrpl_ctrl_pipe_t                               p2_lbrpl_ctrl_pipe_nxt ;
lbrpl_ctrl_pipe_t                               p2_lbrpl_ctrl_pipe_f ;

logic                                           p3_lbrpl_ctrl_pipe_v_f ;

logic                                           lbrpl_input_req_v ;

logic                                           p2_lbrpl_inp_qid_par_chk_en ;
logic                                           p2_lbrpl_inp_qid_par_err_cond ;
logic                                           p3_lbrpl_inp_qid_par_err_nxt ;
logic                                           p3_lbrpl_inp_qid_par_err_f ;
logic                                           p0_lbrpl_inp_frag_cnt_res_chk_en ;
logic                                           p0_lbrpl_inp_frag_cnt_res_err_cond ;
logic                                           p1_lbrpl_inp_frag_cnt_res_err_nxt ;
logic                                           p1_lbrpl_inp_frag_cnt_res_err_f ;

logic                                           p2_lbrpl_enq_cnt_upd_v ;
lsp_lbrpl_enq_cnt_t                             p2_lbrpl_enq_cnt_upd ;
logic [HQM_LSP_LBRPL_ENQ_CNT_WIDTH-1:0]         p2_lbrpl_enq_cnt_pn ;
logic [HQM_LSP_LBRPL_ENQ_CNT_WIDTH-1:0]         p2_lbrpl_enq_cnt_m1 ;
logic                                           p2_lbrpl_enq_cnt_upd_gt0 ;
logic [1:0]                                     p2_lbrpl_enq_cnt_res_pn ;
logic [1:0]                                     p2_lbrpl_enq_cnt_res_m1 ;
logic                                           p2_lbrpl_enq_cnt_pn_carry ;
logic                                           p2_lbrpl_enq_cnt_m1_borrow ;
logic                                           p2_lbrpl_enq_cnt_oflow_cond ;
logic                                           p2_lbrpl_enq_cnt_uflow_cond ;
logic                                           lbrpl_enq_cnt_rmw_pipe_status ;
lbrpl_enq_cnt_rmw_pipe_t                        p0_lbrpl_enq_cnt_rmw_pipe_nxt ;
lbrpl_enq_cnt_rmw_pipe_t                        p0_lbrpl_enq_cnt_rmw_pipe_f_pnc ;
lbrpl_enq_cnt_rmw_pipe_t                        p1_lbrpl_enq_cnt_rmw_pipe_f_pnc ;
lbrpl_enq_cnt_rmw_pipe_t                        p2_lbrpl_enq_cnt_rmw_pipe_f ;
lbrpl_enq_cnt_rmw_pipe_t                        p3_lbrpl_enq_cnt_rmw_pipe_f_nc ;
logic                                           p2_lbrpl_enq_cnt_res_chk_en ;
logic                                           p3_lbrpl_enq_cnt_uflow_err_nxt ;
logic                                           p3_lbrpl_enq_cnt_oflow_err_nxt ;
logic                                           p3_lbrpl_enq_cnt_uflow_err_f ;
logic                                           p3_lbrpl_enq_cnt_oflow_err_f ;
logic                                           p3_lbrpl_enq_cnt_res_err ;
logic                                           p3_lbrpl_enq_cnt_res_chk_en_nxt ;
logic                                           p3_lbrpl_enq_cnt_res_chk_en_f ;
lsp_lbrpl_enq_cnt_t                             p3_lbrpl_enq_cnt_nxt ;
lsp_lbrpl_enq_cnt_t                             p3_lbrpl_enq_cnt_f ;

logic [HQM_NUM_LB_QID-1:0]                      p3_lbrpl_sch_hit ;

logic [HQM_NUM_LB_QID-1:0]                      p3_lbrpl_p2_enq_hit ;

rpl_arb_stat_t                                  p3_lbrpl_arb_stat_nxt [HQM_NUM_LB_QID-1:0] ;
rpl_arb_stat_t                                  p3_lbrpl_arb_stat_f [HQM_NUM_LB_QID-1:0] ;

logic [HQM_NUM_LB_QID-1:0]                      p3_lbrpl_arb_reqs ;
logic                                           p3_lbrpl_arb_update ;
logic                                           p3_lbrpl_arb_winner_pre_v ;
logic                                           p3_lbrpl_arb_winner_v ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_lbrpl_arb_winner ;
logic                                           p3_lbrpl_arb_winner_gp ;
logic                                           p3_lbrpl_sch_req ;
lsp_lb_qid_t                                    p3_lbrpl_sch_req_qid ;
logic                                           p3_lbrpl_sch_stall_smon ;
logic                                           p3_lbrpl_sch_start ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p3_lbrpl_sch_start_qid ;
logic                                           p4_lbrpl_sch_v_nxt ;
logic                                           p4_lbrpl_sch_v_f ;
lsp_lb_qid_t                                    p4_lbrpl_sch_qid_nxt ;
lsp_lb_qid_t                                    p4_lbrpl_sch_qid_f ;
logic                                           p4_lbrpl_sch_hold ;

logic [6:0]                                     rpl_ldb_nalb_db_status_pnc ;
logic                                           rpl_ldb_nalb_db_in_ready ;
logic                                           rpl_ldb_nalb_db_in_valid ;
lsp_nalb_sch_rorply_t                           rpl_ldb_nalb_db_in_data ;

lsp_nalb_sch_rorply_t                           rpl_ldb_nalb_fifo_push_data ;
logic                                           rpl_ldb_nalb_fifo_push ;
logic                                           rpl_ldb_nalb_fifo_afull ;
logic                                           rpl_ldb_nalb_fifo_empty ;
logic                                           rpl_ldb_nalb_fifo_hold ;

//------------------------------------------------------------------------------------------------
// DIRRPL pipe declarations
logic [1:0]                                     dirrpl_input_arb_reqs ;
logic                                           dirrpl_input_arb_winner_pre_v ;
logic                                           dirrpl_input_arb_winner_v ;
logic                                           dirrpl_input_arb_winner ;
logic                                           dirrpl_input_arb_sch ;
lsp_dir_qid_t                                   dirrpl_input_arb_sch_qid ;
logic                                           dirrpl_input_arb_enq ;

lsp_pipe_ctrl_t                                 p0_dirrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p1_dirrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p2_dirrpl_ctrl_pipe ;
lsp_pipe_ctrl_t                                 p3_dirrpl_ctrl_pipe ;

logic                                           p0_dirrpl_ctrl_pipe_v_nxt ;
logic                                           p0_dirrpl_ctrl_pipe_v_nxt_gated ;
logic                                           p0_dirrpl_ctrl_pipe_v_f ;
dirrpl_ctrl_pipe_t                              p0_dirrpl_ctrl_pipe_nxt ;
dirrpl_ctrl_pipe_t                              p0_dirrpl_ctrl_pipe_f ;

logic                                           p1_dirrpl_ctrl_pipe_v_f ;
dirrpl_ctrl_pipe_t                              p1_dirrpl_ctrl_pipe_nxt ;
dirrpl_ctrl_pipe_t                              p1_dirrpl_ctrl_pipe_f ;

logic                                           p2_dirrpl_ctrl_pipe_v_f ;
dirrpl_ctrl_pipe_t                              p2_dirrpl_ctrl_pipe_nxt ;
dirrpl_ctrl_pipe_t                              p2_dirrpl_ctrl_pipe_f ;

logic                                           p3_dirrpl_ctrl_pipe_v_f ;

logic                                           dirrpl_input_req_v ;

logic                                           p0_dirrpl_inp_frag_cnt_res_chk_en ;
logic                                           p0_dirrpl_inp_frag_cnt_res_err_cond ;
logic                                           p1_dirrpl_inp_frag_cnt_res_err_nxt ;
logic                                           p1_dirrpl_inp_frag_cnt_res_err_f ;
logic                                           p2_dirrpl_inp_qid_par_chk_en ;
logic                                           p2_dirrpl_inp_qid_par_err_cond ;
logic                                           p3_dirrpl_inp_qid_par_err_nxt ;
logic                                           p3_dirrpl_inp_qid_par_err_f ;

logic                                           p2_dirrpl_enq_cnt_upd_v ;
lsp_dirrpl_enq_cnt_t                            p2_dirrpl_enq_cnt_upd ;
logic [HQM_LSP_DIRRPL_ENQ_CNT_WIDTH-1:0]        p2_dirrpl_enq_cnt_pn ;
logic [HQM_LSP_DIRRPL_ENQ_CNT_WIDTH-1:0]        p2_dirrpl_enq_cnt_m1 ;
logic                                           p2_dirrpl_enq_cnt_upd_gt0 ;
logic [1:0]                                     p2_dirrpl_enq_cnt_res_pn ;
logic [1:0]                                     p2_dirrpl_enq_cnt_res_m1 ;
logic                                           p2_dirrpl_enq_cnt_pn_carry ;
logic                                           p2_dirrpl_enq_cnt_m1_borrow ;
logic                                           p2_dirrpl_enq_cnt_oflow_cond ;
logic                                           p2_dirrpl_enq_cnt_uflow_cond ;
logic                                           dirrpl_enq_cnt_rmw_pipe_status ;
dirrpl_enq_cnt_rmw_pipe_t                       p0_dirrpl_enq_cnt_rmw_pipe_nxt ;
dirrpl_enq_cnt_rmw_pipe_t                       p0_dirrpl_enq_cnt_rmw_pipe_f_pnc ;
dirrpl_enq_cnt_rmw_pipe_t                       p1_dirrpl_enq_cnt_rmw_pipe_f_pnc ;
dirrpl_enq_cnt_rmw_pipe_t                       p2_dirrpl_enq_cnt_rmw_pipe_f ;
dirrpl_enq_cnt_rmw_pipe_t                       p3_dirrpl_enq_cnt_rmw_pipe_f_nc ;
logic                                           p2_dirrpl_enq_cnt_res_chk_en ;
logic                                           p3_dirrpl_enq_cnt_uflow_err_nxt ;
logic                                           p3_dirrpl_enq_cnt_oflow_err_nxt ;
logic                                           p3_dirrpl_enq_cnt_uflow_err_f ;
logic                                           p3_dirrpl_enq_cnt_oflow_err_f ;
logic                                           p3_dirrpl_enq_cnt_res_err ;
logic                                           p3_dirrpl_enq_cnt_res_chk_en_nxt ;
logic                                           p3_dirrpl_enq_cnt_res_chk_en_f ;
lsp_dirrpl_enq_cnt_t                            p3_dirrpl_enq_cnt_nxt ;
lsp_dirrpl_enq_cnt_t                            p3_dirrpl_enq_cnt_f ;

logic [HQM_NUM_LB_QID-1:0]                      p3_dirrpl_sch_hit ;

logic [HQM_NUM_LB_QID-1:0]                      p3_dirrpl_p2_enq_hit ;

rpl_arb_stat_t                                  p3_dirrpl_arb_stat_nxt [HQM_NUM_LB_QID-1:0] ;
rpl_arb_stat_t                                  p3_dirrpl_arb_stat_f [HQM_NUM_LB_QID-1:0] ;

logic [HQM_NUM_LB_QID-1:0]                      p3_dirrpl_arb_reqs ;
logic                                           p3_dirrpl_arb_update ;
logic                                           p3_dirrpl_arb_winner_pre_v ;
logic                                           p3_dirrpl_arb_winner_v ;
logic [HQM_NUM_LB_QIDB2-1:0]                    p3_dirrpl_arb_winner ;
logic                                           p3_dirrpl_arb_winner_gp ;
logic                                           p3_dirrpl_sch_req ;
lsp_dir_qid_t                                   p3_dirrpl_sch_req_qid ;
logic                                           p3_dirrpl_sch_stall_smon ;
logic                                           p3_dirrpl_sch_start ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           p3_dirrpl_sch_start_qid ;
logic                                           p4_dirrpl_sch_v_nxt ;
logic                                           p4_dirrpl_sch_v_f ;
lsp_dir_qid_t                                   p4_dirrpl_sch_qid_nxt ;
lsp_dir_qid_t                                   p4_dirrpl_sch_qid_f ;
logic                                           p4_dirrpl_sch_hold ;

logic [6:0]                                     rpl_dir_dp_db_status_pnc ;
logic                                           rpl_dir_dp_db_in_ready ;
logic                                           rpl_dir_dp_db_in_valid ;
lsp_dp_sch_rorply_t                             rpl_dir_dp_db_in_data ;

lsp_dp_sch_rorply_t                             rpl_dir_dp_fifo_push_data ;
logic                                           rpl_dir_dp_fifo_push ;
logic                                           rpl_dir_dp_fifo_afull ;
logic                                           rpl_dir_dp_fifo_empty ;
logic                                           rpl_dir_dp_fifo_hold ;

//------------------------------------------------------------------------------------------------
// Error logic declarations
logic                                           lba_cq2qid_rw_pipe_err_nxt ;
logic                                           lba_cq_tok_cnt_rmw_pipe_err_nxt ;
logic                                           lba_qid2cqidix_rw_pipe_err_nxt;
logic                                           atq_enq_cnt_rmw_pipe_err_nxt ;
logic                                           direnq_enq_cnt_rmw_pipe_err_nxt ;
logic                                           lbrpl_enq_cnt_rmw_pipe_err_nxt ;
logic                                           dirrpl_enq_cnt_rmw_pipe_err_nxt ;
logic                                           lba_arbindex_rmw_pipe_err_nxt ;
logic                                           lbwu_cq_wu_cnt_rmw_pipe_err_nxt ;

logic                                           lba_cq2qid_rw_pipe_err_f ;
logic                                           lba_cq_tok_cnt_rmw_pipe_err_f ;
logic                                           lba_qid2cqidix_rw_pipe_err_f ;
logic                                           atq_enq_cnt_rmw_pipe_err_f ;
logic                                           direnq_enq_cnt_rmw_pipe_err_f ;
logic                                           lbrpl_enq_cnt_rmw_pipe_err_f ;
logic                                           dirrpl_enq_cnt_rmw_pipe_err_f ;
logic                                           lba_arbindex_rmw_pipe_err_f ;
logic                                           lbwu_cq_wu_cnt_rmw_pipe_err_f ;

logic                                           atq_fid_if_lim_err_nxt ;
logic                                           atq_fid_if_lim_err_f ;
logic                                           atq_fid_if_lim_err_reported_nxt ;
logic                                           atq_fid_if_lim_err_reported_f ;
logic                                           atq_fid_if_lim_err_v ;

logic                                           atq_tot_act_lim_err_nxt ;
logic                                           atq_tot_act_lim_err_f ;
logic                                           atq_tot_act_lim_err_reported_nxt ;
logic                                           atq_tot_act_lim_err_reported_f ;
logic                                           atq_tot_act_lim_err_v ;

//------------------------------------------------------------------------------------------------
// Memory declarations

logic                                   nalb_sel_nalb_fifo_push ;
logic                                   nalb_sel_nalb_fifo_pop ;
lsp_nalb_sch_unoord_t                   nalb_sel_nalb_fifo_push_data ;
lsp_nalb_sch_unoord_t                   nalb_sel_nalb_fifo_pop_data ;
logic                                   nalb_sel_nalb_fifo_pop_data_v ;
logic                                   nalb_sel_nalb_fifo_afull ;
logic                                   nalb_sel_nalb_fifo_full_nc ;
logic                                   nalb_sel_nalb_fifo_empty ;
logic                                   nalb_sel_nalb_fifo_of ;
logic                                   nalb_sel_nalb_fifo_uf ;
logic [HQM_LSP_NALB_SEL_NALB_FIFO_WMWIDTH-1:0]  nalb_sel_nalb_fifo_hwm ;
logic [31:0]                            nalb_sel_nalb_fifo_status_pnc ;

//------------------------------------------------------------------------------------------------
// AP <> LSP internal interfaces

logic                                   lsp_ap_atm_v ;
logic                                   lsp_ap_atm_ready ;
lsp_ap_atm_t                            lsp_ap_atm_data ;
logic                                   ap_lsp_freeze ;
logic                                   p4_lsp_ap_atm_sched_p ;

logic [1:0]                             credit_fifo_ap_aqed_dec_sch ;
logic                                   credit_fifo_ap_aqed_dec_cmp ;

// Previously used by LSP, still very useful for debug / accounting - used by "_inst" file
logic                                   ap_lsp_enq_v_nc ;
ap_lsp_enq_t                            ap_lsp_enq_data_nc ;

logic                                   ap_lsp_cmd_v ;
logic [1:0]                             ap_lsp_cmd ;

logic [5:0]                             ap_lsp_cq ;
logic                                   ap_lsp_qidix_msb ;
logic [2:0]                             ap_lsp_qidix ;
logic [6:0]                             ap_lsp_qid_nc ;                 // Used in assert
logic [511:0]                           ap_lsp_qid2cqqidix ;

logic                                   ap_lsp_haswork_rlst_v ;
logic                                   ap_lsp_haswork_rlst_func ;

logic                                   ap_lsp_haswork_slst_v ;
logic                                   ap_lsp_haswork_slst_func ;

logic                                   ap_lsp_cmpblast_v ;

logic                                   ap_lsp_dec_fid_cnt_v_nc ;       // Used in assert

// Derived signals
logic [8:0]                             ap_lsp_cq_qidix ;
logic                                   ap_lsp_cmpblast_v_hit ;
logic [15:0]                            ap_lsp_qidixv ;
logic                                   ap_lsp_unblast_slst_v ;
logic                                   ap_lsp_unblast_rlst_v ;
logic                                   ap_lsp_unblast_cmpblast ;
logic                                   ap_lsp_cmd_cmp ;

//------------------------------------------------------------------------------------------------
// smon declarations
logic                                           smon_interrupt_nc ;
logic                                           smon_enabled ;
logic                                           smon_enabled_any ;

logic [HQM_LSP_SMON0_WIDTH-1:0]                 smon0_v ;
logic [(HQM_LSP_SMON0_WIDTH*32)-1:0]            smon0_value ;
logic [(HQM_LSP_SMON0_WIDTH*32)-1:0]            smon0_comp ;

logic                                           smon_qed_lsp_deq_v ;
logic                                           smon_qed_lsp_deq_data_parity_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_qed_lsp_deq_data_cq ;
logic [1:0]                                     smon_qed_lsp_deq_data_qe_wt_nc ;
logic                                           smon_aqed_lsp_deq_v ;
logic                                           smon_aqed_lsp_deq_data_parity_nc ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_aqed_lsp_deq_data_cq ;
logic [1:0]                                     smon_aqed_lsp_deq_data_qe_wt_nc ;

logic                                           smon_lsp_dp_sch_dir_v_nxt ;
logic                                           smon_lsp_dp_sch_dir_rdy_nxt ;
logic [1:0]                                     smon_lsp_dp_sch_dir_cm_nxt ;
logic [1:0]                                     smon_lsp_dp_sch_dir_wbo_nxt ;
logic [7:0]                                     smon_lsp_dp_sch_dir_cq_nxt ;
logic                                           smon_lsp_ap_atm_taken_nxt ;
logic                                           smon_lsp_ap_atm_stall_nxt ;
enum_cmd_lsp_ap_atm_t                           smon_lsp_ap_atm_cmd_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_lsp_ap_atm_cq_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_lsp_ap_atm_qid_nxt ;
logic [HQM_LSP_ARCH_NUM_FIDB2-1:0]              smon_lsp_ap_atm_fid_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_lsp_nalb_sch_unoord_cq_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_lsp_nalb_sch_unoord_qid_nxt ;
logic                                           smon_atq_sel_ap_stall_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_atq_sel_ap_qid_nxt ;
logic                                           smon_rpl_dir_dp_stall_nxt ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          smon_rpl_dir_dp_qid_nxt ;
logic                                           smon_rpl_ldb_nalb_stall_nxt ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_rpl_ldb_nalb_qid_nxt ;
logic [6:0]                                     smon_dp_lsp_enq_dir_data_qid_nxt ;
logic                                           smon_chp_lsp_token_data_is_ldb_nxt ;
logic [7:0]                                     smon_chp_lsp_token_data_cq_nxt ;
logic [12:0]                                    smon_chp_lsp_token_data_count_nxt ;
hqm_pkg::qtype_t                                smon_nalb_lsp_enq_lb_data_qtype_nxt ;
logic [6:0]                                     smon_nalb_lsp_enq_lb_data_qid_nxt ;
logic [6:0]                                     smon_chp_lsp_cmp_data_qid_nxt ;
logic [7:0]                                     smon_chp_lsp_cmp_data_cq_nxt ;
hqm_pkg::qtype_t                                smon_chp_lsp_cmp_data_qtype_nxt ;
logic [11:0]                                    smon_chp_lsp_cmp_data_fid_nxt ;
logic [6:0]                                     smon_rop_lsp_reordercmp_data_qid_nxt ;
logic [7:0]                                     smon_rop_lsp_reordercmp_data_cq_nxt ;
logic [6:0]                                     smon_dp_lsp_enq_rorply_data_qid_nxt ;
logic [6:0]                                     smon_nalb_lsp_enq_rorply_data_qid_nxt ;
logic [12:0]                                    smon_dp_lsp_enq_rorply_data_frag_cnt_nxt ;
logic [14:0]                                    smon_nalb_lsp_enq_rorply_data_frag_cnt_nxt ;
logic [5:0]                                     smon_qed_lsp_deq_data_cq_nxt ;
logic [5:0]                                     smon_aqed_lsp_deq_data_cq_nxt ;

logic                                           smon_chp_lsp_token_v_nxt ;
logic                                           smon_chp_lsp_cmp_v_nxt ;
logic                                           smon_rop_lsp_reordercmp_v_nxt ;
logic                                           smon_nalb_lsp_enq_lb_v_nxt ;
logic                                           smon_dp_lsp_enq_dir_v_nxt ;
logic                                           smon_dp_lsp_enq_rorply_v_nxt ;
logic                                           smon_send_atm_to_cq_v_nxt ;
logic                                           smon_nalb_lsp_enq_rorply_v_nxt ;
logic                                           smon_qed_lsp_deq_v_nxt ;
logic                                           smon_aqed_lsp_deq_v_nxt ;
logic                                           smon_chp_lsp_token_ready_nxt ;
logic                                           smon_chp_lsp_cmp_ready_nxt ;
logic                                           smon_rop_lsp_reordercmp_ready_nxt ;
logic                                           smon_nalb_lsp_enq_lb_ready_nxt ;
logic                                           smon_dp_lsp_enq_dir_ready_nxt ;
logic                                           smon_dp_lsp_enq_rorply_ready_nxt ;
logic                                           smon_send_atm_to_cq_ready_nxt ;
logic                                           smon_nalb_lsp_enq_rorply_ready_nxt ;

logic                                           smon_lsp_dp_sch_dir_v_f ;
logic                                           smon_lsp_dp_sch_dir_rdy_f ;
logic [1:0]                                     smon_lsp_dp_sch_dir_cm_f ;
logic [1:0]                                     smon_lsp_dp_sch_dir_wbo_f ;
logic [7:0]                                     smon_lsp_dp_sch_dir_cq_f ;
logic                                           smon_lsp_dp_sch_dir_taken ;
logic                                           smon_lsp_dp_sch_dir_stalled ;
logic                                           smon_lsp_ap_atm_taken_f ;
logic                                           smon_lsp_ap_atm_stall_f ;
enum_cmd_lsp_ap_atm_t                           smon_lsp_ap_atm_cmd_f ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_lsp_ap_atm_cq_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_lsp_ap_atm_qid_f ;
logic [HQM_LSP_ARCH_NUM_FIDB2-1:0]              smon_lsp_ap_atm_fid_f ;
logic                                           smon_lsp_ap_atm_sch_rlist ;
logic                                           smon_lsp_ap_atm_sch_slist ;
logic                                           smon_lsp_ap_atm_sch_stall ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]            smon_lsp_nalb_sch_unoord_cq_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_lsp_nalb_sch_unoord_qid_f ;
logic                                           smon_atq_sel_ap_stall_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_atq_sel_ap_qid_f ;
logic                                           smon_rpl_dir_dp_stall_f ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]          smon_rpl_dir_dp_qid_f ;
logic                                           smon_rpl_ldb_nalb_stall_f ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]           smon_rpl_ldb_nalb_qid_f ;
logic [6:0]                                     smon_dp_lsp_enq_dir_data_qid_f ;
logic                                           smon_chp_lsp_token_data_is_ldb_f ;
logic [7:0]                                     smon_chp_lsp_token_data_cq_f ;
logic [12:0]                                    smon_chp_lsp_token_data_count_f ;
hqm_pkg::qtype_t                                smon_nalb_lsp_enq_lb_data_qtype_f ;
logic [6:0]                                     smon_nalb_lsp_enq_lb_data_qid_f ;
logic [6:0]                                     smon_chp_lsp_cmp_data_qid_f ;
logic [7:0]                                     smon_chp_lsp_cmp_data_cq_f ;
hqm_pkg::qtype_t                                smon_chp_lsp_cmp_data_qtype_f ;
logic [11:0]                                    smon_chp_lsp_cmp_data_fid_f ;
logic [6:0]                                     smon_rop_lsp_reordercmp_data_qid_f ;
logic [7:0]                                     smon_rop_lsp_reordercmp_data_cq_f ;
logic [6:0]                                     smon_dp_lsp_enq_rorply_data_qid_f ;
logic [6:0]                                     smon_nalb_lsp_enq_rorply_data_qid_f ;
logic [12:0]                                    smon_dp_lsp_enq_rorply_data_frag_cnt_f ;
logic [14:0]                                    smon_nalb_lsp_enq_rorply_data_frag_cnt_f ;
logic [5:0]                                     smon_qed_lsp_deq_data_cq_f ;
logic [5:0]                                     smon_aqed_lsp_deq_data_cq_f ;

logic					        smon_chp_lsp_token_v_f ;
logic					        smon_chp_lsp_cmp_v_f ;
logic					        smon_rop_lsp_reordercmp_v_f ;
logic					        smon_nalb_lsp_enq_lb_v_f ;
logic					        smon_dp_lsp_enq_dir_v_f ;
logic					        smon_dp_lsp_enq_rorply_v_f ;
logic					        smon_send_atm_to_cq_v_f ;
logic					        smon_nalb_lsp_enq_rorply_v_f ;
logic					        smon_qed_lsp_deq_v_f ;
logic					        smon_aqed_lsp_deq_v_f ;
logic					        smon_chp_lsp_token_ready_f ;
logic					        smon_chp_lsp_cmp_ready_f ;
logic					        smon_rop_lsp_reordercmp_ready_f ;
logic					        smon_nalb_lsp_enq_lb_ready_f ;
logic					        smon_dp_lsp_enq_dir_ready_f ;
logic					        smon_dp_lsp_enq_rorply_ready_f ;
logic					        smon_send_atm_to_cq_ready_f ;
logic					        smon_nalb_lsp_enq_rorply_ready_f ;
logic					        smon_chp_lsp_token_taken ;
logic					        smon_chp_lsp_cmp_taken ;
logic					        smon_rop_lsp_reordercmp_taken ;
logic					        smon_nalb_lsp_enq_lb_taken ;
logic					        smon_dp_lsp_enq_dir_taken ;
logic					        smon_dp_lsp_enq_rorply_taken ;
logic					        smon_send_atm_to_cq_taken ;
logic					        smon_nalb_lsp_enq_rorply_taken ;
logic					        smon_chp_lsp_token_stalled ;
logic					        smon_chp_lsp_cmp_stalled ;
logic					        smon_rop_lsp_reordercmp_stalled ;
logic					        smon_nalb_lsp_enq_lb_stalled ;
logic					        smon_dp_lsp_enq_dir_stalled ;
logic					        smon_dp_lsp_enq_rorply_stalled ;
logic					        smon_send_atm_to_cq_stalled ;
logic					        smon_nalb_lsp_enq_rorply_stalled ;

//------------------------------------------------------------------------------------------------
// V2 clock / sync / infrastructure declarations
logic                                           lsp_unit_idle_local ;

logic                                           ap_hqm_proc_clk_en_nc ;
logic                                           atm_clk_idle ;
logic                                           atm_clk_enable ;

//--------
logic                                           aqed_intf_enable_nc ;
logic                                           aqed_intf_idle ;
logic                                           aqed_lsp_dec_fid_cnt_v_idle ;
logic                                           atq_fid_cnt_upd_idle ;
logic                                           atq_stop_atqatm_idle ;
logic                                           chp_lsp_token_rx_sync_enable ;
logic                                           chp_lsp_token_rx_sync_idle ;
logic                                           chp_lsp_cmp_rx_sync_enable ;
logic                                           chp_lsp_cmp_rx_sync_idle ;
logic                                           rop_lsp_reordercmp_rx_sync_enable ;
logic                                           rop_lsp_reordercmp_rx_sync_idle ;
logic                                           nalb_lsp_enq_lb_rx_sync_enable ;
logic                                           nalb_lsp_enq_lb_rx_sync_idle ;
logic                                           dp_lsp_enq_dir_rx_sync_enable ;
logic                                           dp_lsp_enq_dir_rx_sync_idle ;
logic                                           dp_lsp_enq_rorply_rx_sync_enable ;
logic                                           dp_lsp_enq_rorply_rx_sync_idle ;
logic                                           send_atm_to_cq_rx_sync_enable ;
logic                                           send_atm_to_cq_rx_sync_idle ;
logic                                           nalb_lsp_enq_rorply_rx_sync_enable ;
logic                                           nalb_lsp_enq_rorply_rx_sync_idle ;
logic                                           rpl_ldb_nalb_tx_sync_idle ;
logic                                           lsp_nalb_sch_unoord_tx_sync_idle ;
logic                                           atq_sel_ap_tx_sync_idle ;
logic                                           lsp_dp_sch_dir_tx_sync_idle ;
logic                                           rpl_dir_dp_tx_sync_idle ;

logic                                           chp_lsp_token_rx_sync_fifo_of ;
logic                                           chp_lsp_token_rx_sync_fifo_uf ;
logic                                           chp_lsp_cmp_rx_sync_fifo_of ;
logic                                           chp_lsp_cmp_rx_sync_fifo_uf ;
logic                                           qed_lsp_deq_fifo_of ;
logic                                           qed_lsp_deq_fifo_uf ;
logic                                           qed_lsp_deq_fifo_empty ;
logic                                           aqed_lsp_deq_fifo_of ;
logic                                           aqed_lsp_deq_fifo_uf ;
logic                                           aqed_lsp_deq_fifo_empty ;
logic                                           rop_lsp_reordercmp_rx_sync_fifo_of ;
logic                                           rop_lsp_reordercmp_rx_sync_fifo_uf ;
logic                                           nalb_lsp_enq_lb_rx_sync_fifo_of ;
logic                                           nalb_lsp_enq_lb_rx_sync_fifo_uf ;
logic                                           dp_lsp_enq_dir_rx_sync_fifo_of ;
logic                                           dp_lsp_enq_dir_rx_sync_fifo_uf ;
logic                                           dp_lsp_enq_rorply_rx_sync_fifo_of ;
logic                                           dp_lsp_enq_rorply_rx_sync_fifo_uf ;
logic                                           send_atm_to_cq_rx_sync_fifo_of ;
logic                                           send_atm_to_cq_rx_sync_fifo_uf ;
logic                                           nalb_lsp_enq_rorply_rx_sync_fifo_of ;
logic                                           nalb_lsp_enq_rorply_rx_sync_fifo_uf ;
logic                                           rx_sync_fifo_error ;
//--------
logic                                           cfg_rx_enable ;
logic                                           cfg_rx_idle ;
aw_fifo_status_t                                cfg_rx_fifo_status_pnc ;

logic                                           cfg_rx_sync_fifo_of ;
logic                                           cfg_rx_sync_fifo_uf ;
//--------
logic [ HQM_LSP_DIRENQ_ENQ_CNT_MEM_WIDTH-1:0 ] pf_dir_enq_cnt_mem_rdata_nc ;
logic [ HQM_LSP_DIRENQ_TOK_CNT_MEM_WIDTH-1:0 ] pf_dir_tok_cnt_mem_rdata_nc ;
logic [ ( 8 ) - 1 : 0 ] pf_dir_tok_lim_mem_rdata_nc ;
logic [ ( 10 ) - 1 : 0 ] pf_enq_nalb_fifo_mem_rdata_nc ;
logic [ ( 20 ) - 1 : 0 ] pf_uno_atm_cmp_fifo_mem_rdata_nc ;
logic [ ( 18 ) - 1 : 0 ] pf_nalb_cmp_fifo_mem_rdata_nc ;
logic [ ( 55 ) - 1 : 0 ] pf_atm_cmp_fifo_mem_rdata_nc ;
logic [ ( 25 ) - 1 : 0 ] pf_ldb_token_rtn_fifo_mem_rdata_nc ;
logic [ ( 27 ) - 1 : 0 ] pf_nalb_sel_nalb_fifo_mem_rdata_nc ;
logic [ ( 33 ) - 1 : 0 ] pf_cfg_cq2priov_odd_mem_rdata_nc ;
logic [ ( 33 ) - 1 : 0 ] pf_cfg_cq2priov_mem_rdata_nc ;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2priov_odd_mem_raddr_nc;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2priov_mem_raddr_nc;
logic [ ( 29 ) - 1 : 0 ] pf_cfg_cq2qid_0_odd_mem_rdata_nc ;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2qid_0_odd_mem_raddr_nc;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2qid_0_mem_raddr_nc;
logic [ ( 29 ) - 1 : 0 ] pf_cfg_cq2qid_0_mem_rdata_nc ;
logic [ ( 29 ) - 1 : 0 ] pf_cfg_cq2qid_1_odd_mem_rdata_nc ;
logic [ ( 29 ) - 1 : 0 ] pf_cfg_cq2qid_1_mem_rdata_nc ;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2qid_1_odd_mem_raddr_nc;
logic [ ( 5 )  - 1 : 0 ] func_cfg_cq2qid_1_mem_raddr_nc;
logic [ HQM_LSP_LB_QID_ENQ_CNT_MEM_WIDTH-1:0 ] pf_qid_ldb_enqueue_count_mem_rdata_nc ;
logic [ HQM_LSP_LB_QID_IF_CNT_MEM_WIDTH-1:0 ] pf_qid_ldb_inflight_count_mem_rdata_nc ;
logic [ HQM_LSP_LB_QID_IF_LIM_MEM_WIDTH-1:0 ] pf_cfg_qid_ldb_inflight_limit_mem_rdata_nc ;
logic [ ( 528 ) - 1 : 0 ] pf_cfg_qid_ldb_qid2cqidix_mem_rdata_nc ;
logic [ ( 528 ) - 1 : 0 ] pf_cfg_qid_ldb_qid2cqidix2_mem_rdata_nc ;
logic [ ( 13 ) - 1 : 0 ] pf_cq_ldb_token_count_mem_rdata_nc ;
logic [ ( 5 ) - 1 : 0 ] pf_cfg_cq_ldb_token_depth_select_mem_rdata_nc ;
logic [ HQM_LSP_LB_CQ_IF_CNT_MEM_WIDTH-1:0 ] pf_cq_ldb_inflight_count_mem_rdata_nc ;
logic [ HQM_LSP_LB_CQ_IF_LIM_MEM_WIDTH-1:0 ] pf_cfg_cq_ldb_inflight_limit_mem_rdata_nc ;
logic [ HQM_LSP_LB_CQ_IF_THR_MEM_WIDTH-1:0 ] pf_cfg_cq_ldb_inflight_threshold_mem_rdata_nc ;
logic [ HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0 ] pf_cq_nalb_pri_arbindex_mem_rdata_nc ;
logic [ HQM_LSP_LB_ARBINDEX_MEM_WIDTH-1:0 ] pf_cq_atm_pri_arbindex_mem_rdata_nc ;
logic [ HQM_LSP_ATQ_ENQ_CNT_MEM_WIDTH-1:0 ] pf_qid_atq_enqueue_count_mem_rdata_nc ;
logic [ HQM_LSP_ATQ_AQED_ACT_CNT_MEM_WIDTH-1:0 ] pf_qid_aqed_active_count_mem_rdata_nc ;
logic [ HQM_LSP_ATQ_AQED_ACT_LIM_MEM_WIDTH-1:0 ] pf_cfg_qid_aqed_active_limit_mem_rdata_nc ;
logic [ HQM_LSP_LBRPL_ENQ_CNT_MEM_WIDTH-1:0 ] pf_qid_ldb_replay_count_mem_rdata_nc ;
logic [ HQM_LSP_DIRRPL_ENQ_CNT_MEM_WIDTH-1:0 ] pf_qid_dir_replay_count_mem_rdata_nc ;
logic [ ( 66 ) - 1 : 0 ] pf_qid_naldb_tot_enq_cnt_mem_rdata_nc ;
logic [ ( 66 ) - 1 : 0 ] pf_qid_atm_tot_enq_cnt_mem_rdata_nc ;
logic [ ( 66 ) - 1 : 0 ] pf_cq_ldb_tot_sch_cnt_mem_rdata_nc ;
logic [ ( 66 ) - 1 : 0 ] pf_qid_dir_tot_enq_cnt_mem_rdata_nc ;
logic [ ( 66 ) - 1 : 0 ] pf_cq_dir_tot_sch_cnt_mem_rdata_nc ;
logic [ HQM_LSP_LB_QID_ENQ_CNT_WIDTH-1:0 ] pf_qid_naldb_max_depth_mem_rdata_nc ;                // No check bits
logic [ HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1:0 ] pf_qid_dir_max_depth_mem_rdata_nc ;                  // No check bits
logic [ ( 25 ) - 1 : 0 ] pf_chp_lsp_token_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 73 ) - 1 : 0 ] pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 9 ) - 1 : 0 ] pf_qed_lsp_deq_fifo_mem_rdata_nc ;
logic [ ( 9 ) - 1 : 0 ] pf_aqed_lsp_deq_fifo_mem_rdata_nc ;
logic [ ( 17 ) - 1 : 0 ] pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 10 ) - 1 : 0 ] pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 8 ) - 1 : 0 ] pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 23 ) - 1 : 0 ] pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 35 ) - 1 : 0 ] pf_send_atm_to_cq_rx_sync_fifo_mem_rdata_nc ;
logic [ ( 27 ) - 1 : 0 ] pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata_nc ;
logic [ HQM_LSP_ATQ_QID_DPTH_THRSH_MEM_WIDTH-1:0 ] pf_cfg_atm_qid_dpth_thrsh_mem_rdata_nc ;
logic [ HQM_LSP_LB_QID_DPTH_THRSH_MEM_WIDTH-1:0 ] pf_cfg_nalb_qid_dpth_thrsh_mem_rdata_nc ;
logic [ HQM_LSP_DIRENQ_DPTH_THRSH_MEM_WIDTH-1:0 ] pf_cfg_dir_qid_dpth_thrsh_mem_rdata_nc ;
logic [ HQM_LSP_ATQ_ATM_ACTIVE_MEM_WIDTH-1:0 ] pf_qid_atm_active_mem_rdata_nc ;
logic [ ( 19 ) - 1 : 0 ] pf_cq_ldb_wu_count_mem_rdata_nc ;
logic [ ( 17 ) - 1 : 0 ] pf_cfg_cq_ldb_wu_limit_mem_rdata_nc ;
lba_ldb_arb_index2x_t pf_cq_nalb_pri_arbindex_mem_wdata_struct ;
lba_ldb_arb_index2x_t pf_cq_atm_pri_arbindex_mem_wdata_struct ;
logic reset_pf_count_lt_num_dir_qid ;
logic reset_pf_count_lt_num_dir_cq ;
logic reset_pf_count_lt_num_lb_qid ;
logic reset_pf_count_lt_num_lb_cq ;
logic reset_pf_count_lt_num_lb_pcq ;

logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_0_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_1_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_2_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_3_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_4_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_5_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_6_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_ldb_sched_perf_7_count_nc ;
logic [63:0]            hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count_nc ;
logic [31:0]            hqm_lsp_target_cfg_syndrome_hw_syndrome_data_nc ;
logic [31:0]            hqm_lsp_target_cfg_syndrome_sw_syndrome_data_nc ;

logic [31:0]            hqm_lsp_target_cfg_interface_status_reg_f_nc ;

//--------
logic                                   cfgsc_dir_tok_cnt_mem_we ;
lsp_direnq_tok_cnt_t                    cfgsc_dir_tok_cnt_mem_wdata_struct ;
logic [1:0]                             cfgsc_dir_tok_cnt_mem_wdata_struct_cnt_res_nc ;
lsp_direnq_tok_cnt_t                    pf_dir_tok_cnt_mem_wdata_struct ;

logic                                   cfgsc_dir_tok_lim_mem_we ;
lsp_direnq_tok_lim_t                    cfgsc_dir_tok_lim_mem_wdata_struct ;
logic [1:0]                             cfgsc_dir_tok_lim_mem_wdata_struct_spare_nc ;
logic                                   cfgsc_dir_tok_lim_mem_wdata_struct_lim_p_nc ;
lsp_direnq_tok_lim_t                    pf_dir_tok_lim_mem_wdata_struct ;

logic                                           cfgsc_cfg_cq2priov_mem_we ;
logic [32:0]                                    cfgsc_cfg_cq2priov_mem_wdata ;
logic                                           cfgsc_cfg_cq2priov_mem_re ;
logic [32:0]                                    cfgsc_cfg_cq2priov_mem_rdata ;
logic                                           cfgsc_cfg_cq2priov_mem_rdata_nc ;
logic                                           cfgsc_cfg_cq2priov_mem_ack ;
logic                                           cfgsc_func_cfg_cq2priov_mem_we ;
logic [(2*33)-1:0]                              cfgsc_func_cfg_cq2priov_mem_wdata ;
logic                                           cfgsc_func_cfg_cq2priov_mem_re ;
logic [(2*33)-1:0]                              cfgsc_func_cfg_cq2priov_mem_rdata ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2priov_mem_addr ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2priov_mem_raddr_nc ;

logic                                           cfgsc_cfg_cq2qid_0_mem_we ;
logic [28:0]                                    cfgsc_cfg_cq2qid_0_mem_wdata ;
logic                                           cfgsc_cfg_cq2qid_0_mem_re ;
logic [28:0]                                    cfgsc_cfg_cq2qid_0_mem_rdata ;
logic                                           cfgsc_cfg_cq2qid_0_mem_rdata_nc ;
logic                                           cfgsc_cfg_cq2qid_0_mem_ack ;
logic                                           cfgsc_func_cfg_cq2qid_0_mem_we ;
logic [(2*29)-1:0]                              cfgsc_func_cfg_cq2qid_0_mem_wdata ;
logic                                           cfgsc_func_cfg_cq2qid_0_mem_re ;
logic [(2*29)-1:0]                              cfgsc_func_cfg_cq2qid_0_mem_rdata ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2qid_0_mem_addr ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2qid_0_mem_raddr_nc ;

logic                                           cfgsc_cfg_cq2qid_1_mem_we ;
logic [28:0]                                    cfgsc_cfg_cq2qid_1_mem_wdata ;
logic                                           cfgsc_cfg_cq2qid_1_mem_re ;
logic [28:0]                                    cfgsc_cfg_cq2qid_1_mem_rdata ;
logic                                           cfgsc_cfg_cq2qid_1_mem_rdata_nc ;
logic                                           cfgsc_cfg_cq2qid_1_mem_ack ;
logic                                           cfgsc_func_cfg_cq2qid_1_mem_we ;
logic [(2*29)-1:0]                              cfgsc_func_cfg_cq2qid_1_mem_wdata ;
logic                                           cfgsc_func_cfg_cq2qid_1_mem_re ;
logic [(2*29)-1:0]                              cfgsc_func_cfg_cq2qid_1_mem_rdata ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2qid_1_mem_addr ;
logic [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0]        cfgsc_func_cfg_cq2qid_1_mem_raddr_nc ;

logic                                   cfgsc_qid_ldb_inflight_count_mem_we ;
lsp_lb_qid_if_cnt_t                     cfgsc_qid_ldb_inflight_count_mem_wdata_struct ;
logic [1:0]                             cfgsc_qid_ldb_inflight_count_mem_wdata_struct_cnt_res_nc ;
lsp_lb_qid_if_cnt_t                     pf_qid_ldb_inflight_count_mem_wdata_struct ;

logic                                   cfgsc_cfg_qid_ldb_inflight_limit_mem_we ;
lsp_lb_qid_if_lim_t                     cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct ;
logic                                   cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct_lim_p_nc ;
lsp_lb_qid_if_lim_t                     pf_cfg_qid_ldb_inflight_limit_mem_wdata_struct ;

logic                                   cfgsc_cfg_qid_ldb_qid2cqidix_mem_we ;
logic                                   cfgsc_cfg_qid_ldb_qid2cqidix2_mem_we ;

logic                                   cfgsc_cq_ldb_token_count_mem_we ;

logic                                   cfgsc_cfg_cq_ldb_token_depth_select_mem_we ;
lsp_lb_cq_tok_lim_t                     cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct ;
logic                                   cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct_lim_p_nc ;
lsp_lb_cq_tok_lim_t                     pf_cfg_cq_ldb_token_depth_select_mem_wdata_struct ;

logic                                   cfgsc_cq_ldb_inflight_count_mem_we ;
lsp_lb_cq_if_cnt_t                      cfgsc_cq_ldb_inflight_count_mem_wdata_struct ;
logic [1:0]                             cfgsc_cq_ldb_inflight_count_mem_wdata_struct_cnt_res_nc ;
lsp_lb_cq_if_cnt_t                      pf_cq_ldb_inflight_count_mem_wdata_struct ;

logic                                   cfgsc_cfg_cq_ldb_inflight_limit_mem_we ;
lsp_lb_cq_if_lim_t                      cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct ;
logic                                   cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct_lim_p_nc ;
lsp_lb_cq_if_lim_t                      pf_cfg_cq_ldb_inflight_limit_mem_wdata_struct ;

logic                                   cfgsc_cfg_cq_ldb_inflight_threshold_mem_we ;
lsp_lb_cq_if_thr_t                      cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct ;
logic                                   cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct_thr_p_nc ;
lsp_lb_cq_if_thr_t                      pf_cfg_cq_ldb_inflight_threshold_mem_wdata_struct ;

logic                                   cfgsc_cfg_qid_aqed_active_limit_mem_we ;
lsp_atq_aqed_act_lim_t                  cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct ;
logic                                   cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct_lim_p_nc ;
lsp_atq_aqed_act_lim_t                  pf_cfg_qid_aqed_active_limit_mem_wdata_struct ;

logic                                   cfgsc_qid_naldb_tot_enq_cnt_mem_we ;
logic                                   cfgsc_func_qid_naldb_tot_enq_cnt_mem_we ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   cfgsc_func_qid_naldb_tot_enq_cnt_mem_waddr ;
logic [65:0]                            cfgsc_func_qid_naldb_tot_enq_cnt_mem_wdata ;

logic                                   cfgsc_qid_atm_tot_enq_cnt_mem_we ;
logic                                   cfgsc_func_qid_atm_tot_enq_cnt_mem_we ;
logic [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0]   cfgsc_func_qid_atm_tot_enq_cnt_mem_waddr ;
logic [65:0]                            cfgsc_func_qid_atm_tot_enq_cnt_mem_wdata ;

logic                                   cfgsc_cq_ldb_tot_sch_cnt_mem_we ;
logic                                   cfgsc_func_cq_ldb_tot_sch_cnt_mem_we ;
logic [HQM_LSP_ARCH_NUM_LB_CQB2-1:0]    cfgsc_func_cq_ldb_tot_sch_cnt_mem_waddr ;
logic [65:0]                            cfgsc_func_cq_ldb_tot_sch_cnt_mem_wdata ;

logic                                   cfgsc_qid_dir_tot_enq_cnt_mem_we ;
logic                                   cfgsc_func_qid_dir_tot_enq_cnt_mem_we ;
logic [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0]  cfgsc_func_qid_dir_tot_enq_cnt_mem_waddr ;
logic [65:0]                            cfgsc_func_qid_dir_tot_enq_cnt_mem_wdata ;

logic                                   cfgsc_cq_dir_tot_sch_cnt_mem_we ;
logic                                   cfgsc_func_cq_dir_tot_sch_cnt_mem_we ;
logic [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0]   cfgsc_func_cq_dir_tot_sch_cnt_mem_waddr ;
logic [65:0]                            cfgsc_func_cq_dir_tot_sch_cnt_mem_wdata ;

logic                                   cfgsc_qid_naldb_max_depth_mem_we ;

logic                                   cfgsc_qid_dir_max_depth_mem_we ;

logic                                   cfgsc_cfg_atm_qid_dpth_thrsh_mem_we ;

logic                                   cfgsc_cfg_nalb_qid_dpth_thrsh_mem_we ;

logic                                   cfgsc_cfg_dir_qid_dpth_thrsh_mem_we ;

logic                                   cfgsc_cq_ldb_wu_count_mem_re ;
logic                                   cfgsc_cq_ldb_wu_count_mem_we ;

logic                                   cfgsc_cfg_cq_ldb_wu_limit_mem_re ;
logic                                   cfgsc_cfg_cq_ldb_wu_limit_mem_we ;

logic                                   cfgsc_wu_count_wr_ack ;
logic                                   cfgsc_wu_count_rd_ack ;
logic                                   cfgsc_wu_limit_wr_ack ;
logic                                   cfgsc_wu_limit_rd_ack ;
logic [31:0]                            cfgsc_wu_cfg_data_f ;

logic                                   cfgsc_wide_memory_wait_for_write_nxt ;
logic                                   cfgsc_wide_memory_wait_for_write_f ;
logic                                   cfg_mem_ack_qid_naldb_tot_enq_cnt_nxt ;
logic                                   cfg_mem_ack_qid_naldb_tot_enq_cnt_f ;
logic                                   cfg_mem_ack_qid_atm_tot_enq_cnt_nxt ;
logic                                   cfg_mem_ack_qid_atm_tot_enq_cnt_f ;
logic                                   cfg_mem_ack_cq_ldb_tot_sch_cnt_nxt ;
logic                                   cfg_mem_ack_cq_ldb_tot_sch_cnt_f ;
logic                                   cfg_mem_ack_qid_dir_tot_enq_cnt_nxt ;
logic                                   cfg_mem_ack_qid_dir_tot_enq_cnt_f ;
logic                                   cfg_mem_ack_cq_dir_tot_sch_cnt_nxt ;
logic                                   cfg_mem_ack_cq_dir_tot_sch_cnt_f ;

logic                                   cfg_range_reconfig ;

logic                                   mem_access_error_nxt ;
logic                                   mem_access_error_f ;

logic [31:0]                            hqm_lsp_target_cfg_debug_00_reg_nxt ;
logic [31:0]                            hqm_lsp_target_cfg_debug_00_reg_f ;
logic [31:0]                            hqm_lsp_target_cfg_debug_01_reg_nxt ;
logic [31:0]                            hqm_lsp_target_cfg_debug_01_reg_f ;

//------------------------------------------------------------------------------------------------
// Misc logic declarations

//-------------------------------------------------------------------------------------------------
function automatic [1:0] hqm_lsp_calc_thresh_code ;
// Compare enqueue count with cfg threshold, encode with following meaning:
// 00 : <=  0.5  threshold
// 01 : >   0.5  threshold  <= 0.75 threshold
// 10 : >   0.75 threshold  <=      threshold
// 11 : >        threshold
  input logic [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:0] count ;
  input logic [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:0] thresh ;
  logic [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:0] thresh_p25 ;
  logic [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:0] thresh_p50 ;
  logic [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:0] thresh_p75 ;
  logic count_gt_thresh_p50 ;
  logic count_gt_thresh_p75 ;
  logic count_gt_thresh ;
  logic [1:0] code ;
  begin
    thresh_p25          = { 2'h0 , thresh [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:2] } ;
    thresh_p50          = { 1'b0 , thresh [HQM_LSP_MAX_LB_ENQ_COUNT_WIDTH-1:1] } ;

    // Hopefully this will not be a delay issue
    thresh_p75          = thresh_p50 + thresh_p25 ;     // Not possible to overflow

    count_gt_thresh     = ( count > thresh ) ;
    count_gt_thresh_p75 = ( count > thresh_p75 ) ;
    count_gt_thresh_p50 = ( count > thresh_p50 ) ;

    code [0]            = count_gt_thresh | ( count_gt_thresh_p50 & ~ count_gt_thresh_p75 ) ;
    code [1]            = count_gt_thresh_p75 ;
  end
  return code ;
endfunction // hqm_lsp_calc_thresh_code
//-------------------------------------------------------------------------------------------------

logic [ (32) -1 : 0 ]  reset_pf_counter_nxt, reset_pf_counter_f ;
logic hw_init_done_f, hw_init_done_nxt ;
logic reset_pf_active_f , reset_pf_active_nxt ;
logic reset_pf_done_f , reset_pf_done_nxt ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: BEGIN common core interfaces
//*****************************************************************************************************
//*****************************************************************************************************

//---------------------------------------------------------------------------------------------------------
// common core - Reset
logic rst_prep;
logic hqm_gated_rst_n;
logic hqm_inp_gated_rst_n;
assign rst_prep             = hqm_rst_prep_lsp;
assign hqm_gated_rst_n      = hqm_gated_rst_b_lsp;
assign hqm_inp_gated_rst_n  = hqm_inp_gated_rst_b_lsp;

logic hqm_gated_rst_n_start;
logic hqm_gated_rst_n_active;
logic hqm_gated_rst_n_done;
assign hqm_gated_rst_n_start    = hqm_gated_rst_b_start_lsp;
assign hqm_gated_rst_n_active   = hqm_gated_rst_b_active_lsp;
assign hqm_gated_rst_n_done = reset_pf_done_f ;
assign hqm_gated_rst_b_done_lsp = hqm_gated_rst_n_done;

//---------------------------------------------------------------------------------------------------------
// common core - CFG accessible patch & proc registers 
// common core - RFW/SRW RAM gasket
// common core - RAM wrapper for all 2 port RF RAMs
// common core - RAM wrapper for all single PORT SR RAMs
// common core - Interface & clock control
// common core - Configuration Ring, sidecar, interrupt serializer

// The following must be kept in-sync with generated code
// BEGIN HQM_CFG_ACCESS
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] pfcsr_cfg_req_write ; //I CFG
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] pfcsr_cfg_req_read ; //I CFG
cfg_req_t pfcsr_cfg_req ; //I CFG
logic pfcsr_cfg_rsp_ack ; //O CFG
logic pfcsr_cfg_rsp_err ; //O CFG
logic [ ( 32 ) - 1 : 0 ] pfcsr_cfg_rsp_rdata ; //O CFG
 logic [ ( HQM_NUM_DIR_CQ ) - 1 : 0 ] pfcsr_shadow_nxt , pfcsr_shadow_f ;
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_nxt ; //I HQM_LSP_TARGET_CFG_AQED_TOT_ENQUEUE_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_f ; //O HQM_LSP_TARGET_CFG_AQED_TOT_ENQUEUE_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_nxt ; //I HQM_LSP_TARGET_CFG_AQED_TOT_ENQUEUE_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_f ; //O HQM_LSP_TARGET_CFG_AQED_TOT_ENQUEUE_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_nxt ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_f ; //O HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_0
logic hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_v ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_nxt ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_f ; //O HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_1
logic hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_v ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_ATM_NALB_QID_1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_nxt ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_ISSUE_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_f ; //O HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_ISSUE_0
logic hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_v ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_ISSUE_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_nxt ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_f ; //O HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_0
logic hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_v ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_nxt ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_f ; //O HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_1
logic hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_v ; //I HQM_LSP_TARGET_CFG_ARB_WEIGHT_LDB_QID_1
logic hqm_lsp_target_cfg_cnt_win_cos0_en ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS0
logic hqm_lsp_target_cfg_cnt_win_cos0_clr ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS0
logic hqm_lsp_target_cfg_cnt_win_cos0_clrv ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS0
logic hqm_lsp_target_cfg_cnt_win_cos0_inc ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cnt_win_cos0_count ; //O HQM_LSP_TARGET_CFG_CNT_WIN_COS0
logic hqm_lsp_target_cfg_cnt_win_cos1_en ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS1
logic hqm_lsp_target_cfg_cnt_win_cos1_clr ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS1
logic hqm_lsp_target_cfg_cnt_win_cos1_clrv ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS1
logic hqm_lsp_target_cfg_cnt_win_cos1_inc ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cnt_win_cos1_count ; //O HQM_LSP_TARGET_CFG_CNT_WIN_COS1
logic hqm_lsp_target_cfg_cnt_win_cos2_en ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS2
logic hqm_lsp_target_cfg_cnt_win_cos2_clr ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS2
logic hqm_lsp_target_cfg_cnt_win_cos2_clrv ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS2
logic hqm_lsp_target_cfg_cnt_win_cos2_inc ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cnt_win_cos2_count ; //O HQM_LSP_TARGET_CFG_CNT_WIN_COS2
logic hqm_lsp_target_cfg_cnt_win_cos3_en ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS3
logic hqm_lsp_target_cfg_cnt_win_cos3_clr ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS3
logic hqm_lsp_target_cfg_cnt_win_cos3_clrv ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS3
logic hqm_lsp_target_cfg_cnt_win_cos3_inc ; //I HQM_LSP_TARGET_CFG_CNT_WIN_COS3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cnt_win_cos3_count ; //O HQM_LSP_TARGET_CFG_CNT_WIN_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_general_0_reg_nxt ; //I HQM_LSP_TARGET_CFG_CONTROL_GENERAL_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_general_0_reg_f ; //O HQM_LSP_TARGET_CFG_CONTROL_GENERAL_0
logic hqm_lsp_target_cfg_control_general_0_reg_v ; //I HQM_LSP_TARGET_CFG_CONTROL_GENERAL_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_general_1_reg_nxt ; //I HQM_LSP_TARGET_CFG_CONTROL_GENERAL_1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_general_1_reg_f ; //O HQM_LSP_TARGET_CFG_CONTROL_GENERAL_1
logic hqm_lsp_target_cfg_control_general_1_reg_v ; //I HQM_LSP_TARGET_CFG_CONTROL_GENERAL_1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_pipeline_credits_reg_nxt ; //I HQM_LSP_TARGET_CFG_CONTROL_PIPELINE_CREDITS
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_pipeline_credits_reg_f ; //O HQM_LSP_TARGET_CFG_CONTROL_PIPELINE_CREDITS
logic hqm_lsp_target_cfg_control_pipeline_credits_reg_v ; //I HQM_LSP_TARGET_CFG_CONTROL_PIPELINE_CREDITS
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_sched_slot_count_reg_nxt ; //I HQM_LSP_TARGET_CFG_CONTROL_SCHED_SLOT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_control_sched_slot_count_reg_f ; //O HQM_LSP_TARGET_CFG_CONTROL_SCHED_SLOT_COUNT
logic hqm_lsp_target_cfg_control_sched_slot_count_reg_v ; //I HQM_LSP_TARGET_CFG_CONTROL_SCHED_SLOT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cos_ctrl_reg_nxt ; //I HQM_LSP_TARGET_CFG_COS_CTRL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cos_ctrl_reg_f ; //O HQM_LSP_TARGET_CFG_COS_CTRL
logic hqm_lsp_target_cfg_cos_ctrl_reg_v ; //I HQM_LSP_TARGET_CFG_COS_CTRL
logic hqm_lsp_target_cfg_cq_dir_disable_reg_load ; //I HQM_LSP_TARGET_CFG_CQ_DIR_DISABLE
logic [ ( 1 * 1 * 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_dir_disable_reg_nxt ; //I HQM_LSP_TARGET_CFG_CQ_DIR_DISABLE
logic [ ( 1 * 1 * 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_dir_disable_reg_f ; //O HQM_LSP_TARGET_CFG_CQ_DIR_DISABLE
logic hqm_lsp_target_cfg_cq_ldb_disable_reg_load ; //I HQM_LSP_TARGET_CFG_CQ_LDB_DISABLE
logic [ ( 1 * 2 * 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_disable_reg_nxt ; //I HQM_LSP_TARGET_CFG_CQ_LDB_DISABLE
logic [ ( 1 * 2 * 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_disable_reg_f ; //O HQM_LSP_TARGET_CFG_CQ_LDB_DISABLE
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_0
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_0
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_0
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_0
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_1
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_1
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_1
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_1
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_2
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_2
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_2
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_2
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_3
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_3
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_3
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_3
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_4
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_4
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_4
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_4
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_4
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_5
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_5
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_5
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_5
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_5
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_6
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_6
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_6
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_6
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_6
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_en ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_7
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clr ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_7
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clrv ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_7
logic hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_inc ; //I HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_7
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count ; //O HQM_LSP_TARGET_CFG_CQ_LDB_SCHED_SLOT_COUNT_7
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_nxt ; //I HQM_LSP_TARGET_CFG_CQ_LDB_TOT_INFLIGHT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_f ; //O HQM_LSP_TARGET_CFG_CQ_LDB_TOT_INFLIGHT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_nxt ; //I HQM_LSP_TARGET_CFG_CQ_LDB_TOT_INFLIGHT_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_f ; //O HQM_LSP_TARGET_CFG_CQ_LDB_TOT_INFLIGHT_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos0_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_CNT_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos0_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_CNT_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos1_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_CNT_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos1_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_CNT_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos2_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_CNT_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos2_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_CNT_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos3_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_CNT_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_cnt_cos3_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_CNT_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos0_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos0_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_SAT_COS0
logic hqm_lsp_target_cfg_credit_sat_cos0_reg_v ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos1_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos1_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_SAT_COS1
logic hqm_lsp_target_cfg_credit_sat_cos1_reg_v ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos2_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos2_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_SAT_COS2
logic hqm_lsp_target_cfg_credit_sat_cos2_reg_v ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos3_reg_nxt ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_credit_sat_cos3_reg_f ; //O HQM_LSP_TARGET_CFG_CREDIT_SAT_COS3
logic hqm_lsp_target_cfg_credit_sat_cos3_reg_v ; //I HQM_LSP_TARGET_CFG_CREDIT_SAT_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_diagnostic_aw_status_status ; //I HQM_LSP_TARGET_CFG_DIAGNOSTIC_AW_STATUS
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_diagnostic_status_0_status ; //I HQM_LSP_TARGET_CFG_DIAGNOSTIC_STATUS_0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_error_inject_reg_nxt ; //I HQM_LSP_TARGET_CFG_ERROR_INJECT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_error_inject_reg_f ; //O HQM_LSP_TARGET_CFG_ERROR_INJECT
logic hqm_lsp_target_cfg_error_inject_reg_v ; //I HQM_LSP_TARGET_CFG_ERROR_INJECT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_fid_inflight_count_reg_nxt ; //I HQM_LSP_TARGET_CFG_FID_INFLIGHT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_fid_inflight_count_reg_f ; //O HQM_LSP_TARGET_CFG_FID_INFLIGHT_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_fid_inflight_limit_reg_nxt ; //I HQM_LSP_TARGET_CFG_FID_INFLIGHT_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_fid_inflight_limit_reg_f ; //O HQM_LSP_TARGET_CFG_FID_INFLIGHT_LIMIT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_hw_agitate_control_reg_nxt ; //I HQM_LSP_TARGET_CFG_HW_AGITATE_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_hw_agitate_control_reg_f ; //O HQM_LSP_TARGET_CFG_HW_AGITATE_CONTROL
logic hqm_lsp_target_cfg_hw_agitate_control_reg_v ; //I HQM_LSP_TARGET_CFG_HW_AGITATE_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_hw_agitate_select_reg_nxt ; //I HQM_LSP_TARGET_CFG_HW_AGITATE_SELECT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_hw_agitate_select_reg_f ; //O HQM_LSP_TARGET_CFG_HW_AGITATE_SELECT
logic hqm_lsp_target_cfg_hw_agitate_select_reg_v ; //I HQM_LSP_TARGET_CFG_HW_AGITATE_SELECT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_interface_status_reg_nxt ; //I HQM_LSP_TARGET_CFG_INTERFACE_STATUS
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_interface_status_reg_f ; //O HQM_LSP_TARGET_CFG_INTERFACE_STATUS
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_control_reg_nxt ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_control_reg_f ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_CONTROL
logic hqm_lsp_target_cfg_ldb_sched_perf_0_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_0
logic hqm_lsp_target_cfg_ldb_sched_perf_0_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_0
logic hqm_lsp_target_cfg_ldb_sched_perf_0_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_0
logic hqm_lsp_target_cfg_ldb_sched_perf_0_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_0_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_0
logic hqm_lsp_target_cfg_ldb_sched_perf_1_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_1
logic hqm_lsp_target_cfg_ldb_sched_perf_1_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_1
logic hqm_lsp_target_cfg_ldb_sched_perf_1_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_1
logic hqm_lsp_target_cfg_ldb_sched_perf_1_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_1_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_1
logic hqm_lsp_target_cfg_ldb_sched_perf_2_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_2
logic hqm_lsp_target_cfg_ldb_sched_perf_2_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_2
logic hqm_lsp_target_cfg_ldb_sched_perf_2_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_2
logic hqm_lsp_target_cfg_ldb_sched_perf_2_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_2_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_2
logic hqm_lsp_target_cfg_ldb_sched_perf_3_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_3
logic hqm_lsp_target_cfg_ldb_sched_perf_3_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_3
logic hqm_lsp_target_cfg_ldb_sched_perf_3_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_3
logic hqm_lsp_target_cfg_ldb_sched_perf_3_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_3_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_3
logic hqm_lsp_target_cfg_ldb_sched_perf_4_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_4
logic hqm_lsp_target_cfg_ldb_sched_perf_4_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_4
logic hqm_lsp_target_cfg_ldb_sched_perf_4_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_4
logic hqm_lsp_target_cfg_ldb_sched_perf_4_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_4
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_4_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_4
logic hqm_lsp_target_cfg_ldb_sched_perf_5_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_5
logic hqm_lsp_target_cfg_ldb_sched_perf_5_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_5
logic hqm_lsp_target_cfg_ldb_sched_perf_5_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_5
logic hqm_lsp_target_cfg_ldb_sched_perf_5_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_5
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_5_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_5
logic hqm_lsp_target_cfg_ldb_sched_perf_6_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_6
logic hqm_lsp_target_cfg_ldb_sched_perf_6_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_6
logic hqm_lsp_target_cfg_ldb_sched_perf_6_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_6
logic hqm_lsp_target_cfg_ldb_sched_perf_6_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_6
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_6_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_6
logic hqm_lsp_target_cfg_ldb_sched_perf_7_en ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_7
logic hqm_lsp_target_cfg_ldb_sched_perf_7_clr ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_7
logic hqm_lsp_target_cfg_ldb_sched_perf_7_clrv ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_7
logic hqm_lsp_target_cfg_ldb_sched_perf_7_inc ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_7
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_7_count ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_7
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_control_reg_nxt ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f ; //O HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_CONTROL
logic hqm_lsp_target_cfg_ldb_sched_perf_control_reg_v ; //I HQM_LSP_TARGET_CFG_LDB_SCHED_PERF_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_csr_control_reg_nxt ; //I HQM_LSP_TARGET_CFG_LSP_CSR_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_csr_control_reg_f ; //O HQM_LSP_TARGET_CFG_LSP_CSR_CONTROL
logic hqm_lsp_target_cfg_lsp_csr_control_reg_v ; //I HQM_LSP_TARGET_CFG_LSP_CSR_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_nxt ; //I HQM_LSP_TARGET_CFG_LSP_PERF_DIR_SCH_COUNT_H
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_f ; //O HQM_LSP_TARGET_CFG_LSP_PERF_DIR_SCH_COUNT_H
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_nxt ; //I HQM_LSP_TARGET_CFG_LSP_PERF_DIR_SCH_COUNT_L
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_f ; //O HQM_LSP_TARGET_CFG_LSP_PERF_DIR_SCH_COUNT_L
logic hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_en ; //I HQM_LSP_TARGET_CFG_LSP_PERF_LDB_SCH_COUNT
logic hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clr ; //I HQM_LSP_TARGET_CFG_LSP_PERF_LDB_SCH_COUNT
logic hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clrv ; //I HQM_LSP_TARGET_CFG_LSP_PERF_LDB_SCH_COUNT
logic hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_inc ; //I HQM_LSP_TARGET_CFG_LSP_PERF_LDB_SCH_COUNT
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count ; //O HQM_LSP_TARGET_CFG_LSP_PERF_LDB_SCH_COUNT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_patch_control_reg_nxt ; //I HQM_LSP_TARGET_CFG_PATCH_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_patch_control_reg_f ; //O HQM_LSP_TARGET_CFG_PATCH_CONTROL
logic hqm_lsp_target_cfg_patch_control_reg_v ; //I HQM_LSP_TARGET_CFG_PATCH_CONTROL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_pipe_health_hold_00_status ; //I HQM_LSP_TARGET_CFG_PIPE_HEALTH_HOLD_00
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_pipe_health_hold_01_status ; //I HQM_LSP_TARGET_CFG_PIPE_HEALTH_HOLD_01
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_pipe_health_valid_00_status ; //I HQM_LSP_TARGET_CFG_PIPE_HEALTH_VALID_00
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_pipe_health_valid_01_status ; //I HQM_LSP_TARGET_CFG_PIPE_HEALTH_VALID_01
logic hqm_lsp_target_cfg_rdy_cos0_en ; //I HQM_LSP_TARGET_CFG_RDY_COS0
logic hqm_lsp_target_cfg_rdy_cos0_clr ; //I HQM_LSP_TARGET_CFG_RDY_COS0
logic hqm_lsp_target_cfg_rdy_cos0_clrv ; //I HQM_LSP_TARGET_CFG_RDY_COS0
logic hqm_lsp_target_cfg_rdy_cos0_inc ; //I HQM_LSP_TARGET_CFG_RDY_COS0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rdy_cos0_count ; //O HQM_LSP_TARGET_CFG_RDY_COS0
logic hqm_lsp_target_cfg_rdy_cos1_en ; //I HQM_LSP_TARGET_CFG_RDY_COS1
logic hqm_lsp_target_cfg_rdy_cos1_clr ; //I HQM_LSP_TARGET_CFG_RDY_COS1
logic hqm_lsp_target_cfg_rdy_cos1_clrv ; //I HQM_LSP_TARGET_CFG_RDY_COS1
logic hqm_lsp_target_cfg_rdy_cos1_inc ; //I HQM_LSP_TARGET_CFG_RDY_COS1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rdy_cos1_count ; //O HQM_LSP_TARGET_CFG_RDY_COS1
logic hqm_lsp_target_cfg_rdy_cos2_en ; //I HQM_LSP_TARGET_CFG_RDY_COS2
logic hqm_lsp_target_cfg_rdy_cos2_clr ; //I HQM_LSP_TARGET_CFG_RDY_COS2
logic hqm_lsp_target_cfg_rdy_cos2_clrv ; //I HQM_LSP_TARGET_CFG_RDY_COS2
logic hqm_lsp_target_cfg_rdy_cos2_inc ; //I HQM_LSP_TARGET_CFG_RDY_COS2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rdy_cos2_count ; //O HQM_LSP_TARGET_CFG_RDY_COS2
logic hqm_lsp_target_cfg_rdy_cos3_en ; //I HQM_LSP_TARGET_CFG_RDY_COS3
logic hqm_lsp_target_cfg_rdy_cos3_clr ; //I HQM_LSP_TARGET_CFG_RDY_COS3
logic hqm_lsp_target_cfg_rdy_cos3_clrv ; //I HQM_LSP_TARGET_CFG_RDY_COS3
logic hqm_lsp_target_cfg_rdy_cos3_inc ; //I HQM_LSP_TARGET_CFG_RDY_COS3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rdy_cos3_count ; //O HQM_LSP_TARGET_CFG_RDY_COS3
logic hqm_lsp_target_cfg_rnd_loss_cos0_en ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS0
logic hqm_lsp_target_cfg_rnd_loss_cos0_clr ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS0
logic hqm_lsp_target_cfg_rnd_loss_cos0_clrv ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS0
logic hqm_lsp_target_cfg_rnd_loss_cos0_inc ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rnd_loss_cos0_count ; //O HQM_LSP_TARGET_CFG_RND_LOSS_COS0
logic hqm_lsp_target_cfg_rnd_loss_cos1_en ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS1
logic hqm_lsp_target_cfg_rnd_loss_cos1_clr ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS1
logic hqm_lsp_target_cfg_rnd_loss_cos1_clrv ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS1
logic hqm_lsp_target_cfg_rnd_loss_cos1_inc ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rnd_loss_cos1_count ; //O HQM_LSP_TARGET_CFG_RND_LOSS_COS1
logic hqm_lsp_target_cfg_rnd_loss_cos2_en ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS2
logic hqm_lsp_target_cfg_rnd_loss_cos2_clr ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS2
logic hqm_lsp_target_cfg_rnd_loss_cos2_clrv ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS2
logic hqm_lsp_target_cfg_rnd_loss_cos2_inc ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rnd_loss_cos2_count ; //O HQM_LSP_TARGET_CFG_RND_LOSS_COS2
logic hqm_lsp_target_cfg_rnd_loss_cos3_en ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS3
logic hqm_lsp_target_cfg_rnd_loss_cos3_clr ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS3
logic hqm_lsp_target_cfg_rnd_loss_cos3_clrv ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS3
logic hqm_lsp_target_cfg_rnd_loss_cos3_inc ; //I HQM_LSP_TARGET_CFG_RND_LOSS_COS3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_rnd_loss_cos3_count ; //O HQM_LSP_TARGET_CFG_RND_LOSS_COS3
logic hqm_lsp_target_cfg_schd_cos0_en ; //I HQM_LSP_TARGET_CFG_SCHD_COS0
logic hqm_lsp_target_cfg_schd_cos0_clr ; //I HQM_LSP_TARGET_CFG_SCHD_COS0
logic hqm_lsp_target_cfg_schd_cos0_clrv ; //I HQM_LSP_TARGET_CFG_SCHD_COS0
logic hqm_lsp_target_cfg_schd_cos0_inc ; //I HQM_LSP_TARGET_CFG_SCHD_COS0
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_schd_cos0_count ; //O HQM_LSP_TARGET_CFG_SCHD_COS0
logic hqm_lsp_target_cfg_schd_cos1_en ; //I HQM_LSP_TARGET_CFG_SCHD_COS1
logic hqm_lsp_target_cfg_schd_cos1_clr ; //I HQM_LSP_TARGET_CFG_SCHD_COS1
logic hqm_lsp_target_cfg_schd_cos1_clrv ; //I HQM_LSP_TARGET_CFG_SCHD_COS1
logic hqm_lsp_target_cfg_schd_cos1_inc ; //I HQM_LSP_TARGET_CFG_SCHD_COS1
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_schd_cos1_count ; //O HQM_LSP_TARGET_CFG_SCHD_COS1
logic hqm_lsp_target_cfg_schd_cos2_en ; //I HQM_LSP_TARGET_CFG_SCHD_COS2
logic hqm_lsp_target_cfg_schd_cos2_clr ; //I HQM_LSP_TARGET_CFG_SCHD_COS2
logic hqm_lsp_target_cfg_schd_cos2_clrv ; //I HQM_LSP_TARGET_CFG_SCHD_COS2
logic hqm_lsp_target_cfg_schd_cos2_inc ; //I HQM_LSP_TARGET_CFG_SCHD_COS2
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_schd_cos2_count ; //O HQM_LSP_TARGET_CFG_SCHD_COS2
logic hqm_lsp_target_cfg_schd_cos3_en ; //I HQM_LSP_TARGET_CFG_SCHD_COS3
logic hqm_lsp_target_cfg_schd_cos3_clr ; //I HQM_LSP_TARGET_CFG_SCHD_COS3
logic hqm_lsp_target_cfg_schd_cos3_clrv ; //I HQM_LSP_TARGET_CFG_SCHD_COS3
logic hqm_lsp_target_cfg_schd_cos3_inc ; //I HQM_LSP_TARGET_CFG_SCHD_COS3
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_schd_cos3_count ; //O HQM_LSP_TARGET_CFG_SCHD_COS3
logic hqm_lsp_target_cfg_sch_rdy_en ; //I HQM_LSP_TARGET_CFG_SCH_RDY
logic hqm_lsp_target_cfg_sch_rdy_clr ; //I HQM_LSP_TARGET_CFG_SCH_RDY
logic hqm_lsp_target_cfg_sch_rdy_clrv ; //I HQM_LSP_TARGET_CFG_SCH_RDY
logic hqm_lsp_target_cfg_sch_rdy_inc ; //I HQM_LSP_TARGET_CFG_SCH_RDY
logic [ ( 64 ) - 1 : 0] hqm_lsp_target_cfg_sch_rdy_count ; //O HQM_LSP_TARGET_CFG_SCH_RDY
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_ctrl_reg_nxt ; //I HQM_LSP_TARGET_CFG_SHDW_CTRL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_ctrl_reg_f ; //O HQM_LSP_TARGET_CFG_SHDW_CTRL
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos0_reg_nxt ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos0_reg_f ; //O HQM_LSP_TARGET_CFG_SHDW_RANGE_COS0
logic hqm_lsp_target_cfg_shdw_range_cos0_reg_v ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS0
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos1_reg_nxt ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos1_reg_f ; //O HQM_LSP_TARGET_CFG_SHDW_RANGE_COS1
logic hqm_lsp_target_cfg_shdw_range_cos1_reg_v ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS1
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos2_reg_nxt ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos2_reg_f ; //O HQM_LSP_TARGET_CFG_SHDW_RANGE_COS2
logic hqm_lsp_target_cfg_shdw_range_cos2_reg_v ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS2
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos3_reg_nxt ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS3
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_shdw_range_cos3_reg_f ; //O HQM_LSP_TARGET_CFG_SHDW_RANGE_COS3
logic hqm_lsp_target_cfg_shdw_range_cos3_reg_v ; //I HQM_LSP_TARGET_CFG_SHDW_RANGE_COS3
logic hqm_lsp_target_cfg_smon0_disable_smon ; //I HQM_LSP_TARGET_CFG_SMON0
logic [ 24 - 1 : 0 ] hqm_lsp_target_cfg_smon0_smon_v ; //I HQM_LSP_TARGET_CFG_SMON0
logic [ ( 24 * 32 ) - 1 : 0 ] hqm_lsp_target_cfg_smon0_smon_comp ; //I HQM_LSP_TARGET_CFG_SMON0
logic [ ( 24 * 32 ) - 1 : 0 ] hqm_lsp_target_cfg_smon0_smon_val ; //I HQM_LSP_TARGET_CFG_SMON0
logic hqm_lsp_target_cfg_smon0_smon_enabled ; //O HQM_LSP_TARGET_CFG_SMON0
logic hqm_lsp_target_cfg_smon0_smon_interrupt ; //O HQM_LSP_TARGET_CFG_SMON0
logic hqm_lsp_target_cfg_syndrome_hw_capture_v ; //I HQM_LSP_TARGET_CFG_SYNDROME_HW
logic [ ( 31 ) - 1 : 0] hqm_lsp_target_cfg_syndrome_hw_capture_data ; //I HQM_LSP_TARGET_CFG_SYNDROME_HW
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_syndrome_hw_syndrome_data ; //I HQM_LSP_TARGET_CFG_SYNDROME_HW
logic hqm_lsp_target_cfg_syndrome_sw_capture_v ; //I HQM_LSP_TARGET_CFG_SYNDROME_SW
logic [ ( 31 ) - 1 : 0] hqm_lsp_target_cfg_syndrome_sw_capture_data ; //I HQM_LSP_TARGET_CFG_SYNDROME_SW
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_syndrome_sw_syndrome_data ; //I HQM_LSP_TARGET_CFG_SYNDROME_SW
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_unit_idle_reg_nxt ; //I HQM_LSP_TARGET_CFG_UNIT_IDLE
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_unit_idle_reg_f ; //O HQM_LSP_TARGET_CFG_UNIT_IDLE
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_unit_timeout_reg_nxt ; //I HQM_LSP_TARGET_CFG_UNIT_TIMEOUT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_unit_timeout_reg_f ; //O HQM_LSP_TARGET_CFG_UNIT_TIMEOUT
logic [ ( 32 ) - 1 : 0] hqm_lsp_target_cfg_unit_version_status ; //I HQM_LSP_TARGET_CFG_UNIT_VERSION
hqm_lsp_pipe_register_pfcsr i_hqm_lsp_pipe_register_pfcsr (
  .hqm_gated_clk ( hqm_gated_clk ) 
, .hqm_gated_rst_n ( hqm_gated_rst_n ) 
, .rst_prep ( '0 )
, .cfg_req_write ( pfcsr_cfg_req_write )
, .cfg_req_read ( pfcsr_cfg_req_read )
, .cfg_req ( pfcsr_cfg_req )
, .cfg_rsp_ack ( pfcsr_cfg_rsp_ack )
, .cfg_rsp_err ( pfcsr_cfg_rsp_err )
, .cfg_rsp_rdata ( pfcsr_cfg_rsp_rdata )
, .pfcsr_shadow_nxt ( pfcsr_shadow_nxt )
, .pfcsr_shadow_f ( pfcsr_shadow_f )
, .hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_nxt ( hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_nxt )
, .hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_f ( hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_f )
, .hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_nxt ( hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_nxt )
, .hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_f ( hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_f )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_nxt ( hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_nxt )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_f ( hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_f )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_v (  hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_v )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_nxt ( hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_nxt )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_f ( hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_f )
, .hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_v (  hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_v )
, .hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_nxt ( hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_nxt )
, .hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_f ( hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_f )
, .hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_v (  hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_v )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_nxt ( hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_nxt )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_f ( hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_f )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_v (  hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_v )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_nxt ( hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_nxt )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_f ( hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_f )
, .hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_v (  hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_v )
, .hqm_lsp_target_cfg_cnt_win_cos0_en ( hqm_lsp_target_cfg_cnt_win_cos0_en )
, .hqm_lsp_target_cfg_cnt_win_cos0_clr ( hqm_lsp_target_cfg_cnt_win_cos0_clr )
, .hqm_lsp_target_cfg_cnt_win_cos0_clrv ( hqm_lsp_target_cfg_cnt_win_cos0_clrv )
, .hqm_lsp_target_cfg_cnt_win_cos0_inc ( hqm_lsp_target_cfg_cnt_win_cos0_inc )
, .hqm_lsp_target_cfg_cnt_win_cos0_count ( hqm_lsp_target_cfg_cnt_win_cos0_count )
, .hqm_lsp_target_cfg_cnt_win_cos1_en ( hqm_lsp_target_cfg_cnt_win_cos1_en )
, .hqm_lsp_target_cfg_cnt_win_cos1_clr ( hqm_lsp_target_cfg_cnt_win_cos1_clr )
, .hqm_lsp_target_cfg_cnt_win_cos1_clrv ( hqm_lsp_target_cfg_cnt_win_cos1_clrv )
, .hqm_lsp_target_cfg_cnt_win_cos1_inc ( hqm_lsp_target_cfg_cnt_win_cos1_inc )
, .hqm_lsp_target_cfg_cnt_win_cos1_count ( hqm_lsp_target_cfg_cnt_win_cos1_count )
, .hqm_lsp_target_cfg_cnt_win_cos2_en ( hqm_lsp_target_cfg_cnt_win_cos2_en )
, .hqm_lsp_target_cfg_cnt_win_cos2_clr ( hqm_lsp_target_cfg_cnt_win_cos2_clr )
, .hqm_lsp_target_cfg_cnt_win_cos2_clrv ( hqm_lsp_target_cfg_cnt_win_cos2_clrv )
, .hqm_lsp_target_cfg_cnt_win_cos2_inc ( hqm_lsp_target_cfg_cnt_win_cos2_inc )
, .hqm_lsp_target_cfg_cnt_win_cos2_count ( hqm_lsp_target_cfg_cnt_win_cos2_count )
, .hqm_lsp_target_cfg_cnt_win_cos3_en ( hqm_lsp_target_cfg_cnt_win_cos3_en )
, .hqm_lsp_target_cfg_cnt_win_cos3_clr ( hqm_lsp_target_cfg_cnt_win_cos3_clr )
, .hqm_lsp_target_cfg_cnt_win_cos3_clrv ( hqm_lsp_target_cfg_cnt_win_cos3_clrv )
, .hqm_lsp_target_cfg_cnt_win_cos3_inc ( hqm_lsp_target_cfg_cnt_win_cos3_inc )
, .hqm_lsp_target_cfg_cnt_win_cos3_count ( hqm_lsp_target_cfg_cnt_win_cos3_count )
, .hqm_lsp_target_cfg_control_general_0_reg_nxt ( hqm_lsp_target_cfg_control_general_0_reg_nxt )
, .hqm_lsp_target_cfg_control_general_0_reg_f ( hqm_lsp_target_cfg_control_general_0_reg_f )
, .hqm_lsp_target_cfg_control_general_0_reg_v (  hqm_lsp_target_cfg_control_general_0_reg_v )
, .hqm_lsp_target_cfg_control_general_1_reg_nxt ( hqm_lsp_target_cfg_control_general_1_reg_nxt )
, .hqm_lsp_target_cfg_control_general_1_reg_f ( hqm_lsp_target_cfg_control_general_1_reg_f )
, .hqm_lsp_target_cfg_control_general_1_reg_v (  hqm_lsp_target_cfg_control_general_1_reg_v )
, .hqm_lsp_target_cfg_control_pipeline_credits_reg_nxt ( hqm_lsp_target_cfg_control_pipeline_credits_reg_nxt )
, .hqm_lsp_target_cfg_control_pipeline_credits_reg_f ( hqm_lsp_target_cfg_control_pipeline_credits_reg_f )
, .hqm_lsp_target_cfg_control_pipeline_credits_reg_v (  hqm_lsp_target_cfg_control_pipeline_credits_reg_v )
, .hqm_lsp_target_cfg_control_sched_slot_count_reg_nxt ( hqm_lsp_target_cfg_control_sched_slot_count_reg_nxt )
, .hqm_lsp_target_cfg_control_sched_slot_count_reg_f ( hqm_lsp_target_cfg_control_sched_slot_count_reg_f )
, .hqm_lsp_target_cfg_control_sched_slot_count_reg_v (  hqm_lsp_target_cfg_control_sched_slot_count_reg_v )
, .hqm_lsp_target_cfg_cos_ctrl_reg_nxt ( hqm_lsp_target_cfg_cos_ctrl_reg_nxt )
, .hqm_lsp_target_cfg_cos_ctrl_reg_f ( hqm_lsp_target_cfg_cos_ctrl_reg_f )
, .hqm_lsp_target_cfg_cos_ctrl_reg_v (  hqm_lsp_target_cfg_cos_ctrl_reg_v )
, .hqm_lsp_target_cfg_cq_dir_disable_reg_load ( hqm_lsp_target_cfg_cq_dir_disable_reg_load )
, .hqm_lsp_target_cfg_cq_dir_disable_reg_nxt ( hqm_lsp_target_cfg_cq_dir_disable_reg_nxt )
, .hqm_lsp_target_cfg_cq_dir_disable_reg_f ( hqm_lsp_target_cfg_cq_dir_disable_reg_f )
, .hqm_lsp_target_cfg_cq_ldb_disable_reg_load ( hqm_lsp_target_cfg_cq_ldb_disable_reg_load )
, .hqm_lsp_target_cfg_cq_ldb_disable_reg_nxt ( hqm_lsp_target_cfg_cq_ldb_disable_reg_nxt )
, .hqm_lsp_target_cfg_cq_ldb_disable_reg_f ( hqm_lsp_target_cfg_cq_ldb_disable_reg_f )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_en ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_en )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clr ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clr )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clrv ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clrv )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_inc ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_inc )
, .hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count ( hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count )
, .hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_nxt ( hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_nxt )
, .hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_f ( hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_f )
, .hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_nxt ( hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_nxt )
, .hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_f ( hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_f )
, .hqm_lsp_target_cfg_credit_cnt_cos0_reg_nxt ( hqm_lsp_target_cfg_credit_cnt_cos0_reg_nxt )
, .hqm_lsp_target_cfg_credit_cnt_cos0_reg_f ( hqm_lsp_target_cfg_credit_cnt_cos0_reg_f )
, .hqm_lsp_target_cfg_credit_cnt_cos1_reg_nxt ( hqm_lsp_target_cfg_credit_cnt_cos1_reg_nxt )
, .hqm_lsp_target_cfg_credit_cnt_cos1_reg_f ( hqm_lsp_target_cfg_credit_cnt_cos1_reg_f )
, .hqm_lsp_target_cfg_credit_cnt_cos2_reg_nxt ( hqm_lsp_target_cfg_credit_cnt_cos2_reg_nxt )
, .hqm_lsp_target_cfg_credit_cnt_cos2_reg_f ( hqm_lsp_target_cfg_credit_cnt_cos2_reg_f )
, .hqm_lsp_target_cfg_credit_cnt_cos3_reg_nxt ( hqm_lsp_target_cfg_credit_cnt_cos3_reg_nxt )
, .hqm_lsp_target_cfg_credit_cnt_cos3_reg_f ( hqm_lsp_target_cfg_credit_cnt_cos3_reg_f )
, .hqm_lsp_target_cfg_credit_sat_cos0_reg_nxt ( hqm_lsp_target_cfg_credit_sat_cos0_reg_nxt )
, .hqm_lsp_target_cfg_credit_sat_cos0_reg_f ( hqm_lsp_target_cfg_credit_sat_cos0_reg_f )
, .hqm_lsp_target_cfg_credit_sat_cos0_reg_v (  hqm_lsp_target_cfg_credit_sat_cos0_reg_v )
, .hqm_lsp_target_cfg_credit_sat_cos1_reg_nxt ( hqm_lsp_target_cfg_credit_sat_cos1_reg_nxt )
, .hqm_lsp_target_cfg_credit_sat_cos1_reg_f ( hqm_lsp_target_cfg_credit_sat_cos1_reg_f )
, .hqm_lsp_target_cfg_credit_sat_cos1_reg_v (  hqm_lsp_target_cfg_credit_sat_cos1_reg_v )
, .hqm_lsp_target_cfg_credit_sat_cos2_reg_nxt ( hqm_lsp_target_cfg_credit_sat_cos2_reg_nxt )
, .hqm_lsp_target_cfg_credit_sat_cos2_reg_f ( hqm_lsp_target_cfg_credit_sat_cos2_reg_f )
, .hqm_lsp_target_cfg_credit_sat_cos2_reg_v (  hqm_lsp_target_cfg_credit_sat_cos2_reg_v )
, .hqm_lsp_target_cfg_credit_sat_cos3_reg_nxt ( hqm_lsp_target_cfg_credit_sat_cos3_reg_nxt )
, .hqm_lsp_target_cfg_credit_sat_cos3_reg_f ( hqm_lsp_target_cfg_credit_sat_cos3_reg_f )
, .hqm_lsp_target_cfg_credit_sat_cos3_reg_v (  hqm_lsp_target_cfg_credit_sat_cos3_reg_v )
, .hqm_lsp_target_cfg_diagnostic_aw_status_status ( hqm_lsp_target_cfg_diagnostic_aw_status_status )
, .hqm_lsp_target_cfg_diagnostic_status_0_status ( hqm_lsp_target_cfg_diagnostic_status_0_status )
, .hqm_lsp_target_cfg_error_inject_reg_nxt ( hqm_lsp_target_cfg_error_inject_reg_nxt )
, .hqm_lsp_target_cfg_error_inject_reg_f ( hqm_lsp_target_cfg_error_inject_reg_f )
, .hqm_lsp_target_cfg_error_inject_reg_v (  hqm_lsp_target_cfg_error_inject_reg_v )
, .hqm_lsp_target_cfg_fid_inflight_count_reg_nxt ( hqm_lsp_target_cfg_fid_inflight_count_reg_nxt )
, .hqm_lsp_target_cfg_fid_inflight_count_reg_f ( hqm_lsp_target_cfg_fid_inflight_count_reg_f )
, .hqm_lsp_target_cfg_fid_inflight_limit_reg_nxt ( hqm_lsp_target_cfg_fid_inflight_limit_reg_nxt )
, .hqm_lsp_target_cfg_fid_inflight_limit_reg_f ( hqm_lsp_target_cfg_fid_inflight_limit_reg_f )
, .hqm_lsp_target_cfg_hw_agitate_control_reg_nxt ( hqm_lsp_target_cfg_hw_agitate_control_reg_nxt )
, .hqm_lsp_target_cfg_hw_agitate_control_reg_f ( hqm_lsp_target_cfg_hw_agitate_control_reg_f )
, .hqm_lsp_target_cfg_hw_agitate_control_reg_v (  hqm_lsp_target_cfg_hw_agitate_control_reg_v )
, .hqm_lsp_target_cfg_hw_agitate_select_reg_nxt ( hqm_lsp_target_cfg_hw_agitate_select_reg_nxt )
, .hqm_lsp_target_cfg_hw_agitate_select_reg_f ( hqm_lsp_target_cfg_hw_agitate_select_reg_f )
, .hqm_lsp_target_cfg_hw_agitate_select_reg_v (  hqm_lsp_target_cfg_hw_agitate_select_reg_v )
, .hqm_lsp_target_cfg_interface_status_reg_nxt ( hqm_lsp_target_cfg_interface_status_reg_nxt )
, .hqm_lsp_target_cfg_interface_status_reg_f ( hqm_lsp_target_cfg_interface_status_reg_f )
, .hqm_lsp_target_cfg_ldb_sched_control_reg_nxt ( hqm_lsp_target_cfg_ldb_sched_control_reg_nxt )
, .hqm_lsp_target_cfg_ldb_sched_control_reg_f ( hqm_lsp_target_cfg_ldb_sched_control_reg_f )
, .hqm_lsp_target_cfg_ldb_sched_perf_0_en ( hqm_lsp_target_cfg_ldb_sched_perf_0_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_0_clr ( hqm_lsp_target_cfg_ldb_sched_perf_0_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_0_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_0_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_0_inc ( hqm_lsp_target_cfg_ldb_sched_perf_0_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_0_count ( hqm_lsp_target_cfg_ldb_sched_perf_0_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_1_en ( hqm_lsp_target_cfg_ldb_sched_perf_1_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_1_clr ( hqm_lsp_target_cfg_ldb_sched_perf_1_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_1_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_1_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_1_inc ( hqm_lsp_target_cfg_ldb_sched_perf_1_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_1_count ( hqm_lsp_target_cfg_ldb_sched_perf_1_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_2_en ( hqm_lsp_target_cfg_ldb_sched_perf_2_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_2_clr ( hqm_lsp_target_cfg_ldb_sched_perf_2_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_2_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_2_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_2_inc ( hqm_lsp_target_cfg_ldb_sched_perf_2_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_2_count ( hqm_lsp_target_cfg_ldb_sched_perf_2_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_3_en ( hqm_lsp_target_cfg_ldb_sched_perf_3_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_3_clr ( hqm_lsp_target_cfg_ldb_sched_perf_3_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_3_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_3_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_3_inc ( hqm_lsp_target_cfg_ldb_sched_perf_3_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_3_count ( hqm_lsp_target_cfg_ldb_sched_perf_3_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_4_en ( hqm_lsp_target_cfg_ldb_sched_perf_4_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_4_clr ( hqm_lsp_target_cfg_ldb_sched_perf_4_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_4_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_4_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_4_inc ( hqm_lsp_target_cfg_ldb_sched_perf_4_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_4_count ( hqm_lsp_target_cfg_ldb_sched_perf_4_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_5_en ( hqm_lsp_target_cfg_ldb_sched_perf_5_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_5_clr ( hqm_lsp_target_cfg_ldb_sched_perf_5_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_5_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_5_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_5_inc ( hqm_lsp_target_cfg_ldb_sched_perf_5_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_5_count ( hqm_lsp_target_cfg_ldb_sched_perf_5_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_6_en ( hqm_lsp_target_cfg_ldb_sched_perf_6_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_6_clr ( hqm_lsp_target_cfg_ldb_sched_perf_6_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_6_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_6_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_6_inc ( hqm_lsp_target_cfg_ldb_sched_perf_6_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_6_count ( hqm_lsp_target_cfg_ldb_sched_perf_6_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_7_en ( hqm_lsp_target_cfg_ldb_sched_perf_7_en )
, .hqm_lsp_target_cfg_ldb_sched_perf_7_clr ( hqm_lsp_target_cfg_ldb_sched_perf_7_clr )
, .hqm_lsp_target_cfg_ldb_sched_perf_7_clrv ( hqm_lsp_target_cfg_ldb_sched_perf_7_clrv )
, .hqm_lsp_target_cfg_ldb_sched_perf_7_inc ( hqm_lsp_target_cfg_ldb_sched_perf_7_inc )
, .hqm_lsp_target_cfg_ldb_sched_perf_7_count ( hqm_lsp_target_cfg_ldb_sched_perf_7_count )
, .hqm_lsp_target_cfg_ldb_sched_perf_control_reg_nxt ( hqm_lsp_target_cfg_ldb_sched_perf_control_reg_nxt )
, .hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f ( hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f )
, .hqm_lsp_target_cfg_ldb_sched_perf_control_reg_v (  hqm_lsp_target_cfg_ldb_sched_perf_control_reg_v )
, .hqm_lsp_target_cfg_lsp_csr_control_reg_nxt ( hqm_lsp_target_cfg_lsp_csr_control_reg_nxt )
, .hqm_lsp_target_cfg_lsp_csr_control_reg_f ( hqm_lsp_target_cfg_lsp_csr_control_reg_f )
, .hqm_lsp_target_cfg_lsp_csr_control_reg_v (  hqm_lsp_target_cfg_lsp_csr_control_reg_v )
, .hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_nxt ( hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_nxt )
, .hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_f ( hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_f )
, .hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_nxt ( hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_nxt )
, .hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_f ( hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_f )
, .hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_en ( hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_en )
, .hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clr ( hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clr )
, .hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clrv ( hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clrv )
, .hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_inc ( hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_inc )
, .hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count ( hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count )
, .hqm_lsp_target_cfg_patch_control_reg_nxt ( hqm_lsp_target_cfg_patch_control_reg_nxt )
, .hqm_lsp_target_cfg_patch_control_reg_f ( hqm_lsp_target_cfg_patch_control_reg_f )
, .hqm_lsp_target_cfg_patch_control_reg_v (  hqm_lsp_target_cfg_patch_control_reg_v )
, .hqm_lsp_target_cfg_pipe_health_hold_00_status ( hqm_lsp_target_cfg_pipe_health_hold_00_status )
, .hqm_lsp_target_cfg_pipe_health_hold_01_status ( hqm_lsp_target_cfg_pipe_health_hold_01_status )
, .hqm_lsp_target_cfg_pipe_health_valid_00_status ( hqm_lsp_target_cfg_pipe_health_valid_00_status )
, .hqm_lsp_target_cfg_pipe_health_valid_01_status ( hqm_lsp_target_cfg_pipe_health_valid_01_status )
, .hqm_lsp_target_cfg_rdy_cos0_en ( hqm_lsp_target_cfg_rdy_cos0_en )
, .hqm_lsp_target_cfg_rdy_cos0_clr ( hqm_lsp_target_cfg_rdy_cos0_clr )
, .hqm_lsp_target_cfg_rdy_cos0_clrv ( hqm_lsp_target_cfg_rdy_cos0_clrv )
, .hqm_lsp_target_cfg_rdy_cos0_inc ( hqm_lsp_target_cfg_rdy_cos0_inc )
, .hqm_lsp_target_cfg_rdy_cos0_count ( hqm_lsp_target_cfg_rdy_cos0_count )
, .hqm_lsp_target_cfg_rdy_cos1_en ( hqm_lsp_target_cfg_rdy_cos1_en )
, .hqm_lsp_target_cfg_rdy_cos1_clr ( hqm_lsp_target_cfg_rdy_cos1_clr )
, .hqm_lsp_target_cfg_rdy_cos1_clrv ( hqm_lsp_target_cfg_rdy_cos1_clrv )
, .hqm_lsp_target_cfg_rdy_cos1_inc ( hqm_lsp_target_cfg_rdy_cos1_inc )
, .hqm_lsp_target_cfg_rdy_cos1_count ( hqm_lsp_target_cfg_rdy_cos1_count )
, .hqm_lsp_target_cfg_rdy_cos2_en ( hqm_lsp_target_cfg_rdy_cos2_en )
, .hqm_lsp_target_cfg_rdy_cos2_clr ( hqm_lsp_target_cfg_rdy_cos2_clr )
, .hqm_lsp_target_cfg_rdy_cos2_clrv ( hqm_lsp_target_cfg_rdy_cos2_clrv )
, .hqm_lsp_target_cfg_rdy_cos2_inc ( hqm_lsp_target_cfg_rdy_cos2_inc )
, .hqm_lsp_target_cfg_rdy_cos2_count ( hqm_lsp_target_cfg_rdy_cos2_count )
, .hqm_lsp_target_cfg_rdy_cos3_en ( hqm_lsp_target_cfg_rdy_cos3_en )
, .hqm_lsp_target_cfg_rdy_cos3_clr ( hqm_lsp_target_cfg_rdy_cos3_clr )
, .hqm_lsp_target_cfg_rdy_cos3_clrv ( hqm_lsp_target_cfg_rdy_cos3_clrv )
, .hqm_lsp_target_cfg_rdy_cos3_inc ( hqm_lsp_target_cfg_rdy_cos3_inc )
, .hqm_lsp_target_cfg_rdy_cos3_count ( hqm_lsp_target_cfg_rdy_cos3_count )
, .hqm_lsp_target_cfg_rnd_loss_cos0_en ( hqm_lsp_target_cfg_rnd_loss_cos0_en )
, .hqm_lsp_target_cfg_rnd_loss_cos0_clr ( hqm_lsp_target_cfg_rnd_loss_cos0_clr )
, .hqm_lsp_target_cfg_rnd_loss_cos0_clrv ( hqm_lsp_target_cfg_rnd_loss_cos0_clrv )
, .hqm_lsp_target_cfg_rnd_loss_cos0_inc ( hqm_lsp_target_cfg_rnd_loss_cos0_inc )
, .hqm_lsp_target_cfg_rnd_loss_cos0_count ( hqm_lsp_target_cfg_rnd_loss_cos0_count )
, .hqm_lsp_target_cfg_rnd_loss_cos1_en ( hqm_lsp_target_cfg_rnd_loss_cos1_en )
, .hqm_lsp_target_cfg_rnd_loss_cos1_clr ( hqm_lsp_target_cfg_rnd_loss_cos1_clr )
, .hqm_lsp_target_cfg_rnd_loss_cos1_clrv ( hqm_lsp_target_cfg_rnd_loss_cos1_clrv )
, .hqm_lsp_target_cfg_rnd_loss_cos1_inc ( hqm_lsp_target_cfg_rnd_loss_cos1_inc )
, .hqm_lsp_target_cfg_rnd_loss_cos1_count ( hqm_lsp_target_cfg_rnd_loss_cos1_count )
, .hqm_lsp_target_cfg_rnd_loss_cos2_en ( hqm_lsp_target_cfg_rnd_loss_cos2_en )
, .hqm_lsp_target_cfg_rnd_loss_cos2_clr ( hqm_lsp_target_cfg_rnd_loss_cos2_clr )
, .hqm_lsp_target_cfg_rnd_loss_cos2_clrv ( hqm_lsp_target_cfg_rnd_loss_cos2_clrv )
, .hqm_lsp_target_cfg_rnd_loss_cos2_inc ( hqm_lsp_target_cfg_rnd_loss_cos2_inc )
, .hqm_lsp_target_cfg_rnd_loss_cos2_count ( hqm_lsp_target_cfg_rnd_loss_cos2_count )
, .hqm_lsp_target_cfg_rnd_loss_cos3_en ( hqm_lsp_target_cfg_rnd_loss_cos3_en )
, .hqm_lsp_target_cfg_rnd_loss_cos3_clr ( hqm_lsp_target_cfg_rnd_loss_cos3_clr )
, .hqm_lsp_target_cfg_rnd_loss_cos3_clrv ( hqm_lsp_target_cfg_rnd_loss_cos3_clrv )
, .hqm_lsp_target_cfg_rnd_loss_cos3_inc ( hqm_lsp_target_cfg_rnd_loss_cos3_inc )
, .hqm_lsp_target_cfg_rnd_loss_cos3_count ( hqm_lsp_target_cfg_rnd_loss_cos3_count )
, .hqm_lsp_target_cfg_schd_cos0_en ( hqm_lsp_target_cfg_schd_cos0_en )
, .hqm_lsp_target_cfg_schd_cos0_clr ( hqm_lsp_target_cfg_schd_cos0_clr )
, .hqm_lsp_target_cfg_schd_cos0_clrv ( hqm_lsp_target_cfg_schd_cos0_clrv )
, .hqm_lsp_target_cfg_schd_cos0_inc ( hqm_lsp_target_cfg_schd_cos0_inc )
, .hqm_lsp_target_cfg_schd_cos0_count ( hqm_lsp_target_cfg_schd_cos0_count )
, .hqm_lsp_target_cfg_schd_cos1_en ( hqm_lsp_target_cfg_schd_cos1_en )
, .hqm_lsp_target_cfg_schd_cos1_clr ( hqm_lsp_target_cfg_schd_cos1_clr )
, .hqm_lsp_target_cfg_schd_cos1_clrv ( hqm_lsp_target_cfg_schd_cos1_clrv )
, .hqm_lsp_target_cfg_schd_cos1_inc ( hqm_lsp_target_cfg_schd_cos1_inc )
, .hqm_lsp_target_cfg_schd_cos1_count ( hqm_lsp_target_cfg_schd_cos1_count )
, .hqm_lsp_target_cfg_schd_cos2_en ( hqm_lsp_target_cfg_schd_cos2_en )
, .hqm_lsp_target_cfg_schd_cos2_clr ( hqm_lsp_target_cfg_schd_cos2_clr )
, .hqm_lsp_target_cfg_schd_cos2_clrv ( hqm_lsp_target_cfg_schd_cos2_clrv )
, .hqm_lsp_target_cfg_schd_cos2_inc ( hqm_lsp_target_cfg_schd_cos2_inc )
, .hqm_lsp_target_cfg_schd_cos2_count ( hqm_lsp_target_cfg_schd_cos2_count )
, .hqm_lsp_target_cfg_schd_cos3_en ( hqm_lsp_target_cfg_schd_cos3_en )
, .hqm_lsp_target_cfg_schd_cos3_clr ( hqm_lsp_target_cfg_schd_cos3_clr )
, .hqm_lsp_target_cfg_schd_cos3_clrv ( hqm_lsp_target_cfg_schd_cos3_clrv )
, .hqm_lsp_target_cfg_schd_cos3_inc ( hqm_lsp_target_cfg_schd_cos3_inc )
, .hqm_lsp_target_cfg_schd_cos3_count ( hqm_lsp_target_cfg_schd_cos3_count )
, .hqm_lsp_target_cfg_sch_rdy_en ( hqm_lsp_target_cfg_sch_rdy_en )
, .hqm_lsp_target_cfg_sch_rdy_clr ( hqm_lsp_target_cfg_sch_rdy_clr )
, .hqm_lsp_target_cfg_sch_rdy_clrv ( hqm_lsp_target_cfg_sch_rdy_clrv )
, .hqm_lsp_target_cfg_sch_rdy_inc ( hqm_lsp_target_cfg_sch_rdy_inc )
, .hqm_lsp_target_cfg_sch_rdy_count ( hqm_lsp_target_cfg_sch_rdy_count )
, .hqm_lsp_target_cfg_shdw_ctrl_reg_nxt ( hqm_lsp_target_cfg_shdw_ctrl_reg_nxt )
, .hqm_lsp_target_cfg_shdw_ctrl_reg_f ( hqm_lsp_target_cfg_shdw_ctrl_reg_f )
, .hqm_lsp_target_cfg_shdw_range_cos0_reg_nxt ( hqm_lsp_target_cfg_shdw_range_cos0_reg_nxt )
, .hqm_lsp_target_cfg_shdw_range_cos0_reg_f ( hqm_lsp_target_cfg_shdw_range_cos0_reg_f )
, .hqm_lsp_target_cfg_shdw_range_cos0_reg_v (  hqm_lsp_target_cfg_shdw_range_cos0_reg_v )
, .hqm_lsp_target_cfg_shdw_range_cos1_reg_nxt ( hqm_lsp_target_cfg_shdw_range_cos1_reg_nxt )
, .hqm_lsp_target_cfg_shdw_range_cos1_reg_f ( hqm_lsp_target_cfg_shdw_range_cos1_reg_f )
, .hqm_lsp_target_cfg_shdw_range_cos1_reg_v (  hqm_lsp_target_cfg_shdw_range_cos1_reg_v )
, .hqm_lsp_target_cfg_shdw_range_cos2_reg_nxt ( hqm_lsp_target_cfg_shdw_range_cos2_reg_nxt )
, .hqm_lsp_target_cfg_shdw_range_cos2_reg_f ( hqm_lsp_target_cfg_shdw_range_cos2_reg_f )
, .hqm_lsp_target_cfg_shdw_range_cos2_reg_v (  hqm_lsp_target_cfg_shdw_range_cos2_reg_v )
, .hqm_lsp_target_cfg_shdw_range_cos3_reg_nxt ( hqm_lsp_target_cfg_shdw_range_cos3_reg_nxt )
, .hqm_lsp_target_cfg_shdw_range_cos3_reg_f ( hqm_lsp_target_cfg_shdw_range_cos3_reg_f )
, .hqm_lsp_target_cfg_shdw_range_cos3_reg_v (  hqm_lsp_target_cfg_shdw_range_cos3_reg_v )
, .hqm_lsp_target_cfg_smon0_disable_smon ( hqm_lsp_target_cfg_smon0_disable_smon )
, .hqm_lsp_target_cfg_smon0_smon_v ( hqm_lsp_target_cfg_smon0_smon_v )
, .hqm_lsp_target_cfg_smon0_smon_comp ( hqm_lsp_target_cfg_smon0_smon_comp )
, .hqm_lsp_target_cfg_smon0_smon_val ( hqm_lsp_target_cfg_smon0_smon_val )
, .hqm_lsp_target_cfg_smon0_smon_enabled ( hqm_lsp_target_cfg_smon0_smon_enabled )
, .hqm_lsp_target_cfg_smon0_smon_interrupt ( hqm_lsp_target_cfg_smon0_smon_interrupt )
, .hqm_lsp_target_cfg_syndrome_hw_capture_v ( hqm_lsp_target_cfg_syndrome_hw_capture_v )
, .hqm_lsp_target_cfg_syndrome_hw_capture_data ( hqm_lsp_target_cfg_syndrome_hw_capture_data )
, .hqm_lsp_target_cfg_syndrome_hw_syndrome_data ( hqm_lsp_target_cfg_syndrome_hw_syndrome_data )
, .hqm_lsp_target_cfg_syndrome_sw_capture_v ( hqm_lsp_target_cfg_syndrome_sw_capture_v )
, .hqm_lsp_target_cfg_syndrome_sw_capture_data ( hqm_lsp_target_cfg_syndrome_sw_capture_data )
, .hqm_lsp_target_cfg_syndrome_sw_syndrome_data ( hqm_lsp_target_cfg_syndrome_sw_syndrome_data )
, .hqm_lsp_target_cfg_unit_idle_reg_nxt ( hqm_lsp_target_cfg_unit_idle_reg_nxt )
, .hqm_lsp_target_cfg_unit_idle_reg_f ( hqm_lsp_target_cfg_unit_idle_reg_f )
, .hqm_lsp_target_cfg_unit_timeout_reg_nxt ( hqm_lsp_target_cfg_unit_timeout_reg_nxt )
, .hqm_lsp_target_cfg_unit_timeout_reg_f ( hqm_lsp_target_cfg_unit_timeout_reg_f )
, .hqm_lsp_target_cfg_unit_version_status ( hqm_lsp_target_cfg_unit_version_status )
) ;
// END HQM_CFG_ACCESS
//---------------------------------------------------------------------------------------------------------
// BEGIN HQM_RAM_ACCESS
localparam NUM_CFG_ACCESSIBLE_RAM = 34;
localparam CFG_ACCESSIBLE_RAM_CFG_ATM_QID_DPTH_THRSH_MEM = 0; // HQM_LSP_TARGET_CFG_ATM_QID_DPTH_THRSH
localparam CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM = 1; // HQM_LSP_TARGET_CFG_CQ2PRIOV
localparam CFG_ACCESSIBLE_RAM_CFG_QID_AQED_ACTIVE_LIMIT_MEM = 10; // HQM_LSP_TARGET_CFG_QID_AQED_ACTIVE_LIMIT
localparam CFG_ACCESSIBLE_RAM_CFG_QID_LDB_INFLIGHT_LIMIT_MEM = 11; // HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_LIMIT
localparam CFG_ACCESSIBLE_RAM_CFG_QID_LDB_QID2CQIDIX2_MEM = 12; // HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_00 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_01 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_02 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_03 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_04 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_05 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_06 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_07 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_08 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_09 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_10 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_11 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_12 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_13 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_14 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_15
localparam CFG_ACCESSIBLE_RAM_CFG_QID_LDB_QID2CQIDIX_MEM = 13; // HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_00 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_01 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_02 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_03 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_04 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_05 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_06 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_07 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_08 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_09 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_10 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_11 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_12 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_13 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_14 HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_15
localparam CFG_ACCESSIBLE_RAM_CQ_DIR_TOT_SCH_CNT_MEM = 14; // HQM_LSP_TARGET_CFG_CQ_DIR_TOT_SCH_CNTH HQM_LSP_TARGET_CFG_CQ_DIR_TOT_SCH_CNTL
localparam CFG_ACCESSIBLE_RAM_CQ_LDB_INFLIGHT_COUNT_MEM = 15; // HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_COUNT
localparam CFG_ACCESSIBLE_RAM_CQ_LDB_TOKEN_COUNT_MEM = 16; // HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_COUNT
localparam CFG_ACCESSIBLE_RAM_CQ_LDB_TOT_SCH_CNT_MEM = 17; // HQM_LSP_TARGET_CFG_CQ_LDB_TOT_SCH_CNTH HQM_LSP_TARGET_CFG_CQ_LDB_TOT_SCH_CNTL
localparam CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM = 18; // HQM_LSP_TARGET_CFG_CQ_LDB_WU_COUNT
localparam CFG_ACCESSIBLE_RAM_DIR_ENQ_CNT_MEM = 19; // HQM_LSP_TARGET_CFG_QID_DIR_ENQUEUE_COUNT
localparam CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM = 2; // HQM_LSP_TARGET_CFG_CQ2QID0
localparam CFG_ACCESSIBLE_RAM_DIR_TOK_CNT_MEM = 20; // HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_COUNT
localparam CFG_ACCESSIBLE_RAM_DIR_TOK_LIM_MEM = 21; // HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_DEPTH_SELECT_DSI
localparam CFG_ACCESSIBLE_RAM_QID_AQED_ACTIVE_COUNT_MEM = 22; // HQM_LSP_TARGET_CFG_QID_AQED_ACTIVE_COUNT
localparam CFG_ACCESSIBLE_RAM_QID_ATM_ACTIVE_MEM = 23; // HQM_LSP_TARGET_CFG_QID_ATM_ACTIVE
localparam CFG_ACCESSIBLE_RAM_QID_ATM_TOT_ENQ_CNT_MEM = 24; // HQM_LSP_TARGET_CFG_QID_ATM_TOT_ENQ_CNTH HQM_LSP_TARGET_CFG_QID_ATM_TOT_ENQ_CNTL
localparam CFG_ACCESSIBLE_RAM_QID_ATQ_ENQUEUE_COUNT_MEM = 25; // HQM_LSP_TARGET_CFG_QID_ATQ_ENQUEUE_COUNT
localparam CFG_ACCESSIBLE_RAM_QID_DIR_MAX_DEPTH_MEM = 26; // HQM_LSP_TARGET_CFG_QID_DIR_MAX_DEPTH
localparam CFG_ACCESSIBLE_RAM_QID_DIR_REPLAY_COUNT_MEM = 27; // HQM_LSP_TARGET_CFG_QID_DIR_REPLAY_COUNT
localparam CFG_ACCESSIBLE_RAM_QID_DIR_TOT_ENQ_CNT_MEM = 28; // HQM_LSP_TARGET_CFG_QID_DIR_TOT_ENQ_CNTH HQM_LSP_TARGET_CFG_QID_DIR_TOT_ENQ_CNTL
localparam CFG_ACCESSIBLE_RAM_QID_LDB_ENQUEUE_COUNT_MEM = 29; // HQM_LSP_TARGET_CFG_QID_LDB_ENQUEUE_COUNT
localparam CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM = 3; // HQM_LSP_TARGET_CFG_CQ2QID1
localparam CFG_ACCESSIBLE_RAM_QID_LDB_INFLIGHT_COUNT_MEM = 30; // HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_COUNT
localparam CFG_ACCESSIBLE_RAM_QID_LDB_REPLAY_COUNT_MEM = 31; // HQM_LSP_TARGET_CFG_QID_LDB_REPLAY_COUNT
localparam CFG_ACCESSIBLE_RAM_QID_NALDB_MAX_DEPTH_MEM = 32; // HQM_LSP_TARGET_CFG_QID_NALDB_MAX_DEPTH
localparam CFG_ACCESSIBLE_RAM_QID_NALDB_TOT_ENQ_CNT_MEM = 33; // HQM_LSP_TARGET_CFG_QID_NALDB_TOT_ENQ_CNTH HQM_LSP_TARGET_CFG_QID_NALDB_TOT_ENQ_CNTL
localparam CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_INFLIGHT_LIMIT_MEM = 4; // HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_LIMIT
localparam CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_INFLIGHT_THRESHOLD_MEM = 5; // HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_THRESHOLD
localparam CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_TOKEN_DEPTH_SELECT_MEM = 6; // HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_DEPTH_SELECT
localparam CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM = 7; // HQM_LSP_TARGET_CFG_CQ_LDB_WU_LIMIT
localparam CFG_ACCESSIBLE_RAM_CFG_DIR_QID_DPTH_THRSH_MEM = 8; // HQM_LSP_TARGET_CFG_DIR_QID_DPTH_THRSH
localparam CFG_ACCESSIBLE_RAM_CFG_NALB_QID_DPTH_THRSH_MEM = 9; // HQM_LSP_TARGET_CFG_NALB_QID_DPTH_THRSH
logic [( 34 *  1)-1:0] cfg_mem_re;
logic [( 34 *  1)-1:0] cfg_mem_we;
logic [(      20)-1:0] cfg_mem_addr;
logic [(      12)-1:0] cfg_mem_minbit;
logic [(      12)-1:0] cfg_mem_maxbit;
logic [(      32)-1:0] cfg_mem_wdata;
logic [( 34 * 32)-1:0] cfg_mem_rdata;
logic [( 34 *  1)-1:0] cfg_mem_ack;
logic                  cfg_mem_cc_v;
logic [(       8)-1:0] cfg_mem_cc_value;
logic [(       4)-1:0] cfg_mem_cc_width;
logic [(      12)-1:0] cfg_mem_cc_position;


logic                  hqm_list_sel_pipe_rfw_top_ipar_error;

logic                  func_aqed_lsp_deq_fifo_mem_re; //I
logic [(       5)-1:0] func_aqed_lsp_deq_fifo_mem_raddr; //I
logic [(       5)-1:0] func_aqed_lsp_deq_fifo_mem_waddr; //I
logic                  func_aqed_lsp_deq_fifo_mem_we;    //I
logic [(       9)-1:0] func_aqed_lsp_deq_fifo_mem_wdata; //I
logic [(       9)-1:0] func_aqed_lsp_deq_fifo_mem_rdata;

logic                pf_aqed_lsp_deq_fifo_mem_re;    //I
logic [(       5)-1:0] pf_aqed_lsp_deq_fifo_mem_raddr; //I
logic [(       5)-1:0] pf_aqed_lsp_deq_fifo_mem_waddr; //I
logic                  pf_aqed_lsp_deq_fifo_mem_we;    //I
logic [(       9)-1:0] pf_aqed_lsp_deq_fifo_mem_wdata; //I
logic [(       9)-1:0] pf_aqed_lsp_deq_fifo_mem_rdata;

logic                  rf_aqed_lsp_deq_fifo_mem_error;

logic                  func_atm_cmp_fifo_mem_re; //I
logic [(       3)-1:0] func_atm_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] func_atm_cmp_fifo_mem_waddr; //I
logic                  func_atm_cmp_fifo_mem_we;    //I
logic [(      55)-1:0] func_atm_cmp_fifo_mem_wdata; //I
logic [(      55)-1:0] func_atm_cmp_fifo_mem_rdata;

logic                pf_atm_cmp_fifo_mem_re;    //I
logic [(       3)-1:0] pf_atm_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] pf_atm_cmp_fifo_mem_waddr; //I
logic                  pf_atm_cmp_fifo_mem_we;    //I
logic [(      55)-1:0] pf_atm_cmp_fifo_mem_wdata; //I
logic [(      55)-1:0] pf_atm_cmp_fifo_mem_rdata;

logic                  rf_atm_cmp_fifo_mem_error;

logic                  func_cfg_atm_qid_dpth_thrsh_mem_re; //I
logic [(       7)-1:0] func_cfg_atm_qid_dpth_thrsh_mem_addr; //I
logic                  func_cfg_atm_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] func_cfg_atm_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] func_cfg_atm_qid_dpth_thrsh_mem_rdata;

logic                pf_cfg_atm_qid_dpth_thrsh_mem_re;    //I
logic [(       7)-1:0] pf_cfg_atm_qid_dpth_thrsh_mem_addr;  //I
logic                  pf_cfg_atm_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] pf_cfg_atm_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] pf_cfg_atm_qid_dpth_thrsh_mem_rdata;

logic                  rf_cfg_atm_qid_dpth_thrsh_mem_error;

logic                  func_cfg_cq2priov_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2priov_mem_addr; //I
logic                  func_cfg_cq2priov_mem_we;    //I
logic [(      33)-1:0] func_cfg_cq2priov_mem_wdata; //I
logic [(      33)-1:0] func_cfg_cq2priov_mem_rdata;

logic                pf_cfg_cq2priov_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2priov_mem_addr;  //I
logic                  pf_cfg_cq2priov_mem_we;    //I
logic [(      33)-1:0] pf_cfg_cq2priov_mem_wdata; //I
logic [(      33)-1:0] pf_cfg_cq2priov_mem_rdata;

logic                  rf_cfg_cq2priov_mem_error;

logic                  func_cfg_cq2priov_odd_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2priov_odd_mem_addr; //I
logic                  func_cfg_cq2priov_odd_mem_we;    //I
logic [(      33)-1:0] func_cfg_cq2priov_odd_mem_wdata; //I
logic [(      33)-1:0] func_cfg_cq2priov_odd_mem_rdata;

logic                pf_cfg_cq2priov_odd_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2priov_odd_mem_addr;  //I
logic                  pf_cfg_cq2priov_odd_mem_we;    //I
logic [(      33)-1:0] pf_cfg_cq2priov_odd_mem_wdata; //I
logic [(      33)-1:0] pf_cfg_cq2priov_odd_mem_rdata;

logic                  rf_cfg_cq2priov_odd_mem_error;

logic                  func_cfg_cq2qid_0_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2qid_0_mem_addr; //I
logic                  func_cfg_cq2qid_0_mem_we;    //I
logic [(      29)-1:0] func_cfg_cq2qid_0_mem_wdata; //I
logic [(      29)-1:0] func_cfg_cq2qid_0_mem_rdata;

logic                pf_cfg_cq2qid_0_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2qid_0_mem_addr;  //I
logic                  pf_cfg_cq2qid_0_mem_we;    //I
logic [(      29)-1:0] pf_cfg_cq2qid_0_mem_wdata; //I
logic [(      29)-1:0] pf_cfg_cq2qid_0_mem_rdata;

logic                  rf_cfg_cq2qid_0_mem_error;

logic                  func_cfg_cq2qid_0_odd_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2qid_0_odd_mem_addr; //I
logic                  func_cfg_cq2qid_0_odd_mem_we;    //I
logic [(      29)-1:0] func_cfg_cq2qid_0_odd_mem_wdata; //I
logic [(      29)-1:0] func_cfg_cq2qid_0_odd_mem_rdata;

logic                pf_cfg_cq2qid_0_odd_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2qid_0_odd_mem_addr;  //I
logic                  pf_cfg_cq2qid_0_odd_mem_we;    //I
logic [(      29)-1:0] pf_cfg_cq2qid_0_odd_mem_wdata; //I
logic [(      29)-1:0] pf_cfg_cq2qid_0_odd_mem_rdata;

logic                  rf_cfg_cq2qid_0_odd_mem_error;

logic                  func_cfg_cq2qid_1_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2qid_1_mem_addr; //I
logic                  func_cfg_cq2qid_1_mem_we;    //I
logic [(      29)-1:0] func_cfg_cq2qid_1_mem_wdata; //I
logic [(      29)-1:0] func_cfg_cq2qid_1_mem_rdata;

logic                pf_cfg_cq2qid_1_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2qid_1_mem_addr;  //I
logic                  pf_cfg_cq2qid_1_mem_we;    //I
logic [(      29)-1:0] pf_cfg_cq2qid_1_mem_wdata; //I
logic [(      29)-1:0] pf_cfg_cq2qid_1_mem_rdata;

logic                  rf_cfg_cq2qid_1_mem_error;

logic                  func_cfg_cq2qid_1_odd_mem_re; //I
logic [(       5)-1:0] func_cfg_cq2qid_1_odd_mem_addr; //I
logic                  func_cfg_cq2qid_1_odd_mem_we;    //I
logic [(      29)-1:0] func_cfg_cq2qid_1_odd_mem_wdata; //I
logic [(      29)-1:0] func_cfg_cq2qid_1_odd_mem_rdata;

logic                pf_cfg_cq2qid_1_odd_mem_re;    //I
logic [(       5)-1:0] pf_cfg_cq2qid_1_odd_mem_addr;  //I
logic                  pf_cfg_cq2qid_1_odd_mem_we;    //I
logic [(      29)-1:0] pf_cfg_cq2qid_1_odd_mem_wdata; //I
logic [(      29)-1:0] pf_cfg_cq2qid_1_odd_mem_rdata;

logic                  rf_cfg_cq2qid_1_odd_mem_error;

logic                  func_cfg_cq_ldb_inflight_limit_mem_re; //I
logic [(       6)-1:0] func_cfg_cq_ldb_inflight_limit_mem_addr; //I
logic                  func_cfg_cq_ldb_inflight_limit_mem_we;    //I
logic [(      14)-1:0] func_cfg_cq_ldb_inflight_limit_mem_wdata; //I
logic [(      14)-1:0] func_cfg_cq_ldb_inflight_limit_mem_rdata;

logic                pf_cfg_cq_ldb_inflight_limit_mem_re;    //I
logic [(       6)-1:0] pf_cfg_cq_ldb_inflight_limit_mem_addr;  //I
logic                  pf_cfg_cq_ldb_inflight_limit_mem_we;    //I
logic [(      14)-1:0] pf_cfg_cq_ldb_inflight_limit_mem_wdata; //I
logic [(      14)-1:0] pf_cfg_cq_ldb_inflight_limit_mem_rdata;

logic                  rf_cfg_cq_ldb_inflight_limit_mem_error;

logic                  func_cfg_cq_ldb_inflight_threshold_mem_re; //I
logic [(       6)-1:0] func_cfg_cq_ldb_inflight_threshold_mem_addr; //I
logic                  func_cfg_cq_ldb_inflight_threshold_mem_we;    //I
logic [(      14)-1:0] func_cfg_cq_ldb_inflight_threshold_mem_wdata; //I
logic [(      14)-1:0] func_cfg_cq_ldb_inflight_threshold_mem_rdata;

logic                pf_cfg_cq_ldb_inflight_threshold_mem_re;    //I
logic [(       6)-1:0] pf_cfg_cq_ldb_inflight_threshold_mem_addr;  //I
logic                  pf_cfg_cq_ldb_inflight_threshold_mem_we;    //I
logic [(      14)-1:0] pf_cfg_cq_ldb_inflight_threshold_mem_wdata; //I
logic [(      14)-1:0] pf_cfg_cq_ldb_inflight_threshold_mem_rdata;

logic                  rf_cfg_cq_ldb_inflight_threshold_mem_error;

logic                  func_cfg_cq_ldb_token_depth_select_mem_re; //I
logic [(       6)-1:0] func_cfg_cq_ldb_token_depth_select_mem_addr; //I
logic                  func_cfg_cq_ldb_token_depth_select_mem_we;    //I
logic [(       5)-1:0] func_cfg_cq_ldb_token_depth_select_mem_wdata; //I
logic [(       5)-1:0] func_cfg_cq_ldb_token_depth_select_mem_rdata;

logic                pf_cfg_cq_ldb_token_depth_select_mem_re;    //I
logic [(       6)-1:0] pf_cfg_cq_ldb_token_depth_select_mem_addr;  //I
logic                  pf_cfg_cq_ldb_token_depth_select_mem_we;    //I
logic [(       5)-1:0] pf_cfg_cq_ldb_token_depth_select_mem_wdata; //I
logic [(       5)-1:0] pf_cfg_cq_ldb_token_depth_select_mem_rdata;

logic                  rf_cfg_cq_ldb_token_depth_select_mem_error;

logic                  func_cfg_cq_ldb_wu_limit_mem_re; //I
logic [(       6)-1:0] func_cfg_cq_ldb_wu_limit_mem_raddr; //I
logic [(       6)-1:0] func_cfg_cq_ldb_wu_limit_mem_waddr; //I
logic                  func_cfg_cq_ldb_wu_limit_mem_we;    //I
logic [(      17)-1:0] func_cfg_cq_ldb_wu_limit_mem_wdata; //I
logic [(      17)-1:0] func_cfg_cq_ldb_wu_limit_mem_rdata;

logic                pf_cfg_cq_ldb_wu_limit_mem_re;    //I
logic [(       6)-1:0] pf_cfg_cq_ldb_wu_limit_mem_raddr; //I
logic [(       6)-1:0] pf_cfg_cq_ldb_wu_limit_mem_waddr; //I
logic                  pf_cfg_cq_ldb_wu_limit_mem_we;    //I
logic [(      17)-1:0] pf_cfg_cq_ldb_wu_limit_mem_wdata; //I
logic [(      17)-1:0] pf_cfg_cq_ldb_wu_limit_mem_rdata;

logic                  rf_cfg_cq_ldb_wu_limit_mem_error;

logic                  func_cfg_dir_qid_dpth_thrsh_mem_re; //I
logic [(       7)-1:0] func_cfg_dir_qid_dpth_thrsh_mem_addr; //I
logic                  func_cfg_dir_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] func_cfg_dir_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] func_cfg_dir_qid_dpth_thrsh_mem_rdata;

logic                pf_cfg_dir_qid_dpth_thrsh_mem_re;    //I
logic [(       7)-1:0] pf_cfg_dir_qid_dpth_thrsh_mem_addr;  //I
logic                  pf_cfg_dir_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] pf_cfg_dir_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] pf_cfg_dir_qid_dpth_thrsh_mem_rdata;

logic                  rf_cfg_dir_qid_dpth_thrsh_mem_error;

logic                  func_cfg_nalb_qid_dpth_thrsh_mem_re; //I
logic [(       7)-1:0] func_cfg_nalb_qid_dpth_thrsh_mem_addr; //I
logic                  func_cfg_nalb_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] func_cfg_nalb_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] func_cfg_nalb_qid_dpth_thrsh_mem_rdata;

logic                pf_cfg_nalb_qid_dpth_thrsh_mem_re;    //I
logic [(       7)-1:0] pf_cfg_nalb_qid_dpth_thrsh_mem_addr;  //I
logic                  pf_cfg_nalb_qid_dpth_thrsh_mem_we;    //I
logic [(      16)-1:0] pf_cfg_nalb_qid_dpth_thrsh_mem_wdata; //I
logic [(      16)-1:0] pf_cfg_nalb_qid_dpth_thrsh_mem_rdata;

logic                  rf_cfg_nalb_qid_dpth_thrsh_mem_error;

logic                  func_cfg_qid_aqed_active_limit_mem_re; //I
logic [(       7)-1:0] func_cfg_qid_aqed_active_limit_mem_addr; //I
logic                  func_cfg_qid_aqed_active_limit_mem_we;    //I
logic [(      13)-1:0] func_cfg_qid_aqed_active_limit_mem_wdata; //I
logic [(      13)-1:0] func_cfg_qid_aqed_active_limit_mem_rdata;

logic                pf_cfg_qid_aqed_active_limit_mem_re;    //I
logic [(       7)-1:0] pf_cfg_qid_aqed_active_limit_mem_addr;  //I
logic                  pf_cfg_qid_aqed_active_limit_mem_we;    //I
logic [(      13)-1:0] pf_cfg_qid_aqed_active_limit_mem_wdata; //I
logic [(      13)-1:0] pf_cfg_qid_aqed_active_limit_mem_rdata;

logic                  rf_cfg_qid_aqed_active_limit_mem_error;

logic                  func_cfg_qid_ldb_inflight_limit_mem_re; //I
logic [(       7)-1:0] func_cfg_qid_ldb_inflight_limit_mem_addr; //I
logic                  func_cfg_qid_ldb_inflight_limit_mem_we;    //I
logic [(      13)-1:0] func_cfg_qid_ldb_inflight_limit_mem_wdata; //I
logic [(      13)-1:0] func_cfg_qid_ldb_inflight_limit_mem_rdata;

logic                pf_cfg_qid_ldb_inflight_limit_mem_re;    //I
logic [(       7)-1:0] pf_cfg_qid_ldb_inflight_limit_mem_addr;  //I
logic                  pf_cfg_qid_ldb_inflight_limit_mem_we;    //I
logic [(      13)-1:0] pf_cfg_qid_ldb_inflight_limit_mem_wdata; //I
logic [(      13)-1:0] pf_cfg_qid_ldb_inflight_limit_mem_rdata;

logic                  rf_cfg_qid_ldb_inflight_limit_mem_error;

logic                  func_cfg_qid_ldb_qid2cqidix2_mem_re; //I
logic [(       7)-1:0] func_cfg_qid_ldb_qid2cqidix2_mem_addr; //I
logic                  func_cfg_qid_ldb_qid2cqidix2_mem_we;    //I
logic [(     528)-1:0] func_cfg_qid_ldb_qid2cqidix2_mem_wdata; //I
logic [(     528)-1:0] func_cfg_qid_ldb_qid2cqidix2_mem_rdata;

logic                pf_cfg_qid_ldb_qid2cqidix2_mem_re;    //I
logic [(       7)-1:0] pf_cfg_qid_ldb_qid2cqidix2_mem_addr;  //I
logic                  pf_cfg_qid_ldb_qid2cqidix2_mem_we;    //I
logic [(     528)-1:0] pf_cfg_qid_ldb_qid2cqidix2_mem_wdata; //I
logic [(     528)-1:0] pf_cfg_qid_ldb_qid2cqidix2_mem_rdata;

logic                  rf_cfg_qid_ldb_qid2cqidix2_mem_error;

logic                  func_cfg_qid_ldb_qid2cqidix_mem_re; //I
logic [(       7)-1:0] func_cfg_qid_ldb_qid2cqidix_mem_addr; //I
logic                  func_cfg_qid_ldb_qid2cqidix_mem_we;    //I
logic [(     528)-1:0] func_cfg_qid_ldb_qid2cqidix_mem_wdata; //I
logic [(     528)-1:0] func_cfg_qid_ldb_qid2cqidix_mem_rdata;

logic                pf_cfg_qid_ldb_qid2cqidix_mem_re;    //I
logic [(       7)-1:0] pf_cfg_qid_ldb_qid2cqidix_mem_addr;  //I
logic                  pf_cfg_qid_ldb_qid2cqidix_mem_we;    //I
logic [(     528)-1:0] pf_cfg_qid_ldb_qid2cqidix_mem_wdata; //I
logic [(     528)-1:0] pf_cfg_qid_ldb_qid2cqidix_mem_rdata;

logic                  rf_cfg_qid_ldb_qid2cqidix_mem_error;

logic                  func_chp_lsp_cmp_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_chp_lsp_cmp_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_chp_lsp_cmp_rx_sync_fifo_mem_waddr; //I
logic                  func_chp_lsp_cmp_rx_sync_fifo_mem_we;    //I
logic [(      73)-1:0] func_chp_lsp_cmp_rx_sync_fifo_mem_wdata; //I
logic [(      73)-1:0] func_chp_lsp_cmp_rx_sync_fifo_mem_rdata;

logic                pf_chp_lsp_cmp_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_chp_lsp_cmp_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_chp_lsp_cmp_rx_sync_fifo_mem_waddr; //I
logic                  pf_chp_lsp_cmp_rx_sync_fifo_mem_we;    //I
logic [(      73)-1:0] pf_chp_lsp_cmp_rx_sync_fifo_mem_wdata; //I
logic [(      73)-1:0] pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata;

logic                  rf_chp_lsp_cmp_rx_sync_fifo_mem_error;

logic                  func_chp_lsp_token_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_chp_lsp_token_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_chp_lsp_token_rx_sync_fifo_mem_waddr; //I
logic                  func_chp_lsp_token_rx_sync_fifo_mem_we;    //I
logic [(      25)-1:0] func_chp_lsp_token_rx_sync_fifo_mem_wdata; //I
logic [(      25)-1:0] func_chp_lsp_token_rx_sync_fifo_mem_rdata;

logic                pf_chp_lsp_token_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_chp_lsp_token_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_chp_lsp_token_rx_sync_fifo_mem_waddr; //I
logic                  pf_chp_lsp_token_rx_sync_fifo_mem_we;    //I
logic [(      25)-1:0] pf_chp_lsp_token_rx_sync_fifo_mem_wdata; //I
logic [(      25)-1:0] pf_chp_lsp_token_rx_sync_fifo_mem_rdata;

logic                  rf_chp_lsp_token_rx_sync_fifo_mem_error;

logic                  func_cq_atm_pri_arbindex_mem_re; //I
logic [(       5)-1:0] func_cq_atm_pri_arbindex_mem_raddr; //I
logic [(       5)-1:0] func_cq_atm_pri_arbindex_mem_waddr; //I
logic                  func_cq_atm_pri_arbindex_mem_we;    //I
logic [(      96)-1:0] func_cq_atm_pri_arbindex_mem_wdata; //I
logic [(      96)-1:0] func_cq_atm_pri_arbindex_mem_rdata;

logic                pf_cq_atm_pri_arbindex_mem_re;    //I
logic [(       5)-1:0] pf_cq_atm_pri_arbindex_mem_raddr; //I
logic [(       5)-1:0] pf_cq_atm_pri_arbindex_mem_waddr; //I
logic                  pf_cq_atm_pri_arbindex_mem_we;    //I
logic [(      96)-1:0] pf_cq_atm_pri_arbindex_mem_wdata; //I
logic [(      96)-1:0] pf_cq_atm_pri_arbindex_mem_rdata;

logic                  rf_cq_atm_pri_arbindex_mem_error;

logic                  func_cq_dir_tot_sch_cnt_mem_re; //I
logic [(       7)-1:0] func_cq_dir_tot_sch_cnt_mem_raddr; //I
logic [(       7)-1:0] func_cq_dir_tot_sch_cnt_mem_waddr; //I
logic                  func_cq_dir_tot_sch_cnt_mem_we;    //I
logic [(      66)-1:0] func_cq_dir_tot_sch_cnt_mem_wdata; //I
logic [(      66)-1:0] func_cq_dir_tot_sch_cnt_mem_rdata;

logic                pf_cq_dir_tot_sch_cnt_mem_re;    //I
logic [(       7)-1:0] pf_cq_dir_tot_sch_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_cq_dir_tot_sch_cnt_mem_waddr; //I
logic                  pf_cq_dir_tot_sch_cnt_mem_we;    //I
logic [(      66)-1:0] pf_cq_dir_tot_sch_cnt_mem_wdata; //I
logic [(      66)-1:0] pf_cq_dir_tot_sch_cnt_mem_rdata;

logic                  rf_cq_dir_tot_sch_cnt_mem_error;

logic                  func_cq_ldb_inflight_count_mem_re; //I
logic [(       6)-1:0] func_cq_ldb_inflight_count_mem_raddr; //I
logic [(       6)-1:0] func_cq_ldb_inflight_count_mem_waddr; //I
logic                  func_cq_ldb_inflight_count_mem_we;    //I
logic [(      15)-1:0] func_cq_ldb_inflight_count_mem_wdata; //I
logic [(      15)-1:0] func_cq_ldb_inflight_count_mem_rdata;

logic                pf_cq_ldb_inflight_count_mem_re;    //I
logic [(       6)-1:0] pf_cq_ldb_inflight_count_mem_raddr; //I
logic [(       6)-1:0] pf_cq_ldb_inflight_count_mem_waddr; //I
logic                  pf_cq_ldb_inflight_count_mem_we;    //I
logic [(      15)-1:0] pf_cq_ldb_inflight_count_mem_wdata; //I
logic [(      15)-1:0] pf_cq_ldb_inflight_count_mem_rdata;

logic                  rf_cq_ldb_inflight_count_mem_error;

logic                  func_cq_ldb_token_count_mem_re; //I
logic [(       6)-1:0] func_cq_ldb_token_count_mem_raddr; //I
logic [(       6)-1:0] func_cq_ldb_token_count_mem_waddr; //I
logic                  func_cq_ldb_token_count_mem_we;    //I
logic [(      13)-1:0] func_cq_ldb_token_count_mem_wdata; //I
logic [(      13)-1:0] func_cq_ldb_token_count_mem_rdata;

logic                pf_cq_ldb_token_count_mem_re;    //I
logic [(       6)-1:0] pf_cq_ldb_token_count_mem_raddr; //I
logic [(       6)-1:0] pf_cq_ldb_token_count_mem_waddr; //I
logic                  pf_cq_ldb_token_count_mem_we;    //I
logic [(      13)-1:0] pf_cq_ldb_token_count_mem_wdata; //I
logic [(      13)-1:0] pf_cq_ldb_token_count_mem_rdata;

logic                  rf_cq_ldb_token_count_mem_error;

logic                  func_cq_ldb_tot_sch_cnt_mem_re; //I
logic [(       6)-1:0] func_cq_ldb_tot_sch_cnt_mem_raddr; //I
logic [(       6)-1:0] func_cq_ldb_tot_sch_cnt_mem_waddr; //I
logic                  func_cq_ldb_tot_sch_cnt_mem_we;    //I
logic [(      66)-1:0] func_cq_ldb_tot_sch_cnt_mem_wdata; //I
logic [(      66)-1:0] func_cq_ldb_tot_sch_cnt_mem_rdata;

logic                pf_cq_ldb_tot_sch_cnt_mem_re;    //I
logic [(       6)-1:0] pf_cq_ldb_tot_sch_cnt_mem_raddr; //I
logic [(       6)-1:0] pf_cq_ldb_tot_sch_cnt_mem_waddr; //I
logic                  pf_cq_ldb_tot_sch_cnt_mem_we;    //I
logic [(      66)-1:0] pf_cq_ldb_tot_sch_cnt_mem_wdata; //I
logic [(      66)-1:0] pf_cq_ldb_tot_sch_cnt_mem_rdata;

logic                  rf_cq_ldb_tot_sch_cnt_mem_error;

logic                  func_cq_ldb_wu_count_mem_re; //I
logic [(       6)-1:0] func_cq_ldb_wu_count_mem_raddr; //I
logic [(       6)-1:0] func_cq_ldb_wu_count_mem_waddr; //I
logic                  func_cq_ldb_wu_count_mem_we;    //I
logic [(      19)-1:0] func_cq_ldb_wu_count_mem_wdata; //I
logic [(      19)-1:0] func_cq_ldb_wu_count_mem_rdata;

logic                pf_cq_ldb_wu_count_mem_re;    //I
logic [(       6)-1:0] pf_cq_ldb_wu_count_mem_raddr; //I
logic [(       6)-1:0] pf_cq_ldb_wu_count_mem_waddr; //I
logic                  pf_cq_ldb_wu_count_mem_we;    //I
logic [(      19)-1:0] pf_cq_ldb_wu_count_mem_wdata; //I
logic [(      19)-1:0] pf_cq_ldb_wu_count_mem_rdata;

logic                  rf_cq_ldb_wu_count_mem_error;

logic                  func_cq_nalb_pri_arbindex_mem_re; //I
logic [(       5)-1:0] func_cq_nalb_pri_arbindex_mem_raddr; //I
logic [(       5)-1:0] func_cq_nalb_pri_arbindex_mem_waddr; //I
logic                  func_cq_nalb_pri_arbindex_mem_we;    //I
logic [(      96)-1:0] func_cq_nalb_pri_arbindex_mem_wdata; //I
logic [(      96)-1:0] func_cq_nalb_pri_arbindex_mem_rdata;

logic                pf_cq_nalb_pri_arbindex_mem_re;    //I
logic [(       5)-1:0] pf_cq_nalb_pri_arbindex_mem_raddr; //I
logic [(       5)-1:0] pf_cq_nalb_pri_arbindex_mem_waddr; //I
logic                  pf_cq_nalb_pri_arbindex_mem_we;    //I
logic [(      96)-1:0] pf_cq_nalb_pri_arbindex_mem_wdata; //I
logic [(      96)-1:0] pf_cq_nalb_pri_arbindex_mem_rdata;

logic                  rf_cq_nalb_pri_arbindex_mem_error;

logic                  func_dir_enq_cnt_mem_re; //I
logic [(       7)-1:0] func_dir_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] func_dir_enq_cnt_mem_waddr; //I
logic                  func_dir_enq_cnt_mem_we;    //I
logic [(      17)-1:0] func_dir_enq_cnt_mem_wdata; //I
logic [(      17)-1:0] func_dir_enq_cnt_mem_rdata;

logic                pf_dir_enq_cnt_mem_re;    //I
logic [(       7)-1:0] pf_dir_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_dir_enq_cnt_mem_waddr; //I
logic                  pf_dir_enq_cnt_mem_we;    //I
logic [(      17)-1:0] pf_dir_enq_cnt_mem_wdata; //I
logic [(      17)-1:0] pf_dir_enq_cnt_mem_rdata;

logic                  rf_dir_enq_cnt_mem_error;

logic                  func_dir_tok_cnt_mem_re; //I
logic [(       7)-1:0] func_dir_tok_cnt_mem_raddr; //I
logic [(       7)-1:0] func_dir_tok_cnt_mem_waddr; //I
logic                  func_dir_tok_cnt_mem_we;    //I
logic [(      13)-1:0] func_dir_tok_cnt_mem_wdata; //I
logic [(      13)-1:0] func_dir_tok_cnt_mem_rdata;

logic                pf_dir_tok_cnt_mem_re;    //I
logic [(       7)-1:0] pf_dir_tok_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_dir_tok_cnt_mem_waddr; //I
logic                  pf_dir_tok_cnt_mem_we;    //I
logic [(      13)-1:0] pf_dir_tok_cnt_mem_wdata; //I
logic [(      13)-1:0] pf_dir_tok_cnt_mem_rdata;

logic                  rf_dir_tok_cnt_mem_error;

logic                  func_dir_tok_lim_mem_re; //I
logic [(       7)-1:0] func_dir_tok_lim_mem_addr; //I
logic                  func_dir_tok_lim_mem_we;    //I
logic [(       8)-1:0] func_dir_tok_lim_mem_wdata; //I
logic [(       8)-1:0] func_dir_tok_lim_mem_rdata;

logic                pf_dir_tok_lim_mem_re;    //I
logic [(       7)-1:0] pf_dir_tok_lim_mem_addr;  //I
logic                  pf_dir_tok_lim_mem_we;    //I
logic [(       8)-1:0] pf_dir_tok_lim_mem_wdata; //I
logic [(       8)-1:0] pf_dir_tok_lim_mem_rdata;

logic                  rf_dir_tok_lim_mem_error;

logic                  func_dp_lsp_enq_dir_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr; //I
logic                  func_dp_lsp_enq_dir_rx_sync_fifo_mem_we;    //I
logic [(       8)-1:0] func_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata; //I
logic [(       8)-1:0] func_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata;

logic                pf_dp_lsp_enq_dir_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr; //I
logic                  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_we;    //I
logic [(       8)-1:0] pf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata; //I
logic [(       8)-1:0] pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata;

logic                  rf_dp_lsp_enq_dir_rx_sync_fifo_mem_error;

logic                  func_dp_lsp_enq_rorply_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr; //I
logic                  func_dp_lsp_enq_rorply_rx_sync_fifo_mem_we;    //I
logic [(      23)-1:0] func_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata; //I
logic [(      23)-1:0] func_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata;

logic                pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr; //I
logic                  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we;    //I
logic [(      23)-1:0] pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata; //I
logic [(      23)-1:0] pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata;

logic                  rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_error;

logic                  func_enq_nalb_fifo_mem_re; //I
logic [(       2)-1:0] func_enq_nalb_fifo_mem_raddr; //I
logic [(       2)-1:0] func_enq_nalb_fifo_mem_waddr; //I
logic                  func_enq_nalb_fifo_mem_we;    //I
logic [(      10)-1:0] func_enq_nalb_fifo_mem_wdata; //I
logic [(      10)-1:0] func_enq_nalb_fifo_mem_rdata;

logic                pf_enq_nalb_fifo_mem_re;    //I
logic [(       2)-1:0] pf_enq_nalb_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_enq_nalb_fifo_mem_waddr; //I
logic                  pf_enq_nalb_fifo_mem_we;    //I
logic [(      10)-1:0] pf_enq_nalb_fifo_mem_wdata; //I
logic [(      10)-1:0] pf_enq_nalb_fifo_mem_rdata;

logic                  rf_enq_nalb_fifo_mem_error;

logic                  func_ldb_token_rtn_fifo_mem_re; //I
logic [(       3)-1:0] func_ldb_token_rtn_fifo_mem_raddr; //I
logic [(       3)-1:0] func_ldb_token_rtn_fifo_mem_waddr; //I
logic                  func_ldb_token_rtn_fifo_mem_we;    //I
logic [(      25)-1:0] func_ldb_token_rtn_fifo_mem_wdata; //I
logic [(      25)-1:0] func_ldb_token_rtn_fifo_mem_rdata;

logic                pf_ldb_token_rtn_fifo_mem_re;    //I
logic [(       3)-1:0] pf_ldb_token_rtn_fifo_mem_raddr; //I
logic [(       3)-1:0] pf_ldb_token_rtn_fifo_mem_waddr; //I
logic                  pf_ldb_token_rtn_fifo_mem_we;    //I
logic [(      25)-1:0] pf_ldb_token_rtn_fifo_mem_wdata; //I
logic [(      25)-1:0] pf_ldb_token_rtn_fifo_mem_rdata;

logic                  rf_ldb_token_rtn_fifo_mem_error;

logic                  func_nalb_cmp_fifo_mem_re; //I
logic [(       3)-1:0] func_nalb_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] func_nalb_cmp_fifo_mem_waddr; //I
logic                  func_nalb_cmp_fifo_mem_we;    //I
logic [(      18)-1:0] func_nalb_cmp_fifo_mem_wdata; //I
logic [(      18)-1:0] func_nalb_cmp_fifo_mem_rdata;

logic                pf_nalb_cmp_fifo_mem_re;    //I
logic [(       3)-1:0] pf_nalb_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] pf_nalb_cmp_fifo_mem_waddr; //I
logic                  pf_nalb_cmp_fifo_mem_we;    //I
logic [(      18)-1:0] pf_nalb_cmp_fifo_mem_wdata; //I
logic [(      18)-1:0] pf_nalb_cmp_fifo_mem_rdata;

logic                  rf_nalb_cmp_fifo_mem_error;

logic                  func_nalb_lsp_enq_lb_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr; //I
logic                  func_nalb_lsp_enq_lb_rx_sync_fifo_mem_we;    //I
logic [(      10)-1:0] func_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata; //I
logic [(      10)-1:0] func_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata;

logic                pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr; //I
logic                  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we;    //I
logic [(      10)-1:0] pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata; //I
logic [(      10)-1:0] pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata;

logic                  rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_error;

logic                  func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr; //I
logic                  func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we;    //I
logic [(      27)-1:0] func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata; //I
logic [(      27)-1:0] func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata;

logic                pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr; //I
logic                  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we;    //I
logic [(      27)-1:0] pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata; //I
logic [(      27)-1:0] pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata;

logic                  rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_error;

logic                  func_nalb_sel_nalb_fifo_mem_re; //I
logic [(       4)-1:0] func_nalb_sel_nalb_fifo_mem_raddr; //I
logic [(       4)-1:0] func_nalb_sel_nalb_fifo_mem_waddr; //I
logic                  func_nalb_sel_nalb_fifo_mem_we;    //I
logic [(      27)-1:0] func_nalb_sel_nalb_fifo_mem_wdata; //I
logic [(      27)-1:0] func_nalb_sel_nalb_fifo_mem_rdata;

logic                pf_nalb_sel_nalb_fifo_mem_re;    //I
logic [(       4)-1:0] pf_nalb_sel_nalb_fifo_mem_raddr; //I
logic [(       4)-1:0] pf_nalb_sel_nalb_fifo_mem_waddr; //I
logic                  pf_nalb_sel_nalb_fifo_mem_we;    //I
logic [(      27)-1:0] pf_nalb_sel_nalb_fifo_mem_wdata; //I
logic [(      27)-1:0] pf_nalb_sel_nalb_fifo_mem_rdata;

logic                  rf_nalb_sel_nalb_fifo_mem_error;

logic                  func_qed_lsp_deq_fifo_mem_re; //I
logic [(       5)-1:0] func_qed_lsp_deq_fifo_mem_raddr; //I
logic [(       5)-1:0] func_qed_lsp_deq_fifo_mem_waddr; //I
logic                  func_qed_lsp_deq_fifo_mem_we;    //I
logic [(       9)-1:0] func_qed_lsp_deq_fifo_mem_wdata; //I
logic [(       9)-1:0] func_qed_lsp_deq_fifo_mem_rdata;

logic                pf_qed_lsp_deq_fifo_mem_re;    //I
logic [(       5)-1:0] pf_qed_lsp_deq_fifo_mem_raddr; //I
logic [(       5)-1:0] pf_qed_lsp_deq_fifo_mem_waddr; //I
logic                  pf_qed_lsp_deq_fifo_mem_we;    //I
logic [(       9)-1:0] pf_qed_lsp_deq_fifo_mem_wdata; //I
logic [(       9)-1:0] pf_qed_lsp_deq_fifo_mem_rdata;

logic                  rf_qed_lsp_deq_fifo_mem_error;

logic                  func_qid_aqed_active_count_mem_re; //I
logic [(       7)-1:0] func_qid_aqed_active_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_aqed_active_count_mem_waddr; //I
logic                  func_qid_aqed_active_count_mem_we;    //I
logic [(      14)-1:0] func_qid_aqed_active_count_mem_wdata; //I
logic [(      14)-1:0] func_qid_aqed_active_count_mem_rdata;

logic                pf_qid_aqed_active_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_aqed_active_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_aqed_active_count_mem_waddr; //I
logic                  pf_qid_aqed_active_count_mem_we;    //I
logic [(      14)-1:0] pf_qid_aqed_active_count_mem_wdata; //I
logic [(      14)-1:0] pf_qid_aqed_active_count_mem_rdata;

logic                  rf_qid_aqed_active_count_mem_error;

logic                  func_qid_atm_active_mem_re; //I
logic [(       7)-1:0] func_qid_atm_active_mem_raddr; //I
logic [(       7)-1:0] func_qid_atm_active_mem_waddr; //I
logic                  func_qid_atm_active_mem_we;    //I
logic [(      17)-1:0] func_qid_atm_active_mem_wdata; //I
logic [(      17)-1:0] func_qid_atm_active_mem_rdata;

logic                pf_qid_atm_active_mem_re;    //I
logic [(       7)-1:0] pf_qid_atm_active_mem_raddr; //I
logic [(       7)-1:0] pf_qid_atm_active_mem_waddr; //I
logic                  pf_qid_atm_active_mem_we;    //I
logic [(      17)-1:0] pf_qid_atm_active_mem_wdata; //I
logic [(      17)-1:0] pf_qid_atm_active_mem_rdata;

logic                  rf_qid_atm_active_mem_error;

logic                  func_qid_atm_tot_enq_cnt_mem_re; //I
logic [(       7)-1:0] func_qid_atm_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] func_qid_atm_tot_enq_cnt_mem_waddr; //I
logic                  func_qid_atm_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] func_qid_atm_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] func_qid_atm_tot_enq_cnt_mem_rdata;

logic                pf_qid_atm_tot_enq_cnt_mem_re;    //I
logic [(       7)-1:0] pf_qid_atm_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_qid_atm_tot_enq_cnt_mem_waddr; //I
logic                  pf_qid_atm_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] pf_qid_atm_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] pf_qid_atm_tot_enq_cnt_mem_rdata;

logic                  rf_qid_atm_tot_enq_cnt_mem_error;

logic                  func_qid_atq_enqueue_count_mem_re; //I
logic [(       7)-1:0] func_qid_atq_enqueue_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_atq_enqueue_count_mem_waddr; //I
logic                  func_qid_atq_enqueue_count_mem_we;    //I
logic [(      17)-1:0] func_qid_atq_enqueue_count_mem_wdata; //I
logic [(      17)-1:0] func_qid_atq_enqueue_count_mem_rdata;

logic                pf_qid_atq_enqueue_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_atq_enqueue_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_atq_enqueue_count_mem_waddr; //I
logic                  pf_qid_atq_enqueue_count_mem_we;    //I
logic [(      17)-1:0] pf_qid_atq_enqueue_count_mem_wdata; //I
logic [(      17)-1:0] pf_qid_atq_enqueue_count_mem_rdata;

logic                  rf_qid_atq_enqueue_count_mem_error;

logic                  func_qid_dir_max_depth_mem_re; //I
logic [(       7)-1:0] func_qid_dir_max_depth_mem_raddr; //I
logic [(       7)-1:0] func_qid_dir_max_depth_mem_waddr; //I
logic                  func_qid_dir_max_depth_mem_we;    //I
logic [(      15)-1:0] func_qid_dir_max_depth_mem_wdata; //I
logic [(      15)-1:0] func_qid_dir_max_depth_mem_rdata;

logic                pf_qid_dir_max_depth_mem_re;    //I
logic [(       7)-1:0] pf_qid_dir_max_depth_mem_raddr; //I
logic [(       7)-1:0] pf_qid_dir_max_depth_mem_waddr; //I
logic                  pf_qid_dir_max_depth_mem_we;    //I
logic [(      15)-1:0] pf_qid_dir_max_depth_mem_wdata; //I
logic [(      15)-1:0] pf_qid_dir_max_depth_mem_rdata;

logic                  rf_qid_dir_max_depth_mem_error;

logic                  func_qid_dir_replay_count_mem_re; //I
logic [(       7)-1:0] func_qid_dir_replay_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_dir_replay_count_mem_waddr; //I
logic                  func_qid_dir_replay_count_mem_we;    //I
logic [(      17)-1:0] func_qid_dir_replay_count_mem_wdata; //I
logic [(      17)-1:0] func_qid_dir_replay_count_mem_rdata;

logic                pf_qid_dir_replay_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_dir_replay_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_dir_replay_count_mem_waddr; //I
logic                  pf_qid_dir_replay_count_mem_we;    //I
logic [(      17)-1:0] pf_qid_dir_replay_count_mem_wdata; //I
logic [(      17)-1:0] pf_qid_dir_replay_count_mem_rdata;

logic                  rf_qid_dir_replay_count_mem_error;

logic                  func_qid_dir_tot_enq_cnt_mem_re; //I
logic [(       7)-1:0] func_qid_dir_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] func_qid_dir_tot_enq_cnt_mem_waddr; //I
logic                  func_qid_dir_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] func_qid_dir_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] func_qid_dir_tot_enq_cnt_mem_rdata;

logic                pf_qid_dir_tot_enq_cnt_mem_re;    //I
logic [(       7)-1:0] pf_qid_dir_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_qid_dir_tot_enq_cnt_mem_waddr; //I
logic                  pf_qid_dir_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] pf_qid_dir_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] pf_qid_dir_tot_enq_cnt_mem_rdata;

logic                  rf_qid_dir_tot_enq_cnt_mem_error;

logic                  func_qid_ldb_enqueue_count_mem_re; //I
logic [(       7)-1:0] func_qid_ldb_enqueue_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_ldb_enqueue_count_mem_waddr; //I
logic                  func_qid_ldb_enqueue_count_mem_we;    //I
logic [(      17)-1:0] func_qid_ldb_enqueue_count_mem_wdata; //I
logic [(      17)-1:0] func_qid_ldb_enqueue_count_mem_rdata;

logic                pf_qid_ldb_enqueue_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_ldb_enqueue_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_ldb_enqueue_count_mem_waddr; //I
logic                  pf_qid_ldb_enqueue_count_mem_we;    //I
logic [(      17)-1:0] pf_qid_ldb_enqueue_count_mem_wdata; //I
logic [(      17)-1:0] pf_qid_ldb_enqueue_count_mem_rdata;

logic                  rf_qid_ldb_enqueue_count_mem_error;

logic                  func_qid_ldb_inflight_count_mem_re; //I
logic [(       7)-1:0] func_qid_ldb_inflight_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_ldb_inflight_count_mem_waddr; //I
logic                  func_qid_ldb_inflight_count_mem_we;    //I
logic [(      14)-1:0] func_qid_ldb_inflight_count_mem_wdata; //I
logic [(      14)-1:0] func_qid_ldb_inflight_count_mem_rdata;

logic                pf_qid_ldb_inflight_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_ldb_inflight_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_ldb_inflight_count_mem_waddr; //I
logic                  pf_qid_ldb_inflight_count_mem_we;    //I
logic [(      14)-1:0] pf_qid_ldb_inflight_count_mem_wdata; //I
logic [(      14)-1:0] pf_qid_ldb_inflight_count_mem_rdata;

logic                  rf_qid_ldb_inflight_count_mem_error;

logic                  func_qid_ldb_replay_count_mem_re; //I
logic [(       7)-1:0] func_qid_ldb_replay_count_mem_raddr; //I
logic [(       7)-1:0] func_qid_ldb_replay_count_mem_waddr; //I
logic                  func_qid_ldb_replay_count_mem_we;    //I
logic [(      17)-1:0] func_qid_ldb_replay_count_mem_wdata; //I
logic [(      17)-1:0] func_qid_ldb_replay_count_mem_rdata;

logic                pf_qid_ldb_replay_count_mem_re;    //I
logic [(       7)-1:0] pf_qid_ldb_replay_count_mem_raddr; //I
logic [(       7)-1:0] pf_qid_ldb_replay_count_mem_waddr; //I
logic                  pf_qid_ldb_replay_count_mem_we;    //I
logic [(      17)-1:0] pf_qid_ldb_replay_count_mem_wdata; //I
logic [(      17)-1:0] pf_qid_ldb_replay_count_mem_rdata;

logic                  rf_qid_ldb_replay_count_mem_error;

logic                  func_qid_naldb_max_depth_mem_re; //I
logic [(       7)-1:0] func_qid_naldb_max_depth_mem_raddr; //I
logic [(       7)-1:0] func_qid_naldb_max_depth_mem_waddr; //I
logic                  func_qid_naldb_max_depth_mem_we;    //I
logic [(      15)-1:0] func_qid_naldb_max_depth_mem_wdata; //I
logic [(      15)-1:0] func_qid_naldb_max_depth_mem_rdata;

logic                pf_qid_naldb_max_depth_mem_re;    //I
logic [(       7)-1:0] pf_qid_naldb_max_depth_mem_raddr; //I
logic [(       7)-1:0] pf_qid_naldb_max_depth_mem_waddr; //I
logic                  pf_qid_naldb_max_depth_mem_we;    //I
logic [(      15)-1:0] pf_qid_naldb_max_depth_mem_wdata; //I
logic [(      15)-1:0] pf_qid_naldb_max_depth_mem_rdata;

logic                  rf_qid_naldb_max_depth_mem_error;

logic                  func_qid_naldb_tot_enq_cnt_mem_re; //I
logic [(       7)-1:0] func_qid_naldb_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] func_qid_naldb_tot_enq_cnt_mem_waddr; //I
logic                  func_qid_naldb_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] func_qid_naldb_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] func_qid_naldb_tot_enq_cnt_mem_rdata;

logic                pf_qid_naldb_tot_enq_cnt_mem_re;    //I
logic [(       7)-1:0] pf_qid_naldb_tot_enq_cnt_mem_raddr; //I
logic [(       7)-1:0] pf_qid_naldb_tot_enq_cnt_mem_waddr; //I
logic                  pf_qid_naldb_tot_enq_cnt_mem_we;    //I
logic [(      66)-1:0] pf_qid_naldb_tot_enq_cnt_mem_wdata; //I
logic [(      66)-1:0] pf_qid_naldb_tot_enq_cnt_mem_rdata;

logic                  rf_qid_naldb_tot_enq_cnt_mem_error;

logic                  func_rop_lsp_reordercmp_rx_sync_fifo_mem_re; //I
logic [(       3)-1:0] func_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr; //I
logic [(       3)-1:0] func_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr; //I
logic                  func_rop_lsp_reordercmp_rx_sync_fifo_mem_we;    //I
logic [(      17)-1:0] func_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata; //I
logic [(      17)-1:0] func_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata;

logic                pf_rop_lsp_reordercmp_rx_sync_fifo_mem_re;    //I
logic [(       3)-1:0] pf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr; //I
logic [(       3)-1:0] pf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr; //I
logic                  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_we;    //I
logic [(      17)-1:0] pf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata; //I
logic [(      17)-1:0] pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata;

logic                  rf_rop_lsp_reordercmp_rx_sync_fifo_mem_error;

logic                  func_send_atm_to_cq_rx_sync_fifo_mem_re; //I
logic [(       2)-1:0] func_send_atm_to_cq_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] func_send_atm_to_cq_rx_sync_fifo_mem_waddr; //I
logic                  func_send_atm_to_cq_rx_sync_fifo_mem_we;    //I
logic [(      35)-1:0] func_send_atm_to_cq_rx_sync_fifo_mem_wdata; //I
logic [(      35)-1:0] func_send_atm_to_cq_rx_sync_fifo_mem_rdata;

logic                pf_send_atm_to_cq_rx_sync_fifo_mem_re;    //I
logic [(       2)-1:0] pf_send_atm_to_cq_rx_sync_fifo_mem_raddr; //I
logic [(       2)-1:0] pf_send_atm_to_cq_rx_sync_fifo_mem_waddr; //I
logic                  pf_send_atm_to_cq_rx_sync_fifo_mem_we;    //I
logic [(      35)-1:0] pf_send_atm_to_cq_rx_sync_fifo_mem_wdata; //I
logic [(      35)-1:0] pf_send_atm_to_cq_rx_sync_fifo_mem_rdata;

logic                  rf_send_atm_to_cq_rx_sync_fifo_mem_error;

logic                  func_uno_atm_cmp_fifo_mem_re; //I
logic [(       3)-1:0] func_uno_atm_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] func_uno_atm_cmp_fifo_mem_waddr; //I
logic                  func_uno_atm_cmp_fifo_mem_we;    //I
logic [(      20)-1:0] func_uno_atm_cmp_fifo_mem_wdata; //I
logic [(      20)-1:0] func_uno_atm_cmp_fifo_mem_rdata;

logic                pf_uno_atm_cmp_fifo_mem_re;    //I
logic [(       3)-1:0] pf_uno_atm_cmp_fifo_mem_raddr; //I
logic [(       3)-1:0] pf_uno_atm_cmp_fifo_mem_waddr; //I
logic                  pf_uno_atm_cmp_fifo_mem_we;    //I
logic [(      20)-1:0] pf_uno_atm_cmp_fifo_mem_wdata; //I
logic [(      20)-1:0] pf_uno_atm_cmp_fifo_mem_rdata;

logic                  rf_uno_atm_cmp_fifo_mem_error;

hqm_list_sel_pipe_ram_access i_hqm_list_sel_pipe_ram_access (
  .hqm_gated_clk (hqm_gated_clk)
, .hqm_inp_gated_clk (hqm_inp_gated_clk)
, .hqm_gated_rst_n (hqm_gated_rst_n)
, .hqm_inp_gated_rst_n (hqm_inp_gated_rst_n)
,.cfg_mem_re          (cfg_mem_re)
,.cfg_mem_we          (cfg_mem_we)
,.cfg_mem_addr        (cfg_mem_addr)
,.cfg_mem_minbit      (cfg_mem_minbit)
,.cfg_mem_maxbit      (cfg_mem_maxbit)
,.cfg_mem_wdata       (cfg_mem_wdata)
,.cfg_mem_rdata       (cfg_mem_rdata)
,.cfg_mem_ack         (cfg_mem_ack)
,.cfg_mem_cc_v        (cfg_mem_cc_v)
,.cfg_mem_cc_value    (cfg_mem_cc_value)
,.cfg_mem_cc_width    (cfg_mem_cc_width)
,.cfg_mem_cc_position (cfg_mem_cc_position)

,.hqm_list_sel_pipe_rfw_top_ipar_error (hqm_list_sel_pipe_rfw_top_ipar_error)

,.func_aqed_lsp_deq_fifo_mem_re    (func_aqed_lsp_deq_fifo_mem_re)
,.func_aqed_lsp_deq_fifo_mem_raddr (func_aqed_lsp_deq_fifo_mem_raddr)
,.func_aqed_lsp_deq_fifo_mem_waddr (func_aqed_lsp_deq_fifo_mem_waddr)
,.func_aqed_lsp_deq_fifo_mem_we    (func_aqed_lsp_deq_fifo_mem_we)
,.func_aqed_lsp_deq_fifo_mem_wdata (func_aqed_lsp_deq_fifo_mem_wdata)
,.func_aqed_lsp_deq_fifo_mem_rdata (func_aqed_lsp_deq_fifo_mem_rdata)

,.pf_aqed_lsp_deq_fifo_mem_re      (pf_aqed_lsp_deq_fifo_mem_re)
,.pf_aqed_lsp_deq_fifo_mem_raddr (pf_aqed_lsp_deq_fifo_mem_raddr)
,.pf_aqed_lsp_deq_fifo_mem_waddr (pf_aqed_lsp_deq_fifo_mem_waddr)
,.pf_aqed_lsp_deq_fifo_mem_we    (pf_aqed_lsp_deq_fifo_mem_we)
,.pf_aqed_lsp_deq_fifo_mem_wdata (pf_aqed_lsp_deq_fifo_mem_wdata)
,.pf_aqed_lsp_deq_fifo_mem_rdata (pf_aqed_lsp_deq_fifo_mem_rdata)

,.rf_aqed_lsp_deq_fifo_mem_rclk (rf_aqed_lsp_deq_fifo_mem_rclk)
,.rf_aqed_lsp_deq_fifo_mem_rclk_rst_n (rf_aqed_lsp_deq_fifo_mem_rclk_rst_n)
,.rf_aqed_lsp_deq_fifo_mem_re    (rf_aqed_lsp_deq_fifo_mem_re)
,.rf_aqed_lsp_deq_fifo_mem_raddr (rf_aqed_lsp_deq_fifo_mem_raddr)
,.rf_aqed_lsp_deq_fifo_mem_waddr (rf_aqed_lsp_deq_fifo_mem_waddr)
,.rf_aqed_lsp_deq_fifo_mem_wclk (rf_aqed_lsp_deq_fifo_mem_wclk)
,.rf_aqed_lsp_deq_fifo_mem_wclk_rst_n (rf_aqed_lsp_deq_fifo_mem_wclk_rst_n)
,.rf_aqed_lsp_deq_fifo_mem_we    (rf_aqed_lsp_deq_fifo_mem_we)
,.rf_aqed_lsp_deq_fifo_mem_wdata (rf_aqed_lsp_deq_fifo_mem_wdata)
,.rf_aqed_lsp_deq_fifo_mem_rdata (rf_aqed_lsp_deq_fifo_mem_rdata)

,.rf_aqed_lsp_deq_fifo_mem_error (rf_aqed_lsp_deq_fifo_mem_error)

,.func_atm_cmp_fifo_mem_re    (func_atm_cmp_fifo_mem_re)
,.func_atm_cmp_fifo_mem_raddr (func_atm_cmp_fifo_mem_raddr)
,.func_atm_cmp_fifo_mem_waddr (func_atm_cmp_fifo_mem_waddr)
,.func_atm_cmp_fifo_mem_we    (func_atm_cmp_fifo_mem_we)
,.func_atm_cmp_fifo_mem_wdata (func_atm_cmp_fifo_mem_wdata)
,.func_atm_cmp_fifo_mem_rdata (func_atm_cmp_fifo_mem_rdata)

,.pf_atm_cmp_fifo_mem_re      (pf_atm_cmp_fifo_mem_re)
,.pf_atm_cmp_fifo_mem_raddr (pf_atm_cmp_fifo_mem_raddr)
,.pf_atm_cmp_fifo_mem_waddr (pf_atm_cmp_fifo_mem_waddr)
,.pf_atm_cmp_fifo_mem_we    (pf_atm_cmp_fifo_mem_we)
,.pf_atm_cmp_fifo_mem_wdata (pf_atm_cmp_fifo_mem_wdata)
,.pf_atm_cmp_fifo_mem_rdata (pf_atm_cmp_fifo_mem_rdata)

,.rf_atm_cmp_fifo_mem_rclk (rf_atm_cmp_fifo_mem_rclk)
,.rf_atm_cmp_fifo_mem_rclk_rst_n (rf_atm_cmp_fifo_mem_rclk_rst_n)
,.rf_atm_cmp_fifo_mem_re    (rf_atm_cmp_fifo_mem_re)
,.rf_atm_cmp_fifo_mem_raddr (rf_atm_cmp_fifo_mem_raddr)
,.rf_atm_cmp_fifo_mem_waddr (rf_atm_cmp_fifo_mem_waddr)
,.rf_atm_cmp_fifo_mem_wclk (rf_atm_cmp_fifo_mem_wclk)
,.rf_atm_cmp_fifo_mem_wclk_rst_n (rf_atm_cmp_fifo_mem_wclk_rst_n)
,.rf_atm_cmp_fifo_mem_we    (rf_atm_cmp_fifo_mem_we)
,.rf_atm_cmp_fifo_mem_wdata (rf_atm_cmp_fifo_mem_wdata)
,.rf_atm_cmp_fifo_mem_rdata (rf_atm_cmp_fifo_mem_rdata)

,.rf_atm_cmp_fifo_mem_error (rf_atm_cmp_fifo_mem_error)

,.func_cfg_atm_qid_dpth_thrsh_mem_re    (func_cfg_atm_qid_dpth_thrsh_mem_re)
,.func_cfg_atm_qid_dpth_thrsh_mem_addr  (func_cfg_atm_qid_dpth_thrsh_mem_addr)
,.func_cfg_atm_qid_dpth_thrsh_mem_we    (func_cfg_atm_qid_dpth_thrsh_mem_we)
,.func_cfg_atm_qid_dpth_thrsh_mem_wdata (func_cfg_atm_qid_dpth_thrsh_mem_wdata)
,.func_cfg_atm_qid_dpth_thrsh_mem_rdata (func_cfg_atm_qid_dpth_thrsh_mem_rdata)

,.pf_cfg_atm_qid_dpth_thrsh_mem_re      (pf_cfg_atm_qid_dpth_thrsh_mem_re)
,.pf_cfg_atm_qid_dpth_thrsh_mem_addr  (pf_cfg_atm_qid_dpth_thrsh_mem_addr)
,.pf_cfg_atm_qid_dpth_thrsh_mem_we    (pf_cfg_atm_qid_dpth_thrsh_mem_we)
,.pf_cfg_atm_qid_dpth_thrsh_mem_wdata (pf_cfg_atm_qid_dpth_thrsh_mem_wdata)
,.pf_cfg_atm_qid_dpth_thrsh_mem_rdata (pf_cfg_atm_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_atm_qid_dpth_thrsh_mem_rclk (rf_cfg_atm_qid_dpth_thrsh_mem_rclk)
,.rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n (rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n)
,.rf_cfg_atm_qid_dpth_thrsh_mem_re    (rf_cfg_atm_qid_dpth_thrsh_mem_re)
,.rf_cfg_atm_qid_dpth_thrsh_mem_raddr (rf_cfg_atm_qid_dpth_thrsh_mem_raddr)
,.rf_cfg_atm_qid_dpth_thrsh_mem_waddr (rf_cfg_atm_qid_dpth_thrsh_mem_waddr)
,.rf_cfg_atm_qid_dpth_thrsh_mem_wclk (rf_cfg_atm_qid_dpth_thrsh_mem_wclk)
,.rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n (rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n)
,.rf_cfg_atm_qid_dpth_thrsh_mem_we    (rf_cfg_atm_qid_dpth_thrsh_mem_we)
,.rf_cfg_atm_qid_dpth_thrsh_mem_wdata (rf_cfg_atm_qid_dpth_thrsh_mem_wdata)
,.rf_cfg_atm_qid_dpth_thrsh_mem_rdata (rf_cfg_atm_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_atm_qid_dpth_thrsh_mem_error (rf_cfg_atm_qid_dpth_thrsh_mem_error)

,.func_cfg_cq2priov_mem_re    (func_cfg_cq2priov_mem_re)
,.func_cfg_cq2priov_mem_addr  (func_cfg_cq2priov_mem_addr)
,.func_cfg_cq2priov_mem_we    (func_cfg_cq2priov_mem_we)
,.func_cfg_cq2priov_mem_wdata (func_cfg_cq2priov_mem_wdata)
,.func_cfg_cq2priov_mem_rdata (func_cfg_cq2priov_mem_rdata)

,.pf_cfg_cq2priov_mem_re      (pf_cfg_cq2priov_mem_re)
,.pf_cfg_cq2priov_mem_addr  (pf_cfg_cq2priov_mem_addr)
,.pf_cfg_cq2priov_mem_we    (pf_cfg_cq2priov_mem_we)
,.pf_cfg_cq2priov_mem_wdata (pf_cfg_cq2priov_mem_wdata)
,.pf_cfg_cq2priov_mem_rdata (pf_cfg_cq2priov_mem_rdata)

,.rf_cfg_cq2priov_mem_rclk (rf_cfg_cq2priov_mem_rclk)
,.rf_cfg_cq2priov_mem_rclk_rst_n (rf_cfg_cq2priov_mem_rclk_rst_n)
,.rf_cfg_cq2priov_mem_re    (rf_cfg_cq2priov_mem_re)
,.rf_cfg_cq2priov_mem_raddr (rf_cfg_cq2priov_mem_raddr)
,.rf_cfg_cq2priov_mem_waddr (rf_cfg_cq2priov_mem_waddr)
,.rf_cfg_cq2priov_mem_wclk (rf_cfg_cq2priov_mem_wclk)
,.rf_cfg_cq2priov_mem_wclk_rst_n (rf_cfg_cq2priov_mem_wclk_rst_n)
,.rf_cfg_cq2priov_mem_we    (rf_cfg_cq2priov_mem_we)
,.rf_cfg_cq2priov_mem_wdata (rf_cfg_cq2priov_mem_wdata)
,.rf_cfg_cq2priov_mem_rdata (rf_cfg_cq2priov_mem_rdata)

,.rf_cfg_cq2priov_mem_error (rf_cfg_cq2priov_mem_error)

,.func_cfg_cq2priov_odd_mem_re    (func_cfg_cq2priov_odd_mem_re)
,.func_cfg_cq2priov_odd_mem_addr  (func_cfg_cq2priov_odd_mem_addr)
,.func_cfg_cq2priov_odd_mem_we    (func_cfg_cq2priov_odd_mem_we)
,.func_cfg_cq2priov_odd_mem_wdata (func_cfg_cq2priov_odd_mem_wdata)
,.func_cfg_cq2priov_odd_mem_rdata (func_cfg_cq2priov_odd_mem_rdata)

,.pf_cfg_cq2priov_odd_mem_re      (pf_cfg_cq2priov_odd_mem_re)
,.pf_cfg_cq2priov_odd_mem_addr  (pf_cfg_cq2priov_odd_mem_addr)
,.pf_cfg_cq2priov_odd_mem_we    (pf_cfg_cq2priov_odd_mem_we)
,.pf_cfg_cq2priov_odd_mem_wdata (pf_cfg_cq2priov_odd_mem_wdata)
,.pf_cfg_cq2priov_odd_mem_rdata (pf_cfg_cq2priov_odd_mem_rdata)

,.rf_cfg_cq2priov_odd_mem_rclk (rf_cfg_cq2priov_odd_mem_rclk)
,.rf_cfg_cq2priov_odd_mem_rclk_rst_n (rf_cfg_cq2priov_odd_mem_rclk_rst_n)
,.rf_cfg_cq2priov_odd_mem_re    (rf_cfg_cq2priov_odd_mem_re)
,.rf_cfg_cq2priov_odd_mem_raddr (rf_cfg_cq2priov_odd_mem_raddr)
,.rf_cfg_cq2priov_odd_mem_waddr (rf_cfg_cq2priov_odd_mem_waddr)
,.rf_cfg_cq2priov_odd_mem_wclk (rf_cfg_cq2priov_odd_mem_wclk)
,.rf_cfg_cq2priov_odd_mem_wclk_rst_n (rf_cfg_cq2priov_odd_mem_wclk_rst_n)
,.rf_cfg_cq2priov_odd_mem_we    (rf_cfg_cq2priov_odd_mem_we)
,.rf_cfg_cq2priov_odd_mem_wdata (rf_cfg_cq2priov_odd_mem_wdata)
,.rf_cfg_cq2priov_odd_mem_rdata (rf_cfg_cq2priov_odd_mem_rdata)

,.rf_cfg_cq2priov_odd_mem_error (rf_cfg_cq2priov_odd_mem_error)

,.func_cfg_cq2qid_0_mem_re    (func_cfg_cq2qid_0_mem_re)
,.func_cfg_cq2qid_0_mem_addr  (func_cfg_cq2qid_0_mem_addr)
,.func_cfg_cq2qid_0_mem_we    (func_cfg_cq2qid_0_mem_we)
,.func_cfg_cq2qid_0_mem_wdata (func_cfg_cq2qid_0_mem_wdata)
,.func_cfg_cq2qid_0_mem_rdata (func_cfg_cq2qid_0_mem_rdata)

,.pf_cfg_cq2qid_0_mem_re      (pf_cfg_cq2qid_0_mem_re)
,.pf_cfg_cq2qid_0_mem_addr  (pf_cfg_cq2qid_0_mem_addr)
,.pf_cfg_cq2qid_0_mem_we    (pf_cfg_cq2qid_0_mem_we)
,.pf_cfg_cq2qid_0_mem_wdata (pf_cfg_cq2qid_0_mem_wdata)
,.pf_cfg_cq2qid_0_mem_rdata (pf_cfg_cq2qid_0_mem_rdata)

,.rf_cfg_cq2qid_0_mem_rclk (rf_cfg_cq2qid_0_mem_rclk)
,.rf_cfg_cq2qid_0_mem_rclk_rst_n (rf_cfg_cq2qid_0_mem_rclk_rst_n)
,.rf_cfg_cq2qid_0_mem_re    (rf_cfg_cq2qid_0_mem_re)
,.rf_cfg_cq2qid_0_mem_raddr (rf_cfg_cq2qid_0_mem_raddr)
,.rf_cfg_cq2qid_0_mem_waddr (rf_cfg_cq2qid_0_mem_waddr)
,.rf_cfg_cq2qid_0_mem_wclk (rf_cfg_cq2qid_0_mem_wclk)
,.rf_cfg_cq2qid_0_mem_wclk_rst_n (rf_cfg_cq2qid_0_mem_wclk_rst_n)
,.rf_cfg_cq2qid_0_mem_we    (rf_cfg_cq2qid_0_mem_we)
,.rf_cfg_cq2qid_0_mem_wdata (rf_cfg_cq2qid_0_mem_wdata)
,.rf_cfg_cq2qid_0_mem_rdata (rf_cfg_cq2qid_0_mem_rdata)

,.rf_cfg_cq2qid_0_mem_error (rf_cfg_cq2qid_0_mem_error)

,.func_cfg_cq2qid_0_odd_mem_re    (func_cfg_cq2qid_0_odd_mem_re)
,.func_cfg_cq2qid_0_odd_mem_addr  (func_cfg_cq2qid_0_odd_mem_addr)
,.func_cfg_cq2qid_0_odd_mem_we    (func_cfg_cq2qid_0_odd_mem_we)
,.func_cfg_cq2qid_0_odd_mem_wdata (func_cfg_cq2qid_0_odd_mem_wdata)
,.func_cfg_cq2qid_0_odd_mem_rdata (func_cfg_cq2qid_0_odd_mem_rdata)

,.pf_cfg_cq2qid_0_odd_mem_re      (pf_cfg_cq2qid_0_odd_mem_re)
,.pf_cfg_cq2qid_0_odd_mem_addr  (pf_cfg_cq2qid_0_odd_mem_addr)
,.pf_cfg_cq2qid_0_odd_mem_we    (pf_cfg_cq2qid_0_odd_mem_we)
,.pf_cfg_cq2qid_0_odd_mem_wdata (pf_cfg_cq2qid_0_odd_mem_wdata)
,.pf_cfg_cq2qid_0_odd_mem_rdata (pf_cfg_cq2qid_0_odd_mem_rdata)

,.rf_cfg_cq2qid_0_odd_mem_rclk (rf_cfg_cq2qid_0_odd_mem_rclk)
,.rf_cfg_cq2qid_0_odd_mem_rclk_rst_n (rf_cfg_cq2qid_0_odd_mem_rclk_rst_n)
,.rf_cfg_cq2qid_0_odd_mem_re    (rf_cfg_cq2qid_0_odd_mem_re)
,.rf_cfg_cq2qid_0_odd_mem_raddr (rf_cfg_cq2qid_0_odd_mem_raddr)
,.rf_cfg_cq2qid_0_odd_mem_waddr (rf_cfg_cq2qid_0_odd_mem_waddr)
,.rf_cfg_cq2qid_0_odd_mem_wclk (rf_cfg_cq2qid_0_odd_mem_wclk)
,.rf_cfg_cq2qid_0_odd_mem_wclk_rst_n (rf_cfg_cq2qid_0_odd_mem_wclk_rst_n)
,.rf_cfg_cq2qid_0_odd_mem_we    (rf_cfg_cq2qid_0_odd_mem_we)
,.rf_cfg_cq2qid_0_odd_mem_wdata (rf_cfg_cq2qid_0_odd_mem_wdata)
,.rf_cfg_cq2qid_0_odd_mem_rdata (rf_cfg_cq2qid_0_odd_mem_rdata)

,.rf_cfg_cq2qid_0_odd_mem_error (rf_cfg_cq2qid_0_odd_mem_error)

,.func_cfg_cq2qid_1_mem_re    (func_cfg_cq2qid_1_mem_re)
,.func_cfg_cq2qid_1_mem_addr  (func_cfg_cq2qid_1_mem_addr)
,.func_cfg_cq2qid_1_mem_we    (func_cfg_cq2qid_1_mem_we)
,.func_cfg_cq2qid_1_mem_wdata (func_cfg_cq2qid_1_mem_wdata)
,.func_cfg_cq2qid_1_mem_rdata (func_cfg_cq2qid_1_mem_rdata)

,.pf_cfg_cq2qid_1_mem_re      (pf_cfg_cq2qid_1_mem_re)
,.pf_cfg_cq2qid_1_mem_addr  (pf_cfg_cq2qid_1_mem_addr)
,.pf_cfg_cq2qid_1_mem_we    (pf_cfg_cq2qid_1_mem_we)
,.pf_cfg_cq2qid_1_mem_wdata (pf_cfg_cq2qid_1_mem_wdata)
,.pf_cfg_cq2qid_1_mem_rdata (pf_cfg_cq2qid_1_mem_rdata)

,.rf_cfg_cq2qid_1_mem_rclk (rf_cfg_cq2qid_1_mem_rclk)
,.rf_cfg_cq2qid_1_mem_rclk_rst_n (rf_cfg_cq2qid_1_mem_rclk_rst_n)
,.rf_cfg_cq2qid_1_mem_re    (rf_cfg_cq2qid_1_mem_re)
,.rf_cfg_cq2qid_1_mem_raddr (rf_cfg_cq2qid_1_mem_raddr)
,.rf_cfg_cq2qid_1_mem_waddr (rf_cfg_cq2qid_1_mem_waddr)
,.rf_cfg_cq2qid_1_mem_wclk (rf_cfg_cq2qid_1_mem_wclk)
,.rf_cfg_cq2qid_1_mem_wclk_rst_n (rf_cfg_cq2qid_1_mem_wclk_rst_n)
,.rf_cfg_cq2qid_1_mem_we    (rf_cfg_cq2qid_1_mem_we)
,.rf_cfg_cq2qid_1_mem_wdata (rf_cfg_cq2qid_1_mem_wdata)
,.rf_cfg_cq2qid_1_mem_rdata (rf_cfg_cq2qid_1_mem_rdata)

,.rf_cfg_cq2qid_1_mem_error (rf_cfg_cq2qid_1_mem_error)

,.func_cfg_cq2qid_1_odd_mem_re    (func_cfg_cq2qid_1_odd_mem_re)
,.func_cfg_cq2qid_1_odd_mem_addr  (func_cfg_cq2qid_1_odd_mem_addr)
,.func_cfg_cq2qid_1_odd_mem_we    (func_cfg_cq2qid_1_odd_mem_we)
,.func_cfg_cq2qid_1_odd_mem_wdata (func_cfg_cq2qid_1_odd_mem_wdata)
,.func_cfg_cq2qid_1_odd_mem_rdata (func_cfg_cq2qid_1_odd_mem_rdata)

,.pf_cfg_cq2qid_1_odd_mem_re      (pf_cfg_cq2qid_1_odd_mem_re)
,.pf_cfg_cq2qid_1_odd_mem_addr  (pf_cfg_cq2qid_1_odd_mem_addr)
,.pf_cfg_cq2qid_1_odd_mem_we    (pf_cfg_cq2qid_1_odd_mem_we)
,.pf_cfg_cq2qid_1_odd_mem_wdata (pf_cfg_cq2qid_1_odd_mem_wdata)
,.pf_cfg_cq2qid_1_odd_mem_rdata (pf_cfg_cq2qid_1_odd_mem_rdata)

,.rf_cfg_cq2qid_1_odd_mem_rclk (rf_cfg_cq2qid_1_odd_mem_rclk)
,.rf_cfg_cq2qid_1_odd_mem_rclk_rst_n (rf_cfg_cq2qid_1_odd_mem_rclk_rst_n)
,.rf_cfg_cq2qid_1_odd_mem_re    (rf_cfg_cq2qid_1_odd_mem_re)
,.rf_cfg_cq2qid_1_odd_mem_raddr (rf_cfg_cq2qid_1_odd_mem_raddr)
,.rf_cfg_cq2qid_1_odd_mem_waddr (rf_cfg_cq2qid_1_odd_mem_waddr)
,.rf_cfg_cq2qid_1_odd_mem_wclk (rf_cfg_cq2qid_1_odd_mem_wclk)
,.rf_cfg_cq2qid_1_odd_mem_wclk_rst_n (rf_cfg_cq2qid_1_odd_mem_wclk_rst_n)
,.rf_cfg_cq2qid_1_odd_mem_we    (rf_cfg_cq2qid_1_odd_mem_we)
,.rf_cfg_cq2qid_1_odd_mem_wdata (rf_cfg_cq2qid_1_odd_mem_wdata)
,.rf_cfg_cq2qid_1_odd_mem_rdata (rf_cfg_cq2qid_1_odd_mem_rdata)

,.rf_cfg_cq2qid_1_odd_mem_error (rf_cfg_cq2qid_1_odd_mem_error)

,.func_cfg_cq_ldb_inflight_limit_mem_re    (func_cfg_cq_ldb_inflight_limit_mem_re)
,.func_cfg_cq_ldb_inflight_limit_mem_addr  (func_cfg_cq_ldb_inflight_limit_mem_addr)
,.func_cfg_cq_ldb_inflight_limit_mem_we    (func_cfg_cq_ldb_inflight_limit_mem_we)
,.func_cfg_cq_ldb_inflight_limit_mem_wdata (func_cfg_cq_ldb_inflight_limit_mem_wdata)
,.func_cfg_cq_ldb_inflight_limit_mem_rdata (func_cfg_cq_ldb_inflight_limit_mem_rdata)

,.pf_cfg_cq_ldb_inflight_limit_mem_re      (pf_cfg_cq_ldb_inflight_limit_mem_re)
,.pf_cfg_cq_ldb_inflight_limit_mem_addr  (pf_cfg_cq_ldb_inflight_limit_mem_addr)
,.pf_cfg_cq_ldb_inflight_limit_mem_we    (pf_cfg_cq_ldb_inflight_limit_mem_we)
,.pf_cfg_cq_ldb_inflight_limit_mem_wdata (pf_cfg_cq_ldb_inflight_limit_mem_wdata)
,.pf_cfg_cq_ldb_inflight_limit_mem_rdata (pf_cfg_cq_ldb_inflight_limit_mem_rdata)

,.rf_cfg_cq_ldb_inflight_limit_mem_rclk (rf_cfg_cq_ldb_inflight_limit_mem_rclk)
,.rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n (rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n)
,.rf_cfg_cq_ldb_inflight_limit_mem_re    (rf_cfg_cq_ldb_inflight_limit_mem_re)
,.rf_cfg_cq_ldb_inflight_limit_mem_raddr (rf_cfg_cq_ldb_inflight_limit_mem_raddr)
,.rf_cfg_cq_ldb_inflight_limit_mem_waddr (rf_cfg_cq_ldb_inflight_limit_mem_waddr)
,.rf_cfg_cq_ldb_inflight_limit_mem_wclk (rf_cfg_cq_ldb_inflight_limit_mem_wclk)
,.rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n (rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n)
,.rf_cfg_cq_ldb_inflight_limit_mem_we    (rf_cfg_cq_ldb_inflight_limit_mem_we)
,.rf_cfg_cq_ldb_inflight_limit_mem_wdata (rf_cfg_cq_ldb_inflight_limit_mem_wdata)
,.rf_cfg_cq_ldb_inflight_limit_mem_rdata (rf_cfg_cq_ldb_inflight_limit_mem_rdata)

,.rf_cfg_cq_ldb_inflight_limit_mem_error (rf_cfg_cq_ldb_inflight_limit_mem_error)

,.func_cfg_cq_ldb_inflight_threshold_mem_re    (func_cfg_cq_ldb_inflight_threshold_mem_re)
,.func_cfg_cq_ldb_inflight_threshold_mem_addr  (func_cfg_cq_ldb_inflight_threshold_mem_addr)
,.func_cfg_cq_ldb_inflight_threshold_mem_we    (func_cfg_cq_ldb_inflight_threshold_mem_we)
,.func_cfg_cq_ldb_inflight_threshold_mem_wdata (func_cfg_cq_ldb_inflight_threshold_mem_wdata)
,.func_cfg_cq_ldb_inflight_threshold_mem_rdata (func_cfg_cq_ldb_inflight_threshold_mem_rdata)

,.pf_cfg_cq_ldb_inflight_threshold_mem_re      (pf_cfg_cq_ldb_inflight_threshold_mem_re)
,.pf_cfg_cq_ldb_inflight_threshold_mem_addr  (pf_cfg_cq_ldb_inflight_threshold_mem_addr)
,.pf_cfg_cq_ldb_inflight_threshold_mem_we    (pf_cfg_cq_ldb_inflight_threshold_mem_we)
,.pf_cfg_cq_ldb_inflight_threshold_mem_wdata (pf_cfg_cq_ldb_inflight_threshold_mem_wdata)
,.pf_cfg_cq_ldb_inflight_threshold_mem_rdata (pf_cfg_cq_ldb_inflight_threshold_mem_rdata)

,.rf_cfg_cq_ldb_inflight_threshold_mem_rclk (rf_cfg_cq_ldb_inflight_threshold_mem_rclk)
,.rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n (rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n)
,.rf_cfg_cq_ldb_inflight_threshold_mem_re    (rf_cfg_cq_ldb_inflight_threshold_mem_re)
,.rf_cfg_cq_ldb_inflight_threshold_mem_raddr (rf_cfg_cq_ldb_inflight_threshold_mem_raddr)
,.rf_cfg_cq_ldb_inflight_threshold_mem_waddr (rf_cfg_cq_ldb_inflight_threshold_mem_waddr)
,.rf_cfg_cq_ldb_inflight_threshold_mem_wclk (rf_cfg_cq_ldb_inflight_threshold_mem_wclk)
,.rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n (rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n)
,.rf_cfg_cq_ldb_inflight_threshold_mem_we    (rf_cfg_cq_ldb_inflight_threshold_mem_we)
,.rf_cfg_cq_ldb_inflight_threshold_mem_wdata (rf_cfg_cq_ldb_inflight_threshold_mem_wdata)
,.rf_cfg_cq_ldb_inflight_threshold_mem_rdata (rf_cfg_cq_ldb_inflight_threshold_mem_rdata)

,.rf_cfg_cq_ldb_inflight_threshold_mem_error (rf_cfg_cq_ldb_inflight_threshold_mem_error)

,.func_cfg_cq_ldb_token_depth_select_mem_re    (func_cfg_cq_ldb_token_depth_select_mem_re)
,.func_cfg_cq_ldb_token_depth_select_mem_addr  (func_cfg_cq_ldb_token_depth_select_mem_addr)
,.func_cfg_cq_ldb_token_depth_select_mem_we    (func_cfg_cq_ldb_token_depth_select_mem_we)
,.func_cfg_cq_ldb_token_depth_select_mem_wdata (func_cfg_cq_ldb_token_depth_select_mem_wdata)
,.func_cfg_cq_ldb_token_depth_select_mem_rdata (func_cfg_cq_ldb_token_depth_select_mem_rdata)

,.pf_cfg_cq_ldb_token_depth_select_mem_re      (pf_cfg_cq_ldb_token_depth_select_mem_re)
,.pf_cfg_cq_ldb_token_depth_select_mem_addr  (pf_cfg_cq_ldb_token_depth_select_mem_addr)
,.pf_cfg_cq_ldb_token_depth_select_mem_we    (pf_cfg_cq_ldb_token_depth_select_mem_we)
,.pf_cfg_cq_ldb_token_depth_select_mem_wdata (pf_cfg_cq_ldb_token_depth_select_mem_wdata)
,.pf_cfg_cq_ldb_token_depth_select_mem_rdata (pf_cfg_cq_ldb_token_depth_select_mem_rdata)

,.rf_cfg_cq_ldb_token_depth_select_mem_rclk (rf_cfg_cq_ldb_token_depth_select_mem_rclk)
,.rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n (rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n)
,.rf_cfg_cq_ldb_token_depth_select_mem_re    (rf_cfg_cq_ldb_token_depth_select_mem_re)
,.rf_cfg_cq_ldb_token_depth_select_mem_raddr (rf_cfg_cq_ldb_token_depth_select_mem_raddr)
,.rf_cfg_cq_ldb_token_depth_select_mem_waddr (rf_cfg_cq_ldb_token_depth_select_mem_waddr)
,.rf_cfg_cq_ldb_token_depth_select_mem_wclk (rf_cfg_cq_ldb_token_depth_select_mem_wclk)
,.rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n (rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n)
,.rf_cfg_cq_ldb_token_depth_select_mem_we    (rf_cfg_cq_ldb_token_depth_select_mem_we)
,.rf_cfg_cq_ldb_token_depth_select_mem_wdata (rf_cfg_cq_ldb_token_depth_select_mem_wdata)
,.rf_cfg_cq_ldb_token_depth_select_mem_rdata (rf_cfg_cq_ldb_token_depth_select_mem_rdata)

,.rf_cfg_cq_ldb_token_depth_select_mem_error (rf_cfg_cq_ldb_token_depth_select_mem_error)

,.func_cfg_cq_ldb_wu_limit_mem_re    (func_cfg_cq_ldb_wu_limit_mem_re)
,.func_cfg_cq_ldb_wu_limit_mem_raddr (func_cfg_cq_ldb_wu_limit_mem_raddr)
,.func_cfg_cq_ldb_wu_limit_mem_waddr (func_cfg_cq_ldb_wu_limit_mem_waddr)
,.func_cfg_cq_ldb_wu_limit_mem_we    (func_cfg_cq_ldb_wu_limit_mem_we)
,.func_cfg_cq_ldb_wu_limit_mem_wdata (func_cfg_cq_ldb_wu_limit_mem_wdata)
,.func_cfg_cq_ldb_wu_limit_mem_rdata (func_cfg_cq_ldb_wu_limit_mem_rdata)

,.pf_cfg_cq_ldb_wu_limit_mem_re      (pf_cfg_cq_ldb_wu_limit_mem_re)
,.pf_cfg_cq_ldb_wu_limit_mem_raddr (pf_cfg_cq_ldb_wu_limit_mem_raddr)
,.pf_cfg_cq_ldb_wu_limit_mem_waddr (pf_cfg_cq_ldb_wu_limit_mem_waddr)
,.pf_cfg_cq_ldb_wu_limit_mem_we    (pf_cfg_cq_ldb_wu_limit_mem_we)
,.pf_cfg_cq_ldb_wu_limit_mem_wdata (pf_cfg_cq_ldb_wu_limit_mem_wdata)
,.pf_cfg_cq_ldb_wu_limit_mem_rdata (pf_cfg_cq_ldb_wu_limit_mem_rdata)

,.rf_cfg_cq_ldb_wu_limit_mem_rclk (rf_cfg_cq_ldb_wu_limit_mem_rclk)
,.rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n (rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n)
,.rf_cfg_cq_ldb_wu_limit_mem_re    (rf_cfg_cq_ldb_wu_limit_mem_re)
,.rf_cfg_cq_ldb_wu_limit_mem_raddr (rf_cfg_cq_ldb_wu_limit_mem_raddr)
,.rf_cfg_cq_ldb_wu_limit_mem_waddr (rf_cfg_cq_ldb_wu_limit_mem_waddr)
,.rf_cfg_cq_ldb_wu_limit_mem_wclk (rf_cfg_cq_ldb_wu_limit_mem_wclk)
,.rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n (rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n)
,.rf_cfg_cq_ldb_wu_limit_mem_we    (rf_cfg_cq_ldb_wu_limit_mem_we)
,.rf_cfg_cq_ldb_wu_limit_mem_wdata (rf_cfg_cq_ldb_wu_limit_mem_wdata)
,.rf_cfg_cq_ldb_wu_limit_mem_rdata (rf_cfg_cq_ldb_wu_limit_mem_rdata)

,.rf_cfg_cq_ldb_wu_limit_mem_error (rf_cfg_cq_ldb_wu_limit_mem_error)

,.func_cfg_dir_qid_dpth_thrsh_mem_re    (func_cfg_dir_qid_dpth_thrsh_mem_re)
,.func_cfg_dir_qid_dpth_thrsh_mem_addr  (func_cfg_dir_qid_dpth_thrsh_mem_addr)
,.func_cfg_dir_qid_dpth_thrsh_mem_we    (func_cfg_dir_qid_dpth_thrsh_mem_we)
,.func_cfg_dir_qid_dpth_thrsh_mem_wdata (func_cfg_dir_qid_dpth_thrsh_mem_wdata)
,.func_cfg_dir_qid_dpth_thrsh_mem_rdata (func_cfg_dir_qid_dpth_thrsh_mem_rdata)

,.pf_cfg_dir_qid_dpth_thrsh_mem_re      (pf_cfg_dir_qid_dpth_thrsh_mem_re)
,.pf_cfg_dir_qid_dpth_thrsh_mem_addr  (pf_cfg_dir_qid_dpth_thrsh_mem_addr)
,.pf_cfg_dir_qid_dpth_thrsh_mem_we    (pf_cfg_dir_qid_dpth_thrsh_mem_we)
,.pf_cfg_dir_qid_dpth_thrsh_mem_wdata (pf_cfg_dir_qid_dpth_thrsh_mem_wdata)
,.pf_cfg_dir_qid_dpth_thrsh_mem_rdata (pf_cfg_dir_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_dir_qid_dpth_thrsh_mem_rclk (rf_cfg_dir_qid_dpth_thrsh_mem_rclk)
,.rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n (rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n)
,.rf_cfg_dir_qid_dpth_thrsh_mem_re    (rf_cfg_dir_qid_dpth_thrsh_mem_re)
,.rf_cfg_dir_qid_dpth_thrsh_mem_raddr (rf_cfg_dir_qid_dpth_thrsh_mem_raddr)
,.rf_cfg_dir_qid_dpth_thrsh_mem_waddr (rf_cfg_dir_qid_dpth_thrsh_mem_waddr)
,.rf_cfg_dir_qid_dpth_thrsh_mem_wclk (rf_cfg_dir_qid_dpth_thrsh_mem_wclk)
,.rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n (rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n)
,.rf_cfg_dir_qid_dpth_thrsh_mem_we    (rf_cfg_dir_qid_dpth_thrsh_mem_we)
,.rf_cfg_dir_qid_dpth_thrsh_mem_wdata (rf_cfg_dir_qid_dpth_thrsh_mem_wdata)
,.rf_cfg_dir_qid_dpth_thrsh_mem_rdata (rf_cfg_dir_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_dir_qid_dpth_thrsh_mem_error (rf_cfg_dir_qid_dpth_thrsh_mem_error)

,.func_cfg_nalb_qid_dpth_thrsh_mem_re    (func_cfg_nalb_qid_dpth_thrsh_mem_re)
,.func_cfg_nalb_qid_dpth_thrsh_mem_addr  (func_cfg_nalb_qid_dpth_thrsh_mem_addr)
,.func_cfg_nalb_qid_dpth_thrsh_mem_we    (func_cfg_nalb_qid_dpth_thrsh_mem_we)
,.func_cfg_nalb_qid_dpth_thrsh_mem_wdata (func_cfg_nalb_qid_dpth_thrsh_mem_wdata)
,.func_cfg_nalb_qid_dpth_thrsh_mem_rdata (func_cfg_nalb_qid_dpth_thrsh_mem_rdata)

,.pf_cfg_nalb_qid_dpth_thrsh_mem_re      (pf_cfg_nalb_qid_dpth_thrsh_mem_re)
,.pf_cfg_nalb_qid_dpth_thrsh_mem_addr  (pf_cfg_nalb_qid_dpth_thrsh_mem_addr)
,.pf_cfg_nalb_qid_dpth_thrsh_mem_we    (pf_cfg_nalb_qid_dpth_thrsh_mem_we)
,.pf_cfg_nalb_qid_dpth_thrsh_mem_wdata (pf_cfg_nalb_qid_dpth_thrsh_mem_wdata)
,.pf_cfg_nalb_qid_dpth_thrsh_mem_rdata (pf_cfg_nalb_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_nalb_qid_dpth_thrsh_mem_rclk (rf_cfg_nalb_qid_dpth_thrsh_mem_rclk)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n (rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_re    (rf_cfg_nalb_qid_dpth_thrsh_mem_re)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_raddr (rf_cfg_nalb_qid_dpth_thrsh_mem_raddr)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_waddr (rf_cfg_nalb_qid_dpth_thrsh_mem_waddr)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_wclk (rf_cfg_nalb_qid_dpth_thrsh_mem_wclk)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n (rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_we    (rf_cfg_nalb_qid_dpth_thrsh_mem_we)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_wdata (rf_cfg_nalb_qid_dpth_thrsh_mem_wdata)
,.rf_cfg_nalb_qid_dpth_thrsh_mem_rdata (rf_cfg_nalb_qid_dpth_thrsh_mem_rdata)

,.rf_cfg_nalb_qid_dpth_thrsh_mem_error (rf_cfg_nalb_qid_dpth_thrsh_mem_error)

,.func_cfg_qid_aqed_active_limit_mem_re    (func_cfg_qid_aqed_active_limit_mem_re)
,.func_cfg_qid_aqed_active_limit_mem_addr  (func_cfg_qid_aqed_active_limit_mem_addr)
,.func_cfg_qid_aqed_active_limit_mem_we    (func_cfg_qid_aqed_active_limit_mem_we)
,.func_cfg_qid_aqed_active_limit_mem_wdata (func_cfg_qid_aqed_active_limit_mem_wdata)
,.func_cfg_qid_aqed_active_limit_mem_rdata (func_cfg_qid_aqed_active_limit_mem_rdata)

,.pf_cfg_qid_aqed_active_limit_mem_re      (pf_cfg_qid_aqed_active_limit_mem_re)
,.pf_cfg_qid_aqed_active_limit_mem_addr  (pf_cfg_qid_aqed_active_limit_mem_addr)
,.pf_cfg_qid_aqed_active_limit_mem_we    (pf_cfg_qid_aqed_active_limit_mem_we)
,.pf_cfg_qid_aqed_active_limit_mem_wdata (pf_cfg_qid_aqed_active_limit_mem_wdata)
,.pf_cfg_qid_aqed_active_limit_mem_rdata (pf_cfg_qid_aqed_active_limit_mem_rdata)

,.rf_cfg_qid_aqed_active_limit_mem_rclk (rf_cfg_qid_aqed_active_limit_mem_rclk)
,.rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n (rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n)
,.rf_cfg_qid_aqed_active_limit_mem_re    (rf_cfg_qid_aqed_active_limit_mem_re)
,.rf_cfg_qid_aqed_active_limit_mem_raddr (rf_cfg_qid_aqed_active_limit_mem_raddr)
,.rf_cfg_qid_aqed_active_limit_mem_waddr (rf_cfg_qid_aqed_active_limit_mem_waddr)
,.rf_cfg_qid_aqed_active_limit_mem_wclk (rf_cfg_qid_aqed_active_limit_mem_wclk)
,.rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n (rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n)
,.rf_cfg_qid_aqed_active_limit_mem_we    (rf_cfg_qid_aqed_active_limit_mem_we)
,.rf_cfg_qid_aqed_active_limit_mem_wdata (rf_cfg_qid_aqed_active_limit_mem_wdata)
,.rf_cfg_qid_aqed_active_limit_mem_rdata (rf_cfg_qid_aqed_active_limit_mem_rdata)

,.rf_cfg_qid_aqed_active_limit_mem_error (rf_cfg_qid_aqed_active_limit_mem_error)

,.func_cfg_qid_ldb_inflight_limit_mem_re    (func_cfg_qid_ldb_inflight_limit_mem_re)
,.func_cfg_qid_ldb_inflight_limit_mem_addr  (func_cfg_qid_ldb_inflight_limit_mem_addr)
,.func_cfg_qid_ldb_inflight_limit_mem_we    (func_cfg_qid_ldb_inflight_limit_mem_we)
,.func_cfg_qid_ldb_inflight_limit_mem_wdata (func_cfg_qid_ldb_inflight_limit_mem_wdata)
,.func_cfg_qid_ldb_inflight_limit_mem_rdata (func_cfg_qid_ldb_inflight_limit_mem_rdata)

,.pf_cfg_qid_ldb_inflight_limit_mem_re      (pf_cfg_qid_ldb_inflight_limit_mem_re)
,.pf_cfg_qid_ldb_inflight_limit_mem_addr  (pf_cfg_qid_ldb_inflight_limit_mem_addr)
,.pf_cfg_qid_ldb_inflight_limit_mem_we    (pf_cfg_qid_ldb_inflight_limit_mem_we)
,.pf_cfg_qid_ldb_inflight_limit_mem_wdata (pf_cfg_qid_ldb_inflight_limit_mem_wdata)
,.pf_cfg_qid_ldb_inflight_limit_mem_rdata (pf_cfg_qid_ldb_inflight_limit_mem_rdata)

,.rf_cfg_qid_ldb_inflight_limit_mem_rclk (rf_cfg_qid_ldb_inflight_limit_mem_rclk)
,.rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n (rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n)
,.rf_cfg_qid_ldb_inflight_limit_mem_re    (rf_cfg_qid_ldb_inflight_limit_mem_re)
,.rf_cfg_qid_ldb_inflight_limit_mem_raddr (rf_cfg_qid_ldb_inflight_limit_mem_raddr)
,.rf_cfg_qid_ldb_inflight_limit_mem_waddr (rf_cfg_qid_ldb_inflight_limit_mem_waddr)
,.rf_cfg_qid_ldb_inflight_limit_mem_wclk (rf_cfg_qid_ldb_inflight_limit_mem_wclk)
,.rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n (rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n)
,.rf_cfg_qid_ldb_inflight_limit_mem_we    (rf_cfg_qid_ldb_inflight_limit_mem_we)
,.rf_cfg_qid_ldb_inflight_limit_mem_wdata (rf_cfg_qid_ldb_inflight_limit_mem_wdata)
,.rf_cfg_qid_ldb_inflight_limit_mem_rdata (rf_cfg_qid_ldb_inflight_limit_mem_rdata)

,.rf_cfg_qid_ldb_inflight_limit_mem_error (rf_cfg_qid_ldb_inflight_limit_mem_error)

,.func_cfg_qid_ldb_qid2cqidix2_mem_re    (func_cfg_qid_ldb_qid2cqidix2_mem_re)
,.func_cfg_qid_ldb_qid2cqidix2_mem_addr  (func_cfg_qid_ldb_qid2cqidix2_mem_addr)
,.func_cfg_qid_ldb_qid2cqidix2_mem_we    (func_cfg_qid_ldb_qid2cqidix2_mem_we)
,.func_cfg_qid_ldb_qid2cqidix2_mem_wdata (func_cfg_qid_ldb_qid2cqidix2_mem_wdata)
,.func_cfg_qid_ldb_qid2cqidix2_mem_rdata (func_cfg_qid_ldb_qid2cqidix2_mem_rdata)

,.pf_cfg_qid_ldb_qid2cqidix2_mem_re      (pf_cfg_qid_ldb_qid2cqidix2_mem_re)
,.pf_cfg_qid_ldb_qid2cqidix2_mem_addr  (pf_cfg_qid_ldb_qid2cqidix2_mem_addr)
,.pf_cfg_qid_ldb_qid2cqidix2_mem_we    (pf_cfg_qid_ldb_qid2cqidix2_mem_we)
,.pf_cfg_qid_ldb_qid2cqidix2_mem_wdata (pf_cfg_qid_ldb_qid2cqidix2_mem_wdata)
,.pf_cfg_qid_ldb_qid2cqidix2_mem_rdata (pf_cfg_qid_ldb_qid2cqidix2_mem_rdata)

,.rf_cfg_qid_ldb_qid2cqidix2_mem_rclk (rf_cfg_qid_ldb_qid2cqidix2_mem_rclk)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n (rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_re    (rf_cfg_qid_ldb_qid2cqidix2_mem_re)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_raddr (rf_cfg_qid_ldb_qid2cqidix2_mem_raddr)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_waddr (rf_cfg_qid_ldb_qid2cqidix2_mem_waddr)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_wclk (rf_cfg_qid_ldb_qid2cqidix2_mem_wclk)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n (rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_we    (rf_cfg_qid_ldb_qid2cqidix2_mem_we)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_wdata (rf_cfg_qid_ldb_qid2cqidix2_mem_wdata)
,.rf_cfg_qid_ldb_qid2cqidix2_mem_rdata (rf_cfg_qid_ldb_qid2cqidix2_mem_rdata)

,.rf_cfg_qid_ldb_qid2cqidix2_mem_error (rf_cfg_qid_ldb_qid2cqidix2_mem_error)

,.func_cfg_qid_ldb_qid2cqidix_mem_re    (func_cfg_qid_ldb_qid2cqidix_mem_re)
,.func_cfg_qid_ldb_qid2cqidix_mem_addr  (func_cfg_qid_ldb_qid2cqidix_mem_addr)
,.func_cfg_qid_ldb_qid2cqidix_mem_we    (func_cfg_qid_ldb_qid2cqidix_mem_we)
,.func_cfg_qid_ldb_qid2cqidix_mem_wdata (func_cfg_qid_ldb_qid2cqidix_mem_wdata)
,.func_cfg_qid_ldb_qid2cqidix_mem_rdata (func_cfg_qid_ldb_qid2cqidix_mem_rdata)

,.pf_cfg_qid_ldb_qid2cqidix_mem_re      (pf_cfg_qid_ldb_qid2cqidix_mem_re)
,.pf_cfg_qid_ldb_qid2cqidix_mem_addr  (pf_cfg_qid_ldb_qid2cqidix_mem_addr)
,.pf_cfg_qid_ldb_qid2cqidix_mem_we    (pf_cfg_qid_ldb_qid2cqidix_mem_we)
,.pf_cfg_qid_ldb_qid2cqidix_mem_wdata (pf_cfg_qid_ldb_qid2cqidix_mem_wdata)
,.pf_cfg_qid_ldb_qid2cqidix_mem_rdata (pf_cfg_qid_ldb_qid2cqidix_mem_rdata)

,.rf_cfg_qid_ldb_qid2cqidix_mem_rclk (rf_cfg_qid_ldb_qid2cqidix_mem_rclk)
,.rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n (rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n)
,.rf_cfg_qid_ldb_qid2cqidix_mem_re    (rf_cfg_qid_ldb_qid2cqidix_mem_re)
,.rf_cfg_qid_ldb_qid2cqidix_mem_raddr (rf_cfg_qid_ldb_qid2cqidix_mem_raddr)
,.rf_cfg_qid_ldb_qid2cqidix_mem_waddr (rf_cfg_qid_ldb_qid2cqidix_mem_waddr)
,.rf_cfg_qid_ldb_qid2cqidix_mem_wclk (rf_cfg_qid_ldb_qid2cqidix_mem_wclk)
,.rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n (rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n)
,.rf_cfg_qid_ldb_qid2cqidix_mem_we    (rf_cfg_qid_ldb_qid2cqidix_mem_we)
,.rf_cfg_qid_ldb_qid2cqidix_mem_wdata (rf_cfg_qid_ldb_qid2cqidix_mem_wdata)
,.rf_cfg_qid_ldb_qid2cqidix_mem_rdata (rf_cfg_qid_ldb_qid2cqidix_mem_rdata)

,.rf_cfg_qid_ldb_qid2cqidix_mem_error (rf_cfg_qid_ldb_qid2cqidix_mem_error)

,.func_chp_lsp_cmp_rx_sync_fifo_mem_re    (func_chp_lsp_cmp_rx_sync_fifo_mem_re)
,.func_chp_lsp_cmp_rx_sync_fifo_mem_raddr (func_chp_lsp_cmp_rx_sync_fifo_mem_raddr)
,.func_chp_lsp_cmp_rx_sync_fifo_mem_waddr (func_chp_lsp_cmp_rx_sync_fifo_mem_waddr)
,.func_chp_lsp_cmp_rx_sync_fifo_mem_we    (func_chp_lsp_cmp_rx_sync_fifo_mem_we)
,.func_chp_lsp_cmp_rx_sync_fifo_mem_wdata (func_chp_lsp_cmp_rx_sync_fifo_mem_wdata)
,.func_chp_lsp_cmp_rx_sync_fifo_mem_rdata (func_chp_lsp_cmp_rx_sync_fifo_mem_rdata)

,.pf_chp_lsp_cmp_rx_sync_fifo_mem_re      (pf_chp_lsp_cmp_rx_sync_fifo_mem_re)
,.pf_chp_lsp_cmp_rx_sync_fifo_mem_raddr (pf_chp_lsp_cmp_rx_sync_fifo_mem_raddr)
,.pf_chp_lsp_cmp_rx_sync_fifo_mem_waddr (pf_chp_lsp_cmp_rx_sync_fifo_mem_waddr)
,.pf_chp_lsp_cmp_rx_sync_fifo_mem_we    (pf_chp_lsp_cmp_rx_sync_fifo_mem_we)
,.pf_chp_lsp_cmp_rx_sync_fifo_mem_wdata (pf_chp_lsp_cmp_rx_sync_fifo_mem_wdata)
,.pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata (pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata)

,.rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk (rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n (rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_re    (rf_chp_lsp_cmp_rx_sync_fifo_mem_re)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr (rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr (rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk (rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n (rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_we    (rf_chp_lsp_cmp_rx_sync_fifo_mem_we)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata (rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata)
,.rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata (rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata)

,.rf_chp_lsp_cmp_rx_sync_fifo_mem_error (rf_chp_lsp_cmp_rx_sync_fifo_mem_error)

,.func_chp_lsp_token_rx_sync_fifo_mem_re    (func_chp_lsp_token_rx_sync_fifo_mem_re)
,.func_chp_lsp_token_rx_sync_fifo_mem_raddr (func_chp_lsp_token_rx_sync_fifo_mem_raddr)
,.func_chp_lsp_token_rx_sync_fifo_mem_waddr (func_chp_lsp_token_rx_sync_fifo_mem_waddr)
,.func_chp_lsp_token_rx_sync_fifo_mem_we    (func_chp_lsp_token_rx_sync_fifo_mem_we)
,.func_chp_lsp_token_rx_sync_fifo_mem_wdata (func_chp_lsp_token_rx_sync_fifo_mem_wdata)
,.func_chp_lsp_token_rx_sync_fifo_mem_rdata (func_chp_lsp_token_rx_sync_fifo_mem_rdata)

,.pf_chp_lsp_token_rx_sync_fifo_mem_re      (pf_chp_lsp_token_rx_sync_fifo_mem_re)
,.pf_chp_lsp_token_rx_sync_fifo_mem_raddr (pf_chp_lsp_token_rx_sync_fifo_mem_raddr)
,.pf_chp_lsp_token_rx_sync_fifo_mem_waddr (pf_chp_lsp_token_rx_sync_fifo_mem_waddr)
,.pf_chp_lsp_token_rx_sync_fifo_mem_we    (pf_chp_lsp_token_rx_sync_fifo_mem_we)
,.pf_chp_lsp_token_rx_sync_fifo_mem_wdata (pf_chp_lsp_token_rx_sync_fifo_mem_wdata)
,.pf_chp_lsp_token_rx_sync_fifo_mem_rdata (pf_chp_lsp_token_rx_sync_fifo_mem_rdata)

,.rf_chp_lsp_token_rx_sync_fifo_mem_rclk (rf_chp_lsp_token_rx_sync_fifo_mem_rclk)
,.rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n (rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n)
,.rf_chp_lsp_token_rx_sync_fifo_mem_re    (rf_chp_lsp_token_rx_sync_fifo_mem_re)
,.rf_chp_lsp_token_rx_sync_fifo_mem_raddr (rf_chp_lsp_token_rx_sync_fifo_mem_raddr)
,.rf_chp_lsp_token_rx_sync_fifo_mem_waddr (rf_chp_lsp_token_rx_sync_fifo_mem_waddr)
,.rf_chp_lsp_token_rx_sync_fifo_mem_wclk (rf_chp_lsp_token_rx_sync_fifo_mem_wclk)
,.rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n (rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n)
,.rf_chp_lsp_token_rx_sync_fifo_mem_we    (rf_chp_lsp_token_rx_sync_fifo_mem_we)
,.rf_chp_lsp_token_rx_sync_fifo_mem_wdata (rf_chp_lsp_token_rx_sync_fifo_mem_wdata)
,.rf_chp_lsp_token_rx_sync_fifo_mem_rdata (rf_chp_lsp_token_rx_sync_fifo_mem_rdata)

,.rf_chp_lsp_token_rx_sync_fifo_mem_error (rf_chp_lsp_token_rx_sync_fifo_mem_error)

,.func_cq_atm_pri_arbindex_mem_re    (func_cq_atm_pri_arbindex_mem_re)
,.func_cq_atm_pri_arbindex_mem_raddr (func_cq_atm_pri_arbindex_mem_raddr)
,.func_cq_atm_pri_arbindex_mem_waddr (func_cq_atm_pri_arbindex_mem_waddr)
,.func_cq_atm_pri_arbindex_mem_we    (func_cq_atm_pri_arbindex_mem_we)
,.func_cq_atm_pri_arbindex_mem_wdata (func_cq_atm_pri_arbindex_mem_wdata)
,.func_cq_atm_pri_arbindex_mem_rdata (func_cq_atm_pri_arbindex_mem_rdata)

,.pf_cq_atm_pri_arbindex_mem_re      (pf_cq_atm_pri_arbindex_mem_re)
,.pf_cq_atm_pri_arbindex_mem_raddr (pf_cq_atm_pri_arbindex_mem_raddr)
,.pf_cq_atm_pri_arbindex_mem_waddr (pf_cq_atm_pri_arbindex_mem_waddr)
,.pf_cq_atm_pri_arbindex_mem_we    (pf_cq_atm_pri_arbindex_mem_we)
,.pf_cq_atm_pri_arbindex_mem_wdata (pf_cq_atm_pri_arbindex_mem_wdata)
,.pf_cq_atm_pri_arbindex_mem_rdata (pf_cq_atm_pri_arbindex_mem_rdata)

,.rf_cq_atm_pri_arbindex_mem_rclk (rf_cq_atm_pri_arbindex_mem_rclk)
,.rf_cq_atm_pri_arbindex_mem_rclk_rst_n (rf_cq_atm_pri_arbindex_mem_rclk_rst_n)
,.rf_cq_atm_pri_arbindex_mem_re    (rf_cq_atm_pri_arbindex_mem_re)
,.rf_cq_atm_pri_arbindex_mem_raddr (rf_cq_atm_pri_arbindex_mem_raddr)
,.rf_cq_atm_pri_arbindex_mem_waddr (rf_cq_atm_pri_arbindex_mem_waddr)
,.rf_cq_atm_pri_arbindex_mem_wclk (rf_cq_atm_pri_arbindex_mem_wclk)
,.rf_cq_atm_pri_arbindex_mem_wclk_rst_n (rf_cq_atm_pri_arbindex_mem_wclk_rst_n)
,.rf_cq_atm_pri_arbindex_mem_we    (rf_cq_atm_pri_arbindex_mem_we)
,.rf_cq_atm_pri_arbindex_mem_wdata (rf_cq_atm_pri_arbindex_mem_wdata)
,.rf_cq_atm_pri_arbindex_mem_rdata (rf_cq_atm_pri_arbindex_mem_rdata)

,.rf_cq_atm_pri_arbindex_mem_error (rf_cq_atm_pri_arbindex_mem_error)

,.func_cq_dir_tot_sch_cnt_mem_re    (func_cq_dir_tot_sch_cnt_mem_re)
,.func_cq_dir_tot_sch_cnt_mem_raddr (func_cq_dir_tot_sch_cnt_mem_raddr)
,.func_cq_dir_tot_sch_cnt_mem_waddr (func_cq_dir_tot_sch_cnt_mem_waddr)
,.func_cq_dir_tot_sch_cnt_mem_we    (func_cq_dir_tot_sch_cnt_mem_we)
,.func_cq_dir_tot_sch_cnt_mem_wdata (func_cq_dir_tot_sch_cnt_mem_wdata)
,.func_cq_dir_tot_sch_cnt_mem_rdata (func_cq_dir_tot_sch_cnt_mem_rdata)

,.pf_cq_dir_tot_sch_cnt_mem_re      (pf_cq_dir_tot_sch_cnt_mem_re)
,.pf_cq_dir_tot_sch_cnt_mem_raddr (pf_cq_dir_tot_sch_cnt_mem_raddr)
,.pf_cq_dir_tot_sch_cnt_mem_waddr (pf_cq_dir_tot_sch_cnt_mem_waddr)
,.pf_cq_dir_tot_sch_cnt_mem_we    (pf_cq_dir_tot_sch_cnt_mem_we)
,.pf_cq_dir_tot_sch_cnt_mem_wdata (pf_cq_dir_tot_sch_cnt_mem_wdata)
,.pf_cq_dir_tot_sch_cnt_mem_rdata (pf_cq_dir_tot_sch_cnt_mem_rdata)

,.rf_cq_dir_tot_sch_cnt_mem_rclk (rf_cq_dir_tot_sch_cnt_mem_rclk)
,.rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n (rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n)
,.rf_cq_dir_tot_sch_cnt_mem_re    (rf_cq_dir_tot_sch_cnt_mem_re)
,.rf_cq_dir_tot_sch_cnt_mem_raddr (rf_cq_dir_tot_sch_cnt_mem_raddr)
,.rf_cq_dir_tot_sch_cnt_mem_waddr (rf_cq_dir_tot_sch_cnt_mem_waddr)
,.rf_cq_dir_tot_sch_cnt_mem_wclk (rf_cq_dir_tot_sch_cnt_mem_wclk)
,.rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n (rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n)
,.rf_cq_dir_tot_sch_cnt_mem_we    (rf_cq_dir_tot_sch_cnt_mem_we)
,.rf_cq_dir_tot_sch_cnt_mem_wdata (rf_cq_dir_tot_sch_cnt_mem_wdata)
,.rf_cq_dir_tot_sch_cnt_mem_rdata (rf_cq_dir_tot_sch_cnt_mem_rdata)

,.rf_cq_dir_tot_sch_cnt_mem_error (rf_cq_dir_tot_sch_cnt_mem_error)

,.func_cq_ldb_inflight_count_mem_re    (func_cq_ldb_inflight_count_mem_re)
,.func_cq_ldb_inflight_count_mem_raddr (func_cq_ldb_inflight_count_mem_raddr)
,.func_cq_ldb_inflight_count_mem_waddr (func_cq_ldb_inflight_count_mem_waddr)
,.func_cq_ldb_inflight_count_mem_we    (func_cq_ldb_inflight_count_mem_we)
,.func_cq_ldb_inflight_count_mem_wdata (func_cq_ldb_inflight_count_mem_wdata)
,.func_cq_ldb_inflight_count_mem_rdata (func_cq_ldb_inflight_count_mem_rdata)

,.pf_cq_ldb_inflight_count_mem_re      (pf_cq_ldb_inflight_count_mem_re)
,.pf_cq_ldb_inflight_count_mem_raddr (pf_cq_ldb_inflight_count_mem_raddr)
,.pf_cq_ldb_inflight_count_mem_waddr (pf_cq_ldb_inflight_count_mem_waddr)
,.pf_cq_ldb_inflight_count_mem_we    (pf_cq_ldb_inflight_count_mem_we)
,.pf_cq_ldb_inflight_count_mem_wdata (pf_cq_ldb_inflight_count_mem_wdata)
,.pf_cq_ldb_inflight_count_mem_rdata (pf_cq_ldb_inflight_count_mem_rdata)

,.rf_cq_ldb_inflight_count_mem_rclk (rf_cq_ldb_inflight_count_mem_rclk)
,.rf_cq_ldb_inflight_count_mem_rclk_rst_n (rf_cq_ldb_inflight_count_mem_rclk_rst_n)
,.rf_cq_ldb_inflight_count_mem_re    (rf_cq_ldb_inflight_count_mem_re)
,.rf_cq_ldb_inflight_count_mem_raddr (rf_cq_ldb_inflight_count_mem_raddr)
,.rf_cq_ldb_inflight_count_mem_waddr (rf_cq_ldb_inflight_count_mem_waddr)
,.rf_cq_ldb_inflight_count_mem_wclk (rf_cq_ldb_inflight_count_mem_wclk)
,.rf_cq_ldb_inflight_count_mem_wclk_rst_n (rf_cq_ldb_inflight_count_mem_wclk_rst_n)
,.rf_cq_ldb_inflight_count_mem_we    (rf_cq_ldb_inflight_count_mem_we)
,.rf_cq_ldb_inflight_count_mem_wdata (rf_cq_ldb_inflight_count_mem_wdata)
,.rf_cq_ldb_inflight_count_mem_rdata (rf_cq_ldb_inflight_count_mem_rdata)

,.rf_cq_ldb_inflight_count_mem_error (rf_cq_ldb_inflight_count_mem_error)

,.func_cq_ldb_token_count_mem_re    (func_cq_ldb_token_count_mem_re)
,.func_cq_ldb_token_count_mem_raddr (func_cq_ldb_token_count_mem_raddr)
,.func_cq_ldb_token_count_mem_waddr (func_cq_ldb_token_count_mem_waddr)
,.func_cq_ldb_token_count_mem_we    (func_cq_ldb_token_count_mem_we)
,.func_cq_ldb_token_count_mem_wdata (func_cq_ldb_token_count_mem_wdata)
,.func_cq_ldb_token_count_mem_rdata (func_cq_ldb_token_count_mem_rdata)

,.pf_cq_ldb_token_count_mem_re      (pf_cq_ldb_token_count_mem_re)
,.pf_cq_ldb_token_count_mem_raddr (pf_cq_ldb_token_count_mem_raddr)
,.pf_cq_ldb_token_count_mem_waddr (pf_cq_ldb_token_count_mem_waddr)
,.pf_cq_ldb_token_count_mem_we    (pf_cq_ldb_token_count_mem_we)
,.pf_cq_ldb_token_count_mem_wdata (pf_cq_ldb_token_count_mem_wdata)
,.pf_cq_ldb_token_count_mem_rdata (pf_cq_ldb_token_count_mem_rdata)

,.rf_cq_ldb_token_count_mem_rclk (rf_cq_ldb_token_count_mem_rclk)
,.rf_cq_ldb_token_count_mem_rclk_rst_n (rf_cq_ldb_token_count_mem_rclk_rst_n)
,.rf_cq_ldb_token_count_mem_re    (rf_cq_ldb_token_count_mem_re)
,.rf_cq_ldb_token_count_mem_raddr (rf_cq_ldb_token_count_mem_raddr)
,.rf_cq_ldb_token_count_mem_waddr (rf_cq_ldb_token_count_mem_waddr)
,.rf_cq_ldb_token_count_mem_wclk (rf_cq_ldb_token_count_mem_wclk)
,.rf_cq_ldb_token_count_mem_wclk_rst_n (rf_cq_ldb_token_count_mem_wclk_rst_n)
,.rf_cq_ldb_token_count_mem_we    (rf_cq_ldb_token_count_mem_we)
,.rf_cq_ldb_token_count_mem_wdata (rf_cq_ldb_token_count_mem_wdata)
,.rf_cq_ldb_token_count_mem_rdata (rf_cq_ldb_token_count_mem_rdata)

,.rf_cq_ldb_token_count_mem_error (rf_cq_ldb_token_count_mem_error)

,.func_cq_ldb_tot_sch_cnt_mem_re    (func_cq_ldb_tot_sch_cnt_mem_re)
,.func_cq_ldb_tot_sch_cnt_mem_raddr (func_cq_ldb_tot_sch_cnt_mem_raddr)
,.func_cq_ldb_tot_sch_cnt_mem_waddr (func_cq_ldb_tot_sch_cnt_mem_waddr)
,.func_cq_ldb_tot_sch_cnt_mem_we    (func_cq_ldb_tot_sch_cnt_mem_we)
,.func_cq_ldb_tot_sch_cnt_mem_wdata (func_cq_ldb_tot_sch_cnt_mem_wdata)
,.func_cq_ldb_tot_sch_cnt_mem_rdata (func_cq_ldb_tot_sch_cnt_mem_rdata)

,.pf_cq_ldb_tot_sch_cnt_mem_re      (pf_cq_ldb_tot_sch_cnt_mem_re)
,.pf_cq_ldb_tot_sch_cnt_mem_raddr (pf_cq_ldb_tot_sch_cnt_mem_raddr)
,.pf_cq_ldb_tot_sch_cnt_mem_waddr (pf_cq_ldb_tot_sch_cnt_mem_waddr)
,.pf_cq_ldb_tot_sch_cnt_mem_we    (pf_cq_ldb_tot_sch_cnt_mem_we)
,.pf_cq_ldb_tot_sch_cnt_mem_wdata (pf_cq_ldb_tot_sch_cnt_mem_wdata)
,.pf_cq_ldb_tot_sch_cnt_mem_rdata (pf_cq_ldb_tot_sch_cnt_mem_rdata)

,.rf_cq_ldb_tot_sch_cnt_mem_rclk (rf_cq_ldb_tot_sch_cnt_mem_rclk)
,.rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n (rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n)
,.rf_cq_ldb_tot_sch_cnt_mem_re    (rf_cq_ldb_tot_sch_cnt_mem_re)
,.rf_cq_ldb_tot_sch_cnt_mem_raddr (rf_cq_ldb_tot_sch_cnt_mem_raddr)
,.rf_cq_ldb_tot_sch_cnt_mem_waddr (rf_cq_ldb_tot_sch_cnt_mem_waddr)
,.rf_cq_ldb_tot_sch_cnt_mem_wclk (rf_cq_ldb_tot_sch_cnt_mem_wclk)
,.rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n (rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n)
,.rf_cq_ldb_tot_sch_cnt_mem_we    (rf_cq_ldb_tot_sch_cnt_mem_we)
,.rf_cq_ldb_tot_sch_cnt_mem_wdata (rf_cq_ldb_tot_sch_cnt_mem_wdata)
,.rf_cq_ldb_tot_sch_cnt_mem_rdata (rf_cq_ldb_tot_sch_cnt_mem_rdata)

,.rf_cq_ldb_tot_sch_cnt_mem_error (rf_cq_ldb_tot_sch_cnt_mem_error)

,.func_cq_ldb_wu_count_mem_re    (func_cq_ldb_wu_count_mem_re)
,.func_cq_ldb_wu_count_mem_raddr (func_cq_ldb_wu_count_mem_raddr)
,.func_cq_ldb_wu_count_mem_waddr (func_cq_ldb_wu_count_mem_waddr)
,.func_cq_ldb_wu_count_mem_we    (func_cq_ldb_wu_count_mem_we)
,.func_cq_ldb_wu_count_mem_wdata (func_cq_ldb_wu_count_mem_wdata)
,.func_cq_ldb_wu_count_mem_rdata (func_cq_ldb_wu_count_mem_rdata)

,.pf_cq_ldb_wu_count_mem_re      (pf_cq_ldb_wu_count_mem_re)
,.pf_cq_ldb_wu_count_mem_raddr (pf_cq_ldb_wu_count_mem_raddr)
,.pf_cq_ldb_wu_count_mem_waddr (pf_cq_ldb_wu_count_mem_waddr)
,.pf_cq_ldb_wu_count_mem_we    (pf_cq_ldb_wu_count_mem_we)
,.pf_cq_ldb_wu_count_mem_wdata (pf_cq_ldb_wu_count_mem_wdata)
,.pf_cq_ldb_wu_count_mem_rdata (pf_cq_ldb_wu_count_mem_rdata)

,.rf_cq_ldb_wu_count_mem_rclk (rf_cq_ldb_wu_count_mem_rclk)
,.rf_cq_ldb_wu_count_mem_rclk_rst_n (rf_cq_ldb_wu_count_mem_rclk_rst_n)
,.rf_cq_ldb_wu_count_mem_re    (rf_cq_ldb_wu_count_mem_re)
,.rf_cq_ldb_wu_count_mem_raddr (rf_cq_ldb_wu_count_mem_raddr)
,.rf_cq_ldb_wu_count_mem_waddr (rf_cq_ldb_wu_count_mem_waddr)
,.rf_cq_ldb_wu_count_mem_wclk (rf_cq_ldb_wu_count_mem_wclk)
,.rf_cq_ldb_wu_count_mem_wclk_rst_n (rf_cq_ldb_wu_count_mem_wclk_rst_n)
,.rf_cq_ldb_wu_count_mem_we    (rf_cq_ldb_wu_count_mem_we)
,.rf_cq_ldb_wu_count_mem_wdata (rf_cq_ldb_wu_count_mem_wdata)
,.rf_cq_ldb_wu_count_mem_rdata (rf_cq_ldb_wu_count_mem_rdata)

,.rf_cq_ldb_wu_count_mem_error (rf_cq_ldb_wu_count_mem_error)

,.func_cq_nalb_pri_arbindex_mem_re    (func_cq_nalb_pri_arbindex_mem_re)
,.func_cq_nalb_pri_arbindex_mem_raddr (func_cq_nalb_pri_arbindex_mem_raddr)
,.func_cq_nalb_pri_arbindex_mem_waddr (func_cq_nalb_pri_arbindex_mem_waddr)
,.func_cq_nalb_pri_arbindex_mem_we    (func_cq_nalb_pri_arbindex_mem_we)
,.func_cq_nalb_pri_arbindex_mem_wdata (func_cq_nalb_pri_arbindex_mem_wdata)
,.func_cq_nalb_pri_arbindex_mem_rdata (func_cq_nalb_pri_arbindex_mem_rdata)

,.pf_cq_nalb_pri_arbindex_mem_re      (pf_cq_nalb_pri_arbindex_mem_re)
,.pf_cq_nalb_pri_arbindex_mem_raddr (pf_cq_nalb_pri_arbindex_mem_raddr)
,.pf_cq_nalb_pri_arbindex_mem_waddr (pf_cq_nalb_pri_arbindex_mem_waddr)
,.pf_cq_nalb_pri_arbindex_mem_we    (pf_cq_nalb_pri_arbindex_mem_we)
,.pf_cq_nalb_pri_arbindex_mem_wdata (pf_cq_nalb_pri_arbindex_mem_wdata)
,.pf_cq_nalb_pri_arbindex_mem_rdata (pf_cq_nalb_pri_arbindex_mem_rdata)

,.rf_cq_nalb_pri_arbindex_mem_rclk (rf_cq_nalb_pri_arbindex_mem_rclk)
,.rf_cq_nalb_pri_arbindex_mem_rclk_rst_n (rf_cq_nalb_pri_arbindex_mem_rclk_rst_n)
,.rf_cq_nalb_pri_arbindex_mem_re    (rf_cq_nalb_pri_arbindex_mem_re)
,.rf_cq_nalb_pri_arbindex_mem_raddr (rf_cq_nalb_pri_arbindex_mem_raddr)
,.rf_cq_nalb_pri_arbindex_mem_waddr (rf_cq_nalb_pri_arbindex_mem_waddr)
,.rf_cq_nalb_pri_arbindex_mem_wclk (rf_cq_nalb_pri_arbindex_mem_wclk)
,.rf_cq_nalb_pri_arbindex_mem_wclk_rst_n (rf_cq_nalb_pri_arbindex_mem_wclk_rst_n)
,.rf_cq_nalb_pri_arbindex_mem_we    (rf_cq_nalb_pri_arbindex_mem_we)
,.rf_cq_nalb_pri_arbindex_mem_wdata (rf_cq_nalb_pri_arbindex_mem_wdata)
,.rf_cq_nalb_pri_arbindex_mem_rdata (rf_cq_nalb_pri_arbindex_mem_rdata)

,.rf_cq_nalb_pri_arbindex_mem_error (rf_cq_nalb_pri_arbindex_mem_error)

,.func_dir_enq_cnt_mem_re    (func_dir_enq_cnt_mem_re)
,.func_dir_enq_cnt_mem_raddr (func_dir_enq_cnt_mem_raddr)
,.func_dir_enq_cnt_mem_waddr (func_dir_enq_cnt_mem_waddr)
,.func_dir_enq_cnt_mem_we    (func_dir_enq_cnt_mem_we)
,.func_dir_enq_cnt_mem_wdata (func_dir_enq_cnt_mem_wdata)
,.func_dir_enq_cnt_mem_rdata (func_dir_enq_cnt_mem_rdata)

,.pf_dir_enq_cnt_mem_re      (pf_dir_enq_cnt_mem_re)
,.pf_dir_enq_cnt_mem_raddr (pf_dir_enq_cnt_mem_raddr)
,.pf_dir_enq_cnt_mem_waddr (pf_dir_enq_cnt_mem_waddr)
,.pf_dir_enq_cnt_mem_we    (pf_dir_enq_cnt_mem_we)
,.pf_dir_enq_cnt_mem_wdata (pf_dir_enq_cnt_mem_wdata)
,.pf_dir_enq_cnt_mem_rdata (pf_dir_enq_cnt_mem_rdata)

,.rf_dir_enq_cnt_mem_rclk (rf_dir_enq_cnt_mem_rclk)
,.rf_dir_enq_cnt_mem_rclk_rst_n (rf_dir_enq_cnt_mem_rclk_rst_n)
,.rf_dir_enq_cnt_mem_re    (rf_dir_enq_cnt_mem_re)
,.rf_dir_enq_cnt_mem_raddr (rf_dir_enq_cnt_mem_raddr)
,.rf_dir_enq_cnt_mem_waddr (rf_dir_enq_cnt_mem_waddr)
,.rf_dir_enq_cnt_mem_wclk (rf_dir_enq_cnt_mem_wclk)
,.rf_dir_enq_cnt_mem_wclk_rst_n (rf_dir_enq_cnt_mem_wclk_rst_n)
,.rf_dir_enq_cnt_mem_we    (rf_dir_enq_cnt_mem_we)
,.rf_dir_enq_cnt_mem_wdata (rf_dir_enq_cnt_mem_wdata)
,.rf_dir_enq_cnt_mem_rdata (rf_dir_enq_cnt_mem_rdata)

,.rf_dir_enq_cnt_mem_error (rf_dir_enq_cnt_mem_error)

,.func_dir_tok_cnt_mem_re    (func_dir_tok_cnt_mem_re)
,.func_dir_tok_cnt_mem_raddr (func_dir_tok_cnt_mem_raddr)
,.func_dir_tok_cnt_mem_waddr (func_dir_tok_cnt_mem_waddr)
,.func_dir_tok_cnt_mem_we    (func_dir_tok_cnt_mem_we)
,.func_dir_tok_cnt_mem_wdata (func_dir_tok_cnt_mem_wdata)
,.func_dir_tok_cnt_mem_rdata (func_dir_tok_cnt_mem_rdata)

,.pf_dir_tok_cnt_mem_re      (pf_dir_tok_cnt_mem_re)
,.pf_dir_tok_cnt_mem_raddr (pf_dir_tok_cnt_mem_raddr)
,.pf_dir_tok_cnt_mem_waddr (pf_dir_tok_cnt_mem_waddr)
,.pf_dir_tok_cnt_mem_we    (pf_dir_tok_cnt_mem_we)
,.pf_dir_tok_cnt_mem_wdata (pf_dir_tok_cnt_mem_wdata)
,.pf_dir_tok_cnt_mem_rdata (pf_dir_tok_cnt_mem_rdata)

,.rf_dir_tok_cnt_mem_rclk (rf_dir_tok_cnt_mem_rclk)
,.rf_dir_tok_cnt_mem_rclk_rst_n (rf_dir_tok_cnt_mem_rclk_rst_n)
,.rf_dir_tok_cnt_mem_re    (rf_dir_tok_cnt_mem_re)
,.rf_dir_tok_cnt_mem_raddr (rf_dir_tok_cnt_mem_raddr)
,.rf_dir_tok_cnt_mem_waddr (rf_dir_tok_cnt_mem_waddr)
,.rf_dir_tok_cnt_mem_wclk (rf_dir_tok_cnt_mem_wclk)
,.rf_dir_tok_cnt_mem_wclk_rst_n (rf_dir_tok_cnt_mem_wclk_rst_n)
,.rf_dir_tok_cnt_mem_we    (rf_dir_tok_cnt_mem_we)
,.rf_dir_tok_cnt_mem_wdata (rf_dir_tok_cnt_mem_wdata)
,.rf_dir_tok_cnt_mem_rdata (rf_dir_tok_cnt_mem_rdata)

,.rf_dir_tok_cnt_mem_error (rf_dir_tok_cnt_mem_error)

,.func_dir_tok_lim_mem_re    (func_dir_tok_lim_mem_re)
,.func_dir_tok_lim_mem_addr  (func_dir_tok_lim_mem_addr)
,.func_dir_tok_lim_mem_we    (func_dir_tok_lim_mem_we)
,.func_dir_tok_lim_mem_wdata (func_dir_tok_lim_mem_wdata)
,.func_dir_tok_lim_mem_rdata (func_dir_tok_lim_mem_rdata)

,.pf_dir_tok_lim_mem_re      (pf_dir_tok_lim_mem_re)
,.pf_dir_tok_lim_mem_addr  (pf_dir_tok_lim_mem_addr)
,.pf_dir_tok_lim_mem_we    (pf_dir_tok_lim_mem_we)
,.pf_dir_tok_lim_mem_wdata (pf_dir_tok_lim_mem_wdata)
,.pf_dir_tok_lim_mem_rdata (pf_dir_tok_lim_mem_rdata)

,.rf_dir_tok_lim_mem_rclk (rf_dir_tok_lim_mem_rclk)
,.rf_dir_tok_lim_mem_rclk_rst_n (rf_dir_tok_lim_mem_rclk_rst_n)
,.rf_dir_tok_lim_mem_re    (rf_dir_tok_lim_mem_re)
,.rf_dir_tok_lim_mem_raddr (rf_dir_tok_lim_mem_raddr)
,.rf_dir_tok_lim_mem_waddr (rf_dir_tok_lim_mem_waddr)
,.rf_dir_tok_lim_mem_wclk (rf_dir_tok_lim_mem_wclk)
,.rf_dir_tok_lim_mem_wclk_rst_n (rf_dir_tok_lim_mem_wclk_rst_n)
,.rf_dir_tok_lim_mem_we    (rf_dir_tok_lim_mem_we)
,.rf_dir_tok_lim_mem_wdata (rf_dir_tok_lim_mem_wdata)
,.rf_dir_tok_lim_mem_rdata (rf_dir_tok_lim_mem_rdata)

,.rf_dir_tok_lim_mem_error (rf_dir_tok_lim_mem_error)

,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_re    (func_dp_lsp_enq_dir_rx_sync_fifo_mem_re)
,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr (func_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr)
,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr (func_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr)
,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_we    (func_dp_lsp_enq_dir_rx_sync_fifo_mem_we)
,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata (func_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata)
,.func_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata (func_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata)

,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_re      (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_re)
,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr)
,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr)
,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_we    (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_we)
,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata)
,.pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata (pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata)

,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re    (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we    (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata)
,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata)

,.rf_dp_lsp_enq_dir_rx_sync_fifo_mem_error (rf_dp_lsp_enq_dir_rx_sync_fifo_mem_error)

,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_re    (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_we    (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.func_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata (func_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re      (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we    (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata (pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re    (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we    (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_error (rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_error)

,.func_enq_nalb_fifo_mem_re    (func_enq_nalb_fifo_mem_re)
,.func_enq_nalb_fifo_mem_raddr (func_enq_nalb_fifo_mem_raddr)
,.func_enq_nalb_fifo_mem_waddr (func_enq_nalb_fifo_mem_waddr)
,.func_enq_nalb_fifo_mem_we    (func_enq_nalb_fifo_mem_we)
,.func_enq_nalb_fifo_mem_wdata (func_enq_nalb_fifo_mem_wdata)
,.func_enq_nalb_fifo_mem_rdata (func_enq_nalb_fifo_mem_rdata)

,.pf_enq_nalb_fifo_mem_re      (pf_enq_nalb_fifo_mem_re)
,.pf_enq_nalb_fifo_mem_raddr (pf_enq_nalb_fifo_mem_raddr)
,.pf_enq_nalb_fifo_mem_waddr (pf_enq_nalb_fifo_mem_waddr)
,.pf_enq_nalb_fifo_mem_we    (pf_enq_nalb_fifo_mem_we)
,.pf_enq_nalb_fifo_mem_wdata (pf_enq_nalb_fifo_mem_wdata)
,.pf_enq_nalb_fifo_mem_rdata (pf_enq_nalb_fifo_mem_rdata)

,.rf_enq_nalb_fifo_mem_rclk (rf_enq_nalb_fifo_mem_rclk)
,.rf_enq_nalb_fifo_mem_rclk_rst_n (rf_enq_nalb_fifo_mem_rclk_rst_n)
,.rf_enq_nalb_fifo_mem_re    (rf_enq_nalb_fifo_mem_re)
,.rf_enq_nalb_fifo_mem_raddr (rf_enq_nalb_fifo_mem_raddr)
,.rf_enq_nalb_fifo_mem_waddr (rf_enq_nalb_fifo_mem_waddr)
,.rf_enq_nalb_fifo_mem_wclk (rf_enq_nalb_fifo_mem_wclk)
,.rf_enq_nalb_fifo_mem_wclk_rst_n (rf_enq_nalb_fifo_mem_wclk_rst_n)
,.rf_enq_nalb_fifo_mem_we    (rf_enq_nalb_fifo_mem_we)
,.rf_enq_nalb_fifo_mem_wdata (rf_enq_nalb_fifo_mem_wdata)
,.rf_enq_nalb_fifo_mem_rdata (rf_enq_nalb_fifo_mem_rdata)

,.rf_enq_nalb_fifo_mem_error (rf_enq_nalb_fifo_mem_error)

,.func_ldb_token_rtn_fifo_mem_re    (func_ldb_token_rtn_fifo_mem_re)
,.func_ldb_token_rtn_fifo_mem_raddr (func_ldb_token_rtn_fifo_mem_raddr)
,.func_ldb_token_rtn_fifo_mem_waddr (func_ldb_token_rtn_fifo_mem_waddr)
,.func_ldb_token_rtn_fifo_mem_we    (func_ldb_token_rtn_fifo_mem_we)
,.func_ldb_token_rtn_fifo_mem_wdata (func_ldb_token_rtn_fifo_mem_wdata)
,.func_ldb_token_rtn_fifo_mem_rdata (func_ldb_token_rtn_fifo_mem_rdata)

,.pf_ldb_token_rtn_fifo_mem_re      (pf_ldb_token_rtn_fifo_mem_re)
,.pf_ldb_token_rtn_fifo_mem_raddr (pf_ldb_token_rtn_fifo_mem_raddr)
,.pf_ldb_token_rtn_fifo_mem_waddr (pf_ldb_token_rtn_fifo_mem_waddr)
,.pf_ldb_token_rtn_fifo_mem_we    (pf_ldb_token_rtn_fifo_mem_we)
,.pf_ldb_token_rtn_fifo_mem_wdata (pf_ldb_token_rtn_fifo_mem_wdata)
,.pf_ldb_token_rtn_fifo_mem_rdata (pf_ldb_token_rtn_fifo_mem_rdata)

,.rf_ldb_token_rtn_fifo_mem_rclk (rf_ldb_token_rtn_fifo_mem_rclk)
,.rf_ldb_token_rtn_fifo_mem_rclk_rst_n (rf_ldb_token_rtn_fifo_mem_rclk_rst_n)
,.rf_ldb_token_rtn_fifo_mem_re    (rf_ldb_token_rtn_fifo_mem_re)
,.rf_ldb_token_rtn_fifo_mem_raddr (rf_ldb_token_rtn_fifo_mem_raddr)
,.rf_ldb_token_rtn_fifo_mem_waddr (rf_ldb_token_rtn_fifo_mem_waddr)
,.rf_ldb_token_rtn_fifo_mem_wclk (rf_ldb_token_rtn_fifo_mem_wclk)
,.rf_ldb_token_rtn_fifo_mem_wclk_rst_n (rf_ldb_token_rtn_fifo_mem_wclk_rst_n)
,.rf_ldb_token_rtn_fifo_mem_we    (rf_ldb_token_rtn_fifo_mem_we)
,.rf_ldb_token_rtn_fifo_mem_wdata (rf_ldb_token_rtn_fifo_mem_wdata)
,.rf_ldb_token_rtn_fifo_mem_rdata (rf_ldb_token_rtn_fifo_mem_rdata)

,.rf_ldb_token_rtn_fifo_mem_error (rf_ldb_token_rtn_fifo_mem_error)

,.func_nalb_cmp_fifo_mem_re    (func_nalb_cmp_fifo_mem_re)
,.func_nalb_cmp_fifo_mem_raddr (func_nalb_cmp_fifo_mem_raddr)
,.func_nalb_cmp_fifo_mem_waddr (func_nalb_cmp_fifo_mem_waddr)
,.func_nalb_cmp_fifo_mem_we    (func_nalb_cmp_fifo_mem_we)
,.func_nalb_cmp_fifo_mem_wdata (func_nalb_cmp_fifo_mem_wdata)
,.func_nalb_cmp_fifo_mem_rdata (func_nalb_cmp_fifo_mem_rdata)

,.pf_nalb_cmp_fifo_mem_re      (pf_nalb_cmp_fifo_mem_re)
,.pf_nalb_cmp_fifo_mem_raddr (pf_nalb_cmp_fifo_mem_raddr)
,.pf_nalb_cmp_fifo_mem_waddr (pf_nalb_cmp_fifo_mem_waddr)
,.pf_nalb_cmp_fifo_mem_we    (pf_nalb_cmp_fifo_mem_we)
,.pf_nalb_cmp_fifo_mem_wdata (pf_nalb_cmp_fifo_mem_wdata)
,.pf_nalb_cmp_fifo_mem_rdata (pf_nalb_cmp_fifo_mem_rdata)

,.rf_nalb_cmp_fifo_mem_rclk (rf_nalb_cmp_fifo_mem_rclk)
,.rf_nalb_cmp_fifo_mem_rclk_rst_n (rf_nalb_cmp_fifo_mem_rclk_rst_n)
,.rf_nalb_cmp_fifo_mem_re    (rf_nalb_cmp_fifo_mem_re)
,.rf_nalb_cmp_fifo_mem_raddr (rf_nalb_cmp_fifo_mem_raddr)
,.rf_nalb_cmp_fifo_mem_waddr (rf_nalb_cmp_fifo_mem_waddr)
,.rf_nalb_cmp_fifo_mem_wclk (rf_nalb_cmp_fifo_mem_wclk)
,.rf_nalb_cmp_fifo_mem_wclk_rst_n (rf_nalb_cmp_fifo_mem_wclk_rst_n)
,.rf_nalb_cmp_fifo_mem_we    (rf_nalb_cmp_fifo_mem_we)
,.rf_nalb_cmp_fifo_mem_wdata (rf_nalb_cmp_fifo_mem_wdata)
,.rf_nalb_cmp_fifo_mem_rdata (rf_nalb_cmp_fifo_mem_rdata)

,.rf_nalb_cmp_fifo_mem_error (rf_nalb_cmp_fifo_mem_error)

,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_re    (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_re)
,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr)
,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr)
,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_we    (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_we)
,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata)
,.func_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata (func_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata)

,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re      (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re)
,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr)
,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr)
,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we    (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we)
,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata)
,.pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata (pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata)

,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re    (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we    (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata)
,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata)

,.rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_error (rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_error)

,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re    (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we    (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata (func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re      (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we    (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata (pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re    (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we    (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata)
,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata)

,.rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_error (rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_error)

,.func_nalb_sel_nalb_fifo_mem_re    (func_nalb_sel_nalb_fifo_mem_re)
,.func_nalb_sel_nalb_fifo_mem_raddr (func_nalb_sel_nalb_fifo_mem_raddr)
,.func_nalb_sel_nalb_fifo_mem_waddr (func_nalb_sel_nalb_fifo_mem_waddr)
,.func_nalb_sel_nalb_fifo_mem_we    (func_nalb_sel_nalb_fifo_mem_we)
,.func_nalb_sel_nalb_fifo_mem_wdata (func_nalb_sel_nalb_fifo_mem_wdata)
,.func_nalb_sel_nalb_fifo_mem_rdata (func_nalb_sel_nalb_fifo_mem_rdata)

,.pf_nalb_sel_nalb_fifo_mem_re      (pf_nalb_sel_nalb_fifo_mem_re)
,.pf_nalb_sel_nalb_fifo_mem_raddr (pf_nalb_sel_nalb_fifo_mem_raddr)
,.pf_nalb_sel_nalb_fifo_mem_waddr (pf_nalb_sel_nalb_fifo_mem_waddr)
,.pf_nalb_sel_nalb_fifo_mem_we    (pf_nalb_sel_nalb_fifo_mem_we)
,.pf_nalb_sel_nalb_fifo_mem_wdata (pf_nalb_sel_nalb_fifo_mem_wdata)
,.pf_nalb_sel_nalb_fifo_mem_rdata (pf_nalb_sel_nalb_fifo_mem_rdata)

,.rf_nalb_sel_nalb_fifo_mem_rclk (rf_nalb_sel_nalb_fifo_mem_rclk)
,.rf_nalb_sel_nalb_fifo_mem_rclk_rst_n (rf_nalb_sel_nalb_fifo_mem_rclk_rst_n)
,.rf_nalb_sel_nalb_fifo_mem_re    (rf_nalb_sel_nalb_fifo_mem_re)
,.rf_nalb_sel_nalb_fifo_mem_raddr (rf_nalb_sel_nalb_fifo_mem_raddr)
,.rf_nalb_sel_nalb_fifo_mem_waddr (rf_nalb_sel_nalb_fifo_mem_waddr)
,.rf_nalb_sel_nalb_fifo_mem_wclk (rf_nalb_sel_nalb_fifo_mem_wclk)
,.rf_nalb_sel_nalb_fifo_mem_wclk_rst_n (rf_nalb_sel_nalb_fifo_mem_wclk_rst_n)
,.rf_nalb_sel_nalb_fifo_mem_we    (rf_nalb_sel_nalb_fifo_mem_we)
,.rf_nalb_sel_nalb_fifo_mem_wdata (rf_nalb_sel_nalb_fifo_mem_wdata)
,.rf_nalb_sel_nalb_fifo_mem_rdata (rf_nalb_sel_nalb_fifo_mem_rdata)

,.rf_nalb_sel_nalb_fifo_mem_error (rf_nalb_sel_nalb_fifo_mem_error)

,.func_qed_lsp_deq_fifo_mem_re    (func_qed_lsp_deq_fifo_mem_re)
,.func_qed_lsp_deq_fifo_mem_raddr (func_qed_lsp_deq_fifo_mem_raddr)
,.func_qed_lsp_deq_fifo_mem_waddr (func_qed_lsp_deq_fifo_mem_waddr)
,.func_qed_lsp_deq_fifo_mem_we    (func_qed_lsp_deq_fifo_mem_we)
,.func_qed_lsp_deq_fifo_mem_wdata (func_qed_lsp_deq_fifo_mem_wdata)
,.func_qed_lsp_deq_fifo_mem_rdata (func_qed_lsp_deq_fifo_mem_rdata)

,.pf_qed_lsp_deq_fifo_mem_re      (pf_qed_lsp_deq_fifo_mem_re)
,.pf_qed_lsp_deq_fifo_mem_raddr (pf_qed_lsp_deq_fifo_mem_raddr)
,.pf_qed_lsp_deq_fifo_mem_waddr (pf_qed_lsp_deq_fifo_mem_waddr)
,.pf_qed_lsp_deq_fifo_mem_we    (pf_qed_lsp_deq_fifo_mem_we)
,.pf_qed_lsp_deq_fifo_mem_wdata (pf_qed_lsp_deq_fifo_mem_wdata)
,.pf_qed_lsp_deq_fifo_mem_rdata (pf_qed_lsp_deq_fifo_mem_rdata)

,.rf_qed_lsp_deq_fifo_mem_rclk (rf_qed_lsp_deq_fifo_mem_rclk)
,.rf_qed_lsp_deq_fifo_mem_rclk_rst_n (rf_qed_lsp_deq_fifo_mem_rclk_rst_n)
,.rf_qed_lsp_deq_fifo_mem_re    (rf_qed_lsp_deq_fifo_mem_re)
,.rf_qed_lsp_deq_fifo_mem_raddr (rf_qed_lsp_deq_fifo_mem_raddr)
,.rf_qed_lsp_deq_fifo_mem_waddr (rf_qed_lsp_deq_fifo_mem_waddr)
,.rf_qed_lsp_deq_fifo_mem_wclk (rf_qed_lsp_deq_fifo_mem_wclk)
,.rf_qed_lsp_deq_fifo_mem_wclk_rst_n (rf_qed_lsp_deq_fifo_mem_wclk_rst_n)
,.rf_qed_lsp_deq_fifo_mem_we    (rf_qed_lsp_deq_fifo_mem_we)
,.rf_qed_lsp_deq_fifo_mem_wdata (rf_qed_lsp_deq_fifo_mem_wdata)
,.rf_qed_lsp_deq_fifo_mem_rdata (rf_qed_lsp_deq_fifo_mem_rdata)

,.rf_qed_lsp_deq_fifo_mem_error (rf_qed_lsp_deq_fifo_mem_error)

,.func_qid_aqed_active_count_mem_re    (func_qid_aqed_active_count_mem_re)
,.func_qid_aqed_active_count_mem_raddr (func_qid_aqed_active_count_mem_raddr)
,.func_qid_aqed_active_count_mem_waddr (func_qid_aqed_active_count_mem_waddr)
,.func_qid_aqed_active_count_mem_we    (func_qid_aqed_active_count_mem_we)
,.func_qid_aqed_active_count_mem_wdata (func_qid_aqed_active_count_mem_wdata)
,.func_qid_aqed_active_count_mem_rdata (func_qid_aqed_active_count_mem_rdata)

,.pf_qid_aqed_active_count_mem_re      (pf_qid_aqed_active_count_mem_re)
,.pf_qid_aqed_active_count_mem_raddr (pf_qid_aqed_active_count_mem_raddr)
,.pf_qid_aqed_active_count_mem_waddr (pf_qid_aqed_active_count_mem_waddr)
,.pf_qid_aqed_active_count_mem_we    (pf_qid_aqed_active_count_mem_we)
,.pf_qid_aqed_active_count_mem_wdata (pf_qid_aqed_active_count_mem_wdata)
,.pf_qid_aqed_active_count_mem_rdata (pf_qid_aqed_active_count_mem_rdata)

,.rf_qid_aqed_active_count_mem_rclk (rf_qid_aqed_active_count_mem_rclk)
,.rf_qid_aqed_active_count_mem_rclk_rst_n (rf_qid_aqed_active_count_mem_rclk_rst_n)
,.rf_qid_aqed_active_count_mem_re    (rf_qid_aqed_active_count_mem_re)
,.rf_qid_aqed_active_count_mem_raddr (rf_qid_aqed_active_count_mem_raddr)
,.rf_qid_aqed_active_count_mem_waddr (rf_qid_aqed_active_count_mem_waddr)
,.rf_qid_aqed_active_count_mem_wclk (rf_qid_aqed_active_count_mem_wclk)
,.rf_qid_aqed_active_count_mem_wclk_rst_n (rf_qid_aqed_active_count_mem_wclk_rst_n)
,.rf_qid_aqed_active_count_mem_we    (rf_qid_aqed_active_count_mem_we)
,.rf_qid_aqed_active_count_mem_wdata (rf_qid_aqed_active_count_mem_wdata)
,.rf_qid_aqed_active_count_mem_rdata (rf_qid_aqed_active_count_mem_rdata)

,.rf_qid_aqed_active_count_mem_error (rf_qid_aqed_active_count_mem_error)

,.func_qid_atm_active_mem_re    (func_qid_atm_active_mem_re)
,.func_qid_atm_active_mem_raddr (func_qid_atm_active_mem_raddr)
,.func_qid_atm_active_mem_waddr (func_qid_atm_active_mem_waddr)
,.func_qid_atm_active_mem_we    (func_qid_atm_active_mem_we)
,.func_qid_atm_active_mem_wdata (func_qid_atm_active_mem_wdata)
,.func_qid_atm_active_mem_rdata (func_qid_atm_active_mem_rdata)

,.pf_qid_atm_active_mem_re      (pf_qid_atm_active_mem_re)
,.pf_qid_atm_active_mem_raddr (pf_qid_atm_active_mem_raddr)
,.pf_qid_atm_active_mem_waddr (pf_qid_atm_active_mem_waddr)
,.pf_qid_atm_active_mem_we    (pf_qid_atm_active_mem_we)
,.pf_qid_atm_active_mem_wdata (pf_qid_atm_active_mem_wdata)
,.pf_qid_atm_active_mem_rdata (pf_qid_atm_active_mem_rdata)

,.rf_qid_atm_active_mem_rclk (rf_qid_atm_active_mem_rclk)
,.rf_qid_atm_active_mem_rclk_rst_n (rf_qid_atm_active_mem_rclk_rst_n)
,.rf_qid_atm_active_mem_re    (rf_qid_atm_active_mem_re)
,.rf_qid_atm_active_mem_raddr (rf_qid_atm_active_mem_raddr)
,.rf_qid_atm_active_mem_waddr (rf_qid_atm_active_mem_waddr)
,.rf_qid_atm_active_mem_wclk (rf_qid_atm_active_mem_wclk)
,.rf_qid_atm_active_mem_wclk_rst_n (rf_qid_atm_active_mem_wclk_rst_n)
,.rf_qid_atm_active_mem_we    (rf_qid_atm_active_mem_we)
,.rf_qid_atm_active_mem_wdata (rf_qid_atm_active_mem_wdata)
,.rf_qid_atm_active_mem_rdata (rf_qid_atm_active_mem_rdata)

,.rf_qid_atm_active_mem_error (rf_qid_atm_active_mem_error)

,.func_qid_atm_tot_enq_cnt_mem_re    (func_qid_atm_tot_enq_cnt_mem_re)
,.func_qid_atm_tot_enq_cnt_mem_raddr (func_qid_atm_tot_enq_cnt_mem_raddr)
,.func_qid_atm_tot_enq_cnt_mem_waddr (func_qid_atm_tot_enq_cnt_mem_waddr)
,.func_qid_atm_tot_enq_cnt_mem_we    (func_qid_atm_tot_enq_cnt_mem_we)
,.func_qid_atm_tot_enq_cnt_mem_wdata (func_qid_atm_tot_enq_cnt_mem_wdata)
,.func_qid_atm_tot_enq_cnt_mem_rdata (func_qid_atm_tot_enq_cnt_mem_rdata)

,.pf_qid_atm_tot_enq_cnt_mem_re      (pf_qid_atm_tot_enq_cnt_mem_re)
,.pf_qid_atm_tot_enq_cnt_mem_raddr (pf_qid_atm_tot_enq_cnt_mem_raddr)
,.pf_qid_atm_tot_enq_cnt_mem_waddr (pf_qid_atm_tot_enq_cnt_mem_waddr)
,.pf_qid_atm_tot_enq_cnt_mem_we    (pf_qid_atm_tot_enq_cnt_mem_we)
,.pf_qid_atm_tot_enq_cnt_mem_wdata (pf_qid_atm_tot_enq_cnt_mem_wdata)
,.pf_qid_atm_tot_enq_cnt_mem_rdata (pf_qid_atm_tot_enq_cnt_mem_rdata)

,.rf_qid_atm_tot_enq_cnt_mem_rclk (rf_qid_atm_tot_enq_cnt_mem_rclk)
,.rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n (rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n)
,.rf_qid_atm_tot_enq_cnt_mem_re    (rf_qid_atm_tot_enq_cnt_mem_re)
,.rf_qid_atm_tot_enq_cnt_mem_raddr (rf_qid_atm_tot_enq_cnt_mem_raddr)
,.rf_qid_atm_tot_enq_cnt_mem_waddr (rf_qid_atm_tot_enq_cnt_mem_waddr)
,.rf_qid_atm_tot_enq_cnt_mem_wclk (rf_qid_atm_tot_enq_cnt_mem_wclk)
,.rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n (rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n)
,.rf_qid_atm_tot_enq_cnt_mem_we    (rf_qid_atm_tot_enq_cnt_mem_we)
,.rf_qid_atm_tot_enq_cnt_mem_wdata (rf_qid_atm_tot_enq_cnt_mem_wdata)
,.rf_qid_atm_tot_enq_cnt_mem_rdata (rf_qid_atm_tot_enq_cnt_mem_rdata)

,.rf_qid_atm_tot_enq_cnt_mem_error (rf_qid_atm_tot_enq_cnt_mem_error)

,.func_qid_atq_enqueue_count_mem_re    (func_qid_atq_enqueue_count_mem_re)
,.func_qid_atq_enqueue_count_mem_raddr (func_qid_atq_enqueue_count_mem_raddr)
,.func_qid_atq_enqueue_count_mem_waddr (func_qid_atq_enqueue_count_mem_waddr)
,.func_qid_atq_enqueue_count_mem_we    (func_qid_atq_enqueue_count_mem_we)
,.func_qid_atq_enqueue_count_mem_wdata (func_qid_atq_enqueue_count_mem_wdata)
,.func_qid_atq_enqueue_count_mem_rdata (func_qid_atq_enqueue_count_mem_rdata)

,.pf_qid_atq_enqueue_count_mem_re      (pf_qid_atq_enqueue_count_mem_re)
,.pf_qid_atq_enqueue_count_mem_raddr (pf_qid_atq_enqueue_count_mem_raddr)
,.pf_qid_atq_enqueue_count_mem_waddr (pf_qid_atq_enqueue_count_mem_waddr)
,.pf_qid_atq_enqueue_count_mem_we    (pf_qid_atq_enqueue_count_mem_we)
,.pf_qid_atq_enqueue_count_mem_wdata (pf_qid_atq_enqueue_count_mem_wdata)
,.pf_qid_atq_enqueue_count_mem_rdata (pf_qid_atq_enqueue_count_mem_rdata)

,.rf_qid_atq_enqueue_count_mem_rclk (rf_qid_atq_enqueue_count_mem_rclk)
,.rf_qid_atq_enqueue_count_mem_rclk_rst_n (rf_qid_atq_enqueue_count_mem_rclk_rst_n)
,.rf_qid_atq_enqueue_count_mem_re    (rf_qid_atq_enqueue_count_mem_re)
,.rf_qid_atq_enqueue_count_mem_raddr (rf_qid_atq_enqueue_count_mem_raddr)
,.rf_qid_atq_enqueue_count_mem_waddr (rf_qid_atq_enqueue_count_mem_waddr)
,.rf_qid_atq_enqueue_count_mem_wclk (rf_qid_atq_enqueue_count_mem_wclk)
,.rf_qid_atq_enqueue_count_mem_wclk_rst_n (rf_qid_atq_enqueue_count_mem_wclk_rst_n)
,.rf_qid_atq_enqueue_count_mem_we    (rf_qid_atq_enqueue_count_mem_we)
,.rf_qid_atq_enqueue_count_mem_wdata (rf_qid_atq_enqueue_count_mem_wdata)
,.rf_qid_atq_enqueue_count_mem_rdata (rf_qid_atq_enqueue_count_mem_rdata)

,.rf_qid_atq_enqueue_count_mem_error (rf_qid_atq_enqueue_count_mem_error)

,.func_qid_dir_max_depth_mem_re    (func_qid_dir_max_depth_mem_re)
,.func_qid_dir_max_depth_mem_raddr (func_qid_dir_max_depth_mem_raddr)
,.func_qid_dir_max_depth_mem_waddr (func_qid_dir_max_depth_mem_waddr)
,.func_qid_dir_max_depth_mem_we    (func_qid_dir_max_depth_mem_we)
,.func_qid_dir_max_depth_mem_wdata (func_qid_dir_max_depth_mem_wdata)
,.func_qid_dir_max_depth_mem_rdata (func_qid_dir_max_depth_mem_rdata)

,.pf_qid_dir_max_depth_mem_re      (pf_qid_dir_max_depth_mem_re)
,.pf_qid_dir_max_depth_mem_raddr (pf_qid_dir_max_depth_mem_raddr)
,.pf_qid_dir_max_depth_mem_waddr (pf_qid_dir_max_depth_mem_waddr)
,.pf_qid_dir_max_depth_mem_we    (pf_qid_dir_max_depth_mem_we)
,.pf_qid_dir_max_depth_mem_wdata (pf_qid_dir_max_depth_mem_wdata)
,.pf_qid_dir_max_depth_mem_rdata (pf_qid_dir_max_depth_mem_rdata)

,.rf_qid_dir_max_depth_mem_rclk (rf_qid_dir_max_depth_mem_rclk)
,.rf_qid_dir_max_depth_mem_rclk_rst_n (rf_qid_dir_max_depth_mem_rclk_rst_n)
,.rf_qid_dir_max_depth_mem_re    (rf_qid_dir_max_depth_mem_re)
,.rf_qid_dir_max_depth_mem_raddr (rf_qid_dir_max_depth_mem_raddr)
,.rf_qid_dir_max_depth_mem_waddr (rf_qid_dir_max_depth_mem_waddr)
,.rf_qid_dir_max_depth_mem_wclk (rf_qid_dir_max_depth_mem_wclk)
,.rf_qid_dir_max_depth_mem_wclk_rst_n (rf_qid_dir_max_depth_mem_wclk_rst_n)
,.rf_qid_dir_max_depth_mem_we    (rf_qid_dir_max_depth_mem_we)
,.rf_qid_dir_max_depth_mem_wdata (rf_qid_dir_max_depth_mem_wdata)
,.rf_qid_dir_max_depth_mem_rdata (rf_qid_dir_max_depth_mem_rdata)

,.rf_qid_dir_max_depth_mem_error (rf_qid_dir_max_depth_mem_error)

,.func_qid_dir_replay_count_mem_re    (func_qid_dir_replay_count_mem_re)
,.func_qid_dir_replay_count_mem_raddr (func_qid_dir_replay_count_mem_raddr)
,.func_qid_dir_replay_count_mem_waddr (func_qid_dir_replay_count_mem_waddr)
,.func_qid_dir_replay_count_mem_we    (func_qid_dir_replay_count_mem_we)
,.func_qid_dir_replay_count_mem_wdata (func_qid_dir_replay_count_mem_wdata)
,.func_qid_dir_replay_count_mem_rdata (func_qid_dir_replay_count_mem_rdata)

,.pf_qid_dir_replay_count_mem_re      (pf_qid_dir_replay_count_mem_re)
,.pf_qid_dir_replay_count_mem_raddr (pf_qid_dir_replay_count_mem_raddr)
,.pf_qid_dir_replay_count_mem_waddr (pf_qid_dir_replay_count_mem_waddr)
,.pf_qid_dir_replay_count_mem_we    (pf_qid_dir_replay_count_mem_we)
,.pf_qid_dir_replay_count_mem_wdata (pf_qid_dir_replay_count_mem_wdata)
,.pf_qid_dir_replay_count_mem_rdata (pf_qid_dir_replay_count_mem_rdata)

,.rf_qid_dir_replay_count_mem_rclk (rf_qid_dir_replay_count_mem_rclk)
,.rf_qid_dir_replay_count_mem_rclk_rst_n (rf_qid_dir_replay_count_mem_rclk_rst_n)
,.rf_qid_dir_replay_count_mem_re    (rf_qid_dir_replay_count_mem_re)
,.rf_qid_dir_replay_count_mem_raddr (rf_qid_dir_replay_count_mem_raddr)
,.rf_qid_dir_replay_count_mem_waddr (rf_qid_dir_replay_count_mem_waddr)
,.rf_qid_dir_replay_count_mem_wclk (rf_qid_dir_replay_count_mem_wclk)
,.rf_qid_dir_replay_count_mem_wclk_rst_n (rf_qid_dir_replay_count_mem_wclk_rst_n)
,.rf_qid_dir_replay_count_mem_we    (rf_qid_dir_replay_count_mem_we)
,.rf_qid_dir_replay_count_mem_wdata (rf_qid_dir_replay_count_mem_wdata)
,.rf_qid_dir_replay_count_mem_rdata (rf_qid_dir_replay_count_mem_rdata)

,.rf_qid_dir_replay_count_mem_error (rf_qid_dir_replay_count_mem_error)

,.func_qid_dir_tot_enq_cnt_mem_re    (func_qid_dir_tot_enq_cnt_mem_re)
,.func_qid_dir_tot_enq_cnt_mem_raddr (func_qid_dir_tot_enq_cnt_mem_raddr)
,.func_qid_dir_tot_enq_cnt_mem_waddr (func_qid_dir_tot_enq_cnt_mem_waddr)
,.func_qid_dir_tot_enq_cnt_mem_we    (func_qid_dir_tot_enq_cnt_mem_we)
,.func_qid_dir_tot_enq_cnt_mem_wdata (func_qid_dir_tot_enq_cnt_mem_wdata)
,.func_qid_dir_tot_enq_cnt_mem_rdata (func_qid_dir_tot_enq_cnt_mem_rdata)

,.pf_qid_dir_tot_enq_cnt_mem_re      (pf_qid_dir_tot_enq_cnt_mem_re)
,.pf_qid_dir_tot_enq_cnt_mem_raddr (pf_qid_dir_tot_enq_cnt_mem_raddr)
,.pf_qid_dir_tot_enq_cnt_mem_waddr (pf_qid_dir_tot_enq_cnt_mem_waddr)
,.pf_qid_dir_tot_enq_cnt_mem_we    (pf_qid_dir_tot_enq_cnt_mem_we)
,.pf_qid_dir_tot_enq_cnt_mem_wdata (pf_qid_dir_tot_enq_cnt_mem_wdata)
,.pf_qid_dir_tot_enq_cnt_mem_rdata (pf_qid_dir_tot_enq_cnt_mem_rdata)

,.rf_qid_dir_tot_enq_cnt_mem_rclk (rf_qid_dir_tot_enq_cnt_mem_rclk)
,.rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n (rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n)
,.rf_qid_dir_tot_enq_cnt_mem_re    (rf_qid_dir_tot_enq_cnt_mem_re)
,.rf_qid_dir_tot_enq_cnt_mem_raddr (rf_qid_dir_tot_enq_cnt_mem_raddr)
,.rf_qid_dir_tot_enq_cnt_mem_waddr (rf_qid_dir_tot_enq_cnt_mem_waddr)
,.rf_qid_dir_tot_enq_cnt_mem_wclk (rf_qid_dir_tot_enq_cnt_mem_wclk)
,.rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n (rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n)
,.rf_qid_dir_tot_enq_cnt_mem_we    (rf_qid_dir_tot_enq_cnt_mem_we)
,.rf_qid_dir_tot_enq_cnt_mem_wdata (rf_qid_dir_tot_enq_cnt_mem_wdata)
,.rf_qid_dir_tot_enq_cnt_mem_rdata (rf_qid_dir_tot_enq_cnt_mem_rdata)

,.rf_qid_dir_tot_enq_cnt_mem_error (rf_qid_dir_tot_enq_cnt_mem_error)

,.func_qid_ldb_enqueue_count_mem_re    (func_qid_ldb_enqueue_count_mem_re)
,.func_qid_ldb_enqueue_count_mem_raddr (func_qid_ldb_enqueue_count_mem_raddr)
,.func_qid_ldb_enqueue_count_mem_waddr (func_qid_ldb_enqueue_count_mem_waddr)
,.func_qid_ldb_enqueue_count_mem_we    (func_qid_ldb_enqueue_count_mem_we)
,.func_qid_ldb_enqueue_count_mem_wdata (func_qid_ldb_enqueue_count_mem_wdata)
,.func_qid_ldb_enqueue_count_mem_rdata (func_qid_ldb_enqueue_count_mem_rdata)

,.pf_qid_ldb_enqueue_count_mem_re      (pf_qid_ldb_enqueue_count_mem_re)
,.pf_qid_ldb_enqueue_count_mem_raddr (pf_qid_ldb_enqueue_count_mem_raddr)
,.pf_qid_ldb_enqueue_count_mem_waddr (pf_qid_ldb_enqueue_count_mem_waddr)
,.pf_qid_ldb_enqueue_count_mem_we    (pf_qid_ldb_enqueue_count_mem_we)
,.pf_qid_ldb_enqueue_count_mem_wdata (pf_qid_ldb_enqueue_count_mem_wdata)
,.pf_qid_ldb_enqueue_count_mem_rdata (pf_qid_ldb_enqueue_count_mem_rdata)

,.rf_qid_ldb_enqueue_count_mem_rclk (rf_qid_ldb_enqueue_count_mem_rclk)
,.rf_qid_ldb_enqueue_count_mem_rclk_rst_n (rf_qid_ldb_enqueue_count_mem_rclk_rst_n)
,.rf_qid_ldb_enqueue_count_mem_re    (rf_qid_ldb_enqueue_count_mem_re)
,.rf_qid_ldb_enqueue_count_mem_raddr (rf_qid_ldb_enqueue_count_mem_raddr)
,.rf_qid_ldb_enqueue_count_mem_waddr (rf_qid_ldb_enqueue_count_mem_waddr)
,.rf_qid_ldb_enqueue_count_mem_wclk (rf_qid_ldb_enqueue_count_mem_wclk)
,.rf_qid_ldb_enqueue_count_mem_wclk_rst_n (rf_qid_ldb_enqueue_count_mem_wclk_rst_n)
,.rf_qid_ldb_enqueue_count_mem_we    (rf_qid_ldb_enqueue_count_mem_we)
,.rf_qid_ldb_enqueue_count_mem_wdata (rf_qid_ldb_enqueue_count_mem_wdata)
,.rf_qid_ldb_enqueue_count_mem_rdata (rf_qid_ldb_enqueue_count_mem_rdata)

,.rf_qid_ldb_enqueue_count_mem_error (rf_qid_ldb_enqueue_count_mem_error)

,.func_qid_ldb_inflight_count_mem_re    (func_qid_ldb_inflight_count_mem_re)
,.func_qid_ldb_inflight_count_mem_raddr (func_qid_ldb_inflight_count_mem_raddr)
,.func_qid_ldb_inflight_count_mem_waddr (func_qid_ldb_inflight_count_mem_waddr)
,.func_qid_ldb_inflight_count_mem_we    (func_qid_ldb_inflight_count_mem_we)
,.func_qid_ldb_inflight_count_mem_wdata (func_qid_ldb_inflight_count_mem_wdata)
,.func_qid_ldb_inflight_count_mem_rdata (func_qid_ldb_inflight_count_mem_rdata)

,.pf_qid_ldb_inflight_count_mem_re      (pf_qid_ldb_inflight_count_mem_re)
,.pf_qid_ldb_inflight_count_mem_raddr (pf_qid_ldb_inflight_count_mem_raddr)
,.pf_qid_ldb_inflight_count_mem_waddr (pf_qid_ldb_inflight_count_mem_waddr)
,.pf_qid_ldb_inflight_count_mem_we    (pf_qid_ldb_inflight_count_mem_we)
,.pf_qid_ldb_inflight_count_mem_wdata (pf_qid_ldb_inflight_count_mem_wdata)
,.pf_qid_ldb_inflight_count_mem_rdata (pf_qid_ldb_inflight_count_mem_rdata)

,.rf_qid_ldb_inflight_count_mem_rclk (rf_qid_ldb_inflight_count_mem_rclk)
,.rf_qid_ldb_inflight_count_mem_rclk_rst_n (rf_qid_ldb_inflight_count_mem_rclk_rst_n)
,.rf_qid_ldb_inflight_count_mem_re    (rf_qid_ldb_inflight_count_mem_re)
,.rf_qid_ldb_inflight_count_mem_raddr (rf_qid_ldb_inflight_count_mem_raddr)
,.rf_qid_ldb_inflight_count_mem_waddr (rf_qid_ldb_inflight_count_mem_waddr)
,.rf_qid_ldb_inflight_count_mem_wclk (rf_qid_ldb_inflight_count_mem_wclk)
,.rf_qid_ldb_inflight_count_mem_wclk_rst_n (rf_qid_ldb_inflight_count_mem_wclk_rst_n)
,.rf_qid_ldb_inflight_count_mem_we    (rf_qid_ldb_inflight_count_mem_we)
,.rf_qid_ldb_inflight_count_mem_wdata (rf_qid_ldb_inflight_count_mem_wdata)
,.rf_qid_ldb_inflight_count_mem_rdata (rf_qid_ldb_inflight_count_mem_rdata)

,.rf_qid_ldb_inflight_count_mem_error (rf_qid_ldb_inflight_count_mem_error)

,.func_qid_ldb_replay_count_mem_re    (func_qid_ldb_replay_count_mem_re)
,.func_qid_ldb_replay_count_mem_raddr (func_qid_ldb_replay_count_mem_raddr)
,.func_qid_ldb_replay_count_mem_waddr (func_qid_ldb_replay_count_mem_waddr)
,.func_qid_ldb_replay_count_mem_we    (func_qid_ldb_replay_count_mem_we)
,.func_qid_ldb_replay_count_mem_wdata (func_qid_ldb_replay_count_mem_wdata)
,.func_qid_ldb_replay_count_mem_rdata (func_qid_ldb_replay_count_mem_rdata)

,.pf_qid_ldb_replay_count_mem_re      (pf_qid_ldb_replay_count_mem_re)
,.pf_qid_ldb_replay_count_mem_raddr (pf_qid_ldb_replay_count_mem_raddr)
,.pf_qid_ldb_replay_count_mem_waddr (pf_qid_ldb_replay_count_mem_waddr)
,.pf_qid_ldb_replay_count_mem_we    (pf_qid_ldb_replay_count_mem_we)
,.pf_qid_ldb_replay_count_mem_wdata (pf_qid_ldb_replay_count_mem_wdata)
,.pf_qid_ldb_replay_count_mem_rdata (pf_qid_ldb_replay_count_mem_rdata)

,.rf_qid_ldb_replay_count_mem_rclk (rf_qid_ldb_replay_count_mem_rclk)
,.rf_qid_ldb_replay_count_mem_rclk_rst_n (rf_qid_ldb_replay_count_mem_rclk_rst_n)
,.rf_qid_ldb_replay_count_mem_re    (rf_qid_ldb_replay_count_mem_re)
,.rf_qid_ldb_replay_count_mem_raddr (rf_qid_ldb_replay_count_mem_raddr)
,.rf_qid_ldb_replay_count_mem_waddr (rf_qid_ldb_replay_count_mem_waddr)
,.rf_qid_ldb_replay_count_mem_wclk (rf_qid_ldb_replay_count_mem_wclk)
,.rf_qid_ldb_replay_count_mem_wclk_rst_n (rf_qid_ldb_replay_count_mem_wclk_rst_n)
,.rf_qid_ldb_replay_count_mem_we    (rf_qid_ldb_replay_count_mem_we)
,.rf_qid_ldb_replay_count_mem_wdata (rf_qid_ldb_replay_count_mem_wdata)
,.rf_qid_ldb_replay_count_mem_rdata (rf_qid_ldb_replay_count_mem_rdata)

,.rf_qid_ldb_replay_count_mem_error (rf_qid_ldb_replay_count_mem_error)

,.func_qid_naldb_max_depth_mem_re    (func_qid_naldb_max_depth_mem_re)
,.func_qid_naldb_max_depth_mem_raddr (func_qid_naldb_max_depth_mem_raddr)
,.func_qid_naldb_max_depth_mem_waddr (func_qid_naldb_max_depth_mem_waddr)
,.func_qid_naldb_max_depth_mem_we    (func_qid_naldb_max_depth_mem_we)
,.func_qid_naldb_max_depth_mem_wdata (func_qid_naldb_max_depth_mem_wdata)
,.func_qid_naldb_max_depth_mem_rdata (func_qid_naldb_max_depth_mem_rdata)

,.pf_qid_naldb_max_depth_mem_re      (pf_qid_naldb_max_depth_mem_re)
,.pf_qid_naldb_max_depth_mem_raddr (pf_qid_naldb_max_depth_mem_raddr)
,.pf_qid_naldb_max_depth_mem_waddr (pf_qid_naldb_max_depth_mem_waddr)
,.pf_qid_naldb_max_depth_mem_we    (pf_qid_naldb_max_depth_mem_we)
,.pf_qid_naldb_max_depth_mem_wdata (pf_qid_naldb_max_depth_mem_wdata)
,.pf_qid_naldb_max_depth_mem_rdata (pf_qid_naldb_max_depth_mem_rdata)

,.rf_qid_naldb_max_depth_mem_rclk (rf_qid_naldb_max_depth_mem_rclk)
,.rf_qid_naldb_max_depth_mem_rclk_rst_n (rf_qid_naldb_max_depth_mem_rclk_rst_n)
,.rf_qid_naldb_max_depth_mem_re    (rf_qid_naldb_max_depth_mem_re)
,.rf_qid_naldb_max_depth_mem_raddr (rf_qid_naldb_max_depth_mem_raddr)
,.rf_qid_naldb_max_depth_mem_waddr (rf_qid_naldb_max_depth_mem_waddr)
,.rf_qid_naldb_max_depth_mem_wclk (rf_qid_naldb_max_depth_mem_wclk)
,.rf_qid_naldb_max_depth_mem_wclk_rst_n (rf_qid_naldb_max_depth_mem_wclk_rst_n)
,.rf_qid_naldb_max_depth_mem_we    (rf_qid_naldb_max_depth_mem_we)
,.rf_qid_naldb_max_depth_mem_wdata (rf_qid_naldb_max_depth_mem_wdata)
,.rf_qid_naldb_max_depth_mem_rdata (rf_qid_naldb_max_depth_mem_rdata)

,.rf_qid_naldb_max_depth_mem_error (rf_qid_naldb_max_depth_mem_error)

,.func_qid_naldb_tot_enq_cnt_mem_re    (func_qid_naldb_tot_enq_cnt_mem_re)
,.func_qid_naldb_tot_enq_cnt_mem_raddr (func_qid_naldb_tot_enq_cnt_mem_raddr)
,.func_qid_naldb_tot_enq_cnt_mem_waddr (func_qid_naldb_tot_enq_cnt_mem_waddr)
,.func_qid_naldb_tot_enq_cnt_mem_we    (func_qid_naldb_tot_enq_cnt_mem_we)
,.func_qid_naldb_tot_enq_cnt_mem_wdata (func_qid_naldb_tot_enq_cnt_mem_wdata)
,.func_qid_naldb_tot_enq_cnt_mem_rdata (func_qid_naldb_tot_enq_cnt_mem_rdata)

,.pf_qid_naldb_tot_enq_cnt_mem_re      (pf_qid_naldb_tot_enq_cnt_mem_re)
,.pf_qid_naldb_tot_enq_cnt_mem_raddr (pf_qid_naldb_tot_enq_cnt_mem_raddr)
,.pf_qid_naldb_tot_enq_cnt_mem_waddr (pf_qid_naldb_tot_enq_cnt_mem_waddr)
,.pf_qid_naldb_tot_enq_cnt_mem_we    (pf_qid_naldb_tot_enq_cnt_mem_we)
,.pf_qid_naldb_tot_enq_cnt_mem_wdata (pf_qid_naldb_tot_enq_cnt_mem_wdata)
,.pf_qid_naldb_tot_enq_cnt_mem_rdata (pf_qid_naldb_tot_enq_cnt_mem_rdata)

,.rf_qid_naldb_tot_enq_cnt_mem_rclk (rf_qid_naldb_tot_enq_cnt_mem_rclk)
,.rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n (rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n)
,.rf_qid_naldb_tot_enq_cnt_mem_re    (rf_qid_naldb_tot_enq_cnt_mem_re)
,.rf_qid_naldb_tot_enq_cnt_mem_raddr (rf_qid_naldb_tot_enq_cnt_mem_raddr)
,.rf_qid_naldb_tot_enq_cnt_mem_waddr (rf_qid_naldb_tot_enq_cnt_mem_waddr)
,.rf_qid_naldb_tot_enq_cnt_mem_wclk (rf_qid_naldb_tot_enq_cnt_mem_wclk)
,.rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n (rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n)
,.rf_qid_naldb_tot_enq_cnt_mem_we    (rf_qid_naldb_tot_enq_cnt_mem_we)
,.rf_qid_naldb_tot_enq_cnt_mem_wdata (rf_qid_naldb_tot_enq_cnt_mem_wdata)
,.rf_qid_naldb_tot_enq_cnt_mem_rdata (rf_qid_naldb_tot_enq_cnt_mem_rdata)

,.rf_qid_naldb_tot_enq_cnt_mem_error (rf_qid_naldb_tot_enq_cnt_mem_error)

,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_re    (func_rop_lsp_reordercmp_rx_sync_fifo_mem_re)
,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr (func_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr)
,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr (func_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr)
,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_we    (func_rop_lsp_reordercmp_rx_sync_fifo_mem_we)
,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata (func_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata)
,.func_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata (func_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata)

,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_re      (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_re)
,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr)
,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr)
,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_we    (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_we)
,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata)
,.pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata (pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata)

,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re    (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we    (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata)
,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata)

,.rf_rop_lsp_reordercmp_rx_sync_fifo_mem_error (rf_rop_lsp_reordercmp_rx_sync_fifo_mem_error)

,.func_send_atm_to_cq_rx_sync_fifo_mem_re    (func_send_atm_to_cq_rx_sync_fifo_mem_re)
,.func_send_atm_to_cq_rx_sync_fifo_mem_raddr (func_send_atm_to_cq_rx_sync_fifo_mem_raddr)
,.func_send_atm_to_cq_rx_sync_fifo_mem_waddr (func_send_atm_to_cq_rx_sync_fifo_mem_waddr)
,.func_send_atm_to_cq_rx_sync_fifo_mem_we    (func_send_atm_to_cq_rx_sync_fifo_mem_we)
,.func_send_atm_to_cq_rx_sync_fifo_mem_wdata (func_send_atm_to_cq_rx_sync_fifo_mem_wdata)
,.func_send_atm_to_cq_rx_sync_fifo_mem_rdata (func_send_atm_to_cq_rx_sync_fifo_mem_rdata)

,.pf_send_atm_to_cq_rx_sync_fifo_mem_re      (pf_send_atm_to_cq_rx_sync_fifo_mem_re)
,.pf_send_atm_to_cq_rx_sync_fifo_mem_raddr (pf_send_atm_to_cq_rx_sync_fifo_mem_raddr)
,.pf_send_atm_to_cq_rx_sync_fifo_mem_waddr (pf_send_atm_to_cq_rx_sync_fifo_mem_waddr)
,.pf_send_atm_to_cq_rx_sync_fifo_mem_we    (pf_send_atm_to_cq_rx_sync_fifo_mem_we)
,.pf_send_atm_to_cq_rx_sync_fifo_mem_wdata (pf_send_atm_to_cq_rx_sync_fifo_mem_wdata)
,.pf_send_atm_to_cq_rx_sync_fifo_mem_rdata (pf_send_atm_to_cq_rx_sync_fifo_mem_rdata)

,.rf_send_atm_to_cq_rx_sync_fifo_mem_rclk (rf_send_atm_to_cq_rx_sync_fifo_mem_rclk)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n (rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_re    (rf_send_atm_to_cq_rx_sync_fifo_mem_re)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_raddr (rf_send_atm_to_cq_rx_sync_fifo_mem_raddr)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_waddr (rf_send_atm_to_cq_rx_sync_fifo_mem_waddr)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_wclk (rf_send_atm_to_cq_rx_sync_fifo_mem_wclk)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n (rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_we    (rf_send_atm_to_cq_rx_sync_fifo_mem_we)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_wdata (rf_send_atm_to_cq_rx_sync_fifo_mem_wdata)
,.rf_send_atm_to_cq_rx_sync_fifo_mem_rdata (rf_send_atm_to_cq_rx_sync_fifo_mem_rdata)

,.rf_send_atm_to_cq_rx_sync_fifo_mem_error (rf_send_atm_to_cq_rx_sync_fifo_mem_error)

,.func_uno_atm_cmp_fifo_mem_re    (func_uno_atm_cmp_fifo_mem_re)
,.func_uno_atm_cmp_fifo_mem_raddr (func_uno_atm_cmp_fifo_mem_raddr)
,.func_uno_atm_cmp_fifo_mem_waddr (func_uno_atm_cmp_fifo_mem_waddr)
,.func_uno_atm_cmp_fifo_mem_we    (func_uno_atm_cmp_fifo_mem_we)
,.func_uno_atm_cmp_fifo_mem_wdata (func_uno_atm_cmp_fifo_mem_wdata)
,.func_uno_atm_cmp_fifo_mem_rdata (func_uno_atm_cmp_fifo_mem_rdata)

,.pf_uno_atm_cmp_fifo_mem_re      (pf_uno_atm_cmp_fifo_mem_re)
,.pf_uno_atm_cmp_fifo_mem_raddr (pf_uno_atm_cmp_fifo_mem_raddr)
,.pf_uno_atm_cmp_fifo_mem_waddr (pf_uno_atm_cmp_fifo_mem_waddr)
,.pf_uno_atm_cmp_fifo_mem_we    (pf_uno_atm_cmp_fifo_mem_we)
,.pf_uno_atm_cmp_fifo_mem_wdata (pf_uno_atm_cmp_fifo_mem_wdata)
,.pf_uno_atm_cmp_fifo_mem_rdata (pf_uno_atm_cmp_fifo_mem_rdata)

,.rf_uno_atm_cmp_fifo_mem_rclk (rf_uno_atm_cmp_fifo_mem_rclk)
,.rf_uno_atm_cmp_fifo_mem_rclk_rst_n (rf_uno_atm_cmp_fifo_mem_rclk_rst_n)
,.rf_uno_atm_cmp_fifo_mem_re    (rf_uno_atm_cmp_fifo_mem_re)
,.rf_uno_atm_cmp_fifo_mem_raddr (rf_uno_atm_cmp_fifo_mem_raddr)
,.rf_uno_atm_cmp_fifo_mem_waddr (rf_uno_atm_cmp_fifo_mem_waddr)
,.rf_uno_atm_cmp_fifo_mem_wclk (rf_uno_atm_cmp_fifo_mem_wclk)
,.rf_uno_atm_cmp_fifo_mem_wclk_rst_n (rf_uno_atm_cmp_fifo_mem_wclk_rst_n)
,.rf_uno_atm_cmp_fifo_mem_we    (rf_uno_atm_cmp_fifo_mem_we)
,.rf_uno_atm_cmp_fifo_mem_wdata (rf_uno_atm_cmp_fifo_mem_wdata)
,.rf_uno_atm_cmp_fifo_mem_rdata (rf_uno_atm_cmp_fifo_mem_rdata)

,.rf_uno_atm_cmp_fifo_mem_error (rf_uno_atm_cmp_fifo_mem_error)

);
// END HQM_RAM_ACCESS
//---------------------------------------------------------------------------------------------------------
// common core - Interface & clock control

logic wire_lsp_unit_idle ;

assign aqed_intf_idle           = aqed_lsp_dec_fid_cnt_v_idle & atq_fid_cnt_upd_idle & atq_stop_atqatm_idle ;

hqm_AW_module_clock_control # ( .REQS ( 12 ) ) i_hqm_AW_module_clock_control (
          .hqm_inp_gated_clk                    ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n                  ( hqm_inp_gated_rst_n )

        , .hqm_gated_clk                        ( hqm_gated_clk )
        , .hqm_gated_rst_n                      ( hqm_gated_rst_n )

        , .cfg_co_dly                           ( { 2'd0 , hqm_lsp_target_cfg_patch_control_reg_f [ 13 : 0 ] } ) 
        , .cfg_co_disable                       ( hqm_lsp_target_cfg_patch_control_reg_f [ 31 ] ) 

        , .hqm_proc_clk_en                      ( hqm_proc_clk_en_lsp )

        , .unit_idle_local                      ( lsp_unit_idle_local )
        , .unit_idle                            ( wire_lsp_unit_idle )



        , .inp_fifo_empty                       ( {       aqed_intf_idle
                                                        , atm_clk_idle
                                                        , aqed_clk_idle
                                                        , cfg_rx_idle
                                                        , chp_lsp_token_rx_sync_idle
                                                        , chp_lsp_cmp_rx_sync_idle
                                                        , rop_lsp_reordercmp_rx_sync_idle
                                                        , nalb_lsp_enq_lb_rx_sync_idle
                                                        , dp_lsp_enq_dir_rx_sync_idle
                                                        , dp_lsp_enq_rorply_rx_sync_idle
                                                        , send_atm_to_cq_rx_sync_idle 
                                                        , nalb_lsp_enq_rorply_rx_sync_idle
                                                  } )
        , .inp_fifo_en                          ( {       aqed_intf_enable_nc
                                                        , atm_clk_enable
                                                        , aqed_clk_enable
                                                        , cfg_rx_enable
                                                        , chp_lsp_token_rx_sync_enable
                                                        , chp_lsp_cmp_rx_sync_enable
                                                        , rop_lsp_reordercmp_rx_sync_enable
                                                        , nalb_lsp_enq_lb_rx_sync_enable
                                                        , dp_lsp_enq_dir_rx_sync_enable
                                                        , dp_lsp_enq_rorply_rx_sync_enable
                                                        , send_atm_to_cq_rx_sync_enable 
                                                        , nalb_lsp_enq_rorply_rx_sync_enable
                                                  } )
        , .cfg_idle                             ( cfg_idle )
        , .int_idle                             ( int_idle )

        , .rst_prep                             ( rst_prep )
        , .reset_active                         ( hqm_gated_rst_n_active )
) ;

assign cfg_rx_sync_fifo_of              = cfg_rx_fifo_status_pnc.overflow ;
assign cfg_rx_sync_fifo_uf              = cfg_rx_fifo_status_pnc.underflow ;

// Note: The chp_lsp_token_t struct/interface includes a 4-bit cmd field which is unused by LSP and not stored in the rx_sync FIFO memory.
// Since the interfaces are defined in terms of the struct these 4 ms bits (unused by LSP) must be stripped off when referencing the memory.
logic [3:0]             func_chp_lsp_token_rx_sync_fifo_mem_wdata_spare_cmd_nc ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( chp_lsp_token_data ) ) , .SEED ( 32'h0f ) ) i_hqm_AW_rx_sync_chp_lsp_token (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( chp_lsp_token_fifo_status_pnc )

        , .enable                       ( chp_lsp_token_rx_sync_enable )
        , .idle                         ( chp_lsp_token_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( chp_lsp_token_ready )
        , .in_valid                     ( chp_lsp_token_v )
        , .in_data                      ( chp_lsp_token_data )
        , .out_ready                    ( core_chp_lsp_token_ready )
        , .out_valid                    ( core_chp_lsp_token_v )
        , .out_data                     ( core_chp_lsp_token_data )

        , .mem_we                       ( func_chp_lsp_token_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_chp_lsp_token_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( { func_chp_lsp_token_rx_sync_fifo_mem_wdata_spare_cmd_nc , func_chp_lsp_token_rx_sync_fifo_mem_wdata } )    // Truncate unused cmd field
        , .mem_re                       ( func_chp_lsp_token_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_chp_lsp_token_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( { 4'h0 , func_chp_lsp_token_rx_sync_fifo_mem_rdata } )                                                      // Truncate unused cmd field



        , .agit_enable                  ( cfg_agitate_select_f [0] )
        , .agit_control                 ( cfg_agitate_control_f )
) ;

assign chp_lsp_token_rx_sync_fifo_of    = chp_lsp_token_fifo_status_pnc.overflow ;
assign chp_lsp_token_rx_sync_fifo_uf    = chp_lsp_token_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( chp_lsp_cmp_data ) ) , .SEED ( 32'h1e ) ) i_hqm_AW_rx_sync_chp_lsp_cmp (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( chp_lsp_cmp_fifo_status_pnc )

        , .enable                       ( chp_lsp_cmp_rx_sync_enable )
        , .idle                         ( chp_lsp_cmp_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( chp_lsp_cmp_ready )
        , .in_valid                     ( chp_lsp_cmp_v )
        , .in_data                      ( chp_lsp_cmp_data )
        , .out_ready                    ( core_chp_lsp_cmp_ready )
        , .out_valid                    ( core_chp_lsp_cmp_v )
        , .out_data                     ( core_chp_lsp_cmp_data )

        , .mem_we                       ( func_chp_lsp_cmp_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_chp_lsp_cmp_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_chp_lsp_cmp_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_chp_lsp_cmp_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_chp_lsp_cmp_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_chp_lsp_cmp_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [1] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign chp_lsp_cmp_rx_sync_fifo_of      = chp_lsp_cmp_fifo_status_pnc.overflow ;
assign chp_lsp_cmp_rx_sync_fifo_uf      = chp_lsp_cmp_fifo_status_pnc.underflow ;

// Depth increased to 8 to absorb previous 8-deep rop_ord_cmp_fifo functionality
hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( rop_lsp_reordercmp_data ) ) , .DEPTH ( 8 ) , .SEED ( 32'h2d ) ) i_hqm_AW_rx_sync_rop_lsp_reordercmp (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( rop_lsp_reordercmp_fifo_status_pnc )

        , .enable                       ( rop_lsp_reordercmp_rx_sync_enable )
        , .idle                         ( rop_lsp_reordercmp_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( rop_lsp_reordercmp_ready )
        , .in_valid                     ( rop_lsp_reordercmp_v )
        , .in_data                      ( rop_lsp_reordercmp_data )
        , .out_ready                    ( core_rop_lsp_reordercmp_ready )
        , .out_valid                    ( core_rop_lsp_reordercmp_v )
        , .out_data                     ( core_rop_lsp_reordercmp_data )

        , .mem_we                       ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [2] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign rop_lsp_reordercmp_rx_sync_fifo_of       = rop_lsp_reordercmp_fifo_status_pnc.overflow ;
assign rop_lsp_reordercmp_rx_sync_fifo_uf       = rop_lsp_reordercmp_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( nalb_lsp_enq_lb_data ) ) , .SEED ( 32'h3c ) ) i_hqm_AW_rx_sync_nalb_lsp_enq_lb (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( nalb_lsp_enq_lb_fifo_status_pnc )

        , .enable                       ( nalb_lsp_enq_lb_rx_sync_enable )
        , .idle                         ( nalb_lsp_enq_lb_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( nalb_lsp_enq_lb_ready )
        , .in_valid                     ( nalb_lsp_enq_lb_v )
        , .in_data                      ( nalb_lsp_enq_lb_data )
        , .out_ready                    ( core_nalb_lsp_enq_lb_ready )
        , .out_valid                    ( core_nalb_lsp_enq_lb_v )
        , .out_data                     ( core_nalb_lsp_enq_lb_data )

        , .mem_we                       ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [3] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign nalb_lsp_enq_lb_rx_sync_fifo_of  = nalb_lsp_enq_lb_fifo_status_pnc.overflow ;
assign nalb_lsp_enq_lb_rx_sync_fifo_uf  = nalb_lsp_enq_lb_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( dp_lsp_enq_dir_data ) ) , .SEED ( 32'h4b ) ) i_hqm_AW_rx_sync_dp_lsp_enq_dir (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( dp_lsp_enq_dir_fifo_status_pnc )

        , .enable                       ( dp_lsp_enq_dir_rx_sync_enable )
        , .idle                         ( dp_lsp_enq_dir_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( dp_lsp_enq_dir_ready )
        , .in_valid                     ( dp_lsp_enq_dir_v )
        , .in_data                      ( dp_lsp_enq_dir_data )
        , .out_ready                    ( core_dp_lsp_enq_dir_ready )
        , .out_valid                    ( core_dp_lsp_enq_dir_v )
        , .out_data                     ( core_dp_lsp_enq_dir_data )

        , .mem_we                       ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [4] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign dp_lsp_enq_dir_rx_sync_fifo_of   = dp_lsp_enq_dir_fifo_status_pnc.overflow ;
assign dp_lsp_enq_dir_rx_sync_fifo_uf   = dp_lsp_enq_dir_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( dp_lsp_enq_rorply_data ) ) , .SEED ( 32'h5a ) ) i_hqm_AW_rx_sync_dp_lsp_enq_rorply (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( dp_lsp_enq_rorply_fifo_status_pnc )

        , .enable                       ( dp_lsp_enq_rorply_rx_sync_enable )
        , .idle                         ( dp_lsp_enq_rorply_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( dp_lsp_enq_rorply_ready )
        , .in_valid                     ( dp_lsp_enq_rorply_v )
        , .in_data                      ( dp_lsp_enq_rorply_data )
        , .out_ready                    ( core_dp_lsp_enq_rorply_ready )
        , .out_valid                    ( core_dp_lsp_enq_rorply_v )
        , .out_data                     ( core_dp_lsp_enq_rorply_data )

        , .mem_we                       ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [5] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign dp_lsp_enq_rorply_rx_sync_fifo_of        = dp_lsp_enq_rorply_fifo_status_pnc.overflow ;
assign dp_lsp_enq_rorply_rx_sync_fifo_uf        = dp_lsp_enq_rorply_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( aqed_lsp_sch_data ) ) , .SEED ( 32'h69 ) ) i_hqm_AW_rx_sync_send_atm_to_cq (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( send_atm_to_cq_fifo_status_pnc )

        , .enable                       ( send_atm_to_cq_rx_sync_enable )
        , .idle                         ( send_atm_to_cq_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( aqed_lsp_sch_ready )
        , .in_valid                     ( aqed_lsp_sch_v )
        , .in_data                      ( aqed_lsp_sch_data )
        , .out_ready                    ( send_atm_to_cq_ready )
        , .out_valid                    ( send_atm_to_cq_v )
        , .out_data                     ( send_atm_to_cq_data )

        , .mem_we                       ( func_send_atm_to_cq_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_send_atm_to_cq_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_send_atm_to_cq_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_send_atm_to_cq_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_send_atm_to_cq_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_send_atm_to_cq_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [6] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign send_atm_to_cq_rx_sync_fifo_of   = send_atm_to_cq_fifo_status_pnc.overflow ;
assign send_atm_to_cq_rx_sync_fifo_uf   = send_atm_to_cq_fifo_status_pnc.underflow ;

hqm_AW_rx_sync_wagitate # ( .WIDTH ( $bits ( nalb_lsp_enq_rorply_data ) ) , .SEED ( 32'h78 ) ) i_hqm_AW_rx_sync_nalb_lsp_enq_rorply (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )

        , .status                       ( nalb_lsp_enq_rorply_fifo_status_pnc )

        , .enable                       ( nalb_lsp_enq_rorply_rx_sync_enable )
        , .idle                         ( nalb_lsp_enq_rorply_rx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( nalb_lsp_enq_rorply_ready )
        , .in_valid                     ( nalb_lsp_enq_rorply_v )
        , .in_data                      ( nalb_lsp_enq_rorply_data )
        , .out_ready                    ( core_nalb_lsp_enq_rorply_ready )
        , .out_valid                    ( core_nalb_lsp_enq_rorply_v )
        , .out_data                     ( core_nalb_lsp_enq_rorply_data )

        , .mem_we                       ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we )
        , .mem_waddr                    ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr )
        , .mem_wdata                    ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata )
        , .mem_re                       ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re )
        , .mem_raddr                    ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr )
        , .mem_rdata                    ( func_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata )



        , .agit_enable                  ( cfg_agitate_select_f [7] )
        , .agit_control                 ( cfg_agitate_control_f )

) ;

assign nalb_lsp_enq_rorply_rx_sync_fifo_of      = nalb_lsp_enq_rorply_fifo_status_pnc.overflow ;
assign nalb_lsp_enq_rorply_rx_sync_fifo_uf      = nalb_lsp_enq_rorply_fifo_status_pnc.underflow ;

assign rx_sync_fifo_error       = | {   cfg_rx_sync_fifo_of
                                      , cfg_rx_sync_fifo_uf
                                      , chp_lsp_token_rx_sync_fifo_of 
                                      , chp_lsp_token_rx_sync_fifo_uf
                                      , chp_lsp_cmp_rx_sync_fifo_of
                                      , chp_lsp_cmp_rx_sync_fifo_uf
                                      , rop_lsp_reordercmp_rx_sync_fifo_of
                                      , rop_lsp_reordercmp_rx_sync_fifo_uf
                                      , nalb_lsp_enq_lb_rx_sync_fifo_of
                                      , nalb_lsp_enq_lb_rx_sync_fifo_uf
                                      , dp_lsp_enq_dir_rx_sync_fifo_of
                                      , dp_lsp_enq_dir_rx_sync_fifo_uf
                                      , dp_lsp_enq_rorply_rx_sync_fifo_of
                                      , dp_lsp_enq_rorply_rx_sync_fifo_uf
                                      , send_atm_to_cq_rx_sync_fifo_of
                                      , send_atm_to_cq_rx_sync_fifo_uf
                                      , nalb_lsp_enq_rorply_rx_sync_fifo_of
                                      , nalb_lsp_enq_rorply_rx_sync_fifo_uf } ;


hqm_AW_tx_sync # ( .WIDTH ( $bits ( lsp_nalb_sch_rorply_data ) ) ) i_hqm_AW_tx_sync_rpl_ldb_nalb (
          .hqm_gated_clk                ( hqm_gated_clk )
        , .hqm_gated_rst_n              ( hqm_gated_rst_n )

        , .status                       ( rpl_ldb_nalb_db_status_pnc )          // Feeds lsp_nalb_sch_rorplywhich is cfg readable in cfg_interface_status
        , .idle                         ( rpl_ldb_nalb_tx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( rpl_ldb_nalb_db_in_ready )
        , .in_valid                     ( rpl_ldb_nalb_db_in_valid )
        , .in_data                      ( rpl_ldb_nalb_db_in_data )
        , .out_ready                    ( lsp_nalb_sch_rorply_ready )
        , .out_valid                    ( lsp_nalb_sch_rorply_v )
        , .out_data                     ( lsp_nalb_sch_rorply_data )
) ;

hqm_AW_tx_sync # ( .WIDTH ( $bits ( lsp_nalb_sch_unoord_data ) ) ) i_hqm_AW_tx_sync_lsp_nalb_sch_unoord (
          .hqm_gated_clk                ( hqm_gated_clk )
        , .hqm_gated_rst_n              ( hqm_gated_rst_n )

        , .status                       ( lsp_nalb_sch_unoord_status_pnc )      // Feeds lsp_nalb_sch_unoord which is cfg readable in cfg_interface_status
        , .idle                         ( lsp_nalb_sch_unoord_tx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( lsp_nalb_sch_unoord_in_ready )
        , .in_valid                     ( nalb_sel_nalb_fifo_pop_data_v )
        , .in_data                      ( nalb_sel_nalb_fifo_pop_data )
        , .out_ready                    ( lsp_nalb_sch_unoord_ready )
        , .out_valid                    ( lsp_nalb_sch_unoord_v )
        , .out_data                     ( lsp_nalb_sch_unoord_data )
) ;

hqm_AW_tx_sync # ( .WIDTH ( $bits ( lsp_nalb_sch_atq_data ) ) ) i_hqm_AW_tx_sync_atq_sel_ap (
          .hqm_gated_clk                ( hqm_gated_clk )
        , .hqm_gated_rst_n              ( hqm_gated_rst_n )

        , .status                       ( atq_sel_ap_db_status_pnc )            // Feeds lsp_nalb_sch_atq which is cfg readable in cfg_interface_status
        , .idle                         ( atq_sel_ap_tx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( atq_sel_ap_db_in_ready )
        , .in_valid                     ( atq_sel_ap_db_in_valid )
        , .in_data                      ( atq_sel_ap_db_in_data )
        , .out_ready                    ( lsp_nalb_sch_atq_ready )
        , .out_valid                    ( lsp_nalb_sch_atq_v )
        , .out_data                     ( lsp_nalb_sch_atq_data )
) ;

hqm_AW_tx_sync # ( .WIDTH ( $bits ( lsp_dp_sch_dir_pre_data ) ) ) i_hqm_AW_tx_sync_lsp_dp_sch_dir (
          .hqm_gated_clk                ( hqm_gated_clk )
        , .hqm_gated_rst_n              ( hqm_gated_rst_n )

        , .status                       ( dir_sel_dp_db_status_nc )             // Feeds lsp_dp_sch_dir which is cfg readable in cfg_interface_status
        , .idle                         ( lsp_dp_sch_dir_tx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( dir_sel_dp_db_in_ready )
        , .in_valid                     ( dir_sel_dp_db_in_valid )
        , .in_data                      ( dir_sel_dp_db_in_data )
        , .out_ready                    ( lsp_dp_sch_dir_ready )
        , .out_valid                    ( lsp_dp_sch_dir_v )
        , .out_data                     ( lsp_dp_sch_dir_pre_data )
) ;

hqm_AW_tx_sync # ( .WIDTH ( $bits ( lsp_dp_sch_rorply_data ) ) ) i_hqm_AW_tx_sync_rpl_dir_dp (
          .hqm_gated_clk                ( hqm_gated_clk )
        , .hqm_gated_rst_n              ( hqm_gated_rst_n )

        , .status                       ( rpl_dir_dp_db_status_pnc )            // Feeds lsp_dp_sch_rorply which is cfg readable in cfg_interface_status
        , .idle                         ( rpl_dir_dp_tx_sync_idle )
        , .rst_prep                     ( rst_prep )

        , .in_ready                     ( rpl_dir_dp_db_in_ready )
        , .in_valid                     ( rpl_dir_dp_db_in_valid )
        , .in_data                      ( rpl_dir_dp_db_in_data )
        , .out_ready                    ( lsp_dp_sch_rorply_ready )
        , .out_valid                    ( lsp_dp_sch_rorply_v )
        , .out_data                     ( lsp_dp_sch_rorply_data )
) ;


//---------------------------------------------------------------------------------------------------------
// common core - Configuration Ring & config sidecar

cfg_req_t unit_cfg_req ;
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] unit_cfg_req_write ;
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] unit_cfg_req_read ;
logic unit_cfg_rsp_ack ;
logic unit_cfg_rsp_err ;
logic [31:0] unit_cfg_rsp_rdata ;
hqm_AW_cfg_ring_top # (
          .NODE_ID                     ( HQM_LSP_CFG_NODE_ID )
        , .UNIT_ID                     ( HQM_LSP_CFG_UNIT_ID )
        , .UNIT_TGT_MAP                ( HQM_LSP_CFG_UNIT_TGT_MAP )
        , .UNIT_NUM_TGTS               ( HQM_LSP_CFG_UNIT_NUM_TGTS )
) i_hqm_aw_cfg_ring_top (
          .hqm_inp_gated_clk           ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n         ( hqm_inp_gated_rst_n )
        , .hqm_gated_clk               ( hqm_gated_clk )
        , .hqm_gated_rst_n             ( hqm_gated_rst_n )
        , .rst_prep                    ( rst_prep )

        , .cfg_rx_enable               ( cfg_rx_enable )
        , .cfg_rx_idle                 ( cfg_rx_idle )
        , .cfg_rx_fifo_status          ( cfg_rx_fifo_status_pnc )
        , .cfg_idle                    ( cfg_idle )

        , .up_cfg_req_write            ( lsp_cfg_req_up_write )
        , .up_cfg_req_read             ( lsp_cfg_req_up_read )
        , .up_cfg_req                  ( lsp_cfg_req_up )
        , .up_cfg_rsp_ack              ( lsp_cfg_rsp_up_ack )
        , .up_cfg_rsp                  ( lsp_cfg_rsp_up )

        , .down_cfg_req_write          ( lsp_cfg_req_down_write )
        , .down_cfg_req_read           ( lsp_cfg_req_down_read )
        , .down_cfg_req                ( lsp_cfg_req_down )
        , .down_cfg_rsp_ack            ( lsp_cfg_rsp_down_ack )
        , .down_cfg_rsp                ( lsp_cfg_rsp_down )

        , .unit_cfg_req_write          ( unit_cfg_req_write )
        , .unit_cfg_req_read           ( unit_cfg_req_read )
        , .unit_cfg_req                ( unit_cfg_req )
        , .unit_cfg_rsp_ack            ( unit_cfg_rsp_ack )
        , .unit_cfg_rsp_rdata          ( unit_cfg_rsp_rdata )
        , .unit_cfg_rsp_err            ( unit_cfg_rsp_err )
) ;
//------------------------------------------------------------------------------------------------------------------
// Common BCAST/VF Reset logic

logic [15:0] timeout_nc ;
cfg_unit_timeout_t  cfg_unit_timeout;
assign hqm_lsp_target_cfg_unit_timeout_reg_nxt = {hqm_lsp_target_cfg_unit_timeout_reg_f[31:5],5'd31};
assign cfg_unit_timeout = {hqm_lsp_target_cfg_unit_timeout_reg_f[31:5],5'd31};
assign timeout_nc = { cfg_unit_timeout[30:20] , hqm_lsp_target_cfg_unit_timeout_reg_f[4:0] } ;

localparam VERSION = 8'h00 ;
cfg_unit_version_t cfg_unit_version;
assign cfg_unit_version.VERSION = VERSION;
assign cfg_unit_version.SPARE   = '0;
assign hqm_lsp_target_cfg_unit_version_status = cfg_unit_version;

//------------------------------------------------------------------------------------------------------------------

logic cfg_req_idlepipe ;
logic cfg_req_ready ;
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] cfg_req_write_pnc ;
logic [ ( HQM_LSP_CFG_UNIT_NUM_TGTS ) - 1 : 0 ] cfg_req_read_nc ;

logic [31:0]                            cfgsc_cfg_mem_wdata ;
logic                                   cfgsc_cfg_mem_wdata_par ;
logic [1:0]                             cfgsc_cfg_mem_wdata_res ;
logic [NUM_CFG_ACCESSIBLE_RAM-1:0]      cfgsc_cfg_mem_re ;
logic [NUM_CFG_ACCESSIBLE_RAM-1:0]      cfgsc_cfg_mem_we ;
logic [ ( NUM_CFG_ACCESSIBLE_RAM * 32 ) - 1 : 0 ] cfgsc_cfg_mem_rdata ;
logic [NUM_CFG_ACCESSIBLE_RAM-1:0]      cfgsc_cfg_mem_ack ;

hqm_AW_cfg_sc # (
          .MODULE                      ( HQM_LSP_CFG_NODE_ID )
        , .NUM_CFG_TARGETS             ( HQM_LSP_CFG_UNIT_NUM_TGTS )
        , .NUM_CFG_ACCESSIBLE_RAM      ( NUM_CFG_ACCESSIBLE_RAM )
) i_hqm_AW_cfg_sc (
          .hqm_gated_clk               ( hqm_gated_clk )
        , .hqm_gated_rst_n             ( hqm_gated_rst_n )

        , .unit_cfg_req_write          ( unit_cfg_req_write )
        , .unit_cfg_req_read           ( unit_cfg_req_read )
        , .unit_cfg_req                ( unit_cfg_req )
        , .unit_cfg_rsp_ack            ( unit_cfg_rsp_ack )
        , .unit_cfg_rsp_rdata          ( unit_cfg_rsp_rdata )
        , .unit_cfg_rsp_err            ( unit_cfg_rsp_err )

        , .pfcsr_cfg_req_write         ( pfcsr_cfg_req_write )
        , .pfcsr_cfg_req_read          ( pfcsr_cfg_req_read )
        , .pfcsr_cfg_req               ( pfcsr_cfg_req )
        , .pfcsr_cfg_rsp_ack           ( pfcsr_cfg_rsp_ack )
        , .pfcsr_cfg_rsp_err           ( pfcsr_cfg_rsp_err )
        , .pfcsr_cfg_rsp_rdata         ( pfcsr_cfg_rsp_rdata )

        , .cfg_req_write               ( cfg_req_write_pnc )
        , .cfg_req_read                ( cfg_req_read_nc )

        , .cfg_mem_re                  ( cfgsc_cfg_mem_re )
        , .cfg_mem_addr                ( cfg_mem_addr )
        , .cfg_mem_minbit              ( cfg_mem_minbit )
        , .cfg_mem_maxbit              ( cfg_mem_maxbit )
        , .cfg_mem_we                  ( cfgsc_cfg_mem_we )
        , .cfg_mem_wdata               ( cfgsc_cfg_mem_wdata )
        , .cfg_mem_rdata               ( cfgsc_cfg_mem_rdata )
        , .cfg_mem_ack                 ( cfgsc_cfg_mem_ack )
        , .cfg_req_idlepipe            ( cfg_req_idlepipe )
        , .cfg_req_ready               ( cfg_req_ready )

        , .cfg_timout_enable           ( cfg_unit_timeout.ENABLE )
        , .cfg_timout_threshold        ( cfg_unit_timeout.THRESHOLD )
);

//---------------------------------------------------------------------------------------------------------
// common core - Interrupt serializer. Capture all interrutps from unit and send on interrupt ring

hqm_AW_int_serializer # (
          .NUM_INF                      ( HQM_LSP_ALARM_NUM_INF )
        , .NUM_COR                      ( HQM_LSP_ALARM_NUM_COR )
        , .NUM_UNC                      ( HQM_LSP_ALARM_NUM_UNC )
) i_hqm_aw_int_serializer (
          .hqm_inp_gated_clk            ( hqm_inp_gated_clk )
        , .hqm_inp_gated_rst_n          ( hqm_inp_gated_rst_n )
        , .rst_prep                     ( rst_prep )


        , .unit                         ( lsp_uid )

        , .inf_v                        ( int_inf_v )
        , .inf_data                     ( int_inf_data )

        , .cor_v                        ( int_cor_v )
        , .cor_data                     ( int_cor_data )

        , .unc_v                        ( int_unc_v )
        , .unc_data                     ( int_unc_data )

        , .int_up_v                     ( lsp_alarm_up_v )
        , .int_up_data                  ( lsp_alarm_up_data )
        , .int_up_ready                 ( lsp_alarm_up_ready )

        , .int_down_v                   ( lsp_alarm_down_v )
        , .int_down_data                ( lsp_alarm_down_data )
        , .int_down_ready               ( lsp_alarm_down_ready )

        , .status                       ( int_serializer_status_pnc )
        , .int_idle                     ( int_idle )    // Interrupt serializer's contribution to unit idle
) ;

//---------------------------------------------------------------------------------------------------------
// Config sidecar glue logic

hqm_AW_parity_gen #( .WIDTH ( 32 ) ) i_cfgsc_cfg_mem_wdata_par_gen (      // If width < 32, will be zero padded in AW cfg logic
          .d                    ( cfg_mem_wdata )
        , .odd                  ( 1'b1 )
        , .p                    ( cfgsc_cfg_mem_wdata_par )
);

hqm_AW_residue_gen #( .WIDTH ( 32 ) ) i_cfgsc_cfg_mem_wdata_res_gen (
          .a                    ( cfg_mem_wdata )
        , .r                    ( cfgsc_cfg_mem_wdata_res )
) ;

// HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_COUNT
assign cfgsc_dir_tok_cnt_mem_we                 = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_DIR_TOK_CNT_MEM ] ;
assign cfgsc_dir_tok_cnt_mem_wdata_struct       = cfgsc_cfg_mem_wdata [12:0] ;                  // Will get linra warning if size of struct changes
assign cfgsc_dir_tok_cnt_mem_wdata_struct_cnt_res_nc    = cfgsc_dir_tok_cnt_mem_wdata_struct.cnt_res ;

// HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_DEPTH_SELECT_DSI
assign cfgsc_dir_tok_lim_mem_we                 = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_DIR_TOK_LIM_MEM ] ;
assign cfgsc_dir_tok_lim_mem_wdata_struct       = cfgsc_cfg_mem_wdata [7:0] ;                   // Will get linra warning if size of struct changes
assign cfgsc_dir_tok_lim_mem_wdata_struct_spare_nc      = cfgsc_dir_tok_lim_mem_wdata_struct.spare ;
assign cfgsc_dir_tok_lim_mem_wdata_struct_lim_p_nc      = cfgsc_dir_tok_lim_mem_wdata_struct.lim_p ;

// HQM_LSP_TARGET_CFG_CQ2PRIOV
assign cfgsc_cfg_cq2priov_mem_we                = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM ] ;
assign cfgsc_cfg_cq2priov_mem_wdata             = { cfgsc_cfg_mem_wdata_par , cfg_mem_wdata } ;                 // No formatting required
assign cfgsc_cfg_cq2priov_mem_re                = cfgsc_cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM ] ;
// HQM_LSP_TARGET_CFG_CQ2QID0
assign cfgsc_cfg_cq2qid_0_mem_we                = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM ] ;
assign cfgsc_cfg_cq2qid_0_mem_wdata             = { cfgsc_cfg_mem_wdata_par , cfg_mem_wdata [27:0] } ;          // Formatting already done
assign cfgsc_cfg_cq2qid_0_mem_re                = cfgsc_cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM ] ;
// HQM_LSP_TARGET_CFG_CQ2QID1
assign cfgsc_cfg_cq2qid_1_mem_we                = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM ] ;
assign cfgsc_cfg_cq2qid_1_mem_wdata             = { cfgsc_cfg_mem_wdata_par , cfg_mem_wdata [27:0] } ;          // Formatting already done
assign cfgsc_cfg_cq2qid_1_mem_re                = cfgsc_cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM ] ;

// HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_COUNT
assign cfgsc_qid_ldb_inflight_count_mem_we                      = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_LDB_INFLIGHT_COUNT_MEM ] ;
assign cfgsc_qid_ldb_inflight_count_mem_wdata_struct            = cfgsc_cfg_mem_wdata [13:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_qid_ldb_inflight_count_mem_wdata_struct_cnt_res_nc = cfgsc_qid_ldb_inflight_count_mem_wdata_struct.cnt_res ;

// HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_LIMIT
assign cfgsc_cfg_qid_ldb_inflight_limit_mem_we                  = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_QID_LDB_INFLIGHT_LIMIT_MEM ] ;
assign cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct        = cfgsc_cfg_mem_wdata [12:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct_lim_p_nc       = cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct.lim_p ;

// HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_0 .. _15
assign cfgsc_cfg_qid_ldb_qid2cqidix_mem_we      = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_QID_LDB_QID2CQIDIX_MEM ] ;
// HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_0 .. _15
assign cfgsc_cfg_qid_ldb_qid2cqidix2_mem_we     = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_QID_LDB_QID2CQIDIX2_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_COUNT
assign cfgsc_cq_ldb_token_count_mem_we          = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_TOKEN_COUNT_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_DEPTH_SELECT
assign cfgsc_cfg_cq_ldb_token_depth_select_mem_we               = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_TOKEN_DEPTH_SELECT_MEM ] ;
assign cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct     = cfgsc_cfg_mem_wdata [4:0] ;   // Will get linra warning if size of struct changes
assign cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct_lim_p_nc    = cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct.lim_p ;

// HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_COUNT
assign cfgsc_cq_ldb_inflight_count_mem_we                       = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_INFLIGHT_COUNT_MEM ] ;
assign cfgsc_cq_ldb_inflight_count_mem_wdata_struct             = cfgsc_cfg_mem_wdata [13:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_cq_ldb_inflight_count_mem_wdata_struct_cnt_res_nc  = cfgsc_cq_ldb_inflight_count_mem_wdata_struct.cnt_res ;

// HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_LIMIT
assign cfgsc_cfg_cq_ldb_inflight_limit_mem_we                           = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_INFLIGHT_LIMIT_MEM ] ;
assign cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct                 = cfgsc_cfg_mem_wdata [12:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct_lim_p_nc        = cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct.lim_p ;

// HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_THRESHOLD
assign cfgsc_cfg_cq_ldb_inflight_threshold_mem_we                       = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_INFLIGHT_THRESHOLD_MEM ] ;
assign cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct             = cfgsc_cfg_mem_wdata [12:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct_thr_p_nc    = cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct.thr_p ;

// HQM_LSP_TARGET_CFG_QID_AQED_ACTIVE_LIMIT
assign cfgsc_cfg_qid_aqed_active_limit_mem_we                           = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_QID_AQED_ACTIVE_LIMIT_MEM ] ;
assign cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct                 = cfgsc_cfg_mem_wdata [12:0] ;  // Will get linra warning if size of struct changes
assign cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct_lim_p_nc        = cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct.lim_p ;

// HQM_LSP_TARGET_CFG_QID_NALDB_TOT_ENQ_CNTH , CNTL
assign cfgsc_qid_naldb_tot_enq_cnt_mem_we                       = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_NALDB_TOT_ENQ_CNT_MEM ] ;

// HQM_LSP_TARGET_CFG_QID_ATM_TOT_ENQ_CNTH , CNTL
assign cfgsc_qid_atm_tot_enq_cnt_mem_we                         = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_ATM_TOT_ENQ_CNT_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_LDB_TOT_SCH_CNTH , CNTL
assign cfgsc_cq_ldb_tot_sch_cnt_mem_we                          = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_TOT_SCH_CNT_MEM ] ;

// HQM_LSP_TARGET_CFG_QID_DIR_TOT_ENQ_CNTH , CNTL
assign cfgsc_qid_dir_tot_enq_cnt_mem_we                         = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_DIR_TOT_ENQ_CNT_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_DIR_TOT_SCH_CNTH , CNTL
assign cfgsc_cq_dir_tot_sch_cnt_mem_we                          = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_DIR_TOT_SCH_CNT_MEM ] ;

// HQM_LSP_TARGET_CFG_QID_NALDB_MAX_DEPTH
assign cfgsc_qid_naldb_max_depth_mem_we                         = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_NALDB_MAX_DEPTH_MEM ] ;

// HQM_LSP_TARGET_CFG_QID_DIR_MAX_DEPTH
assign cfgsc_qid_dir_max_depth_mem_we                           = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_DIR_MAX_DEPTH_MEM ] ;

// HQM_LSP_TARGET_CFG_ATM_QID_DPTH_THRSH
assign cfgsc_cfg_atm_qid_dpth_thrsh_mem_we                      = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_ATM_QID_DPTH_THRSH_MEM ] ;

// HQM_LSP_TARGET_CFG_NALB_QID_DPTH_THRSH
assign cfgsc_cfg_nalb_qid_dpth_thrsh_mem_we                     = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_NALB_QID_DPTH_THRSH_MEM ] ;

// HQM_LSP_TARGET_CFG_DIR_QID_DPTH_THRSH
assign cfgsc_cfg_dir_qid_dpth_thrsh_mem_we                      = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_DIR_QID_DPTH_THRSH_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_LDB_WU_COUNT
assign cfgsc_cq_ldb_wu_count_mem_re                             = cfgsc_cfg_mem_re [ CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM ] ;
assign cfgsc_cq_ldb_wu_count_mem_we                             = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM ] ;

// HQM_LSP_TARGET_CFG_CQ_LDB_WU_LIMIT
assign cfgsc_cfg_cq_ldb_wu_limit_mem_re                         = cfgsc_cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM ] ;
assign cfgsc_cfg_cq_ldb_wu_limit_mem_we                         = cfgsc_cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM ] ;

assign cfg_range_reconfig                       = cfg_shdw_ctrl_load ;

// Upstream interface to sidecar has the logical depth and width as seen by config
// Downstream interface to ram_access has divided depth and multiplied width based on the splitting FACTOR
hqm_AW_cfg_sc_memsplit #(
          .FACTOR               ( 1 )                                   // odd and even
        , .CFG_MEM_ADDR_WIDTH   ( HQM_LSP_ARCH_NUM_LB_CQB2 )            // f(full logical depth)
        , .MEM_DWIDTH           ( 33 )                                  // width of data which goes to physical memories; includes cc
        , .MEM_AWIDTH           ( HQM_LSP_ARCH_NUM_LB_PCQB2 )           // width of address which goes to physical memories
) i_hqm_AW_cfg_sc_memsplit_cq2priov (
          .clk                          ( hqm_gated_clk )
        , .rst_n                        ( hqm_gated_rst_n )

        // Upstream interface to sidecar
        , .cfgsc_cfg_mem_re             ( cfgsc_cfg_cq2priov_mem_re )
        , .cfgsc_cfg_mem_we             ( cfgsc_cfg_cq2priov_mem_we )
        , .cfgsc_cfg_mem_addr           ( cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] )
        , .cfgsc_cfg_mem_wdata          ( cfgsc_cfg_cq2priov_mem_wdata )                        // after formatting, cc insertion
        , .cfgsc_cfg_mem_rdata          ( cfgsc_cfg_cq2priov_mem_rdata )                        // before formatting
        , .cfgsc_cfg_mem_ack            ( cfgsc_cfg_cq2priov_mem_ack )

        // Upstream interface to functional access (e.g. AW rmw)
        , .mem_read                     ( cfgsc_func_cfg_cq2priov_mem_re )
        , .mem_write                    ( cfgsc_func_cfg_cq2priov_mem_we )                      // Unused - never functionally written
        , .mem_read_addr                ( '0 )                                                  // Single-port memory
        , .mem_write_addr               ( cfgsc_func_cfg_cq2priov_mem_addr )
        , .mem_read_data                ( cfgsc_func_cfg_cq2priov_mem_rdata )
        , .mem_write_data               ( cfgsc_func_cfg_cq2priov_mem_wdata )                   // Unused - never functionally written

        // Downstream interface to ram_access module functional port
        , .func_mem_re                  ( {   func_cfg_cq2priov_odd_mem_re
                                            , func_cfg_cq2priov_mem_re } )
        , .func_mem_we                  ( {   func_cfg_cq2priov_odd_mem_we
                                            , func_cfg_cq2priov_mem_we } )
        , .func_mem_raddr               ( {   func_cfg_cq2priov_odd_mem_raddr_nc                // Single-port memory
                                            , func_cfg_cq2priov_mem_raddr_nc } )
        , .func_mem_waddr               ( {   func_cfg_cq2priov_odd_mem_addr
                                            , func_cfg_cq2priov_mem_addr } )
        , .func_mem_rdata               ( {   func_cfg_cq2priov_odd_mem_rdata
                                            , func_cfg_cq2priov_mem_rdata } )
        , .func_mem_wdata               ( {   func_cfg_cq2priov_odd_mem_wdata
                                            , func_cfg_cq2priov_mem_wdata } )

        // Downstream interface to ram_access module rf port
        , .rf_mem_re                    ( {   rf_cfg_cq2priov_odd_mem_re
                                            , rf_cfg_cq2priov_mem_re } )
        , .rf_mem_we                    ( {   rf_cfg_cq2priov_odd_mem_we
                                            , rf_cfg_cq2priov_mem_we } )
) ;

hqm_AW_cfg_sc_memsplit #(
          .FACTOR               ( 1 )                                   // odd and even
        , .CFG_MEM_ADDR_WIDTH   ( HQM_LSP_ARCH_NUM_LB_CQB2 )            // f(full logical depth)
        , .MEM_DWIDTH           ( 29 )                                  // width of data which goes to physical memories; includes cc
        , .MEM_AWIDTH           ( HQM_LSP_ARCH_NUM_LB_PCQB2 )           // width of address which goes to physical memories
) i_hqm_AW_cfg_sc_memsplit_cq2qid_0 (
          .clk                          ( hqm_gated_clk )
        , .rst_n                        ( hqm_gated_rst_n )

        // Upstream interface to sidecar
        , .cfgsc_cfg_mem_re             ( cfgsc_cfg_cq2qid_0_mem_re )
        , .cfgsc_cfg_mem_we             ( cfgsc_cfg_cq2qid_0_mem_we )
        , .cfgsc_cfg_mem_addr           ( cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] )
        , .cfgsc_cfg_mem_wdata          ( cfgsc_cfg_cq2qid_0_mem_wdata )                        // after formatting, cc insertion
        , .cfgsc_cfg_mem_rdata          ( cfgsc_cfg_cq2qid_0_mem_rdata )                        // before formatting
        , .cfgsc_cfg_mem_ack            ( cfgsc_cfg_cq2qid_0_mem_ack )

        // Upstream interface to functional access (e.g. AW rmw)
        , .mem_read                     ( cfgsc_func_cfg_cq2qid_0_mem_re )
        , .mem_write                    ( cfgsc_func_cfg_cq2qid_0_mem_we )                      // Unused - never functionally written
        , .mem_read_addr                ( '0 )                                                  // Single-port memory
        , .mem_write_addr               ( cfgsc_func_cfg_cq2qid_0_mem_addr )
        , .mem_read_data                ( cfgsc_func_cfg_cq2qid_0_mem_rdata )
        , .mem_write_data               ( cfgsc_func_cfg_cq2qid_0_mem_wdata )                   // Unused - never functionally written

        // Downstream interface to ram_access module functional port
        , .func_mem_re                  ( {   func_cfg_cq2qid_0_odd_mem_re
                                            , func_cfg_cq2qid_0_mem_re } )
        , .func_mem_we                  ( {   func_cfg_cq2qid_0_odd_mem_we
                                            , func_cfg_cq2qid_0_mem_we } )
        , .func_mem_raddr               ( {   func_cfg_cq2qid_0_odd_mem_raddr_nc                // Single-port memory
                                            , func_cfg_cq2qid_0_mem_raddr_nc } )
        , .func_mem_waddr               ( {   func_cfg_cq2qid_0_odd_mem_addr
                                            , func_cfg_cq2qid_0_mem_addr } )
        , .func_mem_rdata               ( {   func_cfg_cq2qid_0_odd_mem_rdata
                                            , func_cfg_cq2qid_0_mem_rdata } )
        , .func_mem_wdata               ( {   func_cfg_cq2qid_0_odd_mem_wdata
                                            , func_cfg_cq2qid_0_mem_wdata } )

        // Downstream interface to ram_access module rf port
        , .rf_mem_re                    ( {   rf_cfg_cq2qid_0_odd_mem_re
                                            , rf_cfg_cq2qid_0_mem_re } )
        , .rf_mem_we                    ( {   rf_cfg_cq2qid_0_odd_mem_we
                                            , rf_cfg_cq2qid_0_mem_we } )
) ;

hqm_AW_cfg_sc_memsplit #(
          .FACTOR               ( 1 )                                   // odd and even
        , .CFG_MEM_ADDR_WIDTH   ( HQM_LSP_ARCH_NUM_LB_CQB2 )            // f(full logical depth)
        , .MEM_DWIDTH           ( 29 )                                  // width of data which goes to physical memories; includes cc
        , .MEM_AWIDTH           ( HQM_LSP_ARCH_NUM_LB_PCQB2 )           // width of address which goes to physical memories
) i_hqm_AW_cfg_sc_memsplit_cq2qid_1 (
          .clk                          ( hqm_gated_clk )
        , .rst_n                        ( hqm_gated_rst_n )

        // Upstream interface to sidecar
        , .cfgsc_cfg_mem_re             ( cfgsc_cfg_cq2qid_1_mem_re )
        , .cfgsc_cfg_mem_we             ( cfgsc_cfg_cq2qid_1_mem_we )
        , .cfgsc_cfg_mem_addr           ( cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] )
        , .cfgsc_cfg_mem_wdata          ( cfgsc_cfg_cq2qid_1_mem_wdata )                        // after formatting, cc insertion
        , .cfgsc_cfg_mem_rdata          ( cfgsc_cfg_cq2qid_1_mem_rdata )                        // before formatting
        , .cfgsc_cfg_mem_ack            ( cfgsc_cfg_cq2qid_1_mem_ack )

        // Upstream interface to functional access (e.g. AW rmw)
        , .mem_read                     ( cfgsc_func_cfg_cq2qid_1_mem_re )
        , .mem_write                    ( cfgsc_func_cfg_cq2qid_1_mem_we )                      // Unused - never functionally written
        , .mem_read_addr                ( '0 )                                                  // Single-port memory
        , .mem_write_addr               ( cfgsc_func_cfg_cq2qid_1_mem_addr )
        , .mem_read_data                ( cfgsc_func_cfg_cq2qid_1_mem_rdata )
        , .mem_write_data               ( cfgsc_func_cfg_cq2qid_1_mem_wdata )                   // Unused - never functionally written

        // Downstream interface to ram_access module functional port
        , .func_mem_re                  ( {   func_cfg_cq2qid_1_odd_mem_re
                                            , func_cfg_cq2qid_1_mem_re } )
        , .func_mem_we                  ( {   func_cfg_cq2qid_1_odd_mem_we
                                            , func_cfg_cq2qid_1_mem_we } )
        , .func_mem_raddr               ( {   func_cfg_cq2qid_1_odd_mem_raddr_nc                // Single-port memory
                                            , func_cfg_cq2qid_1_mem_raddr_nc } )
        , .func_mem_waddr               ( {   func_cfg_cq2qid_1_odd_mem_addr
                                            , func_cfg_cq2qid_1_mem_addr } )
        , .func_mem_rdata               ( {   func_cfg_cq2qid_1_odd_mem_rdata
                                            , func_cfg_cq2qid_1_mem_rdata } )
        , .func_mem_wdata               ( {   func_cfg_cq2qid_1_odd_mem_wdata
                                            , func_cfg_cq2qid_1_mem_wdata } )

        // Downstream interface to ram_access module rf port
        , .rf_mem_re                    ( {   rf_cfg_cq2qid_1_odd_mem_re
                                            , rf_cfg_cq2qid_1_mem_re } )
        , .rf_mem_we                    ( {   rf_cfg_cq2qid_1_odd_mem_we
                                            , rf_cfg_cq2qid_1_mem_we } )
) ;

always_comb begin
  cfg_mem_wdata                                 = cfgsc_cfg_mem_wdata ;
  cfg_mem_we                                    = cfgsc_cfg_mem_we ;
  cfg_mem_re                                    = cfgsc_cfg_mem_re ;
  cfgsc_cfg_mem_rdata                           = cfg_mem_rdata ;
  cfgsc_cfg_mem_ack                             = cfg_mem_ack ;

  cfgsc_wide_memory_wait_for_write_nxt          = cfgsc_wide_memory_wait_for_write_f ;

  // 1-clock pulse
  cfg_mem_ack_qid_naldb_tot_enq_cnt_nxt         = 1'b0 ;
  cfg_mem_ack_qid_atm_tot_enq_cnt_nxt           = 1'b0 ;
  cfg_mem_ack_cq_ldb_tot_sch_cnt_nxt            = 1'b0 ;
  cfg_mem_ack_qid_dir_tot_enq_cnt_nxt           = 1'b0 ;
  cfg_mem_ack_cq_dir_tot_sch_cnt_nxt            = 1'b0 ;

  cfg_mem_cc_v                                  = 1'b0 ;
  cfg_mem_cc_value                              = 8'h0 ;
  cfg_mem_cc_width                              = 4'h1 ;
  cfg_mem_cc_position                           = 12'd0 ;

  func_qid_naldb_tot_enq_cnt_mem_we             = cfgsc_func_qid_naldb_tot_enq_cnt_mem_we ;
  func_qid_naldb_tot_enq_cnt_mem_waddr          = cfgsc_func_qid_naldb_tot_enq_cnt_mem_waddr ;
  func_qid_naldb_tot_enq_cnt_mem_wdata          = cfgsc_func_qid_naldb_tot_enq_cnt_mem_wdata ;

  func_qid_atm_tot_enq_cnt_mem_we               = cfgsc_func_qid_atm_tot_enq_cnt_mem_we ;
  func_qid_atm_tot_enq_cnt_mem_waddr            = cfgsc_func_qid_atm_tot_enq_cnt_mem_waddr ;
  func_qid_atm_tot_enq_cnt_mem_wdata            = cfgsc_func_qid_atm_tot_enq_cnt_mem_wdata ;

  func_cq_ldb_tot_sch_cnt_mem_we                = cfgsc_func_cq_ldb_tot_sch_cnt_mem_we ;
  func_cq_ldb_tot_sch_cnt_mem_waddr             = cfgsc_func_cq_ldb_tot_sch_cnt_mem_waddr ;
  func_cq_ldb_tot_sch_cnt_mem_wdata             = cfgsc_func_cq_ldb_tot_sch_cnt_mem_wdata ;

  func_qid_dir_tot_enq_cnt_mem_we               = cfgsc_func_qid_dir_tot_enq_cnt_mem_we ;
  func_qid_dir_tot_enq_cnt_mem_waddr            = cfgsc_func_qid_dir_tot_enq_cnt_mem_waddr ;
  func_qid_dir_tot_enq_cnt_mem_wdata            = cfgsc_func_qid_dir_tot_enq_cnt_mem_wdata ;

  func_cq_dir_tot_sch_cnt_mem_we                = cfgsc_func_cq_dir_tot_sch_cnt_mem_we ;
  func_cq_dir_tot_sch_cnt_mem_waddr             = cfgsc_func_cq_dir_tot_sch_cnt_mem_waddr ;
  func_cq_dir_tot_sch_cnt_mem_wdata             = cfgsc_func_cq_dir_tot_sch_cnt_mem_wdata ;

  // HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_COUNT
  if ( cfgsc_dir_tok_cnt_mem_we ) begin
    cfg_mem_wdata                                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0]            = cfgsc_dir_tok_cnt_mem_wdata_struct.cnt ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 6'h0 , cfgsc_cfg_mem_wdata_res } ;
    cfg_mem_cc_width                            = 4'h2 ;
    cfg_mem_cc_position                         = HQM_LSP_DIRENQ_TOK_CNT_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_CQ_DIR_TOKEN_DEPTH_SELECT_DSI
  if ( cfgsc_dir_tok_lim_mem_we ) begin
    cfg_mem_wdata                               = {   27'h0             // Don't include spare in parity
                                                    , cfgsc_dir_tok_lim_mem_wdata_struct.disab_opt
                                                    , cfgsc_dir_tok_lim_mem_wdata_struct.lim_sel } ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = 12'd7 ;
  end

  // HQM_LSP_TARGET_CFG_CQ2PRIOV - config write to odd/even memories handled by sc_memsplit

  // HQM_LSP_TARGET_CFG_CQ2QID0 - config write to odd/even memories handled by sc_memsplit, need data formatting for sc and parity gen
  if ( cfgsc_cfg_cq2qid_0_mem_we ) begin
    cfg_mem_wdata                               = {       4'h0                          // RDL has qid fields as 8 bits wide
                                                        , cfgsc_cfg_mem_wdata  [ 24 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [ 16 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [  8 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [  0 +: 7 ] } ;
  end

  // HQM_LSP_TARGET_CFG_CQ2QID1 - config write to odd/even memories handled by sc_memsplit, need data formatting for sc and parity gen
  if ( cfgsc_cfg_cq2qid_1_mem_we ) begin
    cfg_mem_wdata                               = {       4'h0                          // RDL has qid fields as 8 bits wide
                                                        , cfgsc_cfg_mem_wdata  [ 24 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [ 16 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [  8 +: 7 ]
                                                        , cfgsc_cfg_mem_wdata  [  0 +: 7 ] } ;
  end

  // HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_COUNT
  if ( cfgsc_qid_ldb_inflight_count_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_QID_IF_CNT_WIDTH-1:0]     = cfgsc_qid_ldb_inflight_count_mem_wdata_struct.cnt ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 6'h0 , cfgsc_cfg_mem_wdata_res } ;
    cfg_mem_cc_width                            = 4'h2 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_QID_IF_CNT_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_QID_LDB_INFLIGHT_LIMIT
  if ( cfgsc_cfg_qid_ldb_inflight_limit_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_QID_IF_LIM_WIDTH-1:0]     = cfgsc_cfg_qid_ldb_inflight_limit_mem_wdata_struct.lim ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_QID_IF_LIM_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_0 .. _15
  if ( cfgsc_cfg_qid_ldb_qid2cqidix_mem_we ) begin
    cfg_mem_wdata                               = cfgsc_cfg_mem_wdata ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = 12'd512 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_00 ] ) cfg_mem_cc_position   = 12'd512 + 12'd0 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_01 ] ) cfg_mem_cc_position   = 12'd512 + 12'd1 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_02 ] ) cfg_mem_cc_position   = 12'd512 + 12'd2 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_03 ] ) cfg_mem_cc_position   = 12'd512 + 12'd3 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_04 ] ) cfg_mem_cc_position   = 12'd512 + 12'd4 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_05 ] ) cfg_mem_cc_position   = 12'd512 + 12'd5 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_06 ] ) cfg_mem_cc_position   = 12'd512 + 12'd6 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_07 ] ) cfg_mem_cc_position   = 12'd512 + 12'd7 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_08 ] ) cfg_mem_cc_position   = 12'd512 + 12'd8 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_09 ] ) cfg_mem_cc_position   = 12'd512 + 12'd9 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_10 ] ) cfg_mem_cc_position   = 12'd512 + 12'd10 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_11 ] ) cfg_mem_cc_position   = 12'd512 + 12'd11 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_12 ] ) cfg_mem_cc_position   = 12'd512 + 12'd12 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_13 ] ) cfg_mem_cc_position   = 12'd512 + 12'd13 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_14 ] ) cfg_mem_cc_position   = 12'd512 + 12'd14 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX_15 ] ) cfg_mem_cc_position   = 12'd512 + 12'd15 ;
  end

  // HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_0 .. _15
  if ( cfgsc_cfg_qid_ldb_qid2cqidix2_mem_we ) begin
    cfg_mem_wdata                               = cfgsc_cfg_mem_wdata ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = 12'd512 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_00 ] ) cfg_mem_cc_position  = 12'd512 + 12'd0 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_01 ] ) cfg_mem_cc_position  = 12'd512 + 12'd1 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_02 ] ) cfg_mem_cc_position  = 12'd512 + 12'd2 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_03 ] ) cfg_mem_cc_position  = 12'd512 + 12'd3 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_04 ] ) cfg_mem_cc_position  = 12'd512 + 12'd4 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_05 ] ) cfg_mem_cc_position  = 12'd512 + 12'd5 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_06 ] ) cfg_mem_cc_position  = 12'd512 + 12'd6 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_07 ] ) cfg_mem_cc_position  = 12'd512 + 12'd7 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_08 ] ) cfg_mem_cc_position  = 12'd512 + 12'd8 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_09 ] ) cfg_mem_cc_position  = 12'd512 + 12'd9 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_10 ] ) cfg_mem_cc_position  = 12'd512 + 12'd10 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_11 ] ) cfg_mem_cc_position  = 12'd512 + 12'd11 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_12 ] ) cfg_mem_cc_position  = 12'd512 + 12'd12 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_13 ] ) cfg_mem_cc_position  = 12'd512 + 12'd13 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_14 ] ) cfg_mem_cc_position  = 12'd512 + 12'd14 ;
    if ( cfg_req_write_pnc [ HQM_LSP_TARGET_CFG_QID_LDB_QID2CQIDIX2_15 ] ) cfg_mem_cc_position  = 12'd512 + 12'd15 ;
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_COUNT
  if ( cfgsc_cq_ldb_token_count_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ; 
    cfg_mem_wdata [HQM_LSP_LB_CQ_TOK_CNT_WIDTH-1:0]     = cfgsc_cfg_mem_wdata [HQM_LSP_LB_CQ_TOK_CNT_WIDTH-1:0] ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 6'h0 , cfgsc_cfg_mem_wdata_res } ;
    cfg_mem_cc_width                            = 4'h2 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_CQ_TOK_CNT_WIDTH[11:0] ;
  end


  // HQM_LSP_TARGET_CFG_CQ_LDB_TOKEN_DEPTH_SELECT
  if ( cfgsc_cfg_cq_ldb_token_depth_select_mem_we ) begin
    cfg_mem_wdata                               = { 28'h0, cfgsc_cfg_cq_ldb_token_depth_select_mem_wdata_struct.lim_sel } ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = 12'd4 ;
  end

  // HQM_LSP_TARGET_CQ_LDB_INFLIGHT_COUNT
  if ( cfgsc_cq_ldb_inflight_count_mem_we ) begin
    cfg_mem_wdata                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]      = cfgsc_cq_ldb_inflight_count_mem_wdata_struct.cnt ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 6'h0 , cfgsc_cfg_mem_wdata_res } ;
    cfg_mem_cc_width                            = 4'h2 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_CQ_IF_CNT_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_LIMIT
  if ( cfgsc_cfg_cq_ldb_inflight_limit_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_CQ_IF_LIM_WIDTH-1:0]      = { 20'h0, cfgsc_cfg_cq_ldb_inflight_limit_mem_wdata_struct.lim } ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_CQ_IF_LIM_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_INFLIGHT_THRESHOLD
  if ( cfgsc_cfg_cq_ldb_inflight_threshold_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_CQ_IF_THR_WIDTH-1:0]      = { 20'h0, cfgsc_cfg_cq_ldb_inflight_threshold_mem_wdata_struct.thr } ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_CQ_IF_THR_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_QID_AQED_ACTIVE_LIMIT
  if ( cfgsc_cfg_qid_aqed_active_limit_mem_we ) begin
    cfg_mem_wdata                                       = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH-1:0]  = cfgsc_cfg_qid_aqed_active_limit_mem_wdata_struct.lim ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH[11:0] ;
  end

  //*************************************************************************************************************************
  //**** For wide memories (> 32 bits, multiple targets) which require an atomic write capability for the multiple       ****
  //**** targets, intercept the config write (CNTL or CNTH) and transform it into a 66-bit write on the func interface.  ****
  //**** Disable the config write to ram_access, manufacture an ack back to the sc when the actual write has occurred.   ****
  //****   - The sc expects the ack to happen at least 1 clock after it issues the config write                          ****
  //****   - Currently the ram_access module issues the functional write on the same clock that it was requested         ****
  //****   - Therefore, detect when a config write has been requested by the sidecar, and set a target-specific flop     ****
  //****     to generate a 1-clock ack when the write is actually requested by ram_access, which may occur 0..n clocks   ****
  //****     later (current ram_access requests 0 clocks later).                                                         ****

  // HQM_LSP_TARGET_CFG_QID_NALDB_TOT_ENQ_CNTH , CNTL
  if ( cfgsc_qid_naldb_tot_enq_cnt_mem_we ) begin               // Config write of any value writes a 0, use func intf to get all 66 bits
    func_qid_naldb_tot_enq_cnt_mem_we           = 1'b1 ;
    func_qid_naldb_tot_enq_cnt_mem_waddr        = cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    func_qid_naldb_tot_enq_cnt_mem_wdata        = 66'h0 ;

    cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_NALDB_TOT_ENQ_CNT_MEM ] = 1'b0 ;
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b1 ;        // Tentatively set, but override (clear) below if actual mem we is signalled this clock
  end

  // HQM_LSP_TARGET_CFG_QID_ATM_TOT_ENQ_CNTH , CNTL
  if ( cfgsc_qid_atm_tot_enq_cnt_mem_we ) begin               // Config write of any value writes a 0, use func intf to get all 66 bits
    func_qid_atm_tot_enq_cnt_mem_we             = 1'b1 ;
    func_qid_atm_tot_enq_cnt_mem_waddr          = cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    func_qid_atm_tot_enq_cnt_mem_wdata          = 66'h0 ;

    cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_ATM_TOT_ENQ_CNT_MEM ] = 1'b0 ;
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b1 ;        // Tentatively set, but override (clear) below if actual mem we is signalled this clock
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_TOT_SCH_CNTH , CNTL
  if ( cfgsc_cq_ldb_tot_sch_cnt_mem_we ) begin               // Config write of any value writes a 0, use func intf to get all 66 bits
    func_cq_ldb_tot_sch_cnt_mem_we              = 1'b1 ;
    func_cq_ldb_tot_sch_cnt_mem_waddr           = cfg_mem_addr [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
    func_cq_ldb_tot_sch_cnt_mem_wdata           = 66'h0 ;

    cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_TOT_SCH_CNT_MEM ] = 1'b0 ;
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b1 ;        // Tentatively set, but override (clear) below if actual mem we is signalled this clock
  end

  // HQM_LSP_TARGET_CFG_QID_DIR_TOT_ENQ_CNTH , CNTL
  if ( cfgsc_qid_dir_tot_enq_cnt_mem_we ) begin               // Config write of any value writes a 0, use func intf to get all 66 bits
    func_qid_dir_tot_enq_cnt_mem_we             = 1'b1 ;
    func_qid_dir_tot_enq_cnt_mem_waddr          = cfg_mem_addr [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
    func_qid_dir_tot_enq_cnt_mem_wdata          = 66'h0 ;

    cfg_mem_we [ CFG_ACCESSIBLE_RAM_QID_DIR_TOT_ENQ_CNT_MEM ] = 1'b0 ;
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b1 ;        // Tentatively set, but override (clear) below if actual mem we is signalled this clock
  end

  // HQM_LSP_TARGET_CFG_CQ_DIR_TOT_SCH_CNTH , CNTL
  if ( cfgsc_cq_dir_tot_sch_cnt_mem_we ) begin               // Config write of any value writes a 0, use func intf to get all 66 bits
    func_cq_dir_tot_sch_cnt_mem_we              = 1'b1 ;
    func_cq_dir_tot_sch_cnt_mem_waddr           = cfg_mem_addr [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0] ;
    func_cq_dir_tot_sch_cnt_mem_wdata           = 66'h0 ;

    cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_DIR_TOT_SCH_CNT_MEM ] = 1'b0 ;
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b1 ;        // Tentatively set, but override (clear) below if actual mem we is signalled this clock
  end

  // Signal ack on next clock
  if ( rf_qid_naldb_tot_enq_cnt_mem_we ) begin
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b0 ;
    cfg_mem_ack_qid_naldb_tot_enq_cnt_nxt       = cfgsc_wide_memory_wait_for_write_f | cfgsc_qid_naldb_tot_enq_cnt_mem_we ;
  end
  if ( rf_qid_atm_tot_enq_cnt_mem_we ) begin
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b0 ;
    cfg_mem_ack_qid_atm_tot_enq_cnt_nxt         = cfgsc_wide_memory_wait_for_write_f | cfgsc_qid_atm_tot_enq_cnt_mem_we ;
  end
  if ( rf_cq_ldb_tot_sch_cnt_mem_we ) begin
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b0 ;
    cfg_mem_ack_cq_ldb_tot_sch_cnt_nxt          = cfgsc_wide_memory_wait_for_write_f | cfgsc_cq_ldb_tot_sch_cnt_mem_we ;
  end
  if ( rf_qid_dir_tot_enq_cnt_mem_we ) begin
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b0 ;
    cfg_mem_ack_qid_dir_tot_enq_cnt_nxt         = cfgsc_wide_memory_wait_for_write_f | cfgsc_qid_dir_tot_enq_cnt_mem_we ;
  end
  if ( rf_cq_dir_tot_sch_cnt_mem_we ) begin
    cfgsc_wide_memory_wait_for_write_nxt        = 1'b0 ;
    cfg_mem_ack_cq_dir_tot_sch_cnt_nxt          = cfgsc_wide_memory_wait_for_write_f | cfgsc_cq_dir_tot_sch_cnt_mem_we ;
  end

  // Read responses occur conventionally, write responses are generated with glue logic, both must work and are independent
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_NALDB_TOT_ENQ_CNT_MEM ]    = cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_NALDB_TOT_ENQ_CNT_MEM ] | cfg_mem_ack_qid_naldb_tot_enq_cnt_f ;
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_ATM_TOT_ENQ_CNT_MEM ]      = cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_ATM_TOT_ENQ_CNT_MEM ]   | cfg_mem_ack_qid_atm_tot_enq_cnt_f ;
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CQ_LDB_TOT_SCH_CNT_MEM ]       = cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CQ_LDB_TOT_SCH_CNT_MEM ]    | cfg_mem_ack_cq_ldb_tot_sch_cnt_f ;
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_DIR_TOT_ENQ_CNT_MEM ]      = cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_QID_DIR_TOT_ENQ_CNT_MEM ]   | cfg_mem_ack_qid_dir_tot_enq_cnt_f ;
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CQ_DIR_TOT_SCH_CNT_MEM ]       = cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CQ_DIR_TOT_SCH_CNT_MEM ]    | cfg_mem_ack_cq_dir_tot_sch_cnt_f ;
  //****                                                                                                                 ****
  //*************************************************************************************************************************

  // HQM_LSP_TARGET_CFG_QID_NALDB_MAX_DEPTH
  if ( cfgsc_qid_naldb_max_depth_mem_we ) begin
    cfg_mem_wdata                               = 32'h0 ;       // 0 with 0 residue, no need to generate/insert
  end

  // HQM_LSP_TARGET_CFG_QID_DIR_MAX_DEPTH
  if ( cfgsc_qid_dir_max_depth_mem_we ) begin
    cfg_mem_wdata                               = 32'h0 ;       // 0 with 0 residue, no need to generate/insert
  end

  // HQM_LSP_TARGET_CFG_ATM_QID_DPTH_THRSH
  if ( cfgsc_cfg_atm_qid_dpth_thrsh_mem_we ) begin
    cfg_mem_wdata                                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH-1:0]        = cfgsc_cfg_mem_wdata [HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH-1:0] ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_NALB_QID_DPTH_THRSH
  if ( cfgsc_cfg_nalb_qid_dpth_thrsh_mem_we ) begin
    cfg_mem_wdata                                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LB_QID_DPTH_THRSH_WIDTH-1:0]         = cfgsc_cfg_mem_wdata [HQM_LSP_LB_QID_DPTH_THRSH_WIDTH-1:0] ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_LB_QID_DPTH_THRSH_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_DIR_QID_DPTH_THRSH
  if ( cfgsc_cfg_dir_qid_dpth_thrsh_mem_we ) begin
    cfg_mem_wdata                                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH-1:0]         = cfgsc_cfg_mem_wdata [HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH-1:0] ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_WU_COUNT
  if ( cfgsc_cq_ldb_wu_count_mem_we ) begin
    cfg_mem_wdata                               = 32'h0 ;
    cfg_mem_wdata [HQM_LSP_LBWU_CQ_WU_CNT_WIDTH-1:0]            = cfgsc_cfg_mem_wdata [HQM_LSP_LBWU_CQ_WU_CNT_WIDTH-1:0] ;
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 6'h0 , cfgsc_cfg_mem_wdata_res } ;
    cfg_mem_cc_width                            = 4'h2 ;
    cfg_mem_cc_position                         = HQM_LSP_LBWU_CQ_WU_CNT_WIDTH[11:0] ;
  end

  // HQM_LSP_TARGET_CFG_CQ_LDB_WU_LIMIT
  if ( cfgsc_cfg_cq_ldb_wu_limit_mem_we ) begin
    cfg_mem_wdata                               = 32'h0 ;
    cfg_mem_wdata [1+(HQM_LSP_LBWU_CQ_WU_LIM_WIDTH-1):0]        = cfgsc_cfg_mem_wdata [1+(HQM_LSP_LBWU_CQ_WU_LIM_WIDTH-1):0] ;  // lim_v, lim
    cfg_mem_cc_v                                = 1'b1 ;
    cfg_mem_cc_value                            = { 7'h0 , cfgsc_cfg_mem_wdata_par } ;
    cfg_mem_cc_width                            = 4'h1 ;
    cfg_mem_cc_position                         = (HQM_LSP_LBWU_CQ_WU_LIM_WIDTH[11:0] + 12'h1);
  end

  //*************************************************************************************************************************
  //****                                                                                                                 ****
  // Config access to split memories is provided by sc_memsplit
  cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM ]            = 1'b0 ;
  cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM ]            = 1'b0 ;
  cfgsc_cfg_mem_rdata [ ( CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM * 32 ) +: 32 ]    = cfgsc_cfg_cq2priov_mem_rdata [31:0] ;         // strip off parity bit
  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CFG_CQ2PRIOV_MEM ]     = cfgsc_cfg_cq2priov_mem_ack ;

  cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM ]            = 1'b0 ;
  cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM ]            = 1'b0 ;
  cfgsc_cfg_mem_rdata [ ( CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM * 32 ) +: 32 ]    = {   1'b0                                      // strip off parity bit, format
                                                                                    , cfgsc_cfg_cq2qid_0_mem_rdata [27:21]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_0_mem_rdata [20:14]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_0_mem_rdata [13:7]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_0_mem_rdata [6:0] } ;

  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_0_MEM ]     = cfgsc_cfg_cq2qid_0_mem_ack ;

  cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM ]            = 1'b0 ;
  cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM ]            = 1'b0 ;
  cfgsc_cfg_mem_rdata [ ( CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM * 32 ) +: 32 ]    = {   1'b0                                      // strip off parity bit, format
                                                                                    , cfgsc_cfg_cq2qid_1_mem_rdata [27:21]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_1_mem_rdata [20:14]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_1_mem_rdata [13:7]
                                                                                    , 1'b0
                                                                                    , cfgsc_cfg_cq2qid_1_mem_rdata [6:0] } ;

  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CFG_CQ2QID_1_MEM ]     = cfgsc_cfg_cq2qid_1_mem_ack ;

  //****                                                                                                                 ****
  //*************************************************************************************************************************

  //*************************************************************************************************************************
  //****                                                                                                                 ****
  // Config access to wu_count and wu_limit is done through the functional pipe
  cfg_mem_we [ CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM ]         = 1'b0 ;
  cfg_mem_re [ CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM ]         = 1'b0 ;
  cfg_mem_we [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM ]     = 1'b0 ;
  cfg_mem_re [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM ]     = 1'b0 ;

  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM ]                          = cfgsc_wu_count_wr_ack | cfgsc_wu_count_rd_ack ;
  if ( cfgsc_wu_count_rd_ack ) begin
    cfgsc_cfg_mem_rdata [ ( CFG_ACCESSIBLE_RAM_CQ_LDB_WU_COUNT_MEM * 32 ) +: 32 ]       = cfgsc_wu_cfg_data_f ;
  end

  cfgsc_cfg_mem_ack [ CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM ]                      = cfgsc_wu_limit_wr_ack | cfgsc_wu_limit_rd_ack ;
  if ( cfgsc_wu_limit_rd_ack ) begin
    cfgsc_cfg_mem_rdata [ ( CFG_ACCESSIBLE_RAM_CFG_CQ_LDB_WU_LIMIT_MEM * 32 ) +: 32 ]   = cfgsc_wu_cfg_data_f ;
  end
  //****                                                                                                                 ****
  //*************************************************************************************************************************
end // always

assign cfgsc_cfg_cq2priov_mem_rdata_nc          = cfgsc_cfg_cq2priov_mem_rdata [32] ;                   // parity bit not used on cfg read
assign cfgsc_cfg_cq2qid_0_mem_rdata_nc          = cfgsc_cfg_cq2qid_0_mem_rdata [28] ;                   // parity bit not used on cfg read
assign cfgsc_cfg_cq2qid_1_mem_rdata_nc          = cfgsc_cfg_cq2qid_1_mem_rdata [28] ;                   // parity bit not used on cfg read

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfgsc_wide_memory_wait_for_write_f                  <= 1'b0 ;
    cfg_mem_ack_qid_naldb_tot_enq_cnt_f                 <= 1'b0 ;
    cfg_mem_ack_qid_atm_tot_enq_cnt_f                   <= 1'b0 ;
    cfg_mem_ack_cq_ldb_tot_sch_cnt_f                    <= 1'b0 ;
    cfg_mem_ack_qid_dir_tot_enq_cnt_f                   <= 1'b0 ;
    cfg_mem_ack_cq_dir_tot_sch_cnt_f                    <= 1'b0 ;
  end
  else begin
    cfgsc_wide_memory_wait_for_write_f                  <= cfgsc_wide_memory_wait_for_write_nxt ;
    cfg_mem_ack_qid_naldb_tot_enq_cnt_f                 <= cfg_mem_ack_qid_naldb_tot_enq_cnt_nxt ;
    cfg_mem_ack_qid_atm_tot_enq_cnt_f                   <= cfg_mem_ack_qid_atm_tot_enq_cnt_nxt ;
    cfg_mem_ack_cq_ldb_tot_sch_cnt_f                    <= cfg_mem_ack_cq_ldb_tot_sch_cnt_nxt ;
    cfg_mem_ack_qid_dir_tot_enq_cnt_f                   <= cfg_mem_ack_qid_dir_tot_enq_cnt_nxt ;
    cfg_mem_ack_cq_dir_tot_sch_cnt_f                    <= cfg_mem_ack_cq_dir_tot_sch_cnt_nxt ;
  end
end // always

//----
assign pfcsr_shadow_nxt         = {   cfg_dir_tok_lim_disab_opt_nxt    } ;      // Copy of cfg RAM, reset value must match pf reset value

assign {   cfg_dir_tok_lim_disab_opt_f }        = pfcsr_shadow_f ;

//----
assign mem_access_error_nxt     = (   rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_error
                                    | rf_qid_dir_max_depth_mem_error
                                    | rf_cfg_dir_qid_dpth_thrsh_mem_error
                                    | rf_qid_ldb_replay_count_mem_error
                                    | rf_cfg_atm_qid_dpth_thrsh_mem_error
                                    | rf_send_atm_to_cq_rx_sync_fifo_mem_error
                                    | rf_cfg_qid_ldb_inflight_limit_mem_error
                                    | rf_qid_ldb_enqueue_count_mem_error
                                    | rf_qid_dir_tot_enq_cnt_mem_error
                                    | rf_qid_naldb_tot_enq_cnt_mem_error
                                    | rf_atm_cmp_fifo_mem_error
                                    | rf_cfg_qid_ldb_qid2cqidix_mem_error
                                    | rf_qid_atm_tot_enq_cnt_mem_error
                                    | rf_cfg_qid_aqed_active_limit_mem_error
                                    | rf_cq_ldb_tot_sch_cnt_mem_error
                                    | rf_qid_naldb_max_depth_mem_error
                                    | rf_rop_lsp_reordercmp_rx_sync_fifo_mem_error
                                    | rf_dir_enq_cnt_mem_error
                                    | rf_qid_aqed_active_count_mem_error
                                    | rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_error
                                    | rf_qid_ldb_inflight_count_mem_error
                                    | rf_cfg_cq2qid_1_odd_mem_error
                                    | rf_cfg_cq2qid_1_mem_error
                                    | rf_qid_dir_replay_count_mem_error
                                    | rf_dir_tok_cnt_mem_error
                                    | rf_uno_atm_cmp_fifo_mem_error
                                    | rf_nalb_sel_nalb_fifo_mem_error
                                    | rf_chp_lsp_token_rx_sync_fifo_mem_error
                                    | rf_chp_lsp_cmp_rx_sync_fifo_mem_error
                                    | rf_qed_lsp_deq_fifo_mem_error
                                    | rf_aqed_lsp_deq_fifo_mem_error
                                    | rf_cq_dir_tot_sch_cnt_mem_error
                                    | rf_qid_atm_active_mem_error
                                    | rf_cfg_qid_ldb_qid2cqidix2_mem_error
                                    | rf_cq_ldb_token_count_mem_error
                                    | rf_dp_lsp_enq_dir_rx_sync_fifo_mem_error
                                    | rf_ldb_token_rtn_fifo_mem_error
                                    | rf_cfg_nalb_qid_dpth_thrsh_mem_error
                                    | rf_cfg_cq2priov_odd_mem_error
                                    | rf_cfg_cq2priov_mem_error
                                    | rf_cfg_cq2qid_0_odd_mem_error
                                    | rf_cfg_cq2qid_0_mem_error
                                    | rf_cfg_cq_ldb_token_depth_select_mem_error
                                    | rf_enq_nalb_fifo_mem_error
                                    | rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_error
                                    | rf_cq_nalb_pri_arbindex_mem_error
                                    | rf_cq_atm_pri_arbindex_mem_error
                                    | rf_nalb_cmp_fifo_mem_error
                                    | rf_dir_tok_lim_mem_error
                                    | rf_cq_ldb_inflight_count_mem_error
                                    | rf_qid_atq_enqueue_count_mem_error
                                    | rf_cfg_cq_ldb_inflight_threshold_mem_error
                                    | rf_cfg_cq_ldb_inflight_limit_mem_error
                                    | rf_cq_ldb_wu_count_mem_error
                                    | rf_cfg_cq_ldb_wu_limit_mem_error
                                  ) ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: END common core interfaces 
//*****************************************************************************************************
//*****************************************************************************************************















always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    reset_pf_counter_f <= '0 ;
    reset_pf_active_f <= 1'b1 ;
    reset_pf_done_f <= '0 ;
    hw_init_done_f <= '0 ;
  end
  else begin
    reset_pf_counter_f <= reset_pf_counter_nxt ;
    reset_pf_active_f <= reset_pf_active_nxt ;
    reset_pf_done_f <= reset_pf_done_nxt ;
    hw_init_done_f <= hw_init_done_nxt ;
  end
end


//-------------------------------------------------------------------------------------------
// Int Serializer

assign lba_cq2qid_rw_pipe_err_nxt               = lba_cq2qid_rw_pipe_status ;
assign lba_cq_tok_cnt_rmw_pipe_err_nxt          = lba_cq_tok_cnt_rmw_pipe_status ;
assign lba_qid2cqidix_rw_pipe_err_nxt           = lba_qid2cqidix_rw_pipe_status ;
assign atq_enq_cnt_rmw_pipe_err_nxt             = atq_enq_cnt_rmw_pipe_status ;
assign direnq_enq_cnt_rmw_pipe_err_nxt          = direnq_enq_cnt_rmw_pipe_status ;
assign lbrpl_enq_cnt_rmw_pipe_err_nxt           = lbrpl_enq_cnt_rmw_pipe_status ;
assign dirrpl_enq_cnt_rmw_pipe_err_nxt          = dirrpl_enq_cnt_rmw_pipe_status ;
assign lba_arbindex_rmw_pipe_err_nxt            = lba_nalb_pri_arbindex_pipe_status | lba_atm_pri_arbindex_pipe_status ;
assign lbwu_cq_wu_cnt_rmw_pipe_err_nxt          = lbwu_cq_wu_cnt_rmw_pipe_status ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    lba_cq2qid_rw_pipe_err_f            <= 1'b0 ;
    lba_cq_tok_cnt_rmw_pipe_err_f       <= 1'b0 ;
    lba_qid2cqidix_rw_pipe_err_f        <= 1'b0 ;
    atq_enq_cnt_rmw_pipe_err_f          <= 1'b0 ;
    direnq_enq_cnt_rmw_pipe_err_f       <= 1'b0 ;
    lbrpl_enq_cnt_rmw_pipe_err_f        <= 1'b0 ;
    dirrpl_enq_cnt_rmw_pipe_err_f       <= 1'b0 ;
    lba_arbindex_rmw_pipe_err_f         <= 1'b0 ;
    lbwu_cq_wu_cnt_rmw_pipe_err_f       <= 1'b0 ;
  end
  else begin
    lba_cq2qid_rw_pipe_err_f            <= lba_cq2qid_rw_pipe_err_nxt ;
    lba_cq_tok_cnt_rmw_pipe_err_f       <= lba_cq_tok_cnt_rmw_pipe_err_nxt ;
    lba_qid2cqidix_rw_pipe_err_f        <= lba_qid2cqidix_rw_pipe_err_nxt ;
    atq_enq_cnt_rmw_pipe_err_f          <= atq_enq_cnt_rmw_pipe_err_nxt ;
    direnq_enq_cnt_rmw_pipe_err_f       <= direnq_enq_cnt_rmw_pipe_err_nxt ;
    lbrpl_enq_cnt_rmw_pipe_err_f        <= lbrpl_enq_cnt_rmw_pipe_err_nxt ;
    dirrpl_enq_cnt_rmw_pipe_err_f       <= dirrpl_enq_cnt_rmw_pipe_err_nxt ;
    lba_arbindex_rmw_pipe_err_f         <= lba_arbindex_rmw_pipe_err_nxt ;
    lbwu_cq_wu_cnt_rmw_pipe_err_f       <= lbwu_cq_wu_cnt_rmw_pipe_err_nxt ;
  end
end // always


assign atq_fid_if_lim_err_nxt           = p3_atq_qid_v_any & p3_atq_fid_inflight_cnt_gt_lim ;
assign atq_fid_if_lim_err_reported_nxt  = ( atq_fid_if_lim_err_f | atq_fid_if_lim_err_reported_f ) ;    // BCAM corrupted, reset required
assign atq_fid_if_lim_err_v             = atq_fid_if_lim_err_f & ~ atq_fid_if_lim_err_reported_f ;

assign atq_tot_act_lim_err_nxt          = p3_atq_qid_v_any & p3_atq_tot_act_cnt_gt_lim ;
assign atq_tot_act_lim_err_reported_nxt = ( atq_tot_act_lim_err_f | atq_tot_act_lim_err_reported_f ) ;  // LSP hardware failure, reset required
assign atq_tot_act_lim_err_v            = atq_tot_act_lim_err_f & ~ atq_tot_act_lim_err_reported_f ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    atq_fid_if_lim_err_f                <= 1'b0 ;
    atq_fid_if_lim_err_reported_f       <= 1'b0 ;
    atq_tot_act_lim_err_f               <= 1'b0 ;
    atq_tot_act_lim_err_reported_f      <= 1'b0 ;
    mem_access_error_f                  <= 1'b0 ;
  end
  else begin
    atq_fid_if_lim_err_f                <= atq_fid_if_lim_err_nxt ;
    atq_fid_if_lim_err_reported_f       <= atq_fid_if_lim_err_reported_nxt ;
    atq_tot_act_lim_err_f               <= atq_tot_act_lim_err_nxt ;
    atq_tot_act_lim_err_reported_f      <= atq_tot_act_lim_err_reported_nxt ;
    mem_access_error_f                  <= mem_access_error_nxt ;
  end
end // always

always_comb begin
  err_hw_class_01               = '0 ;
  err_hw_class_01 [ 30:28 ]     = 3'h1 ;                                // Class
  err_hw_class_01 [ 27 ]        = 1'b0 ;                                // Spare
  err_hw_class_01 [ 26 ]        = p3_lbrpl_enq_cnt_oflow_err_f ;
  err_hw_class_01 [ 25 ]        = p3_lbrpl_enq_cnt_uflow_err_f ;
  err_hw_class_01 [ 24 ]        = p3_lbrpl_enq_cnt_res_err ;            // Not flopped, but reasonably fast signal
  err_hw_class_01 [ 23 ]        = p1_lbrpl_inp_frag_cnt_res_err_f ;
  err_hw_class_01 [ 22 ]        = p3_dirrpl_enq_cnt_oflow_err_f ;
  err_hw_class_01 [ 21 ]        = p3_dirrpl_enq_cnt_uflow_err_f ;
  err_hw_class_01 [ 20 ]        = p3_dirrpl_enq_cnt_res_err ;           // Not flopped, but reasonably fast signal
  err_hw_class_01 [ 19 ]        = p1_dirrpl_inp_frag_cnt_res_err_f ;
  err_hw_class_01 [ 18 ]        = p3_atq_aqed_act_lim_par_err_f ;
  err_hw_class_01 [ 17 ]        = p3_atq_aqed_act_cnt_oflow_err_f ;
  err_hw_class_01 [ 16 ]        = p3_atq_aqed_act_cnt_uflow_err_f ;
  err_hw_class_01 [ 15 ]        = p3_atq_aqed_act_cnt_res_err_f ;
  err_hw_class_01 [ 14 ]        = 1'b0 ;                                // Spare
  err_hw_class_01 [ 13 ]        = p4_atq_atm_active_res_err_f ;
  err_hw_class_01 [ 12 ]        = p3_atq_enq_cnt_res_err_f ;
  err_hw_class_01 [ 11 ]        = p8_lba_qid_if_lim_par_err_f ;
  err_hw_class_01 [ 10 ]        = p8_lba_qid_if_cnt_oflow_err_f ;
  err_hw_class_01 [  9 ]        = p8_lba_qid_if_cnt_res_err_f ;
  err_hw_class_01 [  8 ]        = p4_atq_qid_dpth_thrsh_par_err_f ;
  err_hw_class_01 [  7 ]        = p3_direnq_dpth_thrsh_par_err_f ;
  err_hw_class_01 [  6 ]        = p8_lba_qid_dpth_thrsh_par_err_f ;
  err_hw_class_01 [  5 ]        = p8_lba_qid_enq_cnt_oflow_err_f ;
  err_hw_class_01 [  4 ]        = p8_lba_qid_enq_cnt_uflow_err_f ;
  err_hw_class_01 [  3 ]        = p8_lba_qid_enq_cnt_res_err_f ;
  err_hw_class_01 [  2 ]        = p3_direnq_enq_cnt_oflow_err_f ;
  err_hw_class_01 [  1 ]        = p3_direnq_enq_cnt_uflow_err_f ;
  err_hw_class_01 [  0 ]        = p3_direnq_enq_cnt_res_err_f ;
  err_hw_class_01_v             = | ( err_hw_class_01 [27:0] ) ;

  err_hw_class_02               = '0 ;
  err_hw_class_02 [ 30:28 ]     = 3'h2 ;                                // Class
  err_hw_class_02 [ 27 ]        = p0_lba_cmpblast_lsp_set_err ;         // Not flopped but fast signal
  err_hw_class_02 [ 26 ]        = p0_lba_cmpblast_ap_rst_err ;          // Not flopped but fast signal
  err_hw_class_02 [ 25 ]        = p8_lba_cq_if_lim_par_err_f ;          // Also includes lba_cq_if_thr parity error
  err_hw_class_02 [ 24 ]        = p8_lba_cq_if_cnt_oflow_err_f ;
  err_hw_class_02 [ 23 ]        = p8_lba_cq_if_cnt_res_err_f ;
  err_hw_class_02 [ 22 ]        = p8_lba_cq_tok_lim_par_err_f ;
  err_hw_class_02 [ 21 ]        = p8_lba_cq_tok_cnt_oflow_err_f ;
  err_hw_class_02 [ 20 ]        = p8_lba_cq_tok_cnt_res_err_f ;
  err_hw_class_02 [ 19 ]        = p3_lba_inp_tok_cnt_res_err_f ;
  err_hw_class_02 [ 18 ]        = p3_direnq_tok_lim_par_err_f ;
  err_hw_class_02 [ 17 ]        = p3_direnq_tok_cnt_oflow_err_f ;
  err_hw_class_02 [ 16 ]        = p3_direnq_tok_cnt_res_err_f ;
  err_hw_class_02 [ 15 ]        = p1_direnq_inp_tok_cnt_res_err_f ;
  err_hw_class_02 [ 14 ]        = rx_sync_fifo_error ;                  // Not flopped but reasonably fast signal
  err_hw_class_02 [ 13 ]        = mem_access_error_f ;
  err_hw_class_02 [ 12 ]        = atq_tot_act_lim_err_v ;               // Not flopped but fast signal
  err_hw_class_02 [ 11 ]        = atq_fid_if_lim_err_v ;                // Not flopped but fast signal
  err_hw_class_02 [ 10 ]        = p4_atq_fid_inflight_cnt_oflow_err_f ;
  err_hw_class_02 [  9 ]        = p4_atq_fid_inflight_cnt_uflow_err_f ;
  err_hw_class_02 [  8 ]        = p3_lbrpl_inp_qid_par_err_f ;
  err_hw_class_02 [  7 ]        = p3_dirrpl_inp_qid_par_err_f ;
  err_hw_class_02 [  6 ]        = p4_atq_tot_act_cnt_oflow_err_f ;
  err_hw_class_02 [  5 ]        = p4_atq_tot_act_cnt_uflow_err_f ;
  err_hw_class_02 [  4 ]        = p3_atq_inp_qid_par_err_f ;
  err_hw_class_02 [  3 ]        = p8_lba_tot_if_cnt_oflow_err_f ;
  err_hw_class_02 [  2 ]        = p8_lba_inp_cq_par_err_f ;
  err_hw_class_02 [  1 ]        = p8_lba_inp_qid_par_err_f ;
  err_hw_class_02 [  0 ]        = p3_direnq_inp_qid_cq_par_err_f ;
  err_hw_class_02_v             = | ( err_hw_class_02 [27:0] ) ;

  err_hw_class_03               = '0 ;
  err_hw_class_03 [ 30:28 ]     = 3'h3 ;                                // Class
  err_hw_class_03 [ 27 ]        = hqm_list_sel_pipe_rfw_top_ipar_error ;
  err_hw_class_03 [ 26 ]        = aqed_deq_credit_error ;               // Flopped by AW
  err_hw_class_03 [ 25 ]        = qed_deq_credit_error ;                // Flopped by AW
  err_hw_class_03 [ 24 ]        = lbwu_cq_wu_cnt_rmw_pipe_err_f ;
  err_hw_class_03 [ 23 ]        = aqed_lsp_deq_fifo_of ;
  err_hw_class_03 [ 22 ]        = aqed_lsp_deq_fifo_uf ;
  err_hw_class_03 [ 21 ]        = qed_lsp_deq_fifo_of ;
  err_hw_class_03 [ 20 ]        = qed_lsp_deq_fifo_uf ;
  err_hw_class_03 [ 19 ]        = p4_lba_cq2qid_priov_par_err_f ;
  err_hw_class_03 [ 18 ]        = p4_lba_cq2qid_qid1_par_err_f ;
  err_hw_class_03 [ 17 ]        = p4_lba_cq2qid_qid0_par_err_f ;
  if ( p8_lba_blast_qid2cqidix_par_err_any ) begin
    err_hw_class_03 [ 16 ]      = 1'b1 ;                                // atm
    err_hw_class_03 [ 15:0 ]    = p8_lba_blast_qid2cqidix_par_err_f ;
  end
  if ( p8_lba_qid2cqidix_par_err_any ) begin
    err_hw_class_03 [ 16 ]      = 1'b0 ;                                // ldb
    err_hw_class_03 [ 15:0 ]    = p8_lba_qid2cqidix_par_err_f ;
  end
  err_hw_class_03_v             = | ( err_hw_class_03 [27:0] ) ;

  err_hw_class_04               = '0 ;
  err_hw_class_04 [ 30:28 ]     = 3'h4 ;                                // Class
  err_hw_class_04 [ 27 ]        = p4_lbwu_inp_par_err_f ;
  err_hw_class_04 [ 26 ]        = p0_lba_cq_arb_error_f ;
  err_hw_class_04 [ 25 ]        = uno_atm_cmp_fifo_of ;
  err_hw_class_04 [ 24 ]        = uno_atm_cmp_fifo_uf ;
  err_hw_class_04 [ 23 ]        = p4_lbwu_cq_wu_lim_par_err_f ;
  err_hw_class_04 [ 22 ]        = p4_lbwu_cq_wu_cnt_res_err_f ;
  err_hw_class_04 [ 21 ]        = ldb_token_rtn_fifo_of ;
  err_hw_class_04 [ 20 ]        = ldb_token_rtn_fifo_uf ;
  err_hw_class_04 [ 19 ]        = atm_cmp_fifo_of ;
  err_hw_class_04 [ 18 ]        = atm_cmp_fifo_uf ;
  err_hw_class_04 [ 17 ]        = enq_nalb_fifo_of ;
  err_hw_class_04 [ 16 ]        = enq_nalb_fifo_uf ;
  err_hw_class_04 [ 15 ]        = nalb_sel_nalb_fifo_of ;
  err_hw_class_04 [ 14 ]        = nalb_sel_nalb_fifo_uf ;
  err_hw_class_04 [ 13 ]        = nalb_cmp_fifo_of ;
  err_hw_class_04 [ 12 ]        = nalb_cmp_fifo_uf ;
  err_hw_class_04 [ 11 ]        = lbrpl_enq_cnt_rmw_pipe_err_f ;
  err_hw_class_04 [ 10 ]        = dirrpl_enq_cnt_rmw_pipe_err_f ;
  err_hw_class_04 [  9 ]        = atq_enq_cnt_rmw_pipe_err_f ;
  err_hw_class_04 [  8 ]        = lba_arbindex_rmw_pipe_err_f ;         // nalb or atm
  err_hw_class_04 [  7 ]        = lba_qid2cqidix_rw_pipe_err_f ;
  err_hw_class_04 [  6 ]        = lba_cq_tok_cnt_rmw_pipe_err_f ;
  err_hw_class_04 [  5 ]        = direnq_enq_cnt_rmw_pipe_err_f ;
  err_hw_class_04 [  4 ]        = lba_cq2qid_rw_pipe_err_f ;
  err_hw_class_04 [  3 ]        = p4_atq_fid_inflight_cnt_res_err_f ;
  err_hw_class_04 [  2 ]        = p4_atq_aqed_tot_enq_cnt_res_err_f ;
  err_hw_class_04 [  1 ]        = p9_lba_nalb_sch_err_f ;
  err_hw_class_04 [  0 ]        = p8_lba_tot_if_cnt_res_err_f ;
  err_hw_class_04_v             = | ( err_hw_class_04 [27:0] ) ;

  err_hw_class_05               = '0 ;
  err_hw_class_05 [ 30:28 ]     = 3'h5 ;                                // Class
  err_hw_class_05 [ 27:5 ]      = '0 ;                                  // spare
  err_hw_class_05 [  4 ]        = p4_atq_tot_enq_cnt_res_err_f ;
  err_hw_class_05 [  3 ]        = p9_lba_tot_enq_cnt_res_err_f ;
  err_hw_class_05 [  2 ]        = p4_direnq_tot_enq_cnt_res_err_f ;
  err_hw_class_05 [  1 ]        = p9_lba_tot_sch_cnt_res_err_f ;
  err_hw_class_05 [  0 ]        = p4_direnq_tot_sch_cnt_res_err_f ;
  err_hw_class_05_v             = | ( err_hw_class_05 [27:0] ) ;
end // always


always_comb begin
  int_inf_v                     = '0 ;
  int_inf_data                  = '0 ;
  int_cor_v                     = '0 ;
  int_cor_data                  = '0 ;
  int_unc_v                     = '0 ;
  int_unc_data                  = '0 ;

  lsp_uid                       = HQM_LSP_CFG_UNIT_ID ;
  cfg_syndrome0_capture_v       = 1'b0 ;
  cfg_syndrome0_capture_data    = 31'h0 ;
  cfg_syndrome1_capture_v       = 1'b0 ;
  cfg_syndrome1_capture_data    = 31'h0 ;

  // Prioritize the interrupts from least serious (sw-caused) to most serious (pf reset required) so that
  // in the unlikely event of simultaneous interrupts, the most important loads the syndrome registers.
  // Keep syndrome for software-causable interrupts separate from hardware errors to avoid confusion.

  // May want to move all "hardware" errors out of cfg_syndrome_1 (cfg_syndrome_sw) for consistency, evolved to this point after token underflow change.
  // token underflow                    : can be caused by sw, CHP screens out so should only get to LSP if CHP hw failure
  // per-CQ completion underflow        : can be caused by sw, CHP screens out so should only get to LSP if CHP hw failure
  // per-QID completion underflow       : can be caused by sw, CHP screens "full" completion but not RELEASE

  // ######################################################################################################
  // This section of code is generated by a script and should not be hand-editted

  //  p8_lba_cq_tok_cnt_uflow_err_f "SW Error" "Load balanced token count underflow
  if ( p8_lba_cq_tok_cnt_uflow_err_f & ~cfg_control_disable_tok_uflow_interrupt  ) begin
    int_inf_v [ 2 ]                                = 1'b1 ;
    int_inf_data [ 2 ].rtype                       = 2'd1 ;
    int_inf_data [ 2 ].rid                         = p8_lba_cq_tok_cnt_uflow_err_rid ;
    int_inf_data [ 2 ].msix_map                    = INGRESS_ERROR ;            // Should be changed to HQM_ALARM : screened by CHP
    cfg_syndrome1_capture_v                        = ~cfg_control_disable_tok_uflow_synd_load ;
    cfg_syndrome1_capture_data                     = 31'h00000001 ;
  end
  //  p3_direnq_tok_cnt_uflow_err_f "SW Error" "Directed token count underflow
  if ( p3_direnq_tok_cnt_uflow_err_f & ~cfg_control_disable_tok_uflow_interrupt  ) begin
    int_inf_v [ 2 ]                                = 1'b1 ;
    int_inf_data [ 2 ].rtype                       = 2'd1 ;
    int_inf_data [ 2 ].rid                         = p3_direnq_tok_cnt_uflow_err_rid ;
    int_inf_data [ 2 ].msix_map                    = INGRESS_ERROR ;            // Should be changed to HQM_ALARM : screened by CHP
    cfg_syndrome1_capture_v                        = ~cfg_control_disable_tok_uflow_synd_load ;
    cfg_syndrome1_capture_data                     = 31'h00000002 ;
  end
  //  p8_lba_tot_if_cnt_uflow_err_f "HW Error" "Total inflight count underflow
  if ( p8_lba_tot_if_cnt_uflow_err_f & ~cfg_control_disable_cq_if_uflow_interrupt  ) begin
    int_inf_v [ 1 ]                                = 1'b1 ;
    int_inf_data [ 1 ].rtype                       = 2'd1 ;
    int_inf_data [ 1 ].rid                         = p8_lba_tot_if_cnt_uflow_err_rid ;
    int_inf_data [ 1 ].msix_map                    = HQM_ALARM ;                // Screened by CHP
    cfg_syndrome1_capture_v                        = ~cfg_control_disable_cq_if_uflow_synd_load ;
    cfg_syndrome1_capture_data                     = 31'h00000004 ;
  end
  //  p8_lba_cq_if_cnt_uflow_err_f "HW Error" "Per-CQ inflight count underflow
  if ( p8_lba_cq_if_cnt_uflow_err_f & ~cfg_control_disable_cq_if_uflow_interrupt  ) begin
    int_inf_v [ 1 ]                                = 1'b1 ;
    int_inf_data [ 1 ].rtype                       = 2'd1 ;
    int_inf_data [ 1 ].rid                         = p8_lba_cq_if_cnt_uflow_err_rid ;
    int_inf_data [ 1 ].msix_map                    = HQM_ALARM ;                // Screened by CHP
    cfg_syndrome1_capture_v                        = ~cfg_control_disable_cq_if_uflow_synd_load ;
    cfg_syndrome1_capture_data                     = 31'h00000008 ;
  end
  //  p8_lba_qid_if_cnt_uflow_err_f "SW Error" "Per-QID inflight count underflow
  if ( p8_lba_qid_if_cnt_uflow_err_f & ~cfg_control_disable_qid_if_uflow_interrupt  ) begin
    int_inf_v [ 0 ]                                = 1'b1 ;
    int_inf_data [ 0 ].rtype                       = 2'd2 ;
    int_inf_data [ 0 ].rid                         = p8_lba_qid_if_cnt_uflow_err_rid ;
    int_inf_data [ 0 ].msix_map                    = INGRESS_ERROR ;            // Possibly caused by sw, much more likely than hw failure in CHP
    cfg_syndrome1_capture_v                        = ~cfg_control_disable_qid_if_uflow_synd_load ;
    cfg_syndrome1_capture_data                     = 31'h00000010 ;
  end
  //  err_hw_class_01_v "HW Error" "Hardware error
  if ( err_hw_class_01_v & ~cfg_control_disable_hwerr_interrupt  ) begin
    int_inf_v [ 3 ]                                = 1'b1 ;
    int_inf_data [ 3 ].rtype                       = 2'd0 ;
    int_inf_data [ 3 ].rid                         = 8'h0 ;
    int_inf_data [ 3 ].msix_map                    = HQM_ALARM ;
    cfg_syndrome0_capture_v                        = ~cfg_control_disable_hwerr_synd_load ;
    cfg_syndrome0_capture_data                     = err_hw_class_01 ;
  end
  //  err_hw_class_02_v "HW Error" "Hardware error
  if ( err_hw_class_02_v & ~cfg_control_disable_hwerr_interrupt  ) begin
    int_inf_v [ 3 ]                                = 1'b1 ;
    int_inf_data [ 3 ].rtype                       = 2'd0 ;
    int_inf_data [ 3 ].rid                         = 8'h0 ;
    int_inf_data [ 3 ].msix_map                    = HQM_ALARM ;
    cfg_syndrome0_capture_v                        = ~cfg_control_disable_hwerr_synd_load ;
    cfg_syndrome0_capture_data                     = err_hw_class_02 ;
  end
  //  err_hw_class_03_v "HW Error" "Hardware error
  if ( err_hw_class_03_v & ~cfg_control_disable_hwerr_interrupt  ) begin
    int_inf_v [ 3 ]                                = 1'b1 ;
    int_inf_data [ 3 ].rtype                       = 2'd0 ;
    int_inf_data [ 3 ].rid                         = 8'h0 ;
    int_inf_data [ 3 ].msix_map                    = HQM_ALARM ;
    cfg_syndrome0_capture_v                        = ~cfg_control_disable_hwerr_synd_load ;
    cfg_syndrome0_capture_data                     = err_hw_class_03 ;
  end
  //  err_hw_class_04_v "HW Error" "Hardware error
  if ( err_hw_class_04_v & ~cfg_control_disable_hwerr_interrupt  ) begin
    int_inf_v [ 3 ]                                = 1'b1 ;
    int_inf_data [ 3 ].rtype                       = 2'd0 ;
    int_inf_data [ 3 ].rid                         = 8'h0 ;
    int_inf_data [ 3 ].msix_map                    = HQM_ALARM ;
    cfg_syndrome0_capture_v                        = ~cfg_control_disable_hwerr_synd_load ;
    cfg_syndrome0_capture_data                     = err_hw_class_04 ;
  end
  //  err_hw_class_05_v "HW Error" Hardware error (non-mission critical)
  if ( err_hw_class_05_v & ~cfg_control_disable_non_mc_interrupt  ) begin
    int_inf_v [ 4 ]                                = 1'b1 ;
    int_inf_data [ 4 ].rtype                       = 2'd0 ;
    int_inf_data [ 4 ].rid                         = 8'h0 ;
    int_inf_data [ 4 ].msix_map                    = HQM_ALARM ;
    cfg_syndrome0_capture_v                        = ~cfg_control_disable_non_mc_synd_load ;
    cfg_syndrome0_capture_data                     = err_hw_class_05 ;
  end
  // ######################################################################################################

end // always


assign int_serializer_status_up         = int_serializer_status_pnc [2:0] ;
assign int_serializer_status_down       = int_serializer_status_pnc [9:7] ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: Unit interfaces and input buffering
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// chp_lsp_token: Used for returning tokens, loads either the LDB TOKRTN FIFO or DIR TOKRTN FIFO, which
// then feed into the LBARB and DIRENQ pipes respectively.

// core_chp_lsp_token_data is sourced by i_hqm_AW_rx_sync_chp_lsp_token

always_comb begin
  if ( core_chp_lsp_token_v & ( core_chp_lsp_token_data.is_ldb == 1'b1 ) )
    core_chp_lsp_token_ready            = ~ ldb_token_rtn_fifo_afull ;
  else
    core_chp_lsp_token_ready            = ~ dir_tokrtn_fifo_afull ;
end // always

assign dir_tokrtn_fifo_push             = core_chp_lsp_token_v & ~ dir_tokrtn_fifo_afull & ( core_chp_lsp_token_data.is_ldb == 1'b0 ) ;
assign dir_tokrtn_fifo_push_data        = core_chp_lsp_token_data ;
assign dir_tokrtn_fifo_afull            = ~ dir_tokrtn_db_in_ready ;

assign ldb_token_rtn_fifo_push          = core_chp_lsp_token_v & ~ ldb_token_rtn_fifo_afull & ( core_chp_lsp_token_data.is_ldb == 1'b1 ) ;
assign ldb_token_rtn_fifo_push_data.cq                  = core_chp_lsp_token_data.cq ;
assign ldb_token_rtn_fifo_push_data.is_ldb              = core_chp_lsp_token_data.is_ldb ;
assign ldb_token_rtn_fifo_push_data.parity              = core_chp_lsp_token_data.parity ;
assign ldb_token_rtn_fifo_push_data.count               = core_chp_lsp_token_data.count ;
assign ldb_token_rtn_fifo_push_data.count_residue       = core_chp_lsp_token_data.count_residue ;

hqm_AW_double_buffer #( .WIDTH ( $bits ( chp_lsp_token_data ) ) ) i_dir_token_rtn_if_db (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( dir_tokrtn_db_status_pnc )
        , .in_ready             ( dir_tokrtn_db_in_ready )
        , .in_valid             ( dir_tokrtn_fifo_push )
        , .in_data              ( dir_tokrtn_fifo_push_data )
        , .out_ready            ( dir_tokrtn_fifo_pop )
        , .out_valid            ( dir_tokrtn_db_out_valid )
        , .out_data             ( dir_tokrtn_fifo_pop_data )
) ;

assign dir_tokrtn_fifo_pop_data_cq      = dir_tokrtn_fifo_pop_data.cq [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0] ;

assign ldb_token_rtn_fifo_hwm           = HQM_LSP_LDB_TOKEN_RTN_FIFO_DEPTH [HQM_LSP_LDB_TOKEN_RTN_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control_latepp #(
          .DEPTH                ( HQM_LSP_LDB_TOKEN_RTN_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_LDB_TOKEN_RTN_FIFO_DWIDTH )
) i_ldb_token_rtn_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( ldb_token_rtn_fifo_push )
        , .push_data            ( ldb_token_rtn_fifo_push_data )
        , .pop                  ( ldb_token_rtn_fifo_pop )
        , .pop_data             ( ldb_token_rtn_fifo_pop_data )

        , .cfg_high_wm          ( ldb_token_rtn_fifo_hwm )

        , .mem_we               ( func_ldb_token_rtn_fifo_mem_we )
        , .mem_waddr            ( func_ldb_token_rtn_fifo_mem_waddr )
        , .mem_wdata            ( func_ldb_token_rtn_fifo_mem_wdata )
        , .mem_re               ( func_ldb_token_rtn_fifo_mem_re )
        , .mem_raddr            ( func_ldb_token_rtn_fifo_mem_raddr )
        , .mem_rdata            ( func_ldb_token_rtn_fifo_mem_rdata )

        , .fifo_status          ( ldb_token_rtn_fifo_status_pnc )
        , .fifo_full            ( ldb_token_rtn_fifo_full_nc )
        , .fifo_afull           ( ldb_token_rtn_fifo_afull )
        , .fifo_empty           ( ldb_token_rtn_fifo_empty )
) ;
assign ldb_token_rtn_fifo_pop_data_nc                   = ldb_token_rtn_fifo_pop_data.cq[7:6] ;

assign ldb_token_rtn_fifo_of                            = ldb_token_rtn_fifo_status_pnc [1] ;
assign ldb_token_rtn_fifo_uf                            = ldb_token_rtn_fifo_status_pnc [0] | cfg_error_inject_f [ 7 ] ;

assign dir_tokrtn_fifo_empty            = ~ dir_tokrtn_db_out_valid ;
assign dir_tokrtn_fifo_pop_data_v       = ~ dir_tokrtn_fifo_empty ;
assign dir_tokrtn_fifo_pop_data_vreq    = dir_tokrtn_fifo_pop_data_v & ~ cause_pipe_idle ;

assign dir_tokrtn_fifo_pop              = direnq_input_arb_tok ;
assign ldb_token_rtn_fifo_pop_data_v    = ~ ldb_token_rtn_fifo_empty ;
assign ldb_token_rtn_fifo_pop_data_vreq = ldb_token_rtn_fifo_pop_data_v & ~ cause_pipe_idle ;

//-----------------------------------------------------------------------------------------------------
// chp_lsp_cmp: Used for returning unordered and atm completions, loads the UNO_ATM_CMP FIFO and
// ATM_CMP FIFO

// core_chp_lsp_cmp_data is sourced by i_hqm_AW_rx_sync_chp_lsp_cmp

// HL parity includes all fields sent to AP, plus fields not used (reord_mode, reord_slot).
// Subtract them out, then derive the other parities that are needed from that.

// Subtract fields not sent to AP and expected to be included in the parity.
// qid parity is sent as part of chp_lsp_cmp.parity so subtract here so not counted twice
hqm_AW_parity_gen #( .WIDTH( 1 + 2 + HQM_LSP_ARCH_NUM_LB_QIDB2 + 3 + 5 ) ) i_atm_ap_par_gen (
          .d            ( {   core_chp_lsp_cmp_data.hist_list_info.parity       // On all of hist_list_info
                            , core_chp_lsp_cmp_data.hist_list_info.qtype
                            , { 1'b0 , core_chp_lsp_cmp_data.hist_list_info.qid }
                            , core_chp_lsp_cmp_data.hist_list_info.reord_mode
                            , core_chp_lsp_cmp_data.hist_list_info.reord_slot } )
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( core_chp_lsp_cmp_data_ap_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 12 ) ) i_atm_fid_par_gen (
          .d            ( {   core_chp_lsp_cmp_data_ap_p
                            , core_chp_lsp_cmp_data.hist_list_info.sn_fid.fid } )
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( core_chp_lsp_cmp_data_cmp_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 3 + 1 + 3 ) ) i_atm_cmp_par_gen (
          .d            ( {   core_chp_lsp_cmp_data_ap_p
                            , core_chp_lsp_cmp_data.hist_list_info.qpri
                            , core_chp_lsp_cmp_data.hist_list_info.qidix_msb
                            , core_chp_lsp_cmp_data.hist_list_info.qidix } )
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( core_chp_lsp_cmp_data_fid_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 2 ) ) i_uno_atm_cmp_cq_qid_par_gen (
          .d            ( {   core_chp_lsp_cmp_data.parity
                            , core_chp_lsp_cmp_data.qe_wt } )
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( core_chp_lsp_cmp_data_cq_qid_p )
) ;

// Only pop from buffer and push to any FIFO if all FIFOs that are needed are available.
// FIFO is "available" if it is not needed, or if it is needed but not afull.

// Note: On a "release" command (user[1:0]=2), the hist_list_info (including qtype) is invalid.
assign core_chp_lsp_cmp_rel_v           = core_chp_lsp_cmp_v & ( core_chp_lsp_cmp_data.user[1:0] == 2'b10 ) ;

assign core_chp_lsp_cmp_uno_v           = core_chp_lsp_cmp_v & ( ~ core_chp_lsp_cmp_rel_v ) & ( core_chp_lsp_cmp_data.hist_list_info.qtype == UNORDERED ) ;
assign core_chp_lsp_cmp_atm_v           = core_chp_lsp_cmp_v & ( ~ core_chp_lsp_cmp_rel_v ) & ( core_chp_lsp_cmp_data.hist_list_info.qtype == ATOMIC ) ;
assign core_chp_lsp_cmp_nalb_v          = core_chp_lsp_cmp_v & ( ~ core_chp_lsp_cmp_rel_v ) & ( ( core_chp_lsp_cmp_data.hist_list_info.qtype == UNORDERED ) |
                                                                                                ( core_chp_lsp_cmp_data.hist_list_info.qtype == ORDERED ) ) ;

assign uno_atm_cmp_fifo_ready           = ~ ( ( core_chp_lsp_cmp_uno_v | core_chp_lsp_cmp_atm_v | core_chp_lsp_cmp_rel_v ) & uno_atm_cmp_fifo_afull ) ;
assign atm_cmp_fifo_ready               = ~ ( core_chp_lsp_cmp_atm_v  & atm_cmp_fifo_afull ) ;
assign nalb_cmp_fifo_ready              = ~ ( core_chp_lsp_cmp_nalb_v & nalb_cmp_fifo_afull ) ;

assign core_chp_lsp_cmp_ready           = uno_atm_cmp_fifo_ready & atm_cmp_fifo_ready & nalb_cmp_fifo_ready ;

assign uno_atm_cmp_fifo_push            = ( core_chp_lsp_cmp_uno_v | core_chp_lsp_cmp_atm_v | core_chp_lsp_cmp_rel_v ) & core_chp_lsp_cmp_ready ;
assign atm_cmp_fifo_push                = core_chp_lsp_cmp_atm_v  & core_chp_lsp_cmp_ready ;
assign nalb_cmp_fifo_push               = core_chp_lsp_cmp_nalb_v & core_chp_lsp_cmp_ready ;

always_comb begin
  uno_atm_cmp_fifo_push_data.cq         = core_chp_lsp_cmp_data.pp ;
  uno_atm_cmp_fifo_push_data.qid        = core_chp_lsp_cmp_data.qid ;
  uno_atm_cmp_fifo_push_data.cq_qid_p   = core_chp_lsp_cmp_data_cq_qid_p ;
  uno_atm_cmp_fifo_push_data.user       = core_chp_lsp_cmp_data.user ;
  uno_atm_cmp_fifo_push_data.spare      = 2'h0 ;
end // always

assign uno_atm_cmp_fifo_hwm             = HQM_LSP_UNO_ATM_CMP_FIFO_DEPTH [HQM_LSP_UNO_ATM_CMP_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control_latepp #(
          .DEPTH                ( HQM_LSP_UNO_ATM_CMP_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_UNO_ATM_CMP_FIFO_DWIDTH )
) i_uno_atm_cmp_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( uno_atm_cmp_fifo_push )
        , .push_data            ( uno_atm_cmp_fifo_push_data )
        , .pop                  ( uno_atm_cmp_fifo_pop )
        , .pop_data             ( uno_atm_cmp_fifo_pop_data )

        , .cfg_high_wm          ( uno_atm_cmp_fifo_hwm )

        , .mem_we               ( func_uno_atm_cmp_fifo_mem_we )
        , .mem_waddr            ( func_uno_atm_cmp_fifo_mem_waddr )
        , .mem_wdata            ( func_uno_atm_cmp_fifo_mem_wdata )
        , .mem_re               ( func_uno_atm_cmp_fifo_mem_re )
        , .mem_raddr            ( func_uno_atm_cmp_fifo_mem_raddr )
        , .mem_rdata            ( func_uno_atm_cmp_fifo_mem_rdata )

        , .fifo_status          ( uno_atm_cmp_fifo_status_pnc )
        , .fifo_full            ( uno_atm_cmp_fifo_full_nc )
        , .fifo_afull           ( uno_atm_cmp_fifo_afull )
        , .fifo_empty           ( uno_atm_cmp_fifo_empty )
) ;
assign uno_atm_cmp_fifo_pop_data_nc                     = uno_atm_cmp_fifo_pop_data.spare ;

assign uno_atm_cmp_fifo_of                              = uno_atm_cmp_fifo_status_pnc [1] ;
assign uno_atm_cmp_fifo_uf                              = uno_atm_cmp_fifo_status_pnc [0] ;

assign uno_atm_cmp_fifo_pop_data_v      = ~ uno_atm_cmp_fifo_empty ;
assign uno_atm_cmp_fifo_pop_data_vreq   = uno_atm_cmp_fifo_pop_data_v & ~ cause_pipe_idle ;

//--------
always_comb begin
  nalb_cmp_fifo_push_data.cq            = core_chp_lsp_cmp_data.pp ;
  nalb_cmp_fifo_push_data.qid           = core_chp_lsp_cmp_data.qid ;
  nalb_cmp_fifo_push_data.qe_wt         = core_chp_lsp_cmp_data.qe_wt ;
  nalb_cmp_fifo_push_data.parity        = core_chp_lsp_cmp_data.parity ;
end // always

assign nalb_cmp_fifo_hwm                = HQM_LSP_NALB_CMP_FIFO_DEPTH [HQM_LSP_NALB_CMP_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control_latepp #(
          .DEPTH                ( HQM_LSP_NALB_CMP_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_NALB_CMP_FIFO_DWIDTH )
) i_nalb_cmp_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( nalb_cmp_fifo_push )
        , .push_data            ( nalb_cmp_fifo_push_data )
        , .pop                  ( nalb_cmp_fifo_pop )
        , .pop_data             ( nalb_cmp_fifo_pop_data )

        , .cfg_high_wm          ( nalb_cmp_fifo_hwm )

        , .mem_we               ( func_nalb_cmp_fifo_mem_we )
        , .mem_waddr            ( func_nalb_cmp_fifo_mem_waddr )
        , .mem_wdata            ( func_nalb_cmp_fifo_mem_wdata )
        , .mem_re               ( func_nalb_cmp_fifo_mem_re )
        , .mem_raddr            ( func_nalb_cmp_fifo_mem_raddr )
        , .mem_rdata            ( func_nalb_cmp_fifo_mem_rdata )

        , .fifo_status          ( nalb_cmp_fifo_status_pnc )
        , .fifo_full            ( nalb_cmp_fifo_full_nc )
        , .fifo_afull           ( nalb_cmp_fifo_afull )
        , .fifo_empty           ( nalb_cmp_fifo_empty )
) ;

assign nalb_cmp_fifo_pop_data_cq_ms_nc                  = nalb_cmp_fifo_pop_data.cq[7:6] ;

assign nalb_cmp_fifo_of                                 = nalb_cmp_fifo_status_pnc [1] ;
assign nalb_cmp_fifo_uf                                 = nalb_cmp_fifo_status_pnc [0] ;

assign nalb_cmp_fifo_pop_data_v         = ~ nalb_cmp_fifo_empty ;
assign nalb_cmp_fifo_pop_data_vreq      = nalb_cmp_fifo_pop_data_v & ~ cause_pipe_idle ;

hqm_AW_parity_gen #( .WIDTH( 1 + HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_nalb_cmp_cq_wt_par_gen (       // Subtract out the qid parity
          .d            ( {   nalb_cmp_fifo_pop_data.parity 
                            , nalb_cmp_fifo_pop_data.qid } )
        , .odd          ( 1'b0 )                                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( nalb_cmp_fifo_pop_data_cq_wt_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 2 ) ) i_nalb_cmp_cq_par_gen (                                  // Subtract out the qe_wt parity
          .d            ( {   nalb_cmp_fifo_pop_data_cq_wt_p
                            , nalb_cmp_fifo_pop_data.qe_wt } )
        , .odd          ( 1'b0 )                                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( nalb_cmp_fifo_pop_data_cq_p )
) ;


//-----------------------------------------------------------------------------------------------------
// qed_lsp_deq, aqed_lsp_deq : Dequeue (sent by QED or AQED to CHP for scheduling) indication

// core_qed_lsp_deq_data and core_aqed_lsp_deq_data are sourced by i_hqm_AW_rx_sync_qed_lsp_deq and i_hqm_AW_rx_sync_aqed_lsp_deq inside i_hqm_lsp_wu_pipe

//-----------------------------------------------------------------------------------------------------
// nalb_lsp_enq_lb : Non-Atomic Load Balanced enqueue requests, loads the enq_nalb and enq_atq FIFOs

// core_nalb_lsp_enq_lb_data is sourced by i_hqm_AW_rx_sync_nalb_lsp_enq_lb

always_comb begin
  if ( core_nalb_lsp_enq_lb_v & ( core_nalb_lsp_enq_lb_data.qtype == ATOMIC ) ) begin
    core_nalb_lsp_enq_lb_ready          = enq_atq_db_in_ready ;
    enq_atq_db_in_valid                 = core_nalb_lsp_enq_lb_v & core_nalb_lsp_enq_lb_ready ;
    enq_nalb_fifo_push                  = 1'b0 ;
  end
  else begin
    core_nalb_lsp_enq_lb_ready          = ~ enq_nalb_fifo_afull ;
    enq_atq_db_in_valid                 = 1'b0  ;
    enq_nalb_fifo_push                  = core_nalb_lsp_enq_lb_v & core_nalb_lsp_enq_lb_ready ;
  end
end // always

assign enq_nalb_fifo_push_data          = core_nalb_lsp_enq_lb_data ;
assign enq_atq_db_in_data               = core_nalb_lsp_enq_lb_data ;

assign enq_nalb_fifo_hwm                = HQM_LSP_ENQ_NALB_FIFO_DEPTH [HQM_LSP_ENQ_NALB_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control_latepp #(
          .DEPTH                ( HQM_LSP_ENQ_NALB_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_ENQ_NALB_FIFO_DWIDTH )
) i_enq_nalb_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( enq_nalb_fifo_push )
        , .push_data            ( enq_nalb_fifo_push_data )
        , .pop                  ( enq_nalb_fifo_pop )
        , .pop_data             ( enq_nalb_fifo_pop_data )

        , .cfg_high_wm          ( enq_nalb_fifo_hwm )

        , .mem_we               ( func_enq_nalb_fifo_mem_we )
        , .mem_waddr            ( func_enq_nalb_fifo_mem_waddr )
        , .mem_wdata            ( func_enq_nalb_fifo_mem_wdata )
        , .mem_re               ( func_enq_nalb_fifo_mem_re )
        , .mem_raddr            ( func_enq_nalb_fifo_mem_raddr )
        , .mem_rdata            ( func_enq_nalb_fifo_mem_rdata )

        , .fifo_status          ( enq_nalb_fifo_status_pnc )
        , .fifo_full            ( enq_nalb_fifo_full_nc )
        , .fifo_afull           ( enq_nalb_fifo_afull )
        , .fifo_empty           ( enq_nalb_fifo_empty )
) ;
assign enq_nalb_fifo_of                         = enq_nalb_fifo_status_pnc [1] ;
assign enq_nalb_fifo_uf                         = enq_nalb_fifo_status_pnc [0] ;

assign enq_nalb_fifo_pop_data_v         = ~ enq_nalb_fifo_empty ;
assign enq_nalb_fifo_pop_data_vreq      = enq_nalb_fifo_pop_data_v & ~ cause_pipe_idle ;

hqm_AW_double_buffer #( .WIDTH ( $bits ( enq_atq_db_in_data ) ) ) i_enq_atq_db (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( enq_atq_db_status_pnc )
        , .in_ready             ( enq_atq_db_in_ready )
        , .in_valid             ( enq_atq_db_in_valid ) 
        , .in_data              ( enq_atq_db_in_data )
        , .out_ready            ( enq_atq_db_out_ready )
        , .out_valid            ( enq_atq_db_out_valid )
        , .out_data             ( enq_atq_db_out_data )
) ;

assign enq_atq_db_out_ready     = enq_atq_fifo_pop ;

assign enq_atq_fifo_pop_data    = enq_atq_db_out_data ;

assign enq_atq_fifo_pop_data_v          = enq_atq_db_out_valid ;
assign enq_atq_fifo_pop_data_vreq       = enq_atq_fifo_pop_data_v & ~ cause_pipe_idle ;

assign enq_atq_fifo_pop         = atq_input_arb_enq ;

//-----------------------------------------------------------------------------------------------------
// nalb_lsp_enq_rorply : Non-Atomic Load Balanced reorder-complete replay requests
// Lower bandwidth, only use double buffer

// core_nalb_lsp_enq_rorply_data is sourced by i_hqm_AW_rx_sync_nalb_lsp_enq_rorply

assign core_nalb_lsp_enq_rorply_ready   = nalbrpl_fifo_pop ;

assign nalbrpl_fifo_pop_data_v          = core_nalb_lsp_enq_rorply_v ;
assign nalbrpl_fifo_pop_data_vreq       = nalbrpl_fifo_pop_data_v & ~ cause_pipe_idle ;

assign nalbrpl_fifo_pop         = lbrpl_input_arb_enq ;
assign nalbrpl_fifo_pop_data    = core_nalb_lsp_enq_rorply_data ;

//-----------------------------------------------------------------------------------------------------
// dp_lsp_enq_rorply : Direct reorder-complete replay requests
// Lower bandwidth, only use double buffer

// core_dp_lsp_enq_rorply_data is sourced by i_hqm_AW_rx_sync_dp_lsp_enq_rorply

assign core_dp_lsp_enq_rorply_ready     = dirrpl_fifo_pop ;

assign dirrpl_fifo_pop_data_v           = core_dp_lsp_enq_rorply_v ;
assign dirrpl_fifo_pop_data_vreq        = dirrpl_fifo_pop_data_v & ~ cause_pipe_idle ;

assign dirrpl_fifo_pop          = dirrpl_input_arb_enq ;
assign dirrpl_fifo_pop_data     = core_dp_lsp_enq_rorply_data ;

//-----------------------------------------------------------------------------------------------------
// send_atm_to_cq : AQED ATM schedule requests - need to decrement AQED Active Count
// send_atm_to_cq_data is sourced by i_hqm_AW_rx_sync_send_atm_to_cq

assign send_atm_to_cq_ready             = send_atm_to_cq_fifo_pop ;

assign send_atm_to_cq_fifo_pop_data_v           = send_atm_to_cq_v ;
assign send_atm_to_cq_fifo_pop_data_vreq        = send_atm_to_cq_fifo_pop_data_v & ~ cause_pipe_idle ;

assign send_atm_to_cq_fifo_pop          = atq_input_arb_cmp ;           // Only asserted if pop_data_v=1
assign send_atm_to_cq_fifo_pop_data     = send_atm_to_cq_data ;
assign send_atm_to_cq_fifo_pop_data_flid_nc     = { send_atm_to_cq_fifo_pop_data.flid_parity , send_atm_to_cq_fifo_pop_data.flid } ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: LBARB pipe - Load Balanced arbitration
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB ATM completions
//-----------------------------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------------------------
assign atm_cmp_fifo_push_data.user              = ( core_chp_lsp_cmp_data.user == 2'b11 ) ;
assign atm_cmp_fifo_push_data.cq                = core_chp_lsp_cmp_data.pp [ 6 : 0 ] ;
assign atm_cmp_fifo_push_data.qid               = core_chp_lsp_cmp_data.qid [ 5 : 0 ] ;
assign atm_cmp_fifo_push_data.qe_wt             = core_chp_lsp_cmp_data.qe_wt ;
assign atm_cmp_fifo_push_data.parity            = core_chp_lsp_cmp_data.parity ;
assign atm_cmp_fifo_push_data.qpri              = core_chp_lsp_cmp_data.hist_list_info.qpri ;
assign atm_cmp_fifo_push_data.qidix_msb         = core_chp_lsp_cmp_data.hist_list_info.qidix_msb ;
assign atm_cmp_fifo_push_data.qidix             = core_chp_lsp_cmp_data.hist_list_info.qidix ;
assign atm_cmp_fifo_push_data.cmp_p             = core_chp_lsp_cmp_data_cmp_p ; // Subtracted out cmp fields not sent to AP, and fid
assign atm_cmp_fifo_push_data.fid               = core_chp_lsp_cmp_data.hist_list_info.sn_fid.fid ;
assign atm_cmp_fifo_push_data.fid_p             = core_chp_lsp_cmp_data_fid_p ;
assign atm_cmp_fifo_push_data.hid               = core_chp_lsp_cmp_data.hid ;
assign atm_cmp_fifo_push_data.hid_p             = core_chp_lsp_cmp_data.hid_parity ;


assign atm_cmp_fifo_hwm                 = HQM_LSP_ATM_CMP_FIFO_DEPTH [HQM_LSP_ATM_CMP_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control_latepp #(
          .DEPTH                ( HQM_LSP_ATM_CMP_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_ATM_CMP_FIFO_DWIDTH )
) i_atm_cmp_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( atm_cmp_fifo_push )
        , .push_data            ( atm_cmp_fifo_push_data )
        , .pop                  ( atm_cmp_fifo_pop )
        , .pop_data             ( atm_cmp_fifo_pop_data )

        , .cfg_high_wm          ( atm_cmp_fifo_hwm )

        , .mem_we               ( func_atm_cmp_fifo_mem_we )
        , .mem_waddr            ( func_atm_cmp_fifo_mem_waddr )
        , .mem_wdata            ( func_atm_cmp_fifo_mem_wdata )
        , .mem_re               ( func_atm_cmp_fifo_mem_re )
        , .mem_raddr            ( func_atm_cmp_fifo_mem_raddr )
        , .mem_rdata            ( func_atm_cmp_fifo_mem_rdata )

        , .fifo_status          ( atm_cmp_fifo_status_pnc )
        , .fifo_full            ( atm_cmp_fifo_full_nc )
        , .fifo_afull           ( atm_cmp_fifo_afull )
        , .fifo_empty           ( atm_cmp_fifo_empty )
) ;

assign atm_cmp_fifo_of                                  = atm_cmp_fifo_status_pnc [1] ;
assign atm_cmp_fifo_uf                                  = atm_cmp_fifo_status_pnc [0] ;

// Can't allow atomic completion if no atm credits - goes to AP
assign atm_cmp_fifo_pop_data_v          = ~ atm_cmp_fifo_empty & ~ p0_lba_atm_credit_hold_cond & ~ atm_cmp_fifo_single_op_hold ;
assign atm_cmp_fifo_pop_data_vreq       = atm_cmp_fifo_pop_data_v & ~ cause_pipe_idle ;

hqm_AW_parity_gen #( .WIDTH( 1 + HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_atm_cmp_cq_wt_par_gen (        // Subtract out the qid parity
          .d            ( {   atm_cmp_fifo_pop_data.parity 
                            , { 1'b0 , atm_cmp_fifo_pop_data.qid } } )
        , .odd          ( 1'b0 )                                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( atm_cmp_fifo_pop_data_cq_wt_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 2 ) ) i_atm_cmp_cq_par_gen (                                   // Subtract out the qe_wt parity
          .d            ( {   atm_cmp_fifo_pop_data_cq_wt_p
                            , atm_cmp_fifo_pop_data.qe_wt } )
        , .odd          ( 1'b0 )                                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( atm_cmp_fifo_pop_data_cq_p )
) ;

hqm_AW_parity_gen #( .WIDTH( 1 + 8 + 2 ) ) i_atm_cmp_qid_par_gen (              // Subtract out the cq and qe_wt parity
          .d            ( {  atm_cmp_fifo_pop_data.parity 
                            , { 1'b0, atm_cmp_fifo_pop_data.cq }
                            , atm_cmp_fifo_pop_data.qe_wt } )
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( atm_cmp_fifo_pop_data_qid_p )
) ;

assign lbi_inp_cmp_qidix_msb            = atm_cmp_fifo_pop_data.qidix_msb ;
assign lbi_inp_cmp_qidix                = atm_cmp_fifo_pop_data.qidix ;
assign lbi_inp_cmp_qpri                 = atm_cmp_fifo_pop_data.qpri ;
assign lbi_inp_cmp_fid                  = atm_cmp_fifo_pop_data.fid ;
assign lbi_inp_cmp_fid_p                = atm_cmp_fifo_pop_data.fid_p ;
assign lbi_inp_cmp_p                    = atm_cmp_fifo_pop_data.cmp_p ;
assign lbi_inp_cmp_hid                  = atm_cmp_fifo_pop_data.hid ;
assign lbi_inp_cmp_hid_p                = atm_cmp_fifo_pop_data.hid_p ;

always_comb begin
  atm_cmp_wait_for_ap_cmp_nxt           = atm_cmp_wait_for_ap_cmp_f ;
  if ( atm_cmp_fifo_pop & cfg_control_single_op_atm_cmp ) begin
    atm_cmp_wait_for_ap_cmp_nxt         = 1'b1 ;
  end
  else if ( ap_lsp_cmd_cmp ) begin
    atm_cmp_wait_for_ap_cmp_nxt         = 1'b0 ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    atm_cmp_wait_for_ap_cmp_f           <= 1'b0 ;
  end
  else begin
    atm_cmp_wait_for_ap_cmp_f           <= atm_cmp_wait_for_ap_cmp_nxt ;
  end
end // always
assign atm_cmp_fifo_single_op_hold      = cfg_control_single_op_atm_cmp & atm_cmp_wait_for_ap_cmp_f ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB CQ selection - ATM , NALB
//-----------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// CQ polling

// Signals derived from AP intf
assign ap_lsp_cq_qidix                  = { ap_lsp_cq , ap_lsp_qidix } ;
assign ap_lsp_cmpblast_v_hit            = ap_lsp_cmpblast_v & p0_lba_cmpblast_chkv_f [ ap_lsp_cq_qidix ] ;
assign ap_lsp_unblast_slst_v            = ap_lsp_cmd_v & ( ap_lsp_cmd == HQM_LSP_AP_LSP_CMD_SCH_SLIST ) ;
assign ap_lsp_unblast_rlst_v            = ap_lsp_cmd_v & ( ap_lsp_cmd == HQM_LSP_AP_LSP_CMD_SCH_RLIST ) ;
assign ap_lsp_unblast_cmpblast          = ap_lsp_cmd_v & ( ap_lsp_cmd == HQM_LSP_AP_LSP_CMD_SCH_SLIST ) & p0_lba_cmpblast_chkv_f [ ap_lsp_cq_qidix ] ;
assign ap_lsp_cmd_cmp                   = ap_lsp_cmd_v & ( ap_lsp_cmd == HQM_LSP_AP_LSP_CMD_CMP ) ;

always_comb begin
  //---------------------------------------------------------------------------------------------------
  // valid vectors indicate that the corresponding traffic type has work to do for the indicated cq/qidix pair
  // All ldb vectors should be correctly adjusted as part of a successful vas reset drain

  // haswork_slst_v indicates whether or not AP has a cqidix on the scheduled list that is ready to be scheduled.
  p0_lba_slist_v_nxt                    =  p0_lba_slist_v_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( ap_lsp_haswork_slst_v & ( ap_lsp_cq_qidix == i ) ) begin
      p0_lba_slist_v_nxt [i]            = ap_lsp_haswork_slst_func ;
    end
    if ( cfg_ldb_sched_control_slist_haswork_v & ( cfg_ldb_sched_control_cq_qidix == i ) ) begin
      p0_lba_slist_v_nxt [ i ]          = cfg_ldb_sched_control_value ;
    end
  end // for i

  // haswork_rlst_v indicates whether or not AP has a qid on the ready list that is ready to be scheduled.
  p0_lba_rlist_v_nxt                    = p0_lba_rlist_v_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( ap_lsp_haswork_rlst_v & ap_lsp_qid2cqqidix [i] ) begin
      p0_lba_rlist_v_nxt [ i ]          = ap_lsp_haswork_rlst_func ;
    end
    if ( cfg_ldb_sched_control_rlist_haswork_v & ( cfg_ldb_sched_control_cq_qidix == i ) ) begin
      p0_lba_rlist_v_nxt [ i ]          = cfg_ldb_sched_control_value ;
    end
  end // for i

  // nalb_v indicates that LSP has a cqidix ready to be scheduled.
  p0_lba_nalb_v_nxt                     = p0_lba_nalb_v_f ;
  if ( p8_lba_qidix_if_v_upd_f | p8_lba_qidix_sch_v_upd_f )
    p0_lba_nalb_v_nxt                   = p8_lba_qidix_has_work ;

  //---------------------------------------------------------------------------------------------------
  // blast vectors prevent the arbiter from looking at the corresponding "has work"/valid vector during
  // the time that it is out of date - from the time the schedule starts (after qid2cqidix lookup) to
  // when LSP/AP updates the corresponding "has work" / valid.
  //
  // For ap_cmpblast, need to conditionally set the cmpblast when indicated by AP.  Do the cmpblast
  // if the slist blast bit is on, or if there is a sched in the pipe for the same {cq,qidix}.  If there
  // is a sched in the pipe, accumulate the cmpblasts that occur while it is in the pipe (match the cq),
  // then when the sched gets to p7 see if the selected qidix got cmpblasted, and if so, do the cmpblast.
  // cmpblasts must be accumulated in the pipe even if the pipe is holding.
  // cmpblast bits are cleared when an slist schedule update comes in from AP.
  p0_lba_slist_blast_nxt                = p0_lba_slist_blast_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( ap_lsp_unblast_slst_v & ap_lsp_qid2cqqidix [i] )
      p0_lba_slist_blast_nxt [i]        = 1'b0 ;
    if ( p7_lba_blast_slist & p7_lba_blast_qid2cqidix_v [i] )
      p0_lba_slist_blast_nxt [i]        = 1'b1 ;
  end // for i

  // cmpblast_chkv is set/cleared similar to slist_blast, but only the specific cq,qidix bit
  p7_lba_ctrl_pipe_sch_cq_qidix = p7_lba_ctrl_pipe_f_pcm ? { p7_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , p7_lba_ctrl_pipe_f.sch_qidix_msb , p7_lba_ctrl_pipe_f.sch_qidix } :
                                                           { p7_lba_ctrl_pipe_f.sch_cq , p7_lba_ctrl_pipe_f.sch_qidix } ;
  p0_lba_cmpblast_chkv_nxt              = p0_lba_cmpblast_chkv_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( ap_lsp_unblast_cmpblast & ( ap_lsp_cq_qidix == i ) )
      p0_lba_cmpblast_chkv_nxt [i]      = 1'b0 ;
    if ( p7_lba_blast_slist & ( { p7_lba_ctrl_pipe_sch_cq_qidix } == i ) )
      p0_lba_cmpblast_chkv_nxt [i]      = 1'b1 ;
  end // for i

  p0_lba_rlist_blast_nxt                = p0_lba_rlist_blast_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( ap_lsp_unblast_rlst_v & ap_lsp_qid2cqqidix [i] )
      p0_lba_rlist_blast_nxt [i]        = 1'b0 ;
    if ( p7_lba_blast_rlist & p7_lba_blast_qid2cqidix_v [i] )
      p0_lba_rlist_blast_nxt [i]        = 1'b1 ;
  end // for i

  p0_lba_nalb_blast_nxt                 = p0_lba_nalb_blast_f ;
  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( p8_lba_ctrl_pipe_v_f & p8_lba_blast_qid2cqidix_v_f [i] & p8_lba_ctrl_pipe_f.sch_nalb_v )
      p0_lba_nalb_blast_nxt [i]         = 1'b0 ;
    if ( p7_lba_blast_nalb & p7_lba_blast_qid2cqidix_v [i] )
      p0_lba_nalb_blast_nxt [i]         = 1'b1 ;
  end // for i

  p0_lba_cmpblast_nxt                   = p0_lba_cmpblast_f ;
  if ( ap_lsp_unblast_cmpblast | ap_lsp_cmpblast_v_hit | p7_lba_set_cmpblast ) begin
    for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
      if ( ap_lsp_unblast_cmpblast & ap_lsp_qid2cqqidix [i] )
        p0_lba_cmpblast_nxt [i]         = 1'b0 ;
      if ( ap_lsp_cmpblast_v_hit & ap_lsp_qid2cqqidix [i] )
        p0_lba_cmpblast_nxt [i]         = 1'b1 ;
      if ( p7_lba_set_cmpblast & p7_lba_blast_qid2cqidix_v [i] )
        p0_lba_cmpblast_nxt [i]         = 1'b1 ;
    end // for i
  end // if

  p0_lba_cmpblast_ap_rst_v_nxt          = ap_lsp_unblast_cmpblast ;
  p0_lba_cmpblast_ap_val_nxt            = p0_lba_cmpblast_chkv_f [ ap_lsp_cq_qidix ] ;
  p0_lba_cmpblast_lsp_set_v_nxt         = p7_lba_blast_slist ;
  p0_lba_cmpblast_lsp_val_nxt           = p0_lba_cmpblast_chkv_f [ p7_lba_ctrl_pipe_sch_cq_qidix ] ;

  //---------------------------------------------------------------------------------------------------
  // lba_cq_has_space indicates that the given cq still has space - satisfies the per-CQ token count,
  // cq-inflight count and total-inflight count checks.  Since the CQs are shared between nalb and ATM
  // the total count and checks include both types.  ATM schedules and token returns must also go down
  // the nalb pipe to support this shared checking.
  p0_lba_cq_has_space_nxt               = p0_lba_cq_has_space_f ;
  if ( p8_lba_cq_if_v_upd_f | p8_lba_cq_tok_v_upd_f | cfgsc_cq_ldb_token_count_mem_we ) begin
    p0_lba_cq_has_space_nxt             = p8_lba_cq_has_space ;
    for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
      if ( cfg_cq_ldb_enable_pcm_f [ i ] & ( ( i & 32'h1 ) == 'h1 ) ) begin
        p0_lba_cq_has_space_nxt [i]     = p0_lba_cq_has_space_nxt [ i - 1 ] ;
      end
      if ( cfgsc_cq_ldb_token_count_mem_we & ( cfg_mem_addr [HQM_NUM_LB_CQB2-1:0] == i ) ) begin        // Should only be done as part of vas reset or cq configuration
        p0_lba_cq_has_space_nxt [i]     = 1'b1 ;
      end
    end // for i
  end // if

  //---------------------------------------------------------------------------------------------------
  // lba_cq_ow indicates that the amount of work scheduled to a given cq is over its configured limit.
  p0_lba_cq_ow_nxt                      = p0_lba_cq_ow_f ;
  if ( p4_lbwu_cq_wu_cnt_upd_v_f | cfgsc_cq_ldb_token_count_mem_we ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
      if ( p4_lbwu_cq_wu_cnt_upd_v_f & ( p4_lbwu_cq_wu_cnt_upd_cq_f == i ) ) begin
        p0_lba_cq_ow_nxt [i]            = p4_lbwu_cq_wu_cnt_upd_gt_lim_f ;
      end
    end // for i

    for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
      if ( cfgsc_cq_ldb_token_count_mem_we & ( cfg_mem_addr [HQM_NUM_LB_CQB2-1:0] == i ) ) begin        // Should only be done as part of vas reset or cq configuration
        p0_lba_cq_ow_nxt [i]            = 1'b0 ;
      end
      if ( cfg_cq_ldb_enable_pcm_f [ i ] & ( ( i & 32'h1 ) == 'h1 ) ) begin
        p0_lba_cq_ow_nxt [i]            = p0_lba_cq_ow_nxt [ i - 1 ] ;
      end
    end // for i
  end // if

  //---------------------------------------------------------------------------------------------------
  // Need ability to limit atomic inflight on a per-qid basis like nalb; separate register to ease PD concerns.
  // On 1 -> 0 transition (sch) qidix should already be blasted so 1 clock delay should not matter.
  // On 0 -> 1 transition (cmp) qidix will be eligible 1 clock later.
  p0_lba_atm_if_v_nxt                   = p0_lba_atm_if_v_f;
  if ( p8_lba_qidix_if_v_upd_f ) begin
    p0_lba_atm_if_v_nxt                 = p8_lba_qidix_if_v_f ;
  end

  //---------------------------------------------------------------------------------------------------
  // lba_cq_busy_sch indicates that the given cq has a scheduling operation (nalb or ATM) active in
  // the LSP pipe.  This prevents the CQ from being prematurely scheduled again before the per-CQ
  // token and inflight statuses have been updated with their correct values from the bottom of the pipe.
  p0_lba_cq_busy_sch_nxt                = p0_lba_cq_busy_sch_f ;
  if ( p8_lba_ctrl_pipe_v_f | p1_lba_issue_sched ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
      if ( p8_lba_ctrl_pipe_v_f & p8_lba_ctrl_pipe_f.sch_v & ( p8_lba_ctrl_pipe_f.sch_cq == i ) ) begin
        p0_lba_cq_busy_sch_nxt [i]        = 1'b0 ;
        if ( cfg_cq_ldb_enable_pcm_f [ i ] | ( ~ ( ( i & 32'h1 ) == 'h1 ) & cfg_cq_ldb_enable_pcm_f [ i + 1 ] ) ) begin
          if ( ( i & 32'h1 ) == 'h1 ) begin
            p0_lba_cq_busy_sch_nxt [ i - 1 ]  = 1'b0 ;
          end
          else begin
            p0_lba_cq_busy_sch_nxt [ i + 1 ]  = 1'b0 ;
          end
        end
      end
      if ( p1_lba_issue_sched & ( p1_lba_ctrl_pipe_f.sch_cq == i ) ) begin      // Since cq vectors aren't looked at until state machine is beyond
        p0_lba_cq_busy_sch_nxt [i]        = 1'b1 ;                              // issue_sched, OK to wait and use p1 cq for delay reasons.
        if ( cfg_cq_ldb_enable_pcm_f [ i ] | ( ~ ( ( i & 32'h1 ) == 'h1 ) & cfg_cq_ldb_enable_pcm_f [ i + 1 ] ) ) begin
          if ( ( i & 32'h1 ) == 'h1 ) begin
            p0_lba_cq_busy_sch_nxt [ i - 1 ]  = 1'b1 ; 
          end
          else begin
            p0_lba_cq_busy_sch_nxt [ i + 1 ]  = 1'b1 ; 
          end
        end
      end
    end // for i
  end // if

end // always

always_comb begin
  ap_lsp_qidixv                         = 16'h0 ;                       //JTC
  ap_lsp_qidixv [ { ap_lsp_qidix_msb , ap_lsp_qidix } ]        = 1'b1 ;
end

// If pop does not occur then OK to not blast; p0 state will be updated by ap_lsp for next clock(s)
assign p0_lba_ctrl_pipe_cmpblast_cond   = p0_lba_pop_cq [0]                               & ap_lsp_cmpblast_v &
                                          ( p1_lba_ctrl_pipe_f_pcm_nxt ?
                                            ( p1_lba_ctrl_pipe_nxt.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p1_lba_ctrl_pipe_nxt.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) ) ;
assign p1_lba_ctrl_pipe_cmpblast_cond   = p1_lba_ctrl_pipe_v_f & p1_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p1_lba_ctrl_pipe_f_pcm ?
                                            ( p1_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p1_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p2_lba_ctrl_pipe_cmpblast_cond   = p2_lba_ctrl_pipe_v_f & p2_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p2_lba_ctrl_pipe_f_pcm ?
                                            ( p2_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p2_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p3_lba_ctrl_pipe_cmpblast_cond   = p3_lba_ctrl_pipe_v_f & p3_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p3_lba_ctrl_pipe_f_pcm ?
                                            ( p3_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p3_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p4_lba_ctrl_pipe_cmpblast_cond   = p4_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p4_lba_ctrl_pipe_f_pcm ?
                                            ( p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p5_lba_ctrl_pipe_cmpblast_cond   = p5_lba_ctrl_pipe_v_f & p5_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p5_lba_ctrl_pipe_f_pcm ?
                                            ( p5_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p5_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p6_lba_ctrl_pipe_cmpblast_cond   = p6_lba_ctrl_pipe_v_f & p6_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p6_lba_ctrl_pipe_f_pcm ?
                                            ( p6_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p6_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;
assign p7_lba_ctrl_pipe_cmpblast_cond   = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.sch_v & ap_lsp_cmpblast_v &
                                          ( p7_lba_ctrl_pipe_f_pcm ?
                                            ( p7_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] ) :
                                            ( p7_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] == ap_lsp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ) ) ;

assign p0_lba_sch_cmpblast_qidixv_blasted       =                                          ap_lsp_qidixv ;              //JTC
assign p1_lba_sch_cmpblast_qidixv_blasted       = p1_lba_sch_cmpblast_qidixv_f           | ap_lsp_qidixv ;
assign p2_lba_sch_cmpblast_qidixv_blasted       = p2_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;
assign p3_lba_sch_cmpblast_qidixv_blasted       = p3_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;
assign p4_lba_sch_cmpblast_qidixv_blasted       = p4_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;
assign p5_lba_sch_cmpblast_qidixv_blasted       = p5_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;
assign p6_lba_sch_cmpblast_qidixv_blasted       = p6_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;
assign p7_lba_sch_cmpblast_qidixv_blasted       = p7_lba_ctrl_pipe_f.sch_cmpblast_qidixv | ap_lsp_qidixv ;

assign p1_lba_ctrl_pipe_f_pcm_nxt = (p1_lba_ctrl_pipe.en & 
                                    ( p0_lba_arb_sch_v | p0_lba_arb_cq_cmp_v )) ? cfg_cq_ldb_enable_pcm_f [ (p0_lba_arb_sch_v) ? p0_lba_cq_arb_winner : lbi_inp_cq_cmp_cq ] : p1_lba_ctrl_pipe_f_pcm ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p0_lba_sch_state_f          <= HQM_LSP_LBA_ARB_STATE_WAIT_FOR_WORK ;
    p1_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p2_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p3_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p4_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p5_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p6_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p7_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
    p8_lba_ctrl_pipe_f_pcm	<= 1'b0 ;
  end
  else begin
    p0_lba_sch_state_f          <= p0_lba_sch_state_nxt ;
    p1_lba_ctrl_pipe_f_pcm	<= p1_lba_ctrl_pipe_f_pcm_nxt ;
    p2_lba_ctrl_pipe_f_pcm	<= p2_lba_ctrl_pipe.en ? p1_lba_ctrl_pipe_f_pcm : p2_lba_ctrl_pipe_f_pcm ;
    p3_lba_ctrl_pipe_f_pcm	<= p3_lba_ctrl_pipe.en ? p2_lba_ctrl_pipe_f_pcm : p3_lba_ctrl_pipe_f_pcm ;
    p4_lba_ctrl_pipe_f_pcm	<= p4_lba_ctrl_pipe.en ? p3_lba_ctrl_pipe_f_pcm : p4_lba_ctrl_pipe_f_pcm ;
    p5_lba_ctrl_pipe_f_pcm	<= p5_lba_ctrl_pipe.en ? p4_lba_ctrl_pipe_f_pcm : p5_lba_ctrl_pipe_f_pcm ;
    p6_lba_ctrl_pipe_f_pcm	<= p6_lba_ctrl_pipe.en ? p5_lba_ctrl_pipe_f_pcm : p6_lba_ctrl_pipe_f_pcm ;
    p7_lba_ctrl_pipe_f_pcm	<= p7_lba_ctrl_pipe.en ? p6_lba_ctrl_pipe_f_pcm : p7_lba_ctrl_pipe_f_pcm ;
    p8_lba_ctrl_pipe_f_pcm	<= p8_lba_ctrl_pipe.en ? p7_lba_ctrl_pipe_f_pcm : p8_lba_ctrl_pipe_f_pcm ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p0_lba_slist_v_f            <= 512'h0 ;
    p0_lba_rlist_v_f            <= 512'h0 ;
    p0_lba_nalb_v_f             <= 512'h0 ;
    p0_lba_slist_blast_f        <= 512'h0 ;
    p0_lba_rlist_blast_f        <= 512'h0 ;
    p0_lba_nalb_blast_f         <= 512'h0 ;
    p0_lba_cmpblast_chkv_f      <= 512'h0 ;
    p0_lba_cmpblast_f           <= 512'h0 ;
    p0_lba_atm_if_v_f           <= { 512 { 1'b1 } } ;
    p0_lba_cq_has_space_f       <= { HQM_NUM_LB_CQ { 1'b1 } } ;
    p0_lba_cq_busy_sch_f        <= { HQM_NUM_LB_CQ { 1'b0 } } ;
    p0_lba_cq_ow_f              <= { HQM_NUM_LB_CQ { 1'b0 } } ;
    p0_lba_cmpblast_ap_val_f    <= 1'b0 ;
    p0_lba_cmpblast_ap_rst_v_f  <= 1'b0 ;
    p0_lba_cmpblast_lsp_set_v_f <= 1'b0 ;
    p0_lba_cmpblast_lsp_val_f   <= 1'b0 ;

    p1_lba_sch_slist_v_f        <= 512'h0 ;
    p1_lba_sch_rlist_v_f        <= 512'h0 ;
    p1_lba_sch_nalb_v_f         <= 512'h0 ;
    p1_lba_sch_cmpblast_qidixv_f        <= 16'h0 ;

    p1_lba_ctrl_pipe_v_f        <= 1'b0 ;
    p2_lba_ctrl_pipe_v_f        <= 1'b0 ;
    p3_lba_ctrl_pipe_v_f        <= 1'b0 ;
    p4_lba_ctrl_pipe_v_f        <= 1'b0 ;
  end
  else begin
    p0_lba_slist_v_f            <= p0_lba_slist_v_nxt ;
    p0_lba_rlist_v_f            <= p0_lba_rlist_v_nxt ;
    p0_lba_nalb_v_f             <= p0_lba_nalb_v_nxt ;
    p0_lba_slist_blast_f        <= p0_lba_slist_blast_nxt ;
    p0_lba_rlist_blast_f        <= p0_lba_rlist_blast_nxt ;
    p0_lba_nalb_blast_f         <= p0_lba_nalb_blast_nxt ;
    p0_lba_cmpblast_chkv_f      <= p0_lba_cmpblast_chkv_nxt ;
    p0_lba_cmpblast_f           <= p0_lba_cmpblast_nxt ;
    p0_lba_atm_if_v_f           <= p0_lba_atm_if_v_nxt ;
    p0_lba_cq_has_space_f       <= p0_lba_cq_has_space_nxt ;
    p0_lba_cq_busy_sch_f        <= p0_lba_cq_busy_sch_nxt ;
    p0_lba_cq_ow_f              <= p0_lba_cq_ow_nxt ;
    p0_lba_cmpblast_ap_val_f    <= p0_lba_cmpblast_ap_val_nxt ;
    p0_lba_cmpblast_ap_rst_v_f  <= p0_lba_cmpblast_ap_rst_v_nxt ;
    p0_lba_cmpblast_lsp_set_v_f <= p0_lba_cmpblast_lsp_set_v_nxt ;
    p0_lba_cmpblast_lsp_val_f   <= p0_lba_cmpblast_lsp_val_nxt ;

    p1_lba_sch_slist_v_f        <= p1_lba_sch_slist_v_nxt ;
    p1_lba_sch_rlist_v_f        <= p1_lba_sch_rlist_v_nxt ;
    p1_lba_sch_nalb_v_f         <= p1_lba_sch_nalb_v_nxt ;
    p1_lba_sch_cmpblast_qidixv_f        <= p1_lba_sch_cmpblast_qidixv_nxt ;

    p1_lba_ctrl_pipe_v_f        <= p1_lba_ctrl_pipe_v_nxt ;
    p2_lba_ctrl_pipe_v_f        <= p2_lba_ctrl_pipe_v_nxt ;
    p3_lba_ctrl_pipe_v_f        <= p3_lba_ctrl_pipe_v_nxt ;
    p4_lba_ctrl_pipe_v_f        <= p4_lba_ctrl_pipe_v_nxt ;
  end
end // always

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
    p1_lba_sch_slist_v_ar [i]   = p1_lba_sch_slist_v_f [ ( i * HQM_QID_PER_CQ ) +: HQM_QID_PER_CQ ] ;             //JTC
    p1_lba_sch_rlist_v_ar [i]   = p1_lba_sch_rlist_v_f [ ( i * HQM_QID_PER_CQ ) +: HQM_QID_PER_CQ ] ;             //JTC
    p1_lba_sch_nalb_v_ar [i]    = p1_lba_sch_nalb_v_f [ ( i * HQM_QID_PER_CQ ) +: HQM_QID_PER_CQ ] ;              //JTC
  end // for
end // always

assign p0_lba_cmpblast_ap_rst_err       = p0_lba_cmpblast_ap_rst_v_f  & ~ p0_lba_cmpblast_ap_val_f ;
assign p0_lba_cmpblast_lsp_set_err      = p0_lba_cmpblast_lsp_set_v_f & p0_lba_cmpblast_lsp_val_f ;

//-----------------------------------------------------------------------------------------------------
// Create the per-CQ vectors for arbitration

// All types of scheduling must be supressed for a CQ which does not have space; space is shared.
// For cqidix vectors OK to just OR all 8 bits; individual ix will be selected below by looking at
// individual bits.

// A given CQ is eligible if any of its 8 qidix's has v=1 and blast=0.
// For slist, depending on mode bit, for a given CQ, if any of its 8 blast bits are 1, that CQ is ineligible.           //JTC

hqm_lsp_cq_sel # (
  .HQM_NUM_LB_CQ ( HQM_NUM_LB_CQ )
, .HQM_QID_PER_CQ ( HQM_QID_PER_CQ )
) i_hqm_lsp_cq_sel_p0 (            //JTC
          .cfg_control_atm_cq_qid_priority_prot         ( cfg_control_atm_cq_qid_priority_prot )
        , .cfg_cq_ldb_disable_f                         ( cfg_cq_ldb_disable_f | core_chp_lsp_ldb_cq_off_f )
        , .slist_v                                      ( p0_lba_slist_v_f )
        , .rlist_v                                      ( p0_lba_rlist_v_f )
        , .nalb_v                                       ( p0_lba_nalb_v_f )
        , .slist_blast                                  ( p0_lba_slist_blast_f )
        , .rlist_blast                                  ( p0_lba_rlist_blast_f )
        , .nalb_blast                                   ( p0_lba_nalb_blast_f )
        , .cmpblast                                     ( p0_lba_cmpblast_f )
        , .atm_if_v                                     ( p0_lba_atm_if_v_f )
        , .cq_has_space                                 ( p0_lba_cq_has_space_f )
        , .cq_busy_sch                                  ( p0_lba_cq_busy_sch_f )
        , .cq_ow                                        ( p0_lba_cq_ow_f )

        , .slist_v_blasted                              ( p0_lba_slist_v_blasted )
        , .rlist_v_blasted                              ( p0_lba_rlist_v_blasted )
        , .nalb_v_blasted                               ( p0_lba_nalb_v_blasted )
        , .slist_has_work                               ( p0_lba_cq_arb_slist_has_work_nc )
        , .rlist_has_work                               ( p0_lba_cq_arb_rlist_has_work_nc )
        , .nalb_has_work                                ( p0_lba_cq_arb_nalb_has_work_nc )
        , .any_has_work                                 ( p0_lba_cq_arb_any_has_work )
        , .cq_arb_reqs                                  ( p0_lba_cq_arb_reqs )
) ;

//*******************************************************************************************************************************************
// Note: since there is a 1-clock delay for the arbiter to produce a valid output, but the rest of the pipe requires (for functional and
// performance reasons) that the output be valid as if there were no latency, the reqs must be derived from the "next" inputs to the
// p0 registers.  Potential static timing / PD issues, but most/all signals are at most a couple of levels removed from
// flop outputs.

// Note: It is possible that cfg_cq_ldb_disable could be changed while there is live traffic because of vas reset.  It doesn't matter on
// exactly which clock the arbiter reacts to such a change, but it does matter that the two instances of hqm_lsp_cq_sel react to it
// consisistently, so theoretically should be using a "nxt" version of cfg_cq_ldb_disable here.  However, it's OK because the only arbiter
// output which cfg_cq_ldb_disabled factors into is cq_arb_reqs, and that is not connected on the one instance, so could actually just wire
// up a constant to the cfg_cq_ldb_disable_f input of that instance and it wouldn't matter.

hqm_lsp_cq_sel #(
  .HQM_NUM_LB_CQ ( HQM_NUM_LB_CQ )
, .HQM_QID_PER_CQ ( HQM_QID_PER_CQ )
) i_hqm_lsp_cq_sel_p0_nxt (                //JTC
          .cfg_control_atm_cq_qid_priority_prot         ( cfg_control_atm_cq_qid_priority_prot )
        , .cfg_cq_ldb_disable_f                         ( cfg_cq_ldb_disable_f | core_chp_lsp_ldb_cq_off_f )
        , .slist_v                                      ( p0_lba_slist_v_nxt )
        , .rlist_v                                      ( p0_lba_rlist_v_nxt )
        , .nalb_v                                       ( p0_lba_nalb_v_nxt )
        , .slist_blast                                  ( p0_lba_slist_blast_nxt )
        , .rlist_blast                                  ( p0_lba_rlist_blast_nxt )
        , .nalb_blast                                   ( p0_lba_nalb_blast_nxt )
        , .cmpblast                                     ( p0_lba_cmpblast_nxt )
        , .atm_if_v                                     ( p0_lba_atm_if_v_nxt )
        , .cq_has_space                                 ( p0_lba_cq_has_space_nxt )
        , .cq_busy_sch                                  ( p0_lba_cq_busy_sch_nxt )
        , .cq_ow                                        ( p0_lba_cq_ow_nxt )

        , .slist_v_blasted                              ( p0_nxt_lba_slist_v_blasted_nc )
        , .rlist_v_blasted                              ( p0_nxt_lba_rlist_v_blasted_nc )
        , .nalb_v_blasted                               ( p0_nxt_lba_nalb_v_blasted_nc )
        , .slist_has_work                               ( p0_nxt_lba_cq_arb_slist_has_work_nc )
        , .rlist_has_work                               ( p0_nxt_lba_cq_arb_rlist_has_work_nc )
        , .nalb_has_work                                ( p0_nxt_lba_cq_arb_nalb_has_work_nc )
        , .any_has_work                                 ( p0_nxt_lba_cq_arb_any_has_work_nc )
        , .cq_arb_reqs                                  ( p0_nxt_lba_cq_arb_reqs )
) ;

//*******************************************************************************************************************************************

assign p0_lba_cq_arb_update             = p0_lba_pop_cq [5] ;

// Note: there is a 1-clock latency inside the arbiter such that when an update occurs, on the next clock
// the output valid is stale.  This should not be an issue since the p0_lba_arb state machine should not
// even look at the schedule requests until the prior schedule/update has made it down to p7.  So there
// should be no need to explicitly mask the arbiter valid output during this "stale clock".

hqm_lsp_cq_cos_arb # (
          .NUM_REQS                     ( HQM_NUM_LB_CQ )
        , .NUM_COS                      ( 4 )
        , .NUM_VAL                      ( HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR )
        , .CNT_WIDTH                    ( 16 )
        , .WEIGHT_WIDTH                 ( 8 )
        , .STARV_AVOID_THRESH_WIDTH     ( 10 )
) i_lba_cq_cos_arb (
          .clk                          ( hqm_gated_clk )
        , .rst_n                        ( hqm_gated_rst_n )

        , .cfg_range                    ( { cfg_range_cos3_f       , cfg_range_cos2_f       , cfg_range_cos1_f       , cfg_range_cos0_f } )
        , .cfg_range_reconfig           ( cfg_range_reconfig )
        , .cfg_credit_sat               ( { cfg_credit_sat_cos3_f  , cfg_credit_sat_cos2_f  , cfg_credit_sat_cos1_f  , cfg_credit_sat_cos0_f } )
        , .cfg_no_extra_credit          ( { cfg_no_extra_credit3_f , cfg_no_extra_credit2_f , cfg_no_extra_credit1_f , cfg_no_extra_credit0_f } )
        , .cfg_starv_avoid_enable       ( cfg_starv_avoid_enable_f )
        , .cfg_starv_avoid_thresh_min   ( cfg_starv_avoid_thresh_min_f )
        , .cfg_starv_avoid_thresh_max   ( cfg_starv_avoid_thresh_max_f )
        , .cfg_credit_cnt               ( { cfg_credit_cnt_cos3    , cfg_credit_cnt_cos2    , cfg_credit_cnt_cos1    , cfg_credit_cnt_cos0   } )
        , .cfg_starv_avoid_cnt          ( { cfg_starv_avoid_cnt_cos3  , cfg_starv_avoid_cnt_cos2  , cfg_starv_avoid_cnt_cos1  , cfg_starv_avoid_cnt_cos0 } )
        , .cfg_schd_cos                 ( cfg_schd_cos )
        , .cfg_rdy_cos                  ( cfg_rdy_cos )
        , .cfg_rnd_loss_cos             ( cfg_rnd_loss_cos )
        , .cfg_cnt_win_cos              ( cfg_cnt_win_cos )

        , .reqs                         ( p0_nxt_lba_cq_arb_reqs )
        , .update                       ( p0_lba_cq_arb_update )
        , .winner_v                     ( p0_lba_cq_arb_winner_pre_v )
        , .winner                       ( p0_lba_cq_arb_winner )
        , .arb_error_f                  ( p0_lba_cq_arb_error_f )
        , .arb_status                   ( p0_lba_cq_arb_status )
) ;

//-----------------------------------------------------------------------------------------------------------------
// If cause_pipe_idle, don't introduce new schedules into the pipe; additional work may accumulate while idle (e.g. from AP)
assign p0_lba_cq_arb_winner_v           = p0_lba_cq_arb_winner_pre_v & { { HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR } { ~ cause_pipe_idle } } ;

// Required performance if different qid is 1/8 clocks.  LSP turns on the blast bit from p7 so scheduling to the same qid must wait until
// the update comes from either the bottom of the LSP pipe (9 clocks) or ATM pipe (13 clocks).
// p0_lba_pop_cq        : sch advances from p0 to p1
// p1_lba_issue_sched   : sch advances from p1 to p2
always_comb begin
  p0_lba_sch_state_nxt                          = p0_lba_sch_state_f ;
  p0_lba_pop_cq                                 = { HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR { 1'b0 } } ;
  p0_lba_sch_state_ready_for_work               = 1'b0 ;
  p1_lba_issue_sched_cond                       = 1'b0 ;
  
  case ( p0_lba_sch_state_f )
    HQM_LSP_LBA_ARB_STATE_WAIT_FOR_WORK : begin
      p0_lba_sch_state_ready_for_work           = 1'b1 ;
      if ( p0_lba_cq_arb_winner_v [0] & ~ p1_lba_ctrl_pipe.hold & ~ p0_lba_ctrl_pipe_sch_hold_cond & ~ cause_pipe_idle &
           p0_lba_sch_state_ready_for_work & ~ p0_lba_restrict_bw_hold_cond ) begin
        p0_lba_sch_state_nxt                    = HQM_LSP_LBA_ARB_STATE_SCHED ;
      end
      p0_lba_pop_cq                             = p0_lba_cq_arb_winner_v &
                                                  { HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR {
                                                      ~ p1_lba_ctrl_pipe.hold & ~ p0_lba_ctrl_pipe_sch_hold_cond &
                                                      ~ cause_pipe_idle & p0_lba_sch_state_ready_for_work & ~ p0_lba_restrict_bw_hold_cond } } ;
    end
    HQM_LSP_LBA_ARB_STATE_SCHED : begin
      if ( ~ p1_lba_ctrl_pipe.hold ) begin
        p0_lba_sch_state_nxt                    = HQM_LSP_LBA_ARB_STATE_WAIT_FOR_BLAST ;
      end
      p1_lba_issue_sched_cond                   = 1'b1 ;
    end
    HQM_LSP_LBA_ARB_STATE_WAIT_FOR_BLAST : begin
      if ( ( ~ cfg_control_single_op_atm_sched &       p7_lba_sched ) |
           (   cfg_control_single_op_atm_sched & ( ( ( p7_lba_sched & ~ p7_lba_ctrl_pipe_f.sch_atm_v ) | ap_lsp_unblast_slst_v | ap_lsp_unblast_rlst_v ) ) ) ) begin
        p0_lba_sch_state_nxt                    = HQM_LSP_LBA_ARB_STATE_WAIT_FOR_WORK ;
      end
    end
    default : begin                     // Same as default assigns above
      p0_lba_sch_state_nxt                      = p0_lba_sch_state_f ;
      p0_lba_pop_cq                             = { HQM_LSP_LBA_CQ_ARB_V_DUP_FACTOR { 1'b0 } } ;
      p0_lba_sch_state_ready_for_work           = 1'b0 ;
      p1_lba_issue_sched_cond                   = 1'b0 ;
    end
  endcase
end // always

assign p1_lba_issue_sched       = p1_lba_issue_sched_cond & ~ p1_lba_ctrl_pipe.hold ;

// p1_lba_sch registers are solely for scheduling info.  If a schedule is
// not selected to move on to p2, they hold.  When a particular CQ arbiter is selected, its
// state is updated as it loads into p1 - we are committed to scheduling that CQ.  It is not possible
// for a CQ to be good for scheduling when it is selected and then go "not good" while it is holding
// in p1.  The has_space bit should have set as it went in to p0, and anything in flight in the lba
// pipe should have been protected by has_space so there should not be any updates in flight that could
// "subtract" from the CQs ability to be scheduled to.
// The p1 sch_cmpblast_qidixv needs to be handled differently than the other pipe levels, because in
// cases where p1 is not holding, but is also not actively popping a CQ, it still needs to do blast
// checking.  So need a dedicated register and control separate from the main pipeline.

always_comb begin
  p1_lba_sch_slist_v_nxt                = p1_lba_sch_slist_v_f ;
  p1_lba_sch_rlist_v_nxt                = p1_lba_sch_rlist_v_f ;
  p1_lba_sch_nalb_v_nxt                 = p1_lba_sch_nalb_v_f ;
  p1_lba_sch_cmpblast_qidixv_nxt        = p1_lba_sch_cmpblast_qidixv_f ;

  if ( p0_lba_pop_cq [0] ) begin    // If state allows pop, p1 sch state registers are available
    if ( p0_lba_ctrl_pipe_cmpblast_cond )
      p1_lba_sch_cmpblast_qidixv_nxt    = p0_lba_sch_cmpblast_qidixv_blasted ;
    else
      p1_lba_sch_cmpblast_qidixv_nxt    = 16'h0 ;
  end
  else begin
    if ( p1_lba_issue_sched ) begin
      p1_lba_sch_cmpblast_qidixv_nxt    = 16'h0 ;
    end
    else begin
      if ( p1_lba_ctrl_pipe_cmpblast_cond ) begin
        p1_lba_sch_cmpblast_qidixv_nxt  = p1_lba_sch_cmpblast_qidixv_blasted ;
      end
    end
  end
  if ( p0_lba_pop_cq [1] ) begin                // If state allows pop, p1 sch state registers are available
    p1_lba_sch_slist_v_nxt              = p0_lba_slist_v_blasted ;
  end
  if ( p0_lba_pop_cq [2] ) begin                // If state allows pop, p1 sch state registers are available
    p1_lba_sch_rlist_v_nxt              = p0_lba_rlist_v_blasted ;
  end
  if ( p0_lba_pop_cq [3] ) begin                // If state allows pop, p1 sch state registers are available
    p1_lba_sch_nalb_v_nxt               = p0_lba_nalb_v_blasted ;
  end
end // always

hqm_AW_parity_gen #( .WIDTH( HQM_NUM_LB_CQB2 ) ) i_lba_sch_cq_par_gen (
          .d            ( p0_lba_cq_arb_winner )                // If delay issue could be done at next pipe level
        , .odd          ( 1'b1 )
        , .p            ( p0_lba_cq_gp )
) ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB Input Request arbitration
//-----------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// Enqueue

assign enq_nalb_fifo_pop                = lbi_enq_req_taken ;

assign lbi_inp_enq_qid                  = enq_nalb_fifo_pop_data.qid ;
assign lbi_inp_enq_qid_p                = enq_nalb_fifo_pop_data.parity ^ ( ^ ( enq_nalb_fifo_pop_data.qtype ) ) ;      // subtract out qtype parity

assign lbi_enq_req_taken                = p0_lba_arb_enq_v & ~ p1_lba_ctrl_pipe.hold ;

//-------------------------------------------------------------------------------------------------
// Token

assign ldb_token_rtn_fifo_pop           = lbi_tok_req_taken ;

assign lbi_inp_tok_cq                   = ldb_token_rtn_fifo_pop_data.cq [HQM_NUM_LB_CQB2-1:0] ;
assign lbi_inp_tok_cq_p                 = ldb_token_rtn_fifo_pop_data.parity ^ ldb_token_rtn_fifo_pop_data.is_ldb ;     // subtract out is_ldb parity

// If ms bits are (erroneously) on, force to a value guaranteed to be detected as underflow when subtracting
assign lbi_inp_tok_cnt_uflow_cond       = | ( ldb_token_rtn_fifo_pop_data.count [12:11] ) ;
assign lbi_inp_tok_cnt                  = { ( ldb_token_rtn_fifo_pop_data.count [10:9] | { 2 { lbi_inp_tok_cnt_uflow_cond } } ) ,
                                                ldb_token_rtn_fifo_pop_data.count [8:0]} ;
assign lbi_inp_tok_cnt_res              = ldb_token_rtn_fifo_pop_data.count_residue ;

assign lbi_tok_req_taken                = p0_lba_arb_tok_v & ~ p1_lba_ctrl_pipe.hold ;

//-------------------------------------------------------------------------------------------------
// QID completions

assign rop_lsp_reordercmp_fifo_pop_data_vreq    = core_rop_lsp_reordercmp_v & ~ cause_pipe_idle ;
assign rop_lsp_reordercmp_fifo_pop_data         = core_rop_lsp_reordercmp_data ;
assign core_rop_lsp_reordercmp_ready            = rop_lsp_reordercmp_fifo_pop ;

assign lbi_qid_cmp_arb_reqs [ HQM_LSP_LBA_QID_ARB_UNO_ATM ]     = uno_atm_cmp_fifo_pop_data_vreq ;              // include RELEASE
assign lbi_qid_cmp_arb_reqs [ HQM_LSP_LBA_QID_ARB_ORD ]         = rop_lsp_reordercmp_fifo_pop_data_vreq ;

hqm_AW_wrand_arb # ( .NUM_REQS ( 2 ) , .SEED ( 1 ) ) i_lbi_qid_cmp_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( lbi_qid_cmp_arb_reqs )
        , .cfg_weight           ( { cfg_lbi_qid_cmp_arb_weight_uno_atm ,                // Equal weights = random
                                    cfg_lbi_qid_cmp_arb_weight_ord } )
        , .winner_v             ( lbi_qid_cmp_arb_winner_v )
        , .winner               ( lbi_qid_cmp_arb_winner )
) ;

assign uno_atm_cmp_fifo_pop_data_qid_p  = uno_atm_cmp_fifo_pop_data.cq_qid_p ^ ( ^ uno_atm_cmp_fifo_pop_data.cq ) ;     // Subtract out the cq parity
assign rop_lsp_reordercmp_fifo_pop_data_qid_p   = rop_lsp_reordercmp_fifo_pop_data.parity ^ ( ^ rop_lsp_reordercmp_fifo_pop_data.cq ) ; // Subtract out the cq parity

always_comb begin
  uno_atm_cmp_fifo_pop                          = 1'b0 ;
  rop_lsp_reordercmp_fifo_pop                   = 1'b0 ;
  lbi_inp_qid_cmp_qid                           = uno_atm_cmp_fifo_pop_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  lbi_inp_qid_cmp_qid_p                         = uno_atm_cmp_fifo_pop_data_qid_p ;
  lbi_inp_qid_cmp_no_dec                        = ( ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b01 ) |
                                                    ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b11 ) ) ;
  lbi_inp_qid_cmp_dec_only                      = ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b10 ) ;
  case ( lbi_qid_cmp_arb_winner )
    HQM_LSP_LBA_QID_ARB_ORD : begin
      rop_lsp_reordercmp_fifo_pop               = lbi_qid_cmp_req_taken ;
      lbi_inp_qid_cmp_qid                       = rop_lsp_reordercmp_fifo_pop_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
      lbi_inp_qid_cmp_qid_p                     = rop_lsp_reordercmp_fifo_pop_data_qid_p ;
      lbi_inp_qid_cmp_no_dec                    = ( rop_lsp_reordercmp_fifo_pop_data.user == 1'b1 ) ;
      lbi_inp_qid_cmp_dec_only                  = 1'b0 ;
    end
    HQM_LSP_LBA_QID_ARB_UNO_ATM : begin
      uno_atm_cmp_fifo_pop                      = lbi_qid_cmp_req_taken ;
      lbi_inp_qid_cmp_qid                       = uno_atm_cmp_fifo_pop_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
      lbi_inp_qid_cmp_qid_p                     = uno_atm_cmp_fifo_pop_data_qid_p ;
      lbi_inp_qid_cmp_no_dec                    = ( ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b01 ) |
                                                    ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b11 ) ) ;
      lbi_inp_qid_cmp_dec_only                  = ( uno_atm_cmp_fifo_pop_data.user[1:0] == 2'b10 ) ;
    end
  endcase
end // always

assign lbi_qid_cmp_req_taken            = p0_lba_arb_qid_cmp_v & ~ p1_lba_ctrl_pipe.hold ;      // includes RELEASE

//-------------------------------------------------------------------------------------------------
// Enqueue vs. QID Completion arbiter
// Requests are not compatible since both must access the qid2cqidix RAM.  Give completions strict priority
// since they are freeing up a resource and not consuming one - avoid starvation.  Support backup mode of toggle
// arbiter in case different starvation issue arises.

assign lbi_ec_arb_reqs [ HQM_LSP_LBA_EC_ARB_CMP ]       = lbi_qid_cmp_arb_winner_v ;    // includes RELEASE
assign lbi_ec_arb_reqs [ HQM_LSP_LBA_EC_ARB_ENQ ]       = enq_nalb_fifo_pop_data_vreq ;
assign lbi_ec_arb_update                                = lbi_enq_req_taken | lbi_qid_cmp_req_taken ;

hqm_AW_strict_arb #( .NUM_REQS ( 2 ) ) i_lbi_ec_arb (
          .reqs                                 ( lbi_ec_arb_reqs )
        , .winner_v                             ( lbi_ec_arb_strict_winner_v )
        , .winner                               ( lbi_ec_arb_strict_winner )
) ;

//----
// Toggle arbiter
assign lbi_ec_arb_tie                           = lbi_ec_arb_reqs [ HQM_LSP_LBA_EC_ARB_CMP ] & lbi_ec_arb_reqs [ HQM_LSP_LBA_EC_ARB_ENQ ] ;
assign lbi_ec_arb_tie_broken                    = lbi_ec_arb_tie & lbi_ec_arb_update & cfg_control_ldb_ce_tog_arb ;

always_comb begin
  lbi_ec_arb_tog_winner_v                       = lbi_ec_arb_strict_winner_v ;
  lbi_ec_arb_tog_nxt                            = lbi_ec_arb_tog_f ;

  if ( lbi_ec_arb_tie ) begin
    if ( lbi_ec_arb_tog_f ) begin
      lbi_ec_arb_tog_winner                     = HQM_LSP_LBA_EC_ARB_ENQ ;
    end
    else begin
      lbi_ec_arb_tog_winner                     = HQM_LSP_LBA_EC_ARB_CMP ;
    end
  end
  else begin
    if ( lbi_ec_arb_reqs [ HQM_LSP_LBA_EC_ARB_CMP ] ) begin
      lbi_ec_arb_tog_winner                     = HQM_LSP_LBA_EC_ARB_CMP ;
    end
    else begin
      lbi_ec_arb_tog_winner                     = HQM_LSP_LBA_EC_ARB_ENQ ;
    end
  end

  if ( lbi_ec_arb_tie_broken ) begin
    lbi_ec_arb_tog_nxt                          = ~ lbi_ec_arb_tog_f ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    lbi_ec_arb_tog_f            <= 1'b0 ;
  end
  else begin
    lbi_ec_arb_tog_f            <= lbi_ec_arb_tog_nxt ;
  end
end // always
//----

always_comb begin
  if ( cfg_control_ldb_ce_tog_arb ) begin
    lbi_ec_arb_winner_v                         = lbi_ec_arb_tog_winner_v ;
    lbi_ec_arb_winner                           = lbi_ec_arb_tog_winner ;
  end
  else begin
    lbi_ec_arb_winner_v                         = lbi_ec_arb_strict_winner_v ;
    lbi_ec_arb_winner                           = lbi_ec_arb_strict_winner   ;
  end

  lbi_ec_arb_enq_v                              = 1'b0 ;
  lbi_ec_arb_cmp_v                              = 1'b0 ;

  case ( lbi_ec_arb_winner )
    HQM_LSP_LBA_EC_ARB_CMP : begin
      lbi_ec_arb_cmp_v                          = lbi_ec_arb_winner_v ;         // includes RELEASE
    end
    HQM_LSP_LBA_EC_ARB_ENQ : begin
      lbi_ec_arb_enq_v                          = lbi_ec_arb_winner_v ;
    end
  endcase
end // always

//-------------------------------------------------------------------------------------------------
// CQ completions

assign lbi_cq_cmp_arb_reqs [ HQM_LSP_LBA_CQ_ARB_ATM ]   = atm_cmp_fifo_pop_data_vreq ;
assign lbi_cq_cmp_arb_reqs [ HQM_LSP_LBA_CQ_ARB_NALB ]  = nalb_cmp_fifo_pop_data_vreq ;

hqm_AW_wrand_arb # ( .NUM_REQS ( 2 ) , .SEED ( 1 ) ) i_lbi_cq_cmp_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( lbi_cq_cmp_arb_reqs )
        , .cfg_weight           ( { cfg_lbi_cq_cmp_arb_weight_nalb ,            // Equal weights = random
                                    cfg_lbi_cq_cmp_arb_weight_atm } )
        , .winner_v             ( lbi_cq_cmp_arb_winner_v )
        , .winner               ( lbi_cq_cmp_arb_winner )
) ;

always_comb begin
  atm_cmp_fifo_pop                              = 1'b0 ;
  nalb_cmp_fifo_pop                             = 1'b0 ;
  lbi_inp_cq_cmp_cq_p                           = atm_cmp_fifo_pop_data_cq_p ;
  lbi_inp_cq_cmp_cq_wt_p                        = atm_cmp_fifo_pop_data_cq_wt_p ;
  lbi_inp_cq_cmp_cq                             = atm_cmp_fifo_pop_data.cq [HQM_NUM_LB_CQB2-1:0] ;
  lbi_inp_cq_cmp_qe_wt                          = atm_cmp_fifo_pop_data.qe_wt ;
  lbi_cq_cmp_arb_atm_v                          = 1'b0 ;
  lbi_inp_cq_cmp_no_dec                         = ( atm_cmp_fifo_pop_data.user == 1'b1) ;
  case ( lbi_cq_cmp_arb_winner )
    HQM_LSP_LBA_CQ_ARB_ATM : begin
      atm_cmp_fifo_pop                          = lbi_cq_cmp_req_taken ;
      lbi_cq_cmp_arb_atm_v                      = lbi_cq_cmp_arb_winner_v ;
      lbi_inp_cq_cmp_cq_p                       = atm_cmp_fifo_pop_data_cq_p ;
      lbi_inp_cq_cmp_cq_wt_p                    = atm_cmp_fifo_pop_data_cq_wt_p ;
      lbi_inp_cq_cmp_cq                         = atm_cmp_fifo_pop_data.cq [HQM_NUM_LB_CQB2-1:0] ;
      lbi_inp_cq_cmp_qe_wt                      = atm_cmp_fifo_pop_data.qe_wt ;
      lbi_inp_cq_cmp_no_dec                     = ( atm_cmp_fifo_pop_data.user == 1'b1) ;
    end
    HQM_LSP_LBA_CQ_ARB_NALB : begin
      nalb_cmp_fifo_pop                         = lbi_cq_cmp_req_taken ;
      lbi_cq_cmp_arb_atm_v                      = 1'b0 ;
      lbi_inp_cq_cmp_cq_p                       = nalb_cmp_fifo_pop_data_cq_p ;
      lbi_inp_cq_cmp_cq_wt_p                    = nalb_cmp_fifo_pop_data_cq_wt_p ;
      lbi_inp_cq_cmp_cq                         = nalb_cmp_fifo_pop_data.cq [HQM_NUM_LB_CQB2-1:0] ;
      lbi_inp_cq_cmp_qe_wt                      = nalb_cmp_fifo_pop_data.qe_wt ;
      lbi_inp_cq_cmp_no_dec                     = 1'b0 ;
    end
  endcase
end // always

assign lbi_cq_cmp_req_taken             = p0_lba_arb_cq_cmp_v & ~ p1_lba_ctrl_pipe.hold ;

//-------------------------------------------------------------------------------------------------
// Manage pipeline credits:
// - don't allow an atomic schedule or completion (go to lsp_ap_atm ) if the atm credit limit is reached
// - don't allow a nalb schedule (goes to nalb_sel_nalb FIFO) if the nalb credit limit is reached

// Need to subtract nalb schedules at p4 from atm_credit_count
// Need to subtract atm schedules at p4 from nalb_credit_count
assign p4_lba_atm_credit_count_dec_miss         = p4_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold & p4_lba_sch_arb_nalb ;
assign p4_lba_nalb_credit_count_dec_miss        = p4_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold & p4_lba_sch_arb_atm ;

// credit counts are at p0 level since that is where it gates off schedule requests, but inc/dec signals
// are controlled by their appropriate enables so that this register must not be under p1 enable control.
assign p0_lba_atm_credit_count_dec_amt          = { 2'h0 , credit_fifo_ap_aqed_dec_sch [0] } +
                                                  { 2'h0 , credit_fifo_ap_aqed_dec_sch [1] } +
                                                  { 2'h0 , credit_fifo_ap_aqed_dec_cmp } +
                                                  { 2'h0 , p4_lba_atm_credit_count_dec_miss } ;

assign p0_lba_atm_credit_count_px               = p0_lba_atm_credit_count_f + { 4'h0 , p0_lba_atm_credit_count_inc } ;
assign p0_lba_atm_credit_count_nxt              = p0_lba_atm_credit_count_px - { 2'h0 , p0_lba_atm_credit_count_dec_amt } ;


assign p0_lba_atm_credit_hold_cond              = ( { 3'h0 , p0_lba_atm_credit_count_f } >= cfg_atm_pipeline_credit_limit ) ;
//--------
assign p0_lba_nalb_credit_count_p1              = p0_lba_nalb_credit_count_f + 5'h1 ;
assign p0_lba_nalb_credit_count_m1              = p0_lba_nalb_credit_count_f - 5'h1 ;
assign p0_lba_nalb_credit_count_m2              = p0_lba_nalb_credit_count_f - 5'h2 ;

assign p0_lba_nalb_credit_count_dec_hit         = nalb_sel_nalb_fifo_pop ;

always_comb begin
  p0_lba_nalb_credit_count_nxt                  = p0_lba_nalb_credit_count_f ;
  case ( { p0_lba_nalb_credit_count_inc , p4_lba_nalb_credit_count_dec_miss , p0_lba_nalb_credit_count_dec_hit } )
    3'b001 ,
    3'b010 ,
    3'b111 : p0_lba_nalb_credit_count_nxt       = p0_lba_nalb_credit_count_m1 ;
    3'b011 : p0_lba_nalb_credit_count_nxt       = p0_lba_nalb_credit_count_m2 ;
    3'b100 : p0_lba_nalb_credit_count_nxt       = p0_lba_nalb_credit_count_p1 ;
    default : begin                     // Same as default assign above
      p0_lba_nalb_credit_count_nxt              = p0_lba_nalb_credit_count_f ;
    end
  endcase
end // always

assign p0_lba_nalb_credit_hold_cond             = ( { 3'h0 , p0_lba_nalb_credit_count_f } >= cfg_lba_pipeline_credit_limit ) ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p0_lba_atm_credit_count_f           <= 5'h0 ;
    p0_lba_nalb_credit_count_f          <= 5'h0 ;
  end
  else begin
    p0_lba_atm_credit_count_f           <= p0_lba_atm_credit_count_nxt ;
    p0_lba_nalb_credit_count_f          <= p0_lba_nalb_credit_count_nxt ;
  end
end // always
assign p0_lba_atm_credit_count_eq_0     = ~ ( | p0_lba_atm_credit_count_f ) ;
assign p0_lba_nalb_credit_count_eq_0    = ~ ( | p0_lba_nalb_credit_count_f ) ;

assign p0_lba_ctrl_pipe_sch_hold_cond   = p0_lba_nalb_credit_hold_cond | p0_lba_atm_credit_hold_cond |  ( ( qed_deq_credit_afull | aqed_deq_credit_afull ) & ~ cfg_control_qe_wt_blk ) ;

//-------------------------------------------------------------------------------------------------
// Final p1 lba arbiter
// The p0_lba_sch_state machine drives the selection, so the "final arbiter" is just a function of what
// that state machine allows.  The state machine determines whether or not a sch is possible; if it
// is not, then any valid combinations of E/T/C are allowed.  If it is possible, the type (slist, rlist,
// nalb) is not determined until later.
// The only need for additional arbitration is between Enqueues and QID completes, because both must
// access the qid2cqidix RAM to calculate the "cq has work" condition for all affected qids.
//
// The compatible actions are:
// schedule: none
// else: T, CQ_C, and either E or QID_C

// Partial conditions, do not include slow pop_cq signal yet
assign p0_lba_arb_pre_enq_v_cond        = lbi_ec_arb_enq_v ;
assign p0_lba_arb_pre_tok_v_cond        = ldb_token_rtn_fifo_pop_data_vreq ;
assign p0_lba_arb_pre_qid_cmp_v_cond    = lbi_ec_arb_cmp_v ;                    // includes RELEASE
assign p0_lba_arb_pre_cq_cmp_v_cond     = lbi_cq_cmp_arb_winner_v & ~ p0_lba_supress_cq_cmp ;

always_comb begin
  p0_lba_arb_winner_pre_v               = 1'b0 ;
  p0_lba_arb_sch_v                      = 1'b0 ;
  p0_lba_arb_pre_enq_v                  = 1'b0 ;
  p0_lba_arb_pre_tok_v                  = 1'b0 ;
  p0_lba_arb_pre_qid_cmp_v              = 1'b0 ;
  p0_lba_arb_pre_cq_cmp_v               = 1'b0 ;

  // Pipe enable included where used
  if ( p0_lba_pop_cq [4] ) begin
    p0_lba_arb_winner_pre_v             = 1'b1 ;        // If pop occurs, winner is not masked - p0_lba_restrict_bw_hold_cond must be 0 if pop allowed
    p0_lba_arb_sch_v                    = 1'b1 ;
  end
  else if ( ( p0_lba_arb_pre_enq_v_cond | p0_lba_arb_pre_tok_v_cond | p0_lba_arb_pre_qid_cmp_v_cond | p0_lba_arb_pre_cq_cmp_v_cond )
            & ~ p0_lba_restrict_bw_hold_cond ) begin
    p0_lba_arb_winner_pre_v             = 1'b1 ;
    p0_lba_arb_pre_enq_v                = p0_lba_arb_pre_enq_v_cond ;
    p0_lba_arb_pre_tok_v                = p0_lba_arb_pre_tok_v_cond ;
    p0_lba_arb_pre_qid_cmp_v            = p0_lba_arb_pre_qid_cmp_v_cond ;               // includes RELEASE
    p0_lba_arb_pre_cq_cmp_v             = p0_lba_arb_pre_cq_cmp_v_cond ;
  end
end // always

// When schedule issued from p0, don't know if it will be nalb or atm.  Increment both counts here, then adjust at
// p4 when it is decided which.

assign p0_lba_atm_credit_count_inc      = p0_lba_arb_winner_v & p1_lba_ctrl_pipe.en &
                                          ( p0_lba_arb_sch_v | p0_lba_arb_cmp_atm_v ) ;                         // Need to subtract nalb schedules at p4
assign p0_lba_nalb_credit_count_inc     = p0_lba_arb_winner_v & p1_lba_ctrl_pipe.en & p0_lba_arb_sch_v ;        // Need to subtract atm schedules at p4

assign p0_lba_restrict_bw_hold_cond     = ( cfg_control_single_op_lba & ( ( ~ lba_pipe_idle_f ) | p1_lba_ctrl_pipe_v_f ) ) |
                                          ( cfg_control_half_bw_lba & p1_lba_ctrl_pipe_v_f ) ;

assign p0_lba_arb_winner_v              = p0_lba_arb_winner_pre_v & ~ p0_lba_restrict_bw_hold_cond ;

// If config is disabling the selection of multiple ops, arbitrate RR to pick which one gets to go
always_comb begin
  if ( cfg_control_disable_multi_op_lba ) begin
    p0_lba_arb_enq_v            = 1'b0 ;
    p0_lba_arb_cq_cmp_v         = 1'b0 ;
    p0_lba_arb_qid_cmp_v        = 1'b0 ;
    p0_lba_arb_tok_v            = 1'b0 ;
    case ( p0_lba_mop_arb_winner )
      2'h0: p0_lba_arb_enq_v            = p0_lba_mop_arb_winner_v ;
      2'h1: p0_lba_arb_cq_cmp_v         = p0_lba_mop_arb_winner_v ;
      2'h2: p0_lba_arb_qid_cmp_v        = p0_lba_mop_arb_winner_v ;
      2'h3: p0_lba_arb_tok_v            = p0_lba_mop_arb_winner_v ;
    endcase
  end
  else begin
    p0_lba_arb_enq_v            = p0_lba_arb_pre_enq_v ;
    p0_lba_arb_cq_cmp_v         = p0_lba_arb_pre_cq_cmp_v ;
    p0_lba_arb_qid_cmp_v        = p0_lba_arb_pre_qid_cmp_v ;
    p0_lba_arb_tok_v            = p0_lba_arb_pre_tok_v ;
  end
end // always

assign p0_lba_mop_arb_reqs [0]  = p0_lba_arb_pre_enq_v_cond ;
assign p0_lba_mop_arb_reqs [1]  = p0_lba_arb_pre_cq_cmp_v_cond ;
assign p0_lba_mop_arb_reqs [2]  = p0_lba_arb_pre_qid_cmp_v_cond ;
assign p0_lba_mop_arb_reqs [3]  = p0_lba_arb_pre_tok_v_cond ;

// Not too picky about the update, don't overburden the "taken" logic, if we're running in this mode we don't care about this
// little extra power or fairness.  Include winner_v in update to avoid AW assertion error.
assign p0_lba_mop_arb_update    = cfg_control_disable_multi_op_lba & p0_lba_mop_arb_winner_pre_v ;

hqm_AW_rr_arb # ( .NUM_REQS ( 4 ) ) i_lba_multi_op_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p0_lba_mop_arb_reqs )
        , .update               ( p0_lba_mop_arb_update )
        , .winner_v             ( p0_lba_mop_arb_winner_pre_v )
        , .winner               ( p0_lba_mop_arb_winner )
) ;

// Defer gating in the slow pop_cq signal until here for static timing reasons
assign p0_lba_mop_arb_winner_v  = p0_lba_mop_arb_winner_pre_v & ~ p0_lba_pop_cq [4] & ~ p0_lba_restrict_bw_hold_cond ;

assign p0_lba_arb_cmp_atm_v     = p0_lba_arb_cq_cmp_v & lbi_cq_cmp_arb_atm_v ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB Scheduling
//-----------------------------------------------------------------------------------------------------

// p0_lba_arb_winner_v is effectively the "pipeline valid" for p0
// If p0 holds for scheduling reasons (credits, blast), still allow p0 valid to progress to p1
// (assuming p1 is not holding) because still may do E/T/C.  If S is being held because of scheduling
// reasons, S input request is gated off, so if arbiter output is still valid must be for E/T/C.
assign p1_lba_ctrl_pipe_v_nxt   = ( p0_lba_arb_winner_v  & ~ p0_lba_ctrl_pipe.hold ) | p1_lba_ctrl_pipe.hold ;
assign p2_lba_ctrl_pipe_v_nxt   = ( p1_lba_ctrl_pipe_v_f & ~ p1_lba_ctrl_pipe.hold ) | p2_lba_ctrl_pipe.hold ;
assign p3_lba_ctrl_pipe_v_nxt   = ( p2_lba_ctrl_pipe_v_f & ~ p2_lba_ctrl_pipe.hold ) | p3_lba_ctrl_pipe.hold ;
assign p4_lba_ctrl_pipe_v_nxt   = ( p3_lba_ctrl_pipe_v_f & ~ p3_lba_ctrl_pipe.hold ) | p4_lba_ctrl_pipe.hold ;
assign p5_lba_ctrl_pipe_v_nxt   = ( p4_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold ) | p5_lba_ctrl_pipe.hold ;

always_comb begin
  p1_lba_ctrl_pipe_nxt                          = p1_lba_ctrl_pipe_f ;
  if ( p1_lba_ctrl_pipe.en ) begin
    p1_lba_ctrl_pipe_nxt                        = '0 ;                          // Safety belt just in case any bits missed
    if ( p0_lba_arb_sch_v ) begin
      p1_lba_ctrl_pipe_nxt.sch_v                = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.sch_cq               = p0_lba_cq_arb_winner ;
      p1_lba_ctrl_pipe_nxt.sch_cq_p             = p0_lba_cq_gp ;
    end
    else begin  // Fields are dont care, but cleaner to avoid x in simulation
      p1_lba_ctrl_pipe_nxt.sch_v                = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.sch_cq               = 6'h0 ;
      p1_lba_ctrl_pipe_nxt.sch_cq_p             = 1'b1 ;
    end
    p1_lba_ctrl_pipe_nxt.sch_rlist_qidixv       = 16'h0 ;                       // Not known until loading p2, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_slist_qidixv       = 16'h0 ;                       // Not known until loading p2, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_nalb_qidixv        = 16'h0 ;                       // Not known until loading p2, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = 16'h0 ;                       // Not known until loading p2, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_nalb_v             = 1'b0 ;                        // Not known until loading p5, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_atm_v              = 1'b0 ;                        // Not known until loading p5, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_atm_rlist          = 1'b0 ;                        // Not known until loading p5, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_qid                = 7'h0 ;                        // Not known until loading p5, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_qidix_msb          = 1'b0 ;                        // Not known until loading p5, not needed yet
    p1_lba_ctrl_pipe_nxt.sch_qidix              = 3'h0 ;                        // Not known until loading p5, not needed yet

    if ( p0_lba_arb_enq_v ) begin
      p1_lba_ctrl_pipe_nxt.enq_v                = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.enq_qid              = lbi_inp_enq_qid ;
      p1_lba_ctrl_pipe_nxt.enq_qid_p            = lbi_inp_enq_qid_p ;
    end
    else begin
      p1_lba_ctrl_pipe_nxt.enq_v                = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.enq_qid              = 7'h0 ;
      p1_lba_ctrl_pipe_nxt.enq_qid_p            = 1'b1 ;
    end

    if ( p0_lba_arb_tok_v ) begin
      p1_lba_ctrl_pipe_nxt.tok_v                = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.tok_cq               = lbi_inp_tok_cq ;
      p1_lba_ctrl_pipe_nxt.tok_cq_p             = lbi_inp_tok_cq_p ;
      p1_lba_ctrl_pipe_nxt.tok_cnt              = lbi_inp_tok_cnt ;
      p1_lba_ctrl_pipe_nxt.tok_cnt_res          = lbi_inp_tok_cnt_res ;
    end
    else begin
      p1_lba_ctrl_pipe_nxt.tok_v                = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.tok_cq               = 6'h0 ;
      p1_lba_ctrl_pipe_nxt.tok_cq_p             = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.tok_cnt              = 11'h0 ;
      p1_lba_ctrl_pipe_nxt.tok_cnt_res          = 2'h0 ;
    end

    if ( p0_lba_arb_qid_cmp_v ) begin                           // include RELEASE - not really a completion
      if ( lbi_inp_qid_cmp_dec_only ) begin                     // RELEASE
        p1_lba_ctrl_pipe_nxt.qid_cmp_v          = 1'b0 ;
        p1_lba_ctrl_pipe_nxt.qid_if_dec_v       = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_qid            = lbi_inp_qid_cmp_qid ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_p          = lbi_inp_qid_cmp_qid_p ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_no_dec     = lbi_inp_qid_cmp_no_dec ;
      end
      else begin
        p1_lba_ctrl_pipe_nxt.qid_cmp_v          = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.qid_if_dec_v       = 1'b0 ;
        p1_lba_ctrl_pipe_nxt.cmp_qid            = lbi_inp_qid_cmp_qid ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_p          = lbi_inp_qid_cmp_qid_p ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_no_dec     = lbi_inp_qid_cmp_no_dec ;
      end
    end
    else begin
      p1_lba_ctrl_pipe_nxt.qid_cmp_v            = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.qid_if_dec_v         = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qid              = 7'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qid_p            = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_qid_no_dec       = 1'b0 ;
    end

    if ( p0_lba_arb_cq_cmp_v ) begin
      p1_lba_ctrl_pipe_nxt.cq_cmp_v             = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_cq               = lbi_inp_cq_cmp_cq ;
      p1_lba_ctrl_pipe_nxt.cmp_cq_p             = lbi_inp_cq_cmp_cq_p ;
      if ( p0_lba_arb_cmp_atm_v ) begin
        p1_lba_ctrl_pipe_nxt.cmp_atm            = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_atm        = { 1'b0 , atm_cmp_fifo_pop_data.qid } ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_atm_p      = atm_cmp_fifo_pop_data_qid_p ;
        p1_lba_ctrl_pipe_nxt.cmp_qidix_msb      = lbi_inp_cmp_qidix_msb ;
        p1_lba_ctrl_pipe_nxt.cmp_qidix          = lbi_inp_cmp_qidix ;
        p1_lba_ctrl_pipe_nxt.cmp_qpri           = lbi_inp_cmp_qpri ;
        p1_lba_ctrl_pipe_nxt.cmp_fid            = lbi_inp_cmp_fid ;
        p1_lba_ctrl_pipe_nxt.cmp_fid_p          = lbi_inp_cmp_fid_p ;
        p1_lba_ctrl_pipe_nxt.cmp_p              = lbi_inp_cmp_p ;
        p1_lba_ctrl_pipe_nxt.cmp_hid            = lbi_inp_cmp_hid ;
        p1_lba_ctrl_pipe_nxt.cmp_hid_p          = lbi_inp_cmp_hid_p ;
        p1_lba_ctrl_pipe_nxt.cmp_cq_no_dec      = lbi_inp_cq_cmp_no_dec ;
      end
      else begin
        p1_lba_ctrl_pipe_nxt.cmp_atm            = 1'b0 ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_atm        = 7'h0 ;
        p1_lba_ctrl_pipe_nxt.cmp_qid_atm_p      = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_qidix_msb      = 1'b0 ;
        p1_lba_ctrl_pipe_nxt.cmp_qidix          = 3'h0 ;
        p1_lba_ctrl_pipe_nxt.cmp_qpri           = 3'h0 ;
        p1_lba_ctrl_pipe_nxt.cmp_fid            = 12'h0 ;
        p1_lba_ctrl_pipe_nxt.cmp_fid_p          = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_p              = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_hid            = 16'h0 ;
        p1_lba_ctrl_pipe_nxt.cmp_hid_p          = 1'b1 ;
        p1_lba_ctrl_pipe_nxt.cmp_cq_no_dec      = lbi_inp_cq_cmp_no_dec ;
      end
    end
    else begin
      p1_lba_ctrl_pipe_nxt.cq_cmp_v             = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.cmp_cq               = 6'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_cq_p             = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_atm              = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qid_atm          = 7'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qid_atm_p        = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_qidix_msb        = 1'b0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qidix            = 3'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_qpri             = 3'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_fid              = 12'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_fid_p            = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_p                = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_hid              = 16'h0 ;
      p1_lba_ctrl_pipe_nxt.cmp_hid_p            = 1'b1 ;
      p1_lba_ctrl_pipe_nxt.cmp_cq_no_dec        = 1'b0 ;
    end
  end
end // always

always_comb begin
  p2_lba_ctrl_pipe_nxt                          = p2_lba_ctrl_pipe_f ;
  if ( p2_lba_ctrl_pipe.en ) begin
    p2_lba_ctrl_pipe_nxt                        = p1_lba_ctrl_pipe_f ;
    if ( p1_lba_ctrl_pipe_f.sch_v ) begin
      if ( p1_lba_ctrl_pipe_f_pcm ) begin
        p2_lba_ctrl_pipe_nxt.sch_rlist_qidixv     = { p1_lba_sch_rlist_v_ar [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b1 } ] , p1_lba_sch_rlist_v_ar [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b0 } ] } ;
        p2_lba_ctrl_pipe_nxt.sch_slist_qidixv     = { p1_lba_sch_slist_v_ar [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b1 } ] , p1_lba_sch_slist_v_ar [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b0 } ] } ;
        p2_lba_ctrl_pipe_nxt.sch_nalb_qidixv      = { p1_lba_sch_nalb_v_ar  [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b1 } ] , p1_lba_sch_nalb_v_ar  [ { p1_lba_ctrl_pipe_f_sch_pcq , 1'b0 } ] } ;
      end
      else begin
        p2_lba_ctrl_pipe_nxt.sch_rlist_qidixv     = { 8'h00 , p1_lba_sch_rlist_v_ar [ p1_lba_ctrl_pipe_f.sch_cq ] } ;
        p2_lba_ctrl_pipe_nxt.sch_slist_qidixv     = { 8'h00 , p1_lba_sch_slist_v_ar [ p1_lba_ctrl_pipe_f.sch_cq ] } ;
        p2_lba_ctrl_pipe_nxt.sch_nalb_qidixv      = { 8'h00 , p1_lba_sch_nalb_v_ar  [ p1_lba_ctrl_pipe_f.sch_cq ] } ;
      end
      if ( p1_lba_ctrl_pipe_cmpblast_cond )
        p2_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv        = p1_lba_sch_cmpblast_qidixv_blasted ;
      else
        p2_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv        = p1_lba_sch_cmpblast_qidixv_f ;
    end
  end
  else if ( p2_lba_ctrl_pipe.hold & p2_lba_ctrl_pipe_cmpblast_cond ) begin
    p2_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p2_lba_sch_cmpblast_qidixv_blasted ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_lba_cq_rpri_f            <= { HQM_QID_PER_CQ_2X { 1'b0 } } ;
    p4_lba_rpri_set_f           <= 1'b0 ;
    p4_lba_rpri_reset_f         <= 1'b0 ;
    p5_lba_rpri_set_f           <= 1'b0 ;
    p5_lba_rpri_reset_f         <= 1'b0 ;
    p6_lba_rpri_f               <= { HQM_LSP_NUM_LB_CQQIDIX { 1'b0 } } ;
  end
  else begin
    p3_lba_cq_rpri_f            <= p3_lba_cq_rpri_nxt ;
    p4_lba_rpri_set_f           <= p4_lba_rpri_set_nxt ;
    p4_lba_rpri_reset_f         <= p4_lba_rpri_reset_nxt ;
    p5_lba_rpri_set_f           <= p5_lba_rpri_set_nxt ;
    p5_lba_rpri_reset_f         <= p5_lba_rpri_reset_nxt ;
    p6_lba_rpri_f               <= p6_lba_rpri_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p1_lba_ctrl_pipe_f            <= p1_lba_ctrl_pipe_nxt ;
  p2_lba_ctrl_pipe_f            <= p2_lba_ctrl_pipe_nxt ;
  p3_lba_ctrl_pipe_f            <= p3_lba_ctrl_pipe_nxt ;
  p4_lba_ctrl_pipe_f            <= p4_lba_ctrl_pipe_nxt ;
  p5_lba_ctrl_pipe_f            <= p5_lba_ctrl_pipe_nxt ;
  p6_lba_ctrl_pipe_f            <= p6_lba_ctrl_pipe_nxt ;
  p7_lba_ctrl_pipe_f            <= p7_lba_ctrl_pipe_nxt ;
  p8_lba_ctrl_pipe_f            <= p8_lba_ctrl_pipe_nxt ;

  p8_lba_sch_pipe_f             <= p8_lba_sch_pipe_nxt ;

end // always

// p0_lba_arb_winner_v is effectively the "pipeline valid" for p0

assign p0_lba_ctrl_pipe.hold    = p0_lba_arb_winner_v  & p1_lba_ctrl_pipe.hold ;
assign p0_lba_ctrl_pipe.en      = 1'b1 ;                                                // State machine always able to advance

assign p1_lba_ctrl_pipe.hold    = p1_lba_ctrl_pipe_v_f & p2_lba_ctrl_pipe.hold ;
assign p1_lba_ctrl_pipe.en      = p0_lba_arb_winner_v  & ~ p1_lba_ctrl_pipe.hold ;

assign p2_lba_ctrl_pipe.hold    = p2_lba_ctrl_pipe_v_f & p3_lba_ctrl_pipe.hold ;
assign p2_lba_ctrl_pipe.en      = p1_lba_ctrl_pipe_v_f & ~ p2_lba_ctrl_pipe.hold ;

assign p3_lba_ctrl_pipe.hold    = p3_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe.hold ;
assign p3_lba_ctrl_pipe.en      = p2_lba_ctrl_pipe_v_f & ~ p3_lba_ctrl_pipe.hold ;

assign p4_from_p5_hold          = p4_lba_ctrl_pipe_v_f & p5_lba_ctrl_pipe.hold ;
assign p4_lba_ctrl_pipe.hold    = p4_from_p5_hold      | p4_lba_atm_sch_hold ;
assign p4_lba_ctrl_pipe.en      = p3_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold ;

assign p5_lba_ctrl_pipe.hold    = p5_lba_ctrl_pipe_v_f & p6_lba_ctrl_pipe.hold ;
assign p5_lba_ctrl_pipe.en      = p4_lba_ctrl_pipe_v_f & ~ p5_lba_ctrl_pipe.hold & ~ p4_lba_atm_sch_hold ;

assign p6_lba_ctrl_pipe.hold    = p6_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe.hold ;
assign p6_lba_ctrl_pipe.en      = p5_lba_ctrl_pipe_v_f & ~ p6_lba_ctrl_pipe.hold ;

assign p7_lba_ctrl_pipe.hold    = p7_lba_ctrl_pipe_v_1_f & p8_lba_ctrl_pipe.hold ;
assign p7_lba_ctrl_pipe.en      = p6_lba_ctrl_pipe_v_f & ~ p7_lba_ctrl_pipe.hold ;

// p8_lba_sch_hold_cond should never occur.
// If the wm and pipeline credits are correctly configured, we will never be attempting to push the nalb FIFO when it is afull/full.
// In theory we could hold the pipe in that case.  However, if we ever do that the LSP and AP pipes will get out of sync
// which opens the window for incorrect functionality (e.g. unblast occurs before blast it is attempting to unblast).
// Also full was "propagating" up through the pipe as a HFN for no good reason.  So just detect as an error and drop
// the push if it occurs (will result in "lost" tokens, inflight).
assign p8_lba_ctrl_pipe.hold    = p8_lba_ctrl_pipe_v_1_f_nnc & p9_lba_ctrl_pipe.hold ;
assign p8_lba_ctrl_pipe.en      = p7_lba_ctrl_pipe_v_f & ~ p8_lba_ctrl_pipe.hold ;

// p9 level is just status registers which are always able to be loaded - no holds
assign p9_lba_ctrl_pipe.hold    = 1'b0 ;
assign p9_lba_ctrl_pipe.en      = p8_lba_ctrl_pipe_v_1_f_nnc & ~ p9_lba_ctrl_pipe.hold ;

always_comb begin
  p3_lba_ctrl_pipe_nxt          = p3_lba_ctrl_pipe_f ;
  p4_lba_ctrl_pipe_nxt          = p4_lba_ctrl_pipe_f ;
  p5_lba_ctrl_pipe_nxt          = p5_lba_ctrl_pipe_f ;
  p6_lba_ctrl_pipe_nxt          = p6_lba_ctrl_pipe_f ;
  p7_lba_ctrl_pipe_nxt          = p7_lba_ctrl_pipe_f ;
  p8_lba_ctrl_pipe_nxt          = p8_lba_ctrl_pipe_f ;

  p3_lba_cq_rpri_nxt            = p3_lba_cq_rpri_f ;
  p4_lba_rpri_set_nxt           = p4_lba_rpri_set_f ;
  p4_lba_rpri_reset_nxt         = p4_lba_rpri_reset_f ;
  p5_lba_rpri_set_nxt           = p5_lba_rpri_set_f ;
  p5_lba_rpri_reset_nxt         = p5_lba_rpri_reset_f ;
  p8_lba_sch_pipe_nxt           = p8_lba_sch_pipe_f ;

  if ( p3_lba_ctrl_pipe.en ) begin
    p3_lba_ctrl_pipe_nxt                        = p2_lba_ctrl_pipe_f ;
    p3_lba_cq_rpri_nxt                          = p2_lba_cq_rpri ;

    if ( p2_lba_ctrl_pipe_cmpblast_cond )
      p3_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p2_lba_sch_cmpblast_qidixv_blasted ;
    else
      p3_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p2_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end
  else if ( p3_lba_ctrl_pipe.hold & p3_lba_ctrl_pipe_cmpblast_cond ) begin
    p3_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p3_lba_sch_cmpblast_qidixv_blasted ;
  end
  //----------------
  if ( p4_lba_ctrl_pipe.en ) begin
    p4_lba_ctrl_pipe_nxt                        = p3_lba_ctrl_pipe_f ;
    p4_lba_rpri_set_nxt                         = p3_lba_rpri_set_cond ;
    p4_lba_rpri_reset_nxt                       = p3_lba_rpri_reset_cond ;

    if ( p3_lba_ctrl_pipe_cmpblast_cond )
      p4_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p3_lba_sch_cmpblast_qidixv_blasted ;
    else
      p4_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p3_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end
  else if ( p4_lba_ctrl_pipe.hold & p4_lba_ctrl_pipe_cmpblast_cond ) begin
    p4_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p4_lba_sch_cmpblast_qidixv_blasted ;
  end
  //----------------
  if ( p5_lba_ctrl_pipe.en ) begin
    p5_lba_ctrl_pipe_nxt                        = p4_lba_ctrl_pipe_f ;
    p5_lba_rpri_set_nxt                         = p4_lba_rpri_set_f ;
    p5_lba_rpri_reset_nxt                       = p4_lba_rpri_reset_f ;

    // Fill in the fields from the schedule arbitration decision
    p5_lba_ctrl_pipe_nxt.sch_nalb_v             = p4_lba_sch_arb_nalb ;
    p5_lba_ctrl_pipe_nxt.sch_atm_v              = p4_lba_sch_arb_atm ;
    p5_lba_ctrl_pipe_nxt.sch_atm_rlist          = p4_lba_sch_atm_rlist_f ;
    p5_lba_ctrl_pipe_nxt.sch_qid                = p4_lba_sch_arb_winner_qid ;
    p5_lba_ctrl_pipe_nxt.sch_qidix_msb          = p4_lba_sch_arb_winner_qidix_msb ;
    p5_lba_ctrl_pipe_nxt.sch_qidix              = p4_lba_sch_arb_winner_qidix ;
    if ( p4_lba_ctrl_pipe_cmpblast_cond )
      p5_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p4_lba_sch_cmpblast_qidixv_blasted ;
    else
      p5_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p4_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end
  else if ( p5_lba_ctrl_pipe.hold & p5_lba_ctrl_pipe_cmpblast_cond ) begin
    p5_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p5_lba_sch_cmpblast_qidixv_blasted ;
  end
  //----------------
  if ( p6_lba_ctrl_pipe.en ) begin
    p6_lba_ctrl_pipe_nxt                        = p5_lba_ctrl_pipe_f ;
    if ( p5_lba_ctrl_pipe_cmpblast_cond )
      p6_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p5_lba_sch_cmpblast_qidixv_blasted ;
    else
      p6_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p5_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end
  else if ( p6_lba_ctrl_pipe.hold & p6_lba_ctrl_pipe_cmpblast_cond ) begin
    p6_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p6_lba_sch_cmpblast_qidixv_blasted ;
  end
  //----------------
  if ( p7_lba_ctrl_pipe.en ) begin
    p7_lba_ctrl_pipe_nxt                        = p6_lba_ctrl_pipe_f ;
    if ( p6_lba_ctrl_pipe_cmpblast_cond )
      p7_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p6_lba_sch_cmpblast_qidixv_blasted ;
    else
      p7_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p6_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end
  else if ( p7_lba_ctrl_pipe.hold & p7_lba_ctrl_pipe_cmpblast_cond ) begin
    p7_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv    = p7_lba_sch_cmpblast_qidixv_blasted ;
  end
  //----------------
  if ( p8_lba_ctrl_pipe.en ) begin
    p8_lba_ctrl_pipe_nxt                        = p7_lba_ctrl_pipe_f ;
    if ( p7_lba_ctrl_pipe_cmpblast_cond )
      p8_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p7_lba_sch_cmpblast_qidixv_blasted ;
    else
      p8_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv  = p7_lba_ctrl_pipe_f.sch_cmpblast_qidixv ;
  end

  // Derive the the sch pipe from the ctrl_pipe
  if ( p8_lba_ctrl_pipe.en ) begin
    p8_lba_sch_pipe_nxt.cq                      = p7_lba_ctrl_pipe_f.sch_cq ;
    p8_lba_sch_pipe_nxt.parity                  = p7_lba_ctrl_pipe_f.sch_cq_p ;  // Add in qid/qidix parity in next stage for delay reasons
    p8_lba_sch_pipe_nxt.slot_msb                = p7_lba_ctrl_pipe_f.sch_qidix_msb ;
    p8_lba_sch_pipe_nxt.slot                    = p7_lba_ctrl_pipe_f.sch_qidix ;
    p8_lba_sch_pipe_nxt.qid                     = p7_lba_ctrl_pipe_f.sch_qid ;
    p8_lba_sch_pipe_nxt.cm_code                 = p7_lba_qid_dpth_thrsh_cm_code ;
  end

end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for per-cq qid, priority and valid.
// p0/1/2/3 for the rw_pipe is lba pipe levels p1/p2/p3/p4
// Separate memories to simplify config access.  Only written by config.

assign p1_lba_ctrl_pipe_v_nxt_gated             = p1_lba_ctrl_pipe_v_nxt & ~ p1_lba_ctrl_pipe.hold ;    // rmw can't handle p0_v_nxt & p0_hold

always_comb begin
  if ( p0_lba_pop_cq [0] ) begin
    p1_lba_cq2qid_rw_pipe_nxt.rw_cmd            = HQM_AW_RWPIPE_READ ;
  end
  else begin
    p1_lba_cq2qid_rw_pipe_nxt.rw_cmd            = HQM_AW_RWPIPE_NOOP ;
  end
  p1_lba_cq2qid_rw_pipe_nxt.pcq                 = ( p1_lba_ctrl_pipe_nxt.sch_cq >> 1 ) ;
  p1_lba_cq2qid_rw_pipe_nxt.data_priov_odd      = { $bits ( lsp_cfg_cq2priov_t ) { 1'b0 } } ;   // Unused - cfg write done elsewhere
  p1_lba_cq2qid_rw_pipe_nxt.data_priov_even     = { $bits ( lsp_cfg_cq2priov_t ) { 1'b0 } } ;   // Unused - cfg write done elsewhere
  p1_lba_cq2qid_rw_pipe_nxt.data_qid_ms_odd     = { $bits ( lsp_cfg_cq2qid_t ) { 1'b0 } } ;     // Unused - cfg write done elsewhere
  p1_lba_cq2qid_rw_pipe_nxt.data_qid_ms_even    = { $bits ( lsp_cfg_cq2qid_t ) { 1'b0 } } ;     // Unused - cfg write done elsewhere
  p1_lba_cq2qid_rw_pipe_nxt.data_qid_ls_odd     = { $bits ( lsp_cfg_cq2qid_t ) { 1'b0 } } ;     // Unused - cfg write done elsewhere
  p1_lba_cq2qid_rw_pipe_nxt.data_qid_ls_even    = { $bits ( lsp_cfg_cq2qid_t ) { 1'b0 } } ;     // Unused - cfg write done elsewhere
end // always

// cq2prio part of this memory stores the full priority without scaling
hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ >> 1 )
        , .WIDTH                ( 2 * ( HQM_LSP_LB_CQ2PRIOV_MEM_WIDTH + ( 2 * HQM_LSP_LB_CQ2QID_MEM_WIDTH ) ) )
) i_cq2qid_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq2qid_rw_pipe_status )

        // cmd input
        , .p0_v_nxt             ( p1_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p1_lba_cq2qid_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p1_lba_cq2qid_rw_pipe_nxt.pcq )
        , .p0_write_data_nxt    ( { p1_lba_cq2qid_rw_pipe_nxt.data_priov_odd ,
                                    p1_lba_cq2qid_rw_pipe_nxt.data_priov_even ,
                                    p1_lba_cq2qid_rw_pipe_nxt.data_qid_ms_odd ,
                                    p1_lba_cq2qid_rw_pipe_nxt.data_qid_ms_even ,
                                    p1_lba_cq2qid_rw_pipe_nxt.data_qid_ls_odd ,
                                    p1_lba_cq2qid_rw_pipe_nxt.data_qid_ls_even } )
        , .p0_hold              ( p1_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p1_lba_cq2qid_rw_pipe_v_f_nc )
        , .p0_rw_f              ( p1_lba_cq2qid_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p1_lba_cq2qid_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p1_lba_cq2qid_rw_pipe_data_f_nc )

        , .p1_hold              ( p2_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p2_lba_cq2qid_rw_pipe_v_f_nc )
        , .p1_rw_f              ( p2_lba_cq2qid_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p2_lba_cq2qid_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p2_lba_cq2qid_rw_pipe_data_f_nc )

        , .p2_hold              ( p3_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p3_lba_cq2qid_rw_pipe_v_f_nc )
        , .p2_rw_f              ( p3_lba_cq2qid_rw_pipe_f_pnc.rw_cmd )      // Unused
        , .p2_addr_f            ( p3_lba_cq2qid_rw_pipe_f_pnc.pcq )         // Same as ctrl_pipe CQ/2
        , .p2_data_f            ( { p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_odd ,
                                    p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_even ,
                                    p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_odd ,
                                    p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_even ,
                                    p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_odd ,
                                    p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_even } )

        , .p3_hold              ( p4_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p4_lba_cq2qid_rw_pipe_v_f_nc )
        , .p3_rw_f              ( p4_lba_cq2qid_rw_pipe_f_nc.rw_cmd )                   // Unused
        , .p3_addr_f            ( p4_lba_cq2qid_rw_pipe_f_nc.pcq )                      // Unused
        , .p3_data_f            ( { p4_lba_cq2qid_rw_pipe_f_nc.data_priov_odd ,         // Unused
                                    p4_lba_cq2qid_rw_pipe_f_nc.data_priov_even ,        // Unused
                                    p4_lba_cq2qid_rw_pipe_f_nc.data_qid_ms_odd ,        // Unused
                                    p4_lba_cq2qid_rw_pipe_f_nc.data_qid_ms_even ,       // Unused
                                    p4_lba_cq2qid_rw_pipe_f_nc.data_qid_ls_odd ,        // Unused
                                    p4_lba_cq2qid_rw_pipe_f_nc.data_qid_ls_even } )     // Unused


        // mem intf
        , .mem_write            ( cfgsc_func_cfg_cq2priov_mem_we )              // Never used - cfg writes done elsewhere, no func write
        , .mem_read             ( cfgsc_func_cfg_cq2priov_mem_re )
        , .mem_addr             ( cfgsc_func_cfg_cq2priov_mem_addr )
        , .mem_write_data       ( {   cfgsc_func_cfg_cq2priov_mem_wdata         // Never used - no func write, cfg writes done elsewhere
                                    , cfgsc_func_cfg_cq2qid_1_mem_wdata         // Never used - no func write, cfg writes done elsewhere
                                    , cfgsc_func_cfg_cq2qid_0_mem_wdata } )     // Never used - no func write, cfg writes done elsewhere
        , .mem_read_data        ( {   cfgsc_func_cfg_cq2priov_mem_rdata
                                    , cfgsc_func_cfg_cq2qid_1_mem_rdata
                                    , cfgsc_func_cfg_cq2qid_0_mem_rdata } )
) ;

assign p3_lba_cq2qid_rw_pipe_rw_cmd_f_nc        = p3_lba_cq2qid_rw_pipe_f_pnc.rw_cmd ;

assign cfgsc_func_cfg_cq2qid_1_mem_we   = cfgsc_func_cfg_cq2priov_mem_we ;      // Never used - cfg writes done elsewhere
assign cfgsc_func_cfg_cq2qid_0_mem_we   = cfgsc_func_cfg_cq2priov_mem_we ;      // Never used - cfg writes done elsewhere

assign cfgsc_func_cfg_cq2qid_1_mem_re   = cfgsc_func_cfg_cq2priov_mem_re ;      // Always functionally read together
assign cfgsc_func_cfg_cq2qid_0_mem_re   = cfgsc_func_cfg_cq2priov_mem_re ;      // Always functionally read together

assign cfgsc_func_cfg_cq2qid_1_mem_addr = cfgsc_func_cfg_cq2priov_mem_addr ;    // Always functionally read together
assign cfgsc_func_cfg_cq2qid_0_mem_addr = cfgsc_func_cfg_cq2priov_mem_addr ;    // Always functionally read together

always_comb begin
  p3_lba_cq2qid_rw_pipe_qid_8_odd       = { p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_odd.qid_4 , p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_odd.qid_4 } ;
  p3_lba_cq2qid_rw_pipe_qid_8_even      = { p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_even.qid_4 , p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_even.qid_4 } ;

  p3_lba_cq2qid_par_chk_en              = p3_lba_ctrl_pipe_v_f & p3_lba_ctrl_pipe_f.sch_v ;

  p3_lba_cq2qid_cq_disable_odd          = cfg_cq_ldb_disable_f [ { p3_lba_cq2qid_rw_pipe_f_pnc.pcq , 1'b1 } ] ;
  p3_lba_cq2qid0_par_chk_en_odd         = p3_lba_cq2qid_par_chk_en &
                                          ( | ( p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_odd.v_8[3:0] ) ) ;
  p3_lba_cq2qid1_par_chk_en_odd         = p3_lba_cq2qid_par_chk_en &
                                          ( | ( p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_odd.v_8[7:4] ) ) ;
  p3_lba_cq2qid_cq_disable_even         = cfg_cq_ldb_disable_f [ { p3_lba_cq2qid_rw_pipe_f_pnc.pcq , 1'b0 } ] ;
  p3_lba_cq2qid0_par_chk_en_even        = p3_lba_cq2qid_par_chk_en &
                                          ( | ( p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_even.v_8[3:0] ) ) ;
  p3_lba_cq2qid1_par_chk_en_even        = p3_lba_cq2qid_par_chk_en &
                                          ( | ( p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_even.v_8[7:4] ) ) ;


  p3_lba_cq2qid_rw_pipe_data_priov_v_16  = { p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_odd.v_8 , p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_even.v_8 } ;

  if ( p3_lba_ctrl_pipe_f.sch_cq[0] ) begin
    p3_lba_cq2qid_rw_pipe_qid_8_x       = p3_lba_cq2qid_rw_pipe_qid_8_odd ;
    p3_lba_cq2qid_rw_pipe_data_priov_x  = p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_odd ;
    p3_lba_cq2qid_rw_pipe_data_qid_ls_x = p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_odd;
    p3_lba_cq2qid_rw_pipe_data_qid_ms_x = p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_odd;
    p3_lba_cq2qid_cq_disable_x          = p3_lba_cq2qid_cq_disable_odd ;
    p3_lba_cq2qid0_par_chk_en_x         = p3_lba_cq2qid0_par_chk_en_odd ;
    p3_lba_cq2qid1_par_chk_en_x         = p3_lba_cq2qid1_par_chk_en_odd ;
  end
  else begin
    p3_lba_cq2qid_rw_pipe_qid_8_x       = p3_lba_cq2qid_rw_pipe_qid_8_even ;
    p3_lba_cq2qid_rw_pipe_data_priov_x  = p3_lba_cq2qid_rw_pipe_f_pnc.data_priov_even ;
    p3_lba_cq2qid_rw_pipe_data_qid_ls_x = p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ls_even;
    p3_lba_cq2qid_rw_pipe_data_qid_ms_x = p3_lba_cq2qid_rw_pipe_f_pnc.data_qid_ms_even;
    p3_lba_cq2qid_cq_disable_x          = p3_lba_cq2qid_cq_disable_even ;
    p3_lba_cq2qid0_par_chk_en_x         = p3_lba_cq2qid0_par_chk_en_even ;
    p3_lba_cq2qid1_par_chk_en_x         = p3_lba_cq2qid1_par_chk_en_even ;
  end
end // always

hqm_AW_parity_check # ( .WIDTH ( 32 ) ) i_lba_cq2qid_priov_par_chk (
          .p                    ( p3_lba_cq2qid_rw_pipe_data_priov_x.p )
        , .d                    ( { p3_lba_cq2qid_rw_pipe_data_priov_x.v_8 ,
                                    p3_lba_cq2qid_rw_pipe_data_priov_x.pri_8 } )
        , .e                    ( p3_lba_cq2qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p3_lba_cq2qid_priov_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( 28 ) ) i_lba_cq2qid_qid0_par_chk (
          .p                    ( p3_lba_cq2qid_rw_pipe_data_qid_ls_x.p )
        , .d                    ( p3_lba_cq2qid_rw_pipe_data_qid_ls_x.qid_4 )
        , .e                    ( p3_lba_cq2qid0_par_chk_en_x )
        , .odd                  ( 1'b1 )
        , .err                  ( p3_lba_cq2qid_qid0_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( 28 ) ) i_lba_cq2qid_qid1_par_chk (
          .p                    ( p3_lba_cq2qid_rw_pipe_data_qid_ms_x.p )
        , .d                    ( p3_lba_cq2qid_rw_pipe_data_qid_ms_x.qid_4 )
        , .e                    ( p3_lba_cq2qid1_par_chk_en_x )
        , .odd                  ( 1'b1 )
        , .err                  ( p3_lba_cq2qid_qid1_par_err_cond )
) ;

assign p3_lba_cq2qid_v_err_cond         = p3_lba_cq2qid_par_chk_en & ~ ( | ( p3_lba_cq2qid_rw_pipe_data_priov_x.v_8[7:0] ) ) ;

//-------------------------------------------------------------------------------------------------
// qid arbiter
// - For slist/rlist and nalb, round robin among eligible qidix's for each priority
// - Pick the highest priority slist/rlist and nalb.  Between slist/rlist, if winner has the
//   same priority, lba_rpri_f toggle vector is used to arbitrate, with slist given preference.
// - Pick either atm (slist/rlist) or nalb based on priority.  If same priority, if one appears to be in the
//   middle of a burst, choose that one (cache locality / cq affinity), else use toggle bit.

always_comb begin
  for ( int i = HQM_QID_PER_CQ ; i < HQM_QID_PER_CQ_2X ; i = i + 1 ) begin              //JTC
    p3_lba_sch_atm_req_upper [i-HQM_QID_PER_CQ]      = ( p3_lba_ctrl_pipe_f_pcm ) &
                                                       ( p3_lba_ctrl_pipe_f.sch_slist_qidixv [i] | p3_lba_ctrl_pipe_f.sch_rlist_qidixv [i] ) &
                                                       p3_lba_cq2qid_rw_pipe_data_priov_v_16 [i] & p3_lba_ctrl_pipe_f.sch_v ;

    p3_lba_sch_nalb_req_upper [i-HQM_QID_PER_CQ]     = p3_lba_ctrl_pipe_f_pcm & p3_lba_ctrl_pipe_f.sch_nalb_qidixv [i] &
                                                       p3_lba_cq2qid_rw_pipe_data_priov_v_16 [i] & p3_lba_ctrl_pipe_f.sch_v ;
  end // for i

  for ( int i = 0 ; i < HQM_QID_PER_CQ ; i = i + 1 ) begin              //JTC
    p3_lba_sch_atm_req [i]      = ( p3_lba_ctrl_pipe_f.sch_slist_qidixv [i] | p3_lba_ctrl_pipe_f.sch_rlist_qidixv [i] ) &
                                  p3_lba_cq2qid_rw_pipe_data_priov_x.v_8[i] & p3_lba_ctrl_pipe_f.sch_v ;

    p3_lba_sch_nalb_req [i]     = p3_lba_ctrl_pipe_f.sch_nalb_qidixv [i] &
                                  p3_lba_cq2qid_rw_pipe_data_priov_x.v_8[i] & p3_lba_ctrl_pipe_f.sch_v ;
  end // for i

  for ( int i = 0 ; i < HQM_LSP_NUM_PRI_BINS ; i = i + 1 ) begin
    // Need to arrange the arbiter requests so that they are:
    // { qidix[7]pri7 , qidix[6]pri7, ... , qidix[0]pri7 ,
    //   qidix[7]pri6 , qidix[6]pri6, ... , qidix[0]pri6 ,
    //   ...
    //   qidix[7]pri0 , qidix[6]pri0, ... , qidix[0]pri0 }
    //
    // p3_lba_sch_atm_arb_pri_reqs and p3_lba_sch_nalb_arb_pri_reqs are organized:
    // pri_reqs[7] = { qidix[7]pri7 , qidix[7]pri6 , ... , qidix[7]pri0 }
    // ...
    // pri_reqs[0] = { qidix[0]pri7 , qidix[0]pri6 , ... , qidix[0]pri0 }
    for ( int j = 0 ; j < HQM_QID_PER_CQ_2X ; j = j + 1 ) begin            //JTC
      p3_lba_sch_atm_arb_reqs [ ( i * HQM_QID_PER_CQ_2X ) + j ]    = ( j >= HQM_QID_PER_CQ ) ? p3_lba_sch_atm_arb_pri_reqs_upper [j-HQM_QID_PER_CQ] [i] : p3_lba_sch_atm_arb_pri_reqs [j] [i] ;
      p3_lba_sch_nalb_arb_reqs [ ( i * HQM_QID_PER_CQ_2X ) + j ]   = ( j >= HQM_QID_PER_CQ ) ? p3_lba_sch_nalb_arb_pri_reqs_upper [j-HQM_QID_PER_CQ] [i] : p3_lba_sch_nalb_arb_pri_reqs [j] [i] ;
    end // for j
  end // for i
end // always

generate
  for ( genvar gi = 0 ; gi < HQM_QID_PER_CQ ; gi = gi + 1 ) begin: gen_lba_sch_dec_pri
    // Create decoded priority/request vector for arbiter.  For the gi'th index, create an 8-bit vector
    // where bit j=1 if the priority for this index = j.
    // If priority binning is done, from this point forward the downstream logic will only see the binned priorities
    assign p3_lba_cq2qid_rw_pipe_pri_scaled [gi]        = p3_lba_cq2qid_rw_pipe_data_priov_x.pri_8 [ (gi * 3) +: 3 ] >> HQM_LSP_PRI_BIN_FACTOR ;
    hqm_AW_bindec #( .WIDTH( HQM_LSP_NUM_PRI_BINSB2 ) ) i_p3_lba_sch_atm_arb_req_upper_bindec (
          .a                            ( p3_lba_cq2qid_rw_pipe_pri_scaled [gi] )
        , .enable                       ( p3_lba_sch_atm_req_upper [gi] )
        , .dec                          ( p3_lba_sch_atm_arb_pri_reqs_upper [gi] )
    ) ;

    hqm_AW_bindec #( .WIDTH( HQM_LSP_NUM_PRI_BINSB2 ) ) i_p3_lba_sch_atm_arb_req_bindec (
          .a                            ( p3_lba_cq2qid_rw_pipe_pri_scaled [gi] )
        , .enable                       ( p3_lba_sch_atm_req [gi] )
        , .dec                          ( p3_lba_sch_atm_arb_pri_reqs [gi] )
    ) ;

    hqm_AW_bindec #( .WIDTH( HQM_LSP_NUM_PRI_BINSB2 ) ) i_p3_lba_sch_nalb_arb_req_upper_bindec (
          .a                            ( p3_lba_cq2qid_rw_pipe_pri_scaled [gi] )
        , .enable                       ( p3_lba_sch_nalb_req_upper [gi] )
        , .dec                          ( p3_lba_sch_nalb_arb_pri_reqs_upper [gi] )
    ) ;
    hqm_AW_bindec #( .WIDTH( HQM_LSP_NUM_PRI_BINSB2 ) ) i_p3_lba_sch_nalb_arb_req_bindec (
          .a                            ( p3_lba_cq2qid_rw_pipe_pri_scaled [gi] )
        , .enable                       ( p3_lba_sch_nalb_req [gi] )
        , .dec                          ( p3_lba_sch_nalb_arb_pri_reqs [gi] )
    ) ;
  end // for
endgenerate

hqm_AW_wrrwrand_arb_windex # (
          .NUM_REQS             ( HQM_QID_PER_CQ_2X )                         //JTC
        , .NUM_PRI              ( HQM_LSP_NUM_PRI_BINS )
        , .WRR_WEIGHT_WIDTH     ( HQM_LSP_NUM_LDB_WRR_COUNTB2 )
        , .SEED                 ( 1 )
) i_p3_lba_sch_atm_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .cfg_weight_wrr       ( cfg_control_ldb_wrr_count_base )
        , .cfg_weight_wrand     ( { cfg_arb_weight_atm_nalb_qid_1_f , cfg_arb_weight_atm_nalb_qid_0_f } )             // Strict (default), or wrand with starvation avoidance
        , .index_f              ( p3_lba_atm_index_rw_pipe_data_pcm.indexes )
        , .count_f              ( p3_lba_atm_index_rw_pipe_data_pcm.counts )
        , .reqs                 ( p3_lba_sch_atm_arb_reqs )
        , .winner_v             ( p3_lba_sch_atm_arb_winner_v )
        , .winner_pri           ( p3_lba_sch_atm_arb_winner_pri )
        , .winner               ( { p3_lba_sch_atm_arb_winner_msb , p3_lba_sch_atm_arb_winner } )
        , .winner_in_seq        ( p3_lba_sch_atm_arb_winner_in_seq )
        , .index_nxt            ( p3_lba_sch_atm_index_upd_pcm )
        , .count_nxt            ( p3_lba_sch_atm_count_upd_pcm )
        , .winner_boosted       ( p3_lba_sch_atm_arb_winner_boosted )
) ;

hqm_AW_wrrwrand_arb_windex # (
          .NUM_REQS             ( HQM_QID_PER_CQ_2X )                         //JTC
        , .NUM_PRI              ( HQM_LSP_NUM_PRI_BINS )
        , .WRR_WEIGHT_WIDTH     ( HQM_LSP_NUM_LDB_WRR_COUNTB2 )
        , .SEED                 ( 2 )
) i_p3_lba_sch_nalb_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .cfg_weight_wrr       ( cfg_control_ldb_wrr_count_base )
        , .cfg_weight_wrand     ( { cfg_arb_weight_atm_nalb_qid_1_f , cfg_arb_weight_atm_nalb_qid_0_f } )             // Strict (default), or wrand with starvation avoidance
        , .index_f              ( p3_lba_nalb_index_rw_pipe_data_pcm.indexes )
        , .count_f              ( p3_lba_nalb_index_rw_pipe_data_pcm.counts )
	, .reqs                 ( p3_lba_sch_nalb_arb_reqs )
        , .winner_v             ( p3_lba_sch_nalb_arb_winner_v )
        , .winner_pri           ( p3_lba_sch_nalb_arb_winner_pri )
        , .winner               ( { p3_lba_sch_nalb_arb_winner_msb , p3_lba_sch_nalb_arb_winner } )
        , .winner_in_seq        ( p3_lba_sch_nalb_arb_winner_in_seq )
        , .index_nxt            ( p3_lba_sch_nalb_index_upd_pcm )
        , .count_nxt            ( p3_lba_sch_nalb_count_upd_pcm )
        , .winner_boosted       ( p3_lba_sch_nalb_arb_winner_boosted )
) ;

always_comb begin
  for ( int i = 0 ; i < HQM_QID_PER_CQ ; i = i + 1 ) begin                      //JTC
    p3_lba_cq2qid_qid_8_upper_ar [i]    = p3_lba_ctrl_pipe_f_pcm ? p3_lba_cq2qid_rw_pipe_qid_8_odd [ (i * 7) +: 7 ] : 8'h00 ;
    p3_lba_cq2qid_qid_8_ar [i]          = p3_lba_ctrl_pipe_f_pcm ? p3_lba_cq2qid_rw_pipe_qid_8_even [ (i * 7) +: 7 ] : p3_lba_cq2qid_rw_pipe_qid_8_x [ (i * 7) +: 7 ] ;
  end // for i
end // always

assign p3_lba_sch_atm_rlist_v           = p3_lba_ctrl_pipe_f.sch_rlist_qidixv [ { p3_lba_sch_atm_arb_winner_msb , p3_lba_sch_atm_arb_winner } ] ;
assign p3_lba_sch_atm_slist_v           = p3_lba_ctrl_pipe_f.sch_slist_qidixv [ { p3_lba_sch_atm_arb_winner_msb , p3_lba_sch_atm_arb_winner } ] ;
assign p3_lba_cq_qidix_rpri             = p3_lba_cq_rpri_f                    [ { p3_lba_sch_atm_arb_winner_msb , p3_lba_sch_atm_arb_winner } ] ;

// Same priority chosen as winner for both slist and rlist (both valid)
assign p3_lba_sch_atm_rlist_slist_collide       = p3_lba_sch_atm_arb_winner_v & p3_lba_sch_atm_slist_v & p3_lba_sch_atm_rlist_v ;

assign p3_lba_rpri_set_cond             = p3_lba_sch_atm_rlist_slist_collide & ~ p3_lba_cq_qidix_rpri & ~ cfg_control_disable_rlist_pri ;
assign p3_lba_rpri_reset_cond           = p3_lba_sch_atm_rlist_v             &   p3_lba_cq_qidix_rpri ;

assign p5_lba_ctrl_pipe_sch_cq_qidix    = p5_lba_ctrl_pipe_f_pcm ? { p5_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , p5_lba_ctrl_pipe_f.sch_qidix_msb , p5_lba_ctrl_pipe_f.sch_qidix } :
                                                                   { p5_lba_ctrl_pipe_f.sch_cq , p5_lba_ctrl_pipe_f.sch_qidix } ;

always_comb begin
  p6_lba_rpri_nxt                       = p6_lba_rpri_f ;

  if ( p6_lba_ctrl_pipe.en & p5_lba_ctrl_pipe_v_f & p5_lba_ctrl_pipe_f.sch_v & p5_lba_ctrl_pipe_f.sch_atm_v ) begin
    for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
      if ( p5_lba_ctrl_pipe_sch_cq_qidix  == i ) begin
        p6_lba_rpri_nxt [i]             = p5_lba_rpri_set_f | ( p6_lba_rpri_f [i] & ~ p5_lba_rpri_reset_f ) ;
      end
    end // for i
  end // if
end // always

// OK to read p6 reg via p2 because of slow sched rate
// Do as much read decoding as possible beforehand to reduce delay at p3
assign p2_lba_cq_rpri                   = p2_lba_ctrl_pipe_f_pcm ? { p6_lba_rpri_f [ { p2_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b1 , 3'h0 } +: 8 ] , 
                                                                     p6_lba_rpri_f [ { p2_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 , 3'h0 } +: 8 ] } :
                                                                   { 8'h00 ,
                                                                     p6_lba_rpri_f [ { p2_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 0 ] ,        3'h0 } +: 8 ] } ;

//--------------------------------------------------------------------
always_comb begin
  p4_lba_sch_atm_v_nxt                  = p4_lba_sch_atm_v_f ;
  p4_lba_sch_atm_qidix_msb_nxt          = p4_lba_sch_atm_qidix_msb_f ;
  p4_lba_sch_atm_qidix_nxt              = p4_lba_sch_atm_qidix_f ;
  p4_lba_sch_atm_pri_nxt                = p4_lba_sch_atm_pri_f ;
  p4_lba_sch_atm_in_seq_nxt             = p4_lba_sch_atm_in_seq_f ;
  p4_lba_sch_atm_qid_nxt                = p4_lba_sch_atm_qid_f ;
  p4_lba_sch_atm_index_upd_pcm_nxt      = p4_lba_sch_atm_index_upd_pcm_f ;
  p4_lba_sch_atm_count_upd_pcm_nxt      = p4_lba_sch_atm_count_upd_pcm_f ;
  p4_lba_sch_atm_rlist_nxt              = p4_lba_sch_atm_rlist_f ;
  p4_lba_atm_index_rw_pipe_data_unch_nxt        = p4_lba_atm_index_rw_pipe_data_unch_f ;
  p4_lba_sch_nalb_v_nxt                 = p4_lba_sch_nalb_v_f ;
  p4_lba_sch_nalb_qidix_msb_nxt         = p4_lba_sch_nalb_qidix_msb_f ;
  p4_lba_sch_nalb_qidix_nxt             = p4_lba_sch_nalb_qidix_f ;
  p4_lba_sch_nalb_pri_nxt               = p4_lba_sch_nalb_pri_f ;
  p4_lba_sch_nalb_in_seq_nxt            = p4_lba_sch_nalb_in_seq_f ;
  p4_lba_sch_nalb_qid_nxt               = p4_lba_sch_nalb_qid_f ;
  p4_lba_sch_nalb_index_upd_pcm_nxt     = p4_lba_sch_nalb_index_upd_pcm_f ;
  p4_lba_sch_nalb_count_upd_pcm_nxt     = p4_lba_sch_nalb_count_upd_pcm_f ;
  p4_lba_sch_arb_tog_nxt                = p4_lba_sch_arb_tog_f ;
  p4_lba_nalb_index_rw_pipe_data_unch_nxt       = p4_lba_nalb_index_rw_pipe_data_unch_f ;

  if ( p4_lba_ctrl_pipe.en ) begin
    p4_lba_sch_atm_v_nxt                = p3_lba_sch_atm_arb_winner_v ;
    p4_lba_sch_atm_qidix_msb_nxt        = p3_lba_sch_atm_arb_winner_msb ;
    p4_lba_sch_atm_qidix_nxt            = p3_lba_sch_atm_arb_winner ;
    case ( { p3_lba_sch_atm_arb_winner_boosted , p3_lba_sch_nalb_arb_winner_boosted } )
      2'b01 : begin
        p4_lba_sch_nalb_pri_nxt         = 3'h0 ;                                // Boost to highest priority
        p4_lba_sch_atm_pri_nxt          = 3'h7 >> HQM_LSP_PRI_BIN_FACTOR ;      // Supress competition to lowest priority
      end
      2'b10 : begin
        p4_lba_sch_atm_pri_nxt          = 3'h0 ;                                // Boost to highest priority
        p4_lba_sch_nalb_pri_nxt         = 3'h7 >> HQM_LSP_PRI_BIN_FACTOR ;      // Supress competition to lowest priority
      end
      2'b11 : begin                                                             // Both boosting, make same, 50/50 chance of getting through
        p4_lba_sch_atm_pri_nxt          = 3'h0 ;
        p4_lba_sch_nalb_pri_nxt         = 3'h0 ;
      end
      default : begin                                                           // No boosting, stick with the original input priorities
        p4_lba_sch_atm_pri_nxt          = p3_lba_sch_atm_arb_winner_pri ;
        p4_lba_sch_nalb_pri_nxt         = p3_lba_sch_nalb_arb_winner_pri ;
      end
    endcase
    p4_lba_sch_atm_in_seq_nxt           = p3_lba_sch_atm_arb_winner_in_seq ;
    p4_lba_sch_atm_qid_nxt              = p3_lba_sch_atm_arb_winner_msb ? p3_lba_cq2qid_qid_8_upper_ar [ p3_lba_sch_atm_arb_winner ] : p3_lba_cq2qid_qid_8_ar [ p3_lba_sch_atm_arb_winner ] ;
    p4_lba_sch_atm_index_upd_pcm_nxt    = p3_lba_sch_atm_index_upd_pcm ;
    p4_lba_sch_atm_count_upd_pcm_nxt    = p3_lba_sch_atm_count_upd_pcm ;
    if ( p3_lba_sch_atm_rlist_slist_collide )
      p4_lba_sch_atm_rlist_nxt          = p3_lba_cq_qidix_rpri ;        // If collision, favor slist but give rlist priority based on history
    else
      p4_lba_sch_atm_rlist_nxt          = p3_lba_sch_atm_rlist_v ;
    p4_lba_atm_index_rw_pipe_data_unch_nxt       = p3_lba_atm_index_rw_pipe_data_unch ;

    p4_lba_sch_nalb_v_nxt               = p3_lba_sch_nalb_arb_winner_v ;
    p4_lba_sch_nalb_qidix_msb_nxt       = p3_lba_sch_nalb_arb_winner_msb ;
    p4_lba_sch_nalb_qidix_nxt           = p3_lba_sch_nalb_arb_winner ;
    p4_lba_sch_nalb_in_seq_nxt          = p3_lba_sch_nalb_arb_winner_in_seq;
    p4_lba_sch_nalb_qid_nxt             = p3_lba_sch_nalb_arb_winner_msb ? p3_lba_cq2qid_qid_8_upper_ar [ p3_lba_sch_nalb_arb_winner ] : p3_lba_cq2qid_qid_8_ar [ p3_lba_sch_nalb_arb_winner ] ;
    p4_lba_sch_nalb_index_upd_pcm_nxt   = p3_lba_sch_nalb_index_upd_pcm ;
    p4_lba_sch_nalb_count_upd_pcm_nxt   = p3_lba_sch_nalb_count_upd_pcm ;
    p4_lba_nalb_index_rw_pipe_data_unch_nxt      = p3_lba_nalb_index_rw_pipe_data_unch ;

    p4_lba_sch_arb_tog_nxt              = ~ p4_lba_sch_arb_tog_f ;                         // free running
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p4_lba_sch_atm_v_f                  <= 1'b0 ;
    p4_lba_sch_nalb_v_f                 <= 1'b0 ;
    p4_lba_sch_arb_tog_f                <= 1'b0 ;
  end
  else begin
    p4_lba_sch_atm_v_f                  <= p4_lba_sch_atm_v_nxt ;
    p4_lba_sch_nalb_v_f                 <= p4_lba_sch_nalb_v_nxt ;
    p4_lba_sch_arb_tog_f                <= p4_lba_sch_arb_tog_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p4_lba_sch_atm_qid_f                  <= p4_lba_sch_atm_qid_nxt ;
  p4_lba_sch_atm_qidix_msb_f            <= p4_lba_sch_atm_qidix_msb_nxt ;
  p4_lba_sch_atm_qidix_f                <= p4_lba_sch_atm_qidix_nxt ;
  p4_lba_sch_atm_pri_f                  <= p4_lba_sch_atm_pri_nxt ;
  p4_lba_sch_atm_in_seq_f               <= p4_lba_sch_atm_in_seq_nxt ;
  p4_lba_sch_atm_index_upd_pcm_f        <= p4_lba_sch_atm_index_upd_pcm_nxt ;
  p4_lba_sch_atm_count_upd_pcm_f        <= p4_lba_sch_atm_count_upd_pcm_nxt ;
  p4_lba_sch_atm_rlist_f                <= p4_lba_sch_atm_rlist_nxt ;
  p4_lba_atm_index_rw_pipe_data_unch_f  <= p4_lba_atm_index_rw_pipe_data_unch_nxt ;
  p4_lba_sch_nalb_qid_f                 <= p4_lba_sch_nalb_qid_nxt ;
  p4_lba_sch_nalb_qidix_msb_f           <= p4_lba_sch_nalb_qidix_msb_nxt ;
  p4_lba_sch_nalb_qidix_f               <= p4_lba_sch_nalb_qidix_nxt ;
  p4_lba_sch_nalb_pri_f                 <= p4_lba_sch_nalb_pri_nxt ;
  p4_lba_sch_nalb_in_seq_f              <= p4_lba_sch_nalb_in_seq_nxt ;
  p4_lba_sch_nalb_index_upd_pcm_f       <= p4_lba_sch_nalb_index_upd_pcm_nxt ;
  p4_lba_sch_nalb_count_upd_pcm_f       <= p4_lba_sch_nalb_count_upd_pcm_nxt ;
  p4_lba_nalb_index_rw_pipe_data_unch_f <= p4_lba_nalb_index_rw_pipe_data_unch_nxt ;
end // always

always_comb begin
  p4_lba_sch_atm_count_upd = p4_lba_sch_atm_count_upd_pcm_f [ 23 : 0 ];
  p4_lba_sch_atm_index_upd = { p4_lba_sch_atm_count_upd_pcm_f [ 30 : 28 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [ 26 : 24 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [ 22 : 20 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [ 18 : 16 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [ 14 : 12 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [ 10 :  8 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [  6 :  4 ]
                             , p4_lba_sch_atm_count_upd_pcm_f [  2 :  0 ]
                             } ;
  p4_lba_sch_nalb_count_upd = p4_lba_sch_nalb_count_upd_pcm_f [ 23 : 0 ];
  p4_lba_sch_nalb_index_upd = { p4_lba_sch_nalb_count_upd_pcm_f [ 30 : 28 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [ 26 : 24 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [ 22 : 20 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [ 18 : 16 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [ 14 : 12 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [ 10 :  8 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [  6 :  4 ]
                              , p4_lba_sch_nalb_count_upd_pcm_f [  2 :  0 ]
                              } ; 
  if ( p4_lba_ctrl_pipe_f.sch_cq[0] ) begin                     // odd CQ has been updated
    p4_lba_atm_index_rw_pipe_data_struct.counts_odd     = p4_lba_sch_atm_count_upd ;
    p4_lba_atm_index_rw_pipe_data_struct.indexes_odd    = p4_lba_sch_atm_index_upd ;
    p4_lba_atm_index_rw_pipe_data_struct.counts_even    = p4_lba_atm_index_rw_pipe_data_unch_f.counts ;
    p4_lba_atm_index_rw_pipe_data_struct.indexes_even   = p4_lba_atm_index_rw_pipe_data_unch_f.indexes ;

    p4_lba_nalb_index_rw_pipe_data_struct.counts_odd    = p4_lba_sch_nalb_count_upd ;
    p4_lba_nalb_index_rw_pipe_data_struct.indexes_odd   = p4_lba_sch_nalb_index_upd ;
    p4_lba_nalb_index_rw_pipe_data_struct.counts_even   = p4_lba_nalb_index_rw_pipe_data_unch_f.counts ;
    p4_lba_nalb_index_rw_pipe_data_struct.indexes_even  = p4_lba_nalb_index_rw_pipe_data_unch_f.indexes ;
  end
  else begin                                                    // even CQ has been updated
    p4_lba_atm_index_rw_pipe_data_struct.counts_odd     = p4_lba_atm_index_rw_pipe_data_unch_f.counts ;
    p4_lba_atm_index_rw_pipe_data_struct.indexes_odd    = p4_lba_atm_index_rw_pipe_data_unch_f.indexes ;
    p4_lba_atm_index_rw_pipe_data_struct.counts_even    = p4_lba_sch_atm_count_upd ;
    p4_lba_atm_index_rw_pipe_data_struct.indexes_even   = p4_lba_sch_atm_index_upd ;

    p4_lba_nalb_index_rw_pipe_data_struct.counts_odd    = p4_lba_nalb_index_rw_pipe_data_unch_f.counts ;
    p4_lba_nalb_index_rw_pipe_data_struct.indexes_odd   = p4_lba_nalb_index_rw_pipe_data_unch_f.indexes ;
    p4_lba_nalb_index_rw_pipe_data_struct.counts_even   = p4_lba_sch_nalb_count_upd ;
    p4_lba_nalb_index_rw_pipe_data_struct.indexes_even  = p4_lba_sch_nalb_index_upd ;
  end
end // always

//--------
assign p4_lba_sch_nalb_in_seq           = p4_lba_sch_nalb_v_f & p4_lba_sch_nalb_in_seq_f ;
assign p4_lba_sch_atm_in_seq            = p4_lba_sch_atm_v_f & p4_lba_sch_atm_in_seq_f ;

// For the selection priority between atm and nalb, the p4 winner priority (possibly boosted) takes precedence.  If they are equal, then
// if one of them is in the middle of a burst sequence that takes precedence.  Otherwise select via toggle.

// Lowest number value priority (0) has highest priority.
assign p4_lba_sch_nalb_sel_pri          = { ~ p4_lba_sch_nalb_v_f , p4_lba_sch_nalb_pri_f , ~ p4_lba_sch_nalb_in_seq } ;
assign p4_lba_sch_atm_sel_pri           = { ~ p4_lba_sch_atm_v_f ,  p4_lba_sch_atm_pri_f ,  ~ p4_lba_sch_atm_in_seq } ;

assign p4_lba_sch_arb_winner_v          = p4_lba_ctrl_pipe_v_f & ( p4_lba_sch_nalb_v_f | p4_lba_sch_atm_v_f ) ;

always_comb begin
  p4_lba_sch_arb_atm_nalb_collide_cond_nc       = 1'b0 ;
  if ( p4_lba_sch_nalb_sel_pri < p4_lba_sch_atm_sel_pri ) begin
    p4_lba_sch_arb_atm_cond     = 1'b0 ;                                // nalb wins
  end
  else if ( p4_lba_sch_nalb_sel_pri > p4_lba_sch_atm_sel_pri ) begin
    p4_lba_sch_arb_atm_cond     = 1'b1 ;                                // atm wins
  end
  else begin                                                            // tie - use toggle to break tie
    p4_lba_sch_arb_atm_cond     = p4_lba_sch_arb_tog_f ;
    p4_lba_sch_arb_atm_nalb_collide_cond_nc     = 1'b1 ;
  end
end // always

assign p4_lba_sch_arb_nalb      = p4_lba_sch_arb_winner_v & ~ p4_lba_sch_arb_atm_cond ;
assign p4_lba_sch_arb_atm       = p4_lba_sch_arb_winner_v &   p4_lba_sch_arb_atm_cond ;

always_comb begin
  if ( p4_lba_sch_arb_atm ) begin       // atm
    p4_lba_sch_arb_winner_qid           = p4_lba_sch_atm_qid_f ;
    p4_lba_sch_arb_winner_qidix_msb     = p4_lba_sch_atm_qidix_msb_f ;
    p4_lba_sch_arb_winner_qidix         = p4_lba_sch_atm_qidix_f ;
  end
  else begin
    p4_lba_sch_arb_winner_qid           = p4_lba_sch_nalb_qid_f ;
    p4_lba_sch_arb_winner_qidix_msb     = p4_lba_sch_nalb_qidix_msb_f ;
    p4_lba_sch_arb_winner_qidix         = p4_lba_sch_nalb_qidix_f ;
  end
end // always

assign p4_lba_sch_arb_winner_cm_code    = p4_atq_cm_code_f [ p4_lba_sch_arb_winner_qid [HQM_NUM_LB_QIDB2-1:0] ] ;       // Coincidental that lba and atq are both p4

//-------------------------------------------------------------------------------------------------
// Update the counts as necessary for the selected qid and cq
assign p7_lba_qid_enq_cnt_upd_v         = p8_lba_ctrl_pipe.en & ( p7_lba_qid_enq_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_qid_if_cnt_upd_v          = p8_lba_ctrl_pipe.en & ( p7_lba_qid_if_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_cq_tok_cnt_upd_v          = p8_lba_ctrl_pipe.en & ( p7_lba_cq_tok_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_cq_if_cnt_upd_v           = p8_lba_ctrl_pipe.en & ( p7_lba_cq_if_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_tot_enq_cnt_upd_v         = p8_lba_ctrl_pipe.en & ( p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_tot_sch_cnt_upd_v         = p8_lba_ctrl_pipe.en & ( p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;
assign p7_lba_max_enq_depth_upd_v       = p8_lba_ctrl_pipe.en & ( p7_lba_max_enq_depth_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_READ ) & p7_lba_enq_cnt_gt_max_depth ;
assign p7_lba_perf_sch_count_upd_v      = p8_lba_ctrl_pipe.en & p7_lba_ctrl_pipe_f.sch_v ;

assign p5_lba_ctrl_pipe_v_nxt_gated     = p5_lba_ctrl_pipe_v_nxt & ~ p5_lba_ctrl_pipe.hold ;    // rmw can't handle p0_v_nxt & p0_hold

assign p7_lba_qid_enq_cnt_res_chk_en            = p7_lba_qid_enq_cnt_upd_v ;
assign p7_lba_qid_dpth_thrsh_par_chk_en         = p7_lba_qid_enq_cnt_res_chk_en ;
assign p7_lba_qid_if_cnt_res_chk_en             = p7_lba_qid_if_cnt_upd_v ;
assign p7_lba_qid_if_lim_par_chk_en             = p7_lba_qid_if_cnt_res_chk_en ;
assign p7_lba_cq_tok_cnt_res_chk_en             = p7_lba_cq_tok_cnt_upd_v ;
assign p7_lba_cq_tok_lim_par_chk_en             = p7_lba_cq_tok_cnt_res_chk_en ;


    //-------------------------------------------------------------------------------------------------
    // Manage storage for per-qid enqueue count, if-count and if-limit.
    // p0/1/2/3 for the rmw_pipe is lba pipe levels p5/p6/p7/p8

    //-------------------------------------------------------------------------------------------------
    // enq_cnt, dpth_thrsh

    always_comb begin
      if ( p4_lba_ctrl_pipe_v_f & ( p4_lba_ctrl_pipe_f.enq_v | p4_lba_sch_arb_nalb ) ) begin    // Don't read/update for atm sch - enq count not maintainted
        p5_lba_qid_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_RMW ;
        p5_lba_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_READ ;
      end
      else begin
        p5_lba_qid_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_NOOP ;
        p5_lba_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_NOOP ;
      end
      if ( p4_lba_sch_arb_nalb ) begin
        p5_lba_qid_enq_cnt_rmw_pipe_nxt.qid         = p4_lba_sch_arb_winner_qid ;
        p5_lba_qid_dpth_thrsh_rw_pipe_nxt.qid       = p4_lba_sch_arb_winner_qid ;
      end
      else begin
        p5_lba_qid_enq_cnt_rmw_pipe_nxt.qid         = p4_lba_ctrl_pipe_f.enq_qid ;
        p5_lba_qid_dpth_thrsh_rw_pipe_nxt.qid       = p4_lba_ctrl_pipe_f.enq_qid ;
      end
      p5_lba_qid_enq_cnt_rmw_pipe_nxt.data          = { $bits ( lsp_lb_qid_enq_cnt_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
      p5_lba_qid_dpth_thrsh_rw_pipe_nxt.data        = { $bits ( lsp_lb_qid_dpth_thrsh_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
    end // always

    hqm_AW_rmw_mem_4pipe_waddr #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID_ENQ_CNT_MEM_WIDTH )
    ) i_lba_qid_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_qid_enq_cnt_rmw_pipe_status_nc )                  // Unused, same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated  )
        , .p0_rw_nxt            ( p5_lba_qid_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_qid_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_qid_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_qid_enq_cnt_rmw_pipe_v_f_nc )                  // Unused, same as cq_tok_cnt pipe
        , .p0_rw_f              ( p5_lba_qid_enq_cnt_rmw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_qid_enq_cnt_rmw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_qid_enq_cnt_rmw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_qid_enq_cnt_rmw_pipe_v_f_nc )                  // Unused, same as cq_tok_cnt pipe
        , .p1_rw_f              ( p6_lba_qid_enq_cnt_rmw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_qid_enq_cnt_rmw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_qid_enq_cnt_rmw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_qid_enq_cnt_rmw_pipe_v_f_nc )                  // Unused, same as cq_tok_cnt pipe
        , .p2_rw_f              ( p7_lba_qid_enq_cnt_rmw_pipe_f.rw_cmd )                // Used to determine upd_v
        , .p2_addr_f            ( p7_lba_qid_enq_cnt_rmw_pipe_f.qid )                   // Used for bypass address
        , .p2_data_f            ( p7_lba_qid_enq_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypdata_sel_nxt   ( p7_lba_qid_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_qid_enq_cnt_upd )
        , .p3_bypaddr_sel_nxt   ( p7_lba_qid_enq_cnt_upd_v )
        , .p3_bypaddr_nxt       ( p7_lba_qid_enq_cnt_rmw_pipe_f.qid )
        , .p3_v_f               ( p8_lba_qid_enq_cnt_rmw_pipe_v_f_nc )                  // Unused, same as cq_tok_cnt pipe
        , .p3_rw_f              ( p8_lba_qid_enq_cnt_rmw_pipe_f_nc.rw_cmd )             // Unused
        , .p3_addr_f            ( p8_lba_qid_enq_cnt_rmw_pipe_f_nc.qid )                // Unused
        , .p3_data_f            ( p8_lba_qid_enq_cnt_rmw_pipe_f_nc.data )               // Unused


        // mem intf
        , .mem_write            ( func_qid_ldb_enqueue_count_mem_we )
        , .mem_read             ( func_qid_ldb_enqueue_count_mem_re )
        , .mem_write_addr       ( func_qid_ldb_enqueue_count_mem_waddr )
        , .mem_read_addr        ( func_qid_ldb_enqueue_count_mem_raddr )
        , .mem_write_data       ( func_qid_ldb_enqueue_count_mem_wdata )
        , .mem_read_data        ( func_qid_ldb_enqueue_count_mem_rdata  )
    ) ;

    hqm_AW_residue_add i_lba_qid_enq_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_qid_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_qid_enq_cnt_res_p1 )
    ) ;

    hqm_AW_residue_sub i_lba_qid_enq_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_qid_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_qid_enq_cnt_res_m1 )
    ) ;

    assign { p7_lba_qid_enq_cnt_p1_carry , p7_lba_qid_enq_cnt_p1 }      = { 1'b0 , p7_lba_qid_enq_cnt_rmw_pipe_f.data.cnt } + {{HQM_LSP_LB_QID_ENQ_CNT_WIDTH{1'b0}}, 1'b1} ;
    assign { p7_lba_qid_enq_cnt_m1_borrow , p7_lba_qid_enq_cnt_m1 }     = { 1'b0 , p7_lba_qid_enq_cnt_rmw_pipe_f.data.cnt } - {{HQM_LSP_LB_QID_ENQ_CNT_WIDTH{1'b0}}, 1'b1} ;

    always_comb begin
      p7_lba_qid_enq_cnt_oflow_cond                 = 1'b0 ;
      p7_lba_qid_enq_cnt_uflow_cond                 = 1'b0 ;
      if ( p7_lba_ctrl_pipe_f.sch_nalb_v ) begin
        if ( p7_lba_qid_enq_cnt_m1_borrow  ) begin
          p7_lba_qid_enq_cnt_upd                    = p7_lba_qid_enq_cnt_rmw_pipe_f.data ;  // Saturate, no residue error
          p7_lba_qid_enq_cnt_uflow_cond             = 1'b1 ;
        end
        else begin
          p7_lba_qid_enq_cnt_upd.cnt               = p7_lba_qid_enq_cnt_m1 ;
          p7_lba_qid_enq_cnt_upd.cnt_res           = p7_lba_qid_enq_cnt_res_m1 ;
        end
      end
      else begin
        if ( p7_lba_ctrl_pipe_f.enq_v & p7_lba_qid_enq_cnt_p1_carry ) begin
          p7_lba_qid_enq_cnt_upd                   = p7_lba_qid_enq_cnt_rmw_pipe_f.data ;  // Saturate, no residue error
          p7_lba_qid_enq_cnt_oflow_cond            = 1'b1 ;
        end
        else begin
          p7_lba_qid_enq_cnt_upd.cnt               = p7_lba_qid_enq_cnt_p1 ;
          p7_lba_qid_enq_cnt_upd.cnt_res           = p7_lba_qid_enq_cnt_res_p1 ;
        end
      end
    end // always

    assign p7_lba_qid_enq_cnt_upd_gt0           = | p7_lba_qid_enq_cnt_upd.cnt ;

    hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LB_QID_ENQ_CNT_WIDTH ) ) i_lba_qid_enq_cnt_res_chk (
          .r                    ( p7_lba_qid_enq_cnt_upd.cnt_res )
        , .d                    ( p7_lba_qid_enq_cnt_upd.cnt )
        , .e                    ( p7_lba_qid_enq_cnt_res_chk_en )
        , .err                  ( p7_lba_qid_enq_cnt_res_err_cond )
    );

    //-------------------------------------------------------------------------------------------------
    // qid_dpth_thrsh
    assign p7_lba_qid_dpth_thrsh_cm_code    = hqm_lsp_calc_thresh_code (   p7_lba_qid_enq_cnt_rmw_pipe_f.data.cnt
                                                                         , p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.data.thrsh ) ;

    hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_LB_QID_DPTH_THRSH_WIDTH ) ) i_lba_qid_dpth_thrsh_par_chk (
          .p                    ( p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.data.thrsh_p )
        , .d                    ( p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.data.thrsh )
        , .e                    ( p7_lba_qid_dpth_thrsh_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_qid_dpth_thrsh_par_err_cond )
    ) ;

    hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID_DPTH_THRSH_MEM_WIDTH )
    ) i_lba_qid_dpth_thrsh_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_qid_dpth_thrsh_rw_pipe_status_nc )                // Unused: same as lba_qid_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_qid_dpth_thrsh_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_qid_dpth_thrsh_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_qid_dpth_thrsh_rw_pipe_v_f_nc )                // Unused: same as cq_tok_cnt_pipe
        , .p0_rw_f              ( p5_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_qid_dpth_thrsh_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_qid_dpth_thrsh_rw_pipe_v_f_nc )                // Unused: same as cq_tok_cnt_pipe
        , .p1_rw_f              ( p6_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_qid_dpth_thrsh_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_qid_dpth_thrsh_rw_pipe_v_f_nc )                // Unused: same as cq_tok_cnt_pipe
        , .p2_rw_f              ( p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.rw_cmd )          // Unused
        , .p2_addr_f            ( p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.qid )             // Unused
        , .p2_data_f            ( p7_lba_qid_dpth_thrsh_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_qid_dpth_thrsh_rw_pipe_v_f_nc )                // Unused: same as cq_tok_cnt_pipe
        , .p3_rw_f              ( p8_lba_qid_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p8_lba_qid_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p8_lba_qid_dpth_thrsh_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cfg_nalb_qid_dpth_thrsh_mem_we )
        , .mem_read             ( func_cfg_nalb_qid_dpth_thrsh_mem_re )
        , .mem_addr             ( func_cfg_nalb_qid_dpth_thrsh_mem_addr )
        , .mem_write_data       ( func_cfg_nalb_qid_dpth_thrsh_mem_wdata )
        , .mem_read_data        ( func_cfg_nalb_qid_dpth_thrsh_mem_rdata )
    ) ;

    //-------------------------------------------------------------------------------------------------
    // qid_if_cnt, qid_if_lim

    always_comb begin
      if ( p4_lba_ctrl_pipe_v_f & ( p4_lba_sch_arb_winner_v | p4_lba_ctrl_pipe_f.qid_cmp_v | p4_lba_ctrl_pipe_f.qid_if_dec_v ) ) begin
        p5_lba_qid_if_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_RMW ;
        p5_lba_qid_if_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_READ ;
      end
      else begin
        p5_lba_qid_if_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_NOOP ;
        p5_lba_qid_if_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_NOOP ;
      end
      if ( p4_lba_sch_arb_winner_v ) begin
        p5_lba_qid_if_cnt_rmw_pipe_nxt.qid          = p4_lba_sch_arb_winner_qid ;
        p5_lba_qid_if_lim_rw_pipe_nxt.qid           = p4_lba_sch_arb_winner_qid ;
      end
      else begin
        p5_lba_qid_if_cnt_rmw_pipe_nxt.qid          = p4_lba_ctrl_pipe_f.cmp_qid ;
        p5_lba_qid_if_lim_rw_pipe_nxt.qid           = p4_lba_ctrl_pipe_f.cmp_qid ;
      end
      p5_lba_qid_if_cnt_rmw_pipe_nxt.data           = { $bits ( lsp_lb_qid_if_cnt_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
      p5_lba_qid_if_lim_rw_pipe_nxt.data            = { $bits ( lsp_lb_qid_if_lim_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
    end // always

    hqm_AW_rmw_mem_4pipe_waddr #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID_IF_CNT_MEM_WIDTH )
    ) i_lba_qid_if_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_qid_if_cnt_rmw_pipe_status_nc )                   // Unused: same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_qid_if_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_qid_if_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_qid_if_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_qid_if_cnt_rmw_pipe_v_f_nc )                   // Unused: same as cq_tok_cnt_pipe
        , .p0_rw_f              ( p5_lba_qid_if_cnt_rmw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_qid_if_cnt_rmw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_qid_if_cnt_rmw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_qid_if_cnt_rmw_pipe_v_f_nc )                   // Unused: same as cq_tok_cnt_pipe
        , .p1_rw_f              ( p6_lba_qid_if_cnt_rmw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_qid_if_cnt_rmw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_qid_if_cnt_rmw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_qid_if_cnt_rmw_pipe_v_f_nc )                   // Unused: same as cq_tok_cnt_pipe
        , .p2_rw_f              ( p7_lba_qid_if_cnt_rmw_pipe_f.rw_cmd )                 // Used to determine upd_v
        , .p2_addr_f            ( p7_lba_qid_if_cnt_rmw_pipe_f.qid )                    // Used for bypass address
        , .p2_data_f            ( p7_lba_qid_if_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypdata_sel_nxt   ( p7_lba_qid_if_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_qid_if_cnt_upd )
        , .p3_bypaddr_sel_nxt   ( p7_lba_qid_if_cnt_upd_v )
        , .p3_bypaddr_nxt       ( p7_lba_qid_if_cnt_rmw_pipe_f.qid )
        , .p3_v_f               ( p8_lba_qid_if_cnt_rmw_pipe_v_f_nc )                   // Unused: same as cq_tok_cnt_pipe
        , .p3_rw_f              ( p8_lba_qid_if_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p3_addr_f            ( p8_lba_qid_if_cnt_rmw_pipe_f_pnc.qid )                // Used for error rid
        , .p3_data_f            ( p8_lba_qid_if_cnt_rmw_pipe_f_pnc.data )               // Unused

        // mem intf
        , .mem_write            ( func_qid_ldb_inflight_count_mem_we  )
        , .mem_read             ( func_qid_ldb_inflight_count_mem_re  )
        , .mem_write_addr       ( func_qid_ldb_inflight_count_mem_waddr  )
        , .mem_read_addr        ( func_qid_ldb_inflight_count_mem_raddr  )
        , .mem_write_data       ( func_qid_ldb_inflight_count_mem_wdata  )
        , .mem_read_data        ( func_qid_ldb_inflight_count_mem_rdata  )
    ) ;

    hqm_AW_residue_add i_lba_qid_if_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_qid_if_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_qid_if_cnt_res_p1 )
    ) ;

    hqm_AW_residue_sub i_lba_qid_if_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_qid_if_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_qid_if_cnt_res_m1 )
    ) ;

    assign { p7_lba_qid_if_cnt_p1_carry , p7_lba_qid_if_cnt_p1 }      = { 1'b0 , p7_lba_qid_if_cnt_rmw_pipe_f.data.cnt } + 13'h1 ;
    assign { p7_lba_qid_if_cnt_m1_borrow , p7_lba_qid_if_cnt_m1 }     = { 1'b0 , p7_lba_qid_if_cnt_rmw_pipe_f.data.cnt } - 13'h1 ;

    always_comb begin
      p7_lba_qid_if_cnt_oflow_cond                      = 1'b0 ;
      p7_lba_qid_if_cnt_uflow_cond                      = 1'b0 ;
      if ( p7_lba_ctrl_pipe_f.sch_v ) begin
        if ( p7_lba_qid_if_cnt_p1_carry  ) begin
          p7_lba_qid_if_cnt_upd                         = p7_lba_qid_if_cnt_rmw_pipe_f.data ;  // Saturate, no residue error
          p7_lba_qid_if_cnt_oflow_cond                  = 1'b1 ;
        end
        else begin
          p7_lba_qid_if_cnt_upd.cnt                     = p7_lba_qid_if_cnt_p1 ;
          p7_lba_qid_if_cnt_upd.cnt_res                 = p7_lba_qid_if_cnt_res_p1 ;
        end
      end
      else if ( p7_lba_ctrl_pipe_f.qid_if_dec_v ) begin // Decrement only, no other qid/cmp action
        if ( p7_lba_qid_if_cnt_m1_borrow  ) begin
          p7_lba_qid_if_cnt_upd                         = p7_lba_qid_if_cnt_rmw_pipe_f.data ;  // Saturate, no residue error
          p7_lba_qid_if_cnt_uflow_cond                  = 1'b1 ;
        end
        else begin
          p7_lba_qid_if_cnt_upd.cnt                     = p7_lba_qid_if_cnt_m1  ;
          p7_lba_qid_if_cnt_upd.cnt_res                 = p7_lba_qid_if_cnt_res_m1  ;
        end
      end
      else begin        // qid_cmp_v
        if ( p7_lba_ctrl_pipe_f.cmp_qid_no_dec ) begin
          p7_lba_qid_if_cnt_upd                         = p7_lba_qid_if_cnt_rmw_pipe_f.data ;  // No change
        end
        else if ( p7_lba_ctrl_pipe_f.qid_cmp_v & p7_lba_qid_if_cnt_m1_borrow  ) begin
          p7_lba_qid_if_cnt_upd                         = p7_lba_qid_if_cnt_rmw_pipe_f.data ;  // Saturate, no residue error
          p7_lba_qid_if_cnt_uflow_cond                  = 1'b1 ;
        end
        else begin
          p7_lba_qid_if_cnt_upd.cnt                     = p7_lba_qid_if_cnt_m1  ;
          p7_lba_qid_if_cnt_upd.cnt_res                 = p7_lba_qid_if_cnt_res_m1  ;
        end
      end
    end // always

    assign p7_lba_qid_if_cnt_upd_lt_lim                 = ( p7_lba_qid_if_cnt_upd.cnt < p7_lba_qid_if_lim_rw_pipe_f_pnc.data.lim ) ;

    hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LB_QID_IF_CNT_WIDTH ) ) i_lba_qid_if_cnt_res_chk (
          .r                    ( p7_lba_qid_if_cnt_upd.cnt_res )
        , .d                    ( p7_lba_qid_if_cnt_upd.cnt )
        , .e                    ( p7_lba_qid_if_cnt_res_chk_en )
        , .err                  ( p7_lba_qid_if_cnt_res_err_cond  )
    );

    hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_LB_QID_IF_LIM_WIDTH ) ) i_lba_qid_if_lim_par_chk (
          .p                    ( p7_lba_qid_if_lim_rw_pipe_f_pnc.data.lim_p )
        , .d                    ( p7_lba_qid_if_lim_rw_pipe_f_pnc.data.lim )
        , .e                    ( p7_lba_qid_if_lim_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_qid_if_lim_par_err_cond )
    ) ;


    hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID_IF_LIM_MEM_WIDTH )
    ) i_lba_qid_if_lim_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_qid_if_lim_rw_pipe_status_nc )                    // Unused: same as lba_qid_if_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_qid_if_lim_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_qid_if_lim_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_qid_if_lim_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_qid_if_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt_pipe
        , .p0_rw_f              ( p5_lba_qid_if_lim_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_qid_if_lim_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_qid_if_lim_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_qid_if_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt_pipe
        , .p1_rw_f              ( p6_lba_qid_if_lim_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_qid_if_lim_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_qid_if_lim_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_qid_if_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt_pipe
        , .p2_rw_f              ( p7_lba_qid_if_lim_rw_pipe_f_pnc.rw_cmd )              // Unused
        , .p2_addr_f            ( p7_lba_qid_if_lim_rw_pipe_f_pnc.qid )                 // Unused
        , .p2_data_f            ( p7_lba_qid_if_lim_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_qid_if_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt_pipe
        , .p3_rw_f              ( p8_lba_qid_if_lim_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p8_lba_qid_if_lim_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p8_lba_qid_if_lim_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cfg_qid_ldb_inflight_limit_mem_we )
        , .mem_read             ( func_cfg_qid_ldb_inflight_limit_mem_re )
        , .mem_addr             ( func_cfg_qid_ldb_inflight_limit_mem_addr )
        , .mem_write_data       ( func_cfg_qid_ldb_inflight_limit_mem_wdata )
        , .mem_read_data        ( func_cfg_qid_ldb_inflight_limit_mem_rdata )
    ) ;


//-------------------------------------------------------------------------------------------------
// For the selected CQ, look up the token count and limit, and inflight count and limit.

// Manage storage for per-cq token count, token limit, inflight count and inflight limit.
// p0/1/2/3 for the rmw_pipe is lba pipe levels p3/p4/p5/p6
//-------------------------------------------------------------------------------------------------
// cq_tok_cnt, cq_tok_lim

always_comb begin
  if ( p4_lba_ctrl_pipe_v_f & ( p4_lba_ctrl_pipe_f.tok_v | p4_lba_ctrl_pipe_f.sch_v ) ) begin
    p5_lba_cq_tok_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_RMW ;          // Only (conditionally) do rmw if tok or sch
    p5_lba_cq_tok_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_READ ;
  end
  else begin
    p5_lba_cq_tok_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_NOOP ;
    p5_lba_cq_tok_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_NOOP ;
  end
  if ( p4_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe_f.enq_v )
    p5_lba_tot_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_RMW ;
  else
    p5_lba_tot_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_NOOP ;
  if ( p4_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe_f.sch_v )
    p5_lba_tot_sch_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_RMW ;
  else
    p5_lba_tot_sch_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_NOOP ;
  if ( p4_lba_ctrl_pipe_v_f & ( p4_lba_ctrl_pipe_f.enq_v | p4_lba_sch_arb_nalb ) ) begin
    p5_lba_max_enq_depth_rmw_pipe_nxt.rw_cmd    = HQM_AW_RMWPIPE_READ ;         // Also check on sch (decrement) in case RW/C (sets to 0) is followed by sch and depth is > 0
                                                                                // Update occurs via bypass going into p8 if curr upd depth > curr max
                                                                                // Stats not maintained for ATM
  end
  else begin
    p5_lba_max_enq_depth_rmw_pipe_nxt.rw_cmd    = HQM_AW_RMWPIPE_NOOP ;
  end
  //----------------------------------------------------------------------------
  if ( p4_lba_ctrl_pipe_f.sch_v ) begin
    p5_lba_cq_tok_cnt_rmw_pipe_nxt.cq           = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
    p5_lba_cq_tok_lim_rw_pipe_nxt.cq            = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
  end
  else begin
    p5_lba_cq_tok_cnt_rmw_pipe_nxt.cq           = p4_lba_ctrl_pipe_f.tok_cq ;
    p5_lba_cq_tok_lim_rw_pipe_nxt.cq            = p4_lba_ctrl_pipe_f.tok_cq ;
  end
  p5_lba_tot_enq_cnt_rmw_pipe_nxt.qid           = p4_lba_ctrl_pipe_f.enq_qid ;
  p5_lba_tot_sch_cnt_rmw_pipe_nxt.cq            = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
  if ( p4_lba_ctrl_pipe_f.enq_v ) begin
    p5_lba_max_enq_depth_rmw_pipe_nxt.qid       = p4_lba_ctrl_pipe_f.enq_qid ;
  end
  else begin
    p5_lba_max_enq_depth_rmw_pipe_nxt.qid       = p4_lba_sch_arb_winner_qid ;
  end
  //----------------------------------------------------------------------------
  p5_lba_cq_tok_cnt_rmw_pipe_nxt.data           = { $bits ( lsp_lb_cq_tok_cnt_t ) { 1'b0 } } ;  // Unused - cfg write done elsewhere
  p5_lba_cq_tok_lim_rw_pipe_nxt.data            = { $bits ( lsp_lb_cq_tok_lim_t ) { 1'b0 } } ;  // Unused - cfg write done elsewhere
  p5_lba_tot_enq_cnt_rmw_pipe_nxt.data          = { $bits ( lsp_arch_cnt_t ) { 1'b0 } } ;       // Unused - cfg write done elsewhere
  p5_lba_tot_sch_cnt_rmw_pipe_nxt.data          = { $bits ( lsp_arch_cnt_t ) { 1'b0 } } ;       // Unused - cfg write done elsewhere
  p5_lba_max_enq_depth_rmw_pipe_nxt.data        = { HQM_LSP_LB_QID_ENQ_CNT_WIDTH { 1'b0 } } ;   // Unused - cfg write done elsewhere
end // always

hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_LB_CQ_TOK_CNT_MEM_WIDTH )
) i_lba_cq_tok_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq_tok_cnt_rmw_pipe_status )

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_cq_tok_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_cq_tok_cnt_rmw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_cq_tok_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_ctrl_pipe_v_f )
        , .p0_rw_f              ( p5_lba_cq_tok_cnt_rmw_pipe_rw_f_nc )                  // Unused
        , .p0_addr_f            ( p5_lba_cq_tok_cnt_rmw_pipe_addr_f_nc )                // Unused
        , .p0_data_f            ( p5_lba_cq_tok_cnt_rmw_pipe_data_f_nc )                // Unused

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_ctrl_pipe_v_f )
        , .p1_rw_f              ( p6_lba_cq_tok_cnt_rmw_pipe_rw_f_nc )                  // Unused
        , .p1_addr_f            ( p6_lba_cq_tok_cnt_rmw_pipe_addr_f_nc )                // Unused
        , .p1_data_f            ( p6_lba_cq_tok_cnt_rmw_pipe_data_f_nc )                // Unused

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_ctrl_pipe_v_f )
        , .p2_rw_f              ( p7_lba_cq_tok_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p7_lba_cq_tok_cnt_rmw_pipe_f.cq )
        , .p2_data_f            ( p7_lba_cq_tok_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p7_lba_cq_tok_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_cq_tok_cnt_upd_cnt )
        , .p3_v_f               ( p8_lba_ctrl_pipe_v_f )
        , .p3_rw_f              ( p8_lba_cq_tok_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p3_addr_f            ( p8_lba_cq_tok_cnt_rmw_pipe_f_pnc.cq )                 // Used for error rid
        , .p3_data_f            ( p8_lba_cq_tok_cnt_rmw_pipe_f_pnc.data )               // Unused


        // mem intf
        , .mem_write            ( func_cq_ldb_token_count_mem_we )
        , .mem_read             ( func_cq_ldb_token_count_mem_re )
        , .mem_write_addr       ( func_cq_ldb_token_count_mem_waddr )
        , .mem_read_addr        ( func_cq_ldb_token_count_mem_raddr )
        , .mem_write_data       ( func_cq_ldb_token_count_mem_wdata )
        , .mem_read_data        ( func_cq_ldb_token_count_mem_rdata )
) ;

hqm_AW_residue_add i_lba_cq_tok_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_cq_tok_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_cq_tok_cnt_res_p1 )
) ;

hqm_AW_residue_sub i_lba_cq_tok_cnt_res_sub (
          .a                    ( p7_lba_ctrl_pipe_f.tok_cnt_res )
        , .b                    ( p7_lba_cq_tok_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_cq_tok_cnt_res_mn )
) ;

assign { p7_lba_cq_tok_cnt_p1_carry , p7_lba_cq_tok_cnt_p1 }    = { 1'b0 , p7_lba_cq_tok_cnt_rmw_pipe_f.data.cnt } + 12'h1 ;
assign { p7_lba_cq_tok_cnt_mn_borrow , p7_lba_cq_tok_cnt_mn }   = { 1'b0 , p7_lba_cq_tok_cnt_rmw_pipe_f.data.cnt } - { 1'b0 , p7_lba_ctrl_pipe_f.tok_cnt } ;

always_comb begin
  p7_lba_cq_tok_cnt_oflow_cond                  = 1'b0 ;
  p7_lba_cq_tok_cnt_uflow_cond                  = 1'b0 ;
  if ( p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.sch_atm_v ) begin
    if ( p7_lba_cq_tok_cnt_p1_carry ) begin
      p7_lba_cq_tok_cnt_upd_cnt                 = p7_lba_cq_tok_cnt_rmw_pipe_f.data ;   // Saturate, no residue error
      p7_lba_cq_tok_cnt_oflow_cond              = 1'b1 ;
    end
    else begin
      p7_lba_cq_tok_cnt_upd_cnt.cnt             = p7_lba_cq_tok_cnt_p1 ;
      p7_lba_cq_tok_cnt_upd_cnt.cnt_res         = p7_lba_cq_tok_cnt_res_p1 ;
    end
  end
  else begin
    if ( p7_lba_cq_tok_cnt_mn_borrow ) begin    // Decrement to 0, no residue error
      p7_lba_cq_tok_cnt_upd_cnt.cnt             = { HQM_LSP_LB_CQ_TOK_CNT_WIDTH { 1'b0 } } ;
      p7_lba_cq_tok_cnt_upd_cnt.cnt_res         = 2'h0 ;
      p7_lba_cq_tok_cnt_uflow_cond              = 1'b1 ;
    end
    else begin
      p7_lba_cq_tok_cnt_upd_cnt.cnt             = p7_lba_cq_tok_cnt_mn ;
      p7_lba_cq_tok_cnt_upd_cnt.cnt_res         = p7_lba_cq_tok_cnt_res_mn ;
    end
  end
end // always

assign p7_lba_cq_tok_cnt_upd_lt_lim_next        = ( p7_lba_cq_tok_cnt_upd_cnt.cnt < p7_lba_cq_tok_limit ) ;
assign p7_lba_cq_tok_cnt_upd_gt_0               = | p7_lba_cq_tok_cnt_upd_cnt.cnt ;

assign p2_lba_inp_tok_cnt_res_chk_en            = p2_lba_ctrl_pipe_v_f & p3_lba_ctrl_pipe.en & p2_lba_ctrl_pipe_f.tok_v ;

hqm_AW_residue_check #( .WIDTH ( 11 ) ) i_lba_inp_tok_cnt_res_chk (
          .r                    ( p2_lba_ctrl_pipe_f.tok_cnt_res )
        , .d                    ( p2_lba_ctrl_pipe_f.tok_cnt )
        , .e                    ( p2_lba_inp_tok_cnt_res_chk_en )
        , .err                  ( p2_lba_inp_tok_cnt_res_err_cond )
) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LB_CQ_TOK_CNT_WIDTH ) ) i_lba_cq_tok_cnt_res_chk (
          .r                    ( p7_lba_cq_tok_cnt_upd_cnt.cnt_res )
        , .d                    ( p7_lba_cq_tok_cnt_upd_cnt.cnt )
        , .e                    ( p7_lba_cq_tok_cnt_res_chk_en )
        , .err                  ( p7_lba_cq_tok_cnt_res_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_LB_CQ_TOK_LIM_SEL_WIDTH ) ) i_lba_cq_tok_lim_par_chk (
          .p                    ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.data.lim_p )
        , .d                    ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.data.lim_sel )
        , .e                    ( p7_lba_cq_tok_lim_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_cq_tok_lim_par_err_cond )
) ;

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_LB_CQ_TOK_LIM_SEL_MEM_WIDTH )
    ) i_lba_cq_tok_lim_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq_tok_lim_rw_pipe_status_nc )                    // Unused: same as lba_cq_tok_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_cq_tok_lim_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_cq_tok_lim_rw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_cq_tok_lim_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_cq_tok_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt pipe
        , .p0_rw_f              ( p5_lba_cq_tok_lim_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_cq_tok_lim_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_cq_tok_lim_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_cq_tok_lim_rw_pipe_v_f_nc )                    // Unused: same as cq_tok_cnt pipe
        , .p1_rw_f              ( p6_lba_cq_tok_lim_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_cq_tok_lim_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_cq_tok_lim_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_ctrl_pipe_v_1_f )                              // Same as cq_tok_cnt pipe, replicated to reduce transitive fanout
        , .p2_rw_f              ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.rw_cmd )          // Unused
        , .p2_addr_f            ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.cq )              // Unused
        , .p2_data_f            ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_ctrl_pipe_v_1_f_nnc )                          // Same as cq_tok_cnt pipe,  replicated to reduce transitive fanout
        , .p3_rw_f              ( p8_lba_cq_tok_lim_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p8_lba_cq_tok_lim_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p8_lba_cq_tok_lim_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cfg_cq_ldb_token_depth_select_mem_we )
        , .mem_read             ( func_cfg_cq_ldb_token_depth_select_mem_re )
        , .mem_addr             ( func_cfg_cq_ldb_token_depth_select_mem_addr )
        , .mem_write_data       ( func_cfg_cq_ldb_token_depth_select_mem_wdata )
        , .mem_read_data        ( func_cfg_cq_ldb_token_depth_select_mem_rdata )
) ;

always_comb begin
  case ( p7_lba_cq_tok_lim_rw_pipe_f_pnc.data.lim_sel )
    4'h0 :      begin p7_lba_cq_tok_limit       = 11'h004 ;     end
    4'h1 :      begin p7_lba_cq_tok_limit       = 11'h008 ;     end
    4'h2 :      begin p7_lba_cq_tok_limit       = 11'h010 ;     end
    4'h3 :      begin p7_lba_cq_tok_limit       = 11'h020 ;     end
    4'h4 :      begin p7_lba_cq_tok_limit       = 11'h040 ;     end
    4'h5 :      begin p7_lba_cq_tok_limit       = 11'h080 ;     end
    4'h6 :      begin p7_lba_cq_tok_limit       = 11'h100 ;     end
    4'h7 :      begin p7_lba_cq_tok_limit       = 11'h200 ;     end
    4'h8 :      begin p7_lba_cq_tok_limit       = 11'h400 ;     end
    default :   begin p7_lba_cq_tok_limit       = 11'h000 ;     end
  endcase
end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for lba total enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ARCH_CNT_MEM_WIDTH )
) i_lba_tot_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_tot_enq_cnt_rmw_pipe_status_nc )                  // Unused, same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_tot_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_tot_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_tot_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_tot_enq_cnt_rmw_pipe_v_f_nc )                  // Unused
        , .p0_rw_f              ( p5_lba_tot_enq_cnt_rmw_pipe_rw_f_nc )                 // Unused
        , .p0_addr_f            ( p5_lba_tot_enq_cnt_rmw_pipe_addr_f_nc )               // Unused
        , .p0_data_f            ( p5_lba_tot_enq_cnt_rmw_pipe_data_f_nc )               // Unused

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_tot_enq_cnt_rmw_pipe_v_f_nc )                  // Unused
        , .p1_rw_f              ( p6_lba_tot_enq_cnt_rmw_pipe_rw_f_nc )                 // Unused
        , .p1_addr_f            ( p6_lba_tot_enq_cnt_rmw_pipe_addr_f_nc )               // Unused
        , .p1_data_f            ( p6_lba_tot_enq_cnt_rmw_pipe_data_f_nc )               // Unused

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_tot_enq_cnt_rmw_pipe_v_f_nc )                  // Unused
        , .p2_rw_f              ( p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd )            // Used to determine upd_v
        , .p2_addr_f            ( p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.qid )               // Unused
        , .p2_data_f            ( p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p7_lba_tot_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_tot_enq_cnt_upd )
        , .p3_v_f               ( p8_lba_tot_enq_cnt_rmw_pipe_v_f_nc )                  // Unused
        , .p3_rw_f              ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd )            // Used for res_chk_en
        , .p3_addr_f            ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.qid )               // Unused
        , .p3_data_f            ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.data )              // Used for res_chk

        // mem intf
        , .mem_write            ( cfgsc_func_qid_naldb_tot_enq_cnt_mem_we )
        , .mem_read             ( func_qid_naldb_tot_enq_cnt_mem_re )
        , .mem_write_addr       ( cfgsc_func_qid_naldb_tot_enq_cnt_mem_waddr )
        , .mem_read_addr        ( func_qid_naldb_tot_enq_cnt_mem_raddr )
        , .mem_write_data       ( cfgsc_func_qid_naldb_tot_enq_cnt_mem_wdata )
        , .mem_read_data        ( func_qid_naldb_tot_enq_cnt_mem_rdata )
    ) ;

hqm_AW_residue_add i_lba_tot_enq_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .r                    ( p7_lba_tot_enq_cnt_res_p1 )
) ;

assign p7_lba_tot_enq_cnt_p1            = p7_lba_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt + 64'h1 ;          // wrap

assign p7_lba_tot_enq_cnt_upd.cnt       = p7_lba_tot_enq_cnt_p1 ;
assign p7_lba_tot_enq_cnt_upd.cnt_res   = p7_lba_tot_enq_cnt_res_p1 ;

assign p8_lba_tot_enq_cnt_res_chk_en    = p9_lba_ctrl_pipe.en & ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ARCH_CNT_WIDTH ) ) i_lba_tot_enq_cnt_res_chk (
          .r                    ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .d                    ( p8_lba_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt )
        , .e                    ( p8_lba_tot_enq_cnt_res_chk_en )
        , .err                  ( p9_lba_tot_enq_cnt_res_err_nxt )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for lba total schedule count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_ARCH_CNT_MEM_WIDTH )
) i_lba_tot_sch_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_tot_sch_cnt_rmw_pipe_status_nc )                          // Unused, same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_tot_sch_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_tot_sch_cnt_rmw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_tot_sch_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_tot_sch_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p0_rw_f              ( p5_lba_tot_sch_cnt_rmw_pipe_rw_f_nc )         // Unused
        , .p0_addr_f            ( p5_lba_tot_sch_cnt_rmw_pipe_addr_f_nc )       // Unused
        , .p0_data_f            ( p5_lba_tot_sch_cnt_rmw_pipe_datav_f_nc )      // Unused

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_tot_sch_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p1_rw_f              ( p6_lba_tot_sch_cnt_rmw_pipe_rw_f_nc )         // Unused
        , .p1_addr_f            ( p6_lba_tot_sch_cnt_rmw_pipe_addr_f_nc )       // Unused
        , .p1_data_f            ( p6_lba_tot_sch_cnt_rmw_pipe_datav_f_nc )      // Unused

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_tot_sch_cnt_rmw_pipe_v_f_nc )
        , .p2_rw_f              ( p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd )    // Used to determine upd_v
        , .p2_addr_f            ( p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.cq )        // Unused
        , .p2_data_f            ( p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p6_lba_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p7_lba_tot_sch_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_tot_sch_cnt_upd )
        , .p3_v_f               ( p8_lba_tot_sch_cnt_rmw_pipe_v_f_nc )
        , .p3_rw_f              ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd )    // Used for res_chk_en
        , .p3_addr_f            ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.cq )        // Unused
        , .p3_data_f            ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.data )      // Used for res_chk

        // mem intf
        , .mem_write            ( cfgsc_func_cq_ldb_tot_sch_cnt_mem_we )
        , .mem_read             ( func_cq_ldb_tot_sch_cnt_mem_re )
        , .mem_write_addr       ( cfgsc_func_cq_ldb_tot_sch_cnt_mem_waddr )
        , .mem_read_addr        ( func_cq_ldb_tot_sch_cnt_mem_raddr )
        , .mem_write_data       ( cfgsc_func_cq_ldb_tot_sch_cnt_mem_wdata )
        , .mem_read_data        ( func_cq_ldb_tot_sch_cnt_mem_rdata )
    ) ;

hqm_AW_residue_add i_lba_tot_sch_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .r                    ( p7_lba_tot_sch_cnt_res_p1 )
) ;

assign p7_lba_tot_sch_cnt_p1                    = p7_lba_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt + 64'h1 ;          // wrap

assign p7_lba_tot_sch_cnt_upd.cnt       = p7_lba_tot_sch_cnt_p1 ;
assign p7_lba_tot_sch_cnt_upd.cnt_res   = p7_lba_tot_sch_cnt_res_p1 ;

assign p8_lba_tot_sch_cnt_res_chk_en    = p9_lba_ctrl_pipe.en & ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ARCH_CNT_WIDTH ) ) i_lba_tot_sch_cnt_res_chk (
          .r                    ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .d                    ( p8_lba_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt )
        , .e                    ( p8_lba_tot_sch_cnt_res_chk_en )
        , .err                  ( p9_lba_tot_sch_cnt_res_err_nxt )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for lba total enqueue count
hqm_AW_rmw_mem_4pipe_waddr #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID_ENQ_CNT_WIDTH )
) i_lba_max_enq_depth_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_max_enq_depth_rmw_pipe_status_nc )                        // Unused, same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_max_enq_depth_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_max_enq_depth_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_max_enq_depth_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_max_enq_depth_rmw_pipe_v_f_nc )                // Unused
        , .p0_rw_f              ( p5_lba_max_enq_depth_rmw_pipe_rw_f_nc )               // Unused
        , .p0_addr_f            ( p5_lba_max_enq_depth_rmw_pipe_addr_f_nc )             // Unused
        , .p0_data_f            ( p5_lba_max_enq_depth_rmw_pipe_data_f_nc )             // Unused

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_max_enq_depth_rmw_pipe_v_f_nc )                // Unused
        , .p1_rw_f              ( p6_lba_max_enq_depth_rmw_pipe_rw_f_nc )               // Unused
        , .p1_addr_f            ( p6_lba_max_enq_depth_rmw_pipe_addr_f_nc )             // Unused
        , .p1_data_f            ( p6_lba_max_enq_depth_rmw_pipe_data_f_nc )             // Unused

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_max_enq_depth_rmw_pipe_v_f_nc )                // Unused
        , .p2_rw_f              ( p7_lba_max_enq_depth_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p7_lba_max_enq_depth_rmw_pipe_f.qid )
        , .p2_data_f            ( p7_lba_max_enq_depth_rmw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypdata_sel_nxt   ( p7_lba_max_enq_depth_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_max_enq_depth_upd )
        , .p3_bypaddr_sel_nxt   ( p7_lba_max_enq_depth_upd_v )
        , .p3_bypaddr_nxt       ( p7_lba_max_enq_depth_rmw_pipe_f.qid )
        , .p3_v_f               ( p8_lba_max_enq_depth_rmw_pipe_v_f_nc )                // Unused
        , .p3_rw_f              ( p8_lba_max_enq_depth_rmw_pipe_f_nc.rw_cmd )           // Unused
        , .p3_addr_f            ( p8_lba_max_enq_depth_rmw_pipe_f_nc.qid )              // Unused
        , .p3_data_f            ( p8_lba_max_enq_depth_rmw_pipe_f_nc.data )             // Unused

        // mem intf
        , .mem_write            ( func_qid_naldb_max_depth_mem_we )
        , .mem_read             ( func_qid_naldb_max_depth_mem_re )
        , .mem_write_addr       ( func_qid_naldb_max_depth_mem_waddr )
        , .mem_read_addr        ( func_qid_naldb_max_depth_mem_raddr )
        , .mem_write_data       ( func_qid_naldb_max_depth_mem_wdata )
        , .mem_read_data        ( func_qid_naldb_max_depth_mem_rdata )
) ;

assign p7_lba_enq_cnt_gt_max_depth           = ( p7_lba_qid_enq_cnt_upd.cnt > p7_lba_max_enq_depth_rmw_pipe_f.data ) ;
assign p7_lba_max_enq_depth_upd              = p7_lba_qid_enq_cnt_upd.cnt ;

//-------------------------------------------------------------------------------------------------
// cq_if_cnt, cq_if_lim, cq_if_thr, tot_if_cnt

always_comb begin
  if ( p4_lba_ctrl_pipe_v_f & ( p4_lba_ctrl_pipe_f.cq_cmp_v | p4_lba_ctrl_pipe_f.sch_v ) ) begin
    p5_lba_cq_if_cnt_rmw_pipe_nxt.rw_cmd        = HQM_AW_RMWPIPE_RMW ;          // Only (conditionally) do rmw if cmp or sch
    p5_lba_cq_if_lim_rw_pipe_nxt.rw_cmd         = HQM_AW_RWPIPE_READ ;
    p5_lba_cq_if_thr_rw_pipe_nxt.rw_cmd         = HQM_AW_RWPIPE_READ ;
  end
  else begin
    p5_lba_cq_if_cnt_rmw_pipe_nxt.rw_cmd        = HQM_AW_RMWPIPE_NOOP ;
    p5_lba_cq_if_lim_rw_pipe_nxt.rw_cmd         = HQM_AW_RWPIPE_NOOP ;
    p5_lba_cq_if_thr_rw_pipe_nxt.rw_cmd         = HQM_AW_RWPIPE_NOOP ;
  end
  if ( p4_lba_ctrl_pipe_f.sch_v ) begin
    p5_lba_cq_if_cnt_rmw_pipe_nxt.cq            = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
    p5_lba_cq_if_lim_rw_pipe_nxt.cq             = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
    p5_lba_cq_if_thr_rw_pipe_nxt.cq             = p4_lba_ctrl_pipe_f_pcm ? { p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0 } : p4_lba_ctrl_pipe_f.sch_cq ;
  end
  else begin
    p5_lba_cq_if_cnt_rmw_pipe_nxt.cq            = p4_lba_ctrl_pipe_f.cmp_cq ;
    p5_lba_cq_if_lim_rw_pipe_nxt.cq             = p4_lba_ctrl_pipe_f.cmp_cq ;
    p5_lba_cq_if_thr_rw_pipe_nxt.cq             = p4_lba_ctrl_pipe_f.cmp_cq ;
  end
  p5_lba_cq_if_cnt_rmw_pipe_nxt.data            = { $bits ( lsp_lb_cq_if_cnt_t ) { 1'b0 } } ;   // Unused - cfg write done elsewhere
  p5_lba_cq_if_lim_rw_pipe_nxt.data             = { $bits ( lsp_lb_cq_if_lim_t ) { 1'b0 } } ;   // Unused - cfg write done elsewhere
  p5_lba_cq_if_thr_rw_pipe_nxt.data             = { $bits ( lsp_lb_cq_if_lim_t ) { 1'b0 } } ;   // Unused - cfg write done elsewhere
end // always

hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_LB_CQ_IF_CNT_MEM_WIDTH )
) i_lba_cq_if_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq_if_cnt_rmw_pipe_status_nc )            // Unused, same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_cq_if_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_cq_if_cnt_rmw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_cq_if_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p5_lba_cq_if_cnt_rmw_pipe_v_f_nc )            // Unused, same as cq_tok_cnt pipe
        , .p0_rw_f              ( p5_lba_cq_if_cnt_rmw_pipe_rw_f_nc )           // Unused
        , .p0_addr_f            ( p5_lba_cq_if_cnt_rmw_pipe_addr_f_nc )         // Unused
        , .p0_data_f            ( p5_lba_cq_if_cnt_rmw_pipe_data_f_nc )         // Unused

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_cq_if_cnt_rmw_pipe_v_f_nc )            // Unused, same as cq_tok_cnt pipe
        , .p1_rw_f              ( p6_lba_cq_if_cnt_rmw_pipe_rw_f_nc )           // Unused
        , .p1_addr_f            ( p6_lba_cq_if_cnt_rmw_pipe_addr_f_nc )         // Unused
        , .p1_data_f            ( p6_lba_cq_if_cnt_rmw_pipe_data_f_nc )         // Unused

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_cq_if_cnt_rmw_pipe_v_f_nc )            // Unused, same as cq_tok_cnt pipe
        , .p2_rw_f              ( p7_lba_cq_if_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p7_lba_cq_if_cnt_rmw_pipe_f.cq )
        , .p2_data_f            ( p7_lba_cq_if_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p7_lba_cq_if_cnt_upd_v )
        , .p3_bypdata_nxt       ( p7_lba_cq_if_cnt_upd_cnt )
        , .p3_v_f               ( p8_lba_cq_if_cnt_rmw_pipe_v_f_nc )
        , .p3_rw_f              ( p8_lba_cq_if_cnt_rmw_pipe_f_pnc.rw_cmd )      // Unused
        , .p3_addr_f            ( p8_lba_cq_if_cnt_rmw_pipe_f_pnc.cq )          // Used for error rid
        , .p3_data_f            ( p8_lba_cq_if_cnt_rmw_pipe_f_pnc.data )        // Unused


        // mem intf
        , .mem_write            ( func_cq_ldb_inflight_count_mem_we )
        , .mem_read             ( func_cq_ldb_inflight_count_mem_re )
        , .mem_write_addr       ( func_cq_ldb_inflight_count_mem_waddr )
        , .mem_read_addr        ( func_cq_ldb_inflight_count_mem_raddr )
        , .mem_write_data       ( func_cq_ldb_inflight_count_mem_wdata )
        , .mem_read_data        ( func_cq_ldb_inflight_count_mem_rdata )
) ;

hqm_AW_residue_add i_lba_cq_if_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_cq_if_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_cq_if_cnt_res_p1 )
) ;
hqm_AW_residue_add i_lba_tot_if_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_tot_if_cnt_f.cnt_res )
        , .r                    ( p7_lba_tot_if_cnt_res_p1 )
) ;

hqm_AW_residue_sub i_lba_cq_if_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_cq_if_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p7_lba_cq_if_cnt_res_m1 )
) ;
hqm_AW_residue_sub i_lba_tot_if_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p7_lba_tot_if_cnt_f.cnt_res )
        , .r                    ( p7_lba_tot_if_cnt_res_m1 )
) ;


assign { p7_lba_cq_if_cnt_p1_carry , p7_lba_cq_if_cnt_p1 }      = { 1'b0 , p7_lba_cq_if_cnt_rmw_pipe_f.data.cnt } + 13'h1 ;
assign { p7_lba_cq_if_cnt_m1_borrow , p7_lba_cq_if_cnt_m1 }     = { 1'b0 , p7_lba_cq_if_cnt_rmw_pipe_f.data.cnt } - 13'h1 ;

assign { p7_lba_tot_if_cnt_p1_carry , p7_lba_tot_if_cnt_p1 }    = { 1'b0 , p7_lba_tot_if_cnt_f.cnt } + 13'h1 ;
assign { p7_lba_tot_if_cnt_m1_borrow , p7_lba_tot_if_cnt_m1 }   = { 1'b0 , p7_lba_tot_if_cnt_f.cnt } - 13'h1 ;

always_comb begin
  p7_lba_cq_if_cnt_oflow_cond                   = 1'b0 ;
  p7_lba_cq_if_cnt_uflow_cond                   = 1'b0 ;
  p7_lba_tot_if_cnt_oflow_cond                  = 1'b0 ;
  p7_lba_tot_if_cnt_uflow_cond                  = 1'b0 ;
  if ( p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.sch_atm_v ) begin
    if ( p7_lba_cq_if_cnt_p1_carry ) begin
      p7_lba_cq_if_cnt_upd_cnt                  = p7_lba_cq_if_cnt_rmw_pipe_f.data ;    // Saturate, no residue error
      p7_lba_cq_if_cnt_oflow_cond               = 1'b1 ;
    end
    else begin
      p7_lba_cq_if_cnt_upd_cnt.cnt              = p7_lba_cq_if_cnt_p1 ;
      p7_lba_cq_if_cnt_upd_cnt.cnt_res          = p7_lba_cq_if_cnt_res_p1 ;
    end
    if ( p7_lba_tot_if_cnt_p1_carry ) begin
      p7_lba_tot_if_cnt_upd_cnt                 = p7_lba_tot_if_cnt_f ;                 // Saturate, no residue error
      p7_lba_tot_if_cnt_oflow_cond              = 1'b1 ;
    end
    else begin
      p7_lba_tot_if_cnt_upd_cnt.cnt             = p7_lba_tot_if_cnt_p1 ;
      p7_lba_tot_if_cnt_upd_cnt.cnt_res         = p7_lba_tot_if_cnt_res_p1 ;
    end
  end
  else begin
    if ( p7_lba_ctrl_pipe_f.cmp_cq_no_dec ) begin
      p7_lba_cq_if_cnt_upd_cnt                  = p7_lba_cq_if_cnt_rmw_pipe_f.data ;    // No change 
    end
    else if ( p7_lba_cq_if_cnt_m1_borrow ) begin
      p7_lba_cq_if_cnt_upd_cnt                  = p7_lba_cq_if_cnt_rmw_pipe_f.data ;    // Saturate, no residue error
      p7_lba_cq_if_cnt_uflow_cond               = 1'b1 ;
    end
    else begin
      p7_lba_cq_if_cnt_upd_cnt.cnt              = p7_lba_cq_if_cnt_m1 ;
      p7_lba_cq_if_cnt_upd_cnt.cnt_res          = p7_lba_cq_if_cnt_res_m1 ;
    end
    if ( p7_lba_ctrl_pipe_f.cmp_cq_no_dec ) begin
      p7_lba_tot_if_cnt_upd_cnt                 = p7_lba_tot_if_cnt_f ;                 // Saturate, no residue error
    end
    else if ( p7_lba_tot_if_cnt_m1_borrow ) begin
      p7_lba_tot_if_cnt_upd_cnt                 = p7_lba_tot_if_cnt_f ;                 // Saturate, no residue error
      p7_lba_tot_if_cnt_uflow_cond              = 1'b1 ;
    end
    else begin
      p7_lba_tot_if_cnt_upd_cnt.cnt             = p7_lba_tot_if_cnt_m1 ;
      p7_lba_tot_if_cnt_upd_cnt.cnt_res         = p7_lba_tot_if_cnt_res_m1 ;
    end
  end
end // always

assign p7_lba_cq_if_cnt_upd_lt_lim              = ( p7_lba_cq_if_cnt_upd_cnt.cnt         <  p7_lba_cq_if_lim_rw_pipe_f_pnc.data.lim ) ;
assign p7_lba_cq_if_cnt_upd_le_thr              = ( p7_lba_cq_if_cnt_upd_cnt.cnt         <= p7_lba_cq_if_thr_rw_pipe_f_pnc.data.thr ) ;
assign p7_lba_cq_if_cnt_upd_gt_0                = | p7_lba_cq_if_cnt_upd_cnt.cnt ;

assign p7_lba_tot_if_cnt_upd_lt_lim             = ( p7_lba_tot_if_cnt_upd_cnt.cnt  < cfg_cq_ldb_tot_inflight_limit_f ) ;

// Should be correctly adjusted as part of a successful vas reset drain
always_comb begin
  cfg_cq_ldb_tot_inflight_count_nxt             = cfg_cq_ldb_tot_inflight_count_f ;
  if ( p7_lba_cq_if_cnt_upd_v ) begin
    cfg_cq_ldb_tot_inflight_count_nxt           = p7_lba_tot_if_cnt_upd_cnt ;
  end
end // always

assign p7_lba_tot_if_cnt_f                      = cfg_cq_ldb_tot_inflight_count_f ;


assign p7_lba_cq_if_cnt_res_chk_en              = p7_lba_cq_if_cnt_upd_v ;
assign p7_lba_cq_if_lim_par_chk_en              = p7_lba_cq_if_cnt_res_chk_en ;
assign p7_lba_cq_if_thr_par_chk_en              = p7_lba_cq_if_cnt_res_chk_en ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LB_CQ_IF_CNT_WIDTH ) ) i_lba_tot_if_cnt_res_chk (
          .r                    ( cfg_cq_ldb_tot_inflight_count_f.cnt_res )
        , .d                    ( cfg_cq_ldb_tot_inflight_count_f.cnt )
        , .e                    ( p7_lba_cq_if_cnt_upd_v )
        , .err                  ( p7_lba_tot_if_cnt_res_err_cond )
) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LB_CQ_IF_CNT_WIDTH ) ) i_lba_cq_if_cnt_res_chk (
          .r                    ( p7_lba_cq_if_cnt_upd_cnt.cnt_res )
        , .d                    ( p7_lba_cq_if_cnt_upd_cnt.cnt )
        , .e                    ( p7_lba_cq_if_cnt_res_chk_en )
        , .err                  ( p7_lba_cq_if_cnt_res_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_LB_CQ_IF_LIM_WIDTH ) ) i_lba_cq_if_lim_par_chk (
          .p                    ( p7_lba_cq_if_lim_rw_pipe_f_pnc.data.lim_p )
        , .d                    ( p7_lba_cq_if_lim_rw_pipe_f_pnc.data.lim )
        , .e                    ( p7_lba_cq_if_lim_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_cq_if_lim_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_LB_CQ_IF_THR_WIDTH ) ) i_lba_cq_if_thr_par_chk (
          .p                    ( p7_lba_cq_if_thr_rw_pipe_f_pnc.data.thr_p )
        , .d                    ( p7_lba_cq_if_thr_rw_pipe_f_pnc.data.thr )
        , .e                    ( p7_lba_cq_if_thr_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_cq_if_thr_par_err_cond )
) ;

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_LB_CQ_IF_LIM_MEM_WIDTH )
    ) i_lba_cq_if_lim_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq_if_lim_rw_pipe_status_nc )             // Unused: same as lba_cq_if_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_cq_if_lim_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_cq_if_lim_rw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_cq_if_lim_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_cq_if_lim_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p0_rw_f              ( p5_lba_cq_if_lim_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_cq_if_lim_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_cq_if_lim_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_cq_if_lim_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p1_rw_f              ( p6_lba_cq_if_lim_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_cq_if_lim_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_cq_if_lim_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_cq_if_lim_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe 
        , .p2_rw_f              ( p7_lba_cq_if_lim_rw_pipe_f_pnc.rw_cmd )       // Unused
        , .p2_addr_f            ( p7_lba_cq_if_lim_rw_pipe_f_pnc.cq )           // Unused
        , .p2_data_f            ( p7_lba_cq_if_lim_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_cq_if_lim_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p3_rw_f              ( p8_lba_cq_if_lim_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p8_lba_cq_if_lim_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p8_lba_cq_if_lim_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cfg_cq_ldb_inflight_limit_mem_we )
        , .mem_read             ( func_cfg_cq_ldb_inflight_limit_mem_re )
        , .mem_addr             ( func_cfg_cq_ldb_inflight_limit_mem_addr )
        , .mem_write_data       ( func_cfg_cq_ldb_inflight_limit_mem_wdata )
        , .mem_read_data        ( func_cfg_cq_ldb_inflight_limit_mem_rdata )
) ;

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WIDTH                ( HQM_LSP_LB_CQ_IF_THR_MEM_WIDTH )
    ) i_lba_cq_if_thr_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_cq_if_thr_rw_pipe_status_nc )             // Unused: same as lba_cq_if_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_cq_if_thr_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_cq_if_thr_rw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p5_lba_cq_if_thr_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_cq_if_thr_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p0_rw_f              ( p5_lba_cq_if_thr_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_cq_if_thr_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_cq_if_thr_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_cq_if_thr_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p1_rw_f              ( p6_lba_cq_if_thr_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_cq_if_thr_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_cq_if_thr_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_cq_if_thr_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe 
        , .p2_rw_f              ( p7_lba_cq_if_thr_rw_pipe_f_pnc.rw_cmd )       // Unused
        , .p2_addr_f            ( p7_lba_cq_if_thr_rw_pipe_f_pnc.cq )           // Unused
        , .p2_data_f            ( p7_lba_cq_if_thr_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_cq_if_thr_rw_pipe_v_f_nc )             // Unused: same as cq_tok_cnt pipe
        , .p3_rw_f              ( p8_lba_cq_if_thr_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p8_lba_cq_if_thr_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p8_lba_cq_if_thr_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cfg_cq_ldb_inflight_threshold_mem_we )
        , .mem_read             ( func_cfg_cq_ldb_inflight_threshold_mem_re )
        , .mem_addr             ( func_cfg_cq_ldb_inflight_threshold_mem_addr )
        , .mem_write_data       ( func_cfg_cq_ldb_inflight_threshold_mem_wdata )
        , .mem_read_data        ( func_cfg_cq_ldb_inflight_threshold_mem_rdata )
) ;

// Purpose of qid parity checking is just to check the input qid.  Just use the copy in rmw pipe for qid[0].

assign p7_lba_inp_enq_qid_par_chk_en    = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.enq_v ;
assign p7_lba_inp_cmp_qid_par_chk_en    = p7_lba_ctrl_pipe_v_f & ( p7_lba_ctrl_pipe_f.qid_cmp_v | p7_lba_ctrl_pipe_f.qid_if_dec_v ) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_lba_inp_enq_qid_par_chk (
          .p                    ( p7_lba_ctrl_pipe_f.enq_qid_p )
        , .d                    ( p7_lba_qid_enq_cnt_rmw_pipe_f.qid )
        , .e                    ( p7_lba_inp_enq_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_inp_enq_qid_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_lba_inp_cmp_qid_par_chk (
          .p                    ( p7_lba_ctrl_pipe_f.cmp_qid_p )
        , .d                    ( p7_lba_qid_if_cnt_rmw_pipe_f.qid )
        , .e                    ( p7_lba_inp_cmp_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_inp_cmp_qid_par_err_cond )
) ;

assign p7_lba_inp_qid_par_err_cond      = p7_lba_inp_enq_qid_par_err_cond | p7_lba_inp_cmp_qid_par_err_cond ;


// Purpose of cq parity checking is just to check the input cq.

assign p7_lba_inp_tok_cq_par_chk_en     = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.tok_v ;
assign p7_lba_inp_cmp_cq_par_chk_en     = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.cq_cmp_v ;

hqm_AW_parity_check # ( .WIDTH ( HQM_NUM_LB_CQB2 ) ) i_lba_inp_tok_cq_par_chk (
          .p                    ( p7_lba_ctrl_pipe_f.tok_cq_p )
        , .d                    ( p7_lba_cq_tok_cnt_rmw_pipe_f.cq )
        , .e                    ( p7_lba_inp_tok_cq_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_inp_tok_cq_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_NUM_LB_CQB2 ) ) i_lba_inp_cmp_cq_par_chk (
          .p                    ( p7_lba_ctrl_pipe_f.cmp_cq_p )
        , .d                    ( p7_lba_cq_if_cnt_rmw_pipe_f.cq )
        , .e                    ( p7_lba_inp_cmp_cq_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_inp_cmp_cq_par_err_cond )
) ;

assign p7_lba_inp_cq_par_err_cond       = p7_lba_inp_tok_cq_par_err_cond | p7_lba_inp_cmp_cq_par_err_cond ;

//-------------------------------------------------------------------------------------------------
// qid2cqidix  Needed for updating per qidix-based vectors for "has work",
// for (nalb) enqueues, lb schedules and qid completions.
// p0/1/2/3 for the rw_pipe is lba pipe levels p5/p6/p7/p8
// Only written by config.

always_comb begin
  if ( p4_lba_sch_arb_winner_v | p4_lba_ctrl_pipe_f.enq_v | p4_lba_ctrl_pipe_f.qid_cmp_v | p4_lba_ctrl_pipe_f.qid_if_dec_v ) begin
    p5_lba_qid2cqidix_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_READ ;                          // Don't do lookup unless necessary
  end
  else begin
    p5_lba_qid2cqidix_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_NOOP ;
  end
  // Note: this is (only reason) why can't simultaneously do enq and cmp
  if ( p4_lba_sch_arb_winner_v )
    p5_lba_qid2cqidix_rw_pipe_nxt.qid             = p4_lba_sch_arb_winner_qid ;
  else if ( p4_lba_ctrl_pipe_f.enq_v )
    p5_lba_qid2cqidix_rw_pipe_nxt.qid             = p4_lba_ctrl_pipe_f.enq_qid ;
  else
    p5_lba_qid2cqidix_rw_pipe_nxt.qid             = p4_lba_ctrl_pipe_f.cmp_qid ;
  p5_lba_qid2cqidix_rw_pipe_nxt.data            = { $bits ( lsp_cfg_qid2cqidix_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
end // always

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID2CQIDIX_MEM_WIDTH )
) i_lba_qid2cqidix_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_qid2cqidix_rw_pipe_status )

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_qid2cqidix_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_qid2cqidix_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_qid2cqidix_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_qid2cqidix_rw_pipe_v_f_nc )                    // Unused: same as lba_cq_tok_cnt
        , .p0_rw_f              ( p5_lba_qid2cqidix_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_qid2cqidix_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_qid2cqidix_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_qid2cqidix_rw_pipe_v_f_nc )                    // Unused: same as lba_cq_tok_cnt
        , .p1_rw_f              ( p6_lba_qid2cqidix_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_qid2cqidix_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_qid2cqidix_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_qid2cqidix_rw_pipe_v_f_nc )
        , .p2_rw_f              ( p7_lba_qid2cqidix_rw_pipe_f.rw_cmd )                  // Used to distinguish parity check
        , .p2_addr_f            ( p7_lba_qid2cqidix_rw_pipe_f.qid )                     // Unused by hw, used by non-synth checking code
        , .p2_data_f            ( p7_lba_qid2cqidix_rw_pipe_f.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_qid2cqidix_rw_pipe_v_f_nc )
        , .p3_rw_f              ( p8_lba_qid2cqidix_rw_pipe_f_nc.rw_cmd )               // Unused
        , .p3_addr_f            ( p8_lba_qid2cqidix_rw_pipe_f_nc.qid )                  // Unused
        , .p3_data_f            ( p8_lba_qid2cqidix_rw_pipe_f_nc.data )                 // Unused


        // mem intf
        , .mem_write            ( func_cfg_qid_ldb_qid2cqidix_mem_we )                  // Never used - cfg writes done elsewhere
        , .mem_read             ( func_cfg_qid_ldb_qid2cqidix_mem_re )
        , .mem_addr             ( func_cfg_qid_ldb_qid2cqidix_mem_addr )
        , .mem_write_data       ( func_cfg_qid_ldb_qid2cqidix_mem_wdata )               // Never used - cfg writes done elsewhere
        , .mem_read_data        ( func_cfg_qid_ldb_qid2cqidix_mem_rdata )
) ;

assign p7_lba_qid2cqidix_v              = p7_lba_qid2cqidix_rw_pipe_f.data.qidixv ;

assign p7_lba_qid2cqidix_p              = p7_lba_qid2cqidix_rw_pipe_f.data.parity ;     // 16 bits

assign p7_lba_qid2cqidix_par_chk_en     = p7_lba_ctrl_pipe_v_f & ( p7_lba_qid2cqidix_rw_pipe_f.rw_cmd == HQM_AW_RWPIPE_READ ) ;

// Configuration error: cq2qid config inconsistent with qid2cqidix - if a qid was selected for scheduling, at least one of the
// qidix for that cq must = 1.
assign p7_lba_qid2cqidix_ix             = p7_lba_ctrl_pipe_f_pcm ? { p7_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , p7_lba_ctrl_pipe_f.sch_qidix_msb , 3'h0 } : { p7_lba_ctrl_pipe_f.sch_cq , 3'h0 } ;
assign p7_lba_qid2cqidix_v_qidix        = p7_lba_qid2cqidix_v [ p7_lba_qid2cqidix_ix +: 8 ] ; 
assign p7_lba_qid2cqidix_sch_v_err_cond = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.sch_v & ~ ( | p7_lba_qid2cqidix_v_qidix ) ;
assign p7_lba_qid2cqidix_enq_v_err_cond = p7_lba_ctrl_pipe_v_f & p7_lba_ctrl_pipe_f.enq_v & ~ ( | p7_lba_qid2cqidix_v ) ;       // 512-bit OR

generate
  for ( genvar gi = 0 ; gi < 16 ; gi = gi + 1 ) begin: gen_qid2cqidix_par_chk
    hqm_AW_parity_check # ( .WIDTH ( 32 ) ) i_lba_qid2cqidix_par_chk (
          .p                    ( p7_lba_qid2cqidix_p [gi] )
        , .d                    ( p7_lba_qid2cqidix_v [ ( gi * 32 ) +: 32 ] )
        , .e                    ( p7_lba_qid2cqidix_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_qid2cqidix_par_err_cond [gi] )
    ) ;
  end
endgenerate

always_comb begin
  // Don't hold - 1-clock pulse to report
  p8_lba_qid2cqidix_par_err_nxt        = 16'h0 ;
  if ( p7_lba_ctrl_pipe_v_f & ~ p8_lba_ctrl_pipe.hold ) begin
    p8_lba_qid2cqidix_par_err_nxt      = p7_lba_qid2cqidix_par_err_cond ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p8_lba_qid2cqidix_par_err_f        <= 16'h0 ;
  end
  else begin
    p8_lba_qid2cqidix_par_err_f        <= p8_lba_qid2cqidix_par_err_nxt ;
  end
end // always

assign p8_lba_qid2cqidix_par_err_any  = ( | p8_lba_qid2cqidix_par_err_f ) | cfg_error_inject_f [ 4 ] ;

//-------------------------------------------------------------------------------------------------
// RR arbiter index state for atm, nalb and ldb arbiters.  For each CQ, 3-bit index per priority bin,
// plus 3-bit count per qidix (weight).  Separate storage for nalb and atm - want to support the ability
// for a particular type to burst without interrupting each other.
// p0/1/2 for the rw_pipe is lba pipe levels p1/p2/p3 for atm and nalb.

assign p4_lba_nalb_sch_arb_update               = p4_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe_f.sch_v & ~ p4_lba_ctrl_pipe.hold & ~ p4_lba_sch_arb_atm ;
assign p4_lba_atm_sch_arb_update                = p4_lba_ctrl_pipe_v_f & p4_lba_ctrl_pipe_f.sch_v & ~ p4_lba_ctrl_pipe.hold &   p4_lba_sch_arb_atm ;

assign p1_lba_ctrl_pipe_nxt_sch_pcq             = p1_lba_ctrl_pipe_nxt.sch_cq >> 1 ;
assign p1_lba_ctrl_pipe_f_sch_pcq               = p1_lba_ctrl_pipe_f.sch_cq >> 1 ;
assign p4_lba_ctrl_pipe_f_sch_pcq               = p4_lba_ctrl_pipe_f.sch_cq >> 1 ;

// Max 1 schedule per 8 clocks, no need for internal bypasses, better static timing with rf pipe.
hqm_AW_rf_mem_3pipe_core #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ >> 1 )
        , .WIDTH                ( HQM_LSP_LB_ARBINDEX_MEM_WIDTH )
) i_cq_nalb_pri_arbindex_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_nalb_pri_arbindex_pipe_status )

        // Read pipe
        , .p0_v_nxt             ( p1_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rd_v_nxt          ( p0_lba_pop_cq [0] )
        , .p0_addr_nxt          ( p1_lba_ctrl_pipe_nxt_sch_pcq )
        , .p0_hold              ( p1_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p1_lba_nalb_index_v_f_nc )
        , .p0_addr_f            ( p1_lba_nalb_index_rw_pipe_addr_f_nc )

        , .p1_hold              ( p2_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p2_lba_nalb_index_v_f_nc )
        , .p1_addr_f            ( p2_lba_nalb_index_rw_pipe_addr_f_nc )

        , .p2_hold              ( p3_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p3_lba_nalb_index_v_f_nc )
        , .p2_addr_f            ( p3_lba_nalb_index_rw_pipe_addr_f_nc )
        , .p2_data_f            ( p3_lba_nalb_index_rw_pipe_data_f )
        , .p2_data_nobyp_f      ( p3_lba_nalb_index_rw_pipe_data_nobyp_f_nc )   // Unused
        , .p2_byp_v_nxt         ( 1'b0 )                                        // Unused
        , .p2_bypdata_nxt       ( { HQM_LSP_LB_ARBINDEX_MEM_WIDTH { 1'b0 } } )  // Unused

        // Write pipe
        , .pw_v_nxt             ( p4_lba_nalb_sch_arb_update )
        , .pw_addr_nxt          ( p4_lba_ctrl_pipe_f_sch_pcq )
        , .pw_data_nxt          ( p4_lba_nalb_index_rw_pipe_data_struct )
        , .pw_v_f               ( pw_lba_nalb_index_v_f_nc )
        , .pw_addr_f            ( pw_lba_nalb_index_rw_pipe_addr_f_nc )
        , .pw_data_f            ( pw_lba_nalb_index_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cq_nalb_pri_arbindex_mem_we )
        , .mem_read             ( func_cq_nalb_pri_arbindex_mem_re )
        , .mem_write_addr       ( func_cq_nalb_pri_arbindex_mem_waddr )
        , .mem_read_addr        ( func_cq_nalb_pri_arbindex_mem_raddr )
        , .mem_write_data       ( func_cq_nalb_pri_arbindex_mem_wdata )
        , .mem_read_data        ( func_cq_nalb_pri_arbindex_mem_rdata )
) ;

always_comb begin
  p3_lba_nalb_index_rw_pipe_data_struct         = p3_lba_nalb_index_rw_pipe_data_f ;
  p3_lba_nalb_index_rw_pipe_data_odd.counts     = p3_lba_nalb_index_rw_pipe_data_struct.counts_odd ;
  p3_lba_nalb_index_rw_pipe_data_odd.indexes    = p3_lba_nalb_index_rw_pipe_data_struct.indexes_odd ;
  p3_lba_nalb_index_rw_pipe_data_even.counts    = p3_lba_nalb_index_rw_pipe_data_struct.counts_even ;
  p3_lba_nalb_index_rw_pipe_data_even.indexes   = p3_lba_nalb_index_rw_pipe_data_struct.indexes_even ;

  if ( p3_lba_ctrl_pipe_f.sch_cq[0] ) begin
    p3_lba_nalb_index_rw_pipe_data_x.counts     = p3_lba_nalb_index_rw_pipe_data_odd.counts ;
    p3_lba_nalb_index_rw_pipe_data_x.indexes    = p3_lba_nalb_index_rw_pipe_data_odd.indexes ;
    p3_lba_nalb_index_rw_pipe_data_unch.counts  = p3_lba_nalb_index_rw_pipe_data_even.counts ;
    p3_lba_nalb_index_rw_pipe_data_unch.indexes = p3_lba_nalb_index_rw_pipe_data_even.indexes ;
  end
  else begin
    p3_lba_nalb_index_rw_pipe_data_x.counts     = p3_lba_nalb_index_rw_pipe_data_even.counts ;
    p3_lba_nalb_index_rw_pipe_data_x.indexes    = p3_lba_nalb_index_rw_pipe_data_even.indexes ;
    p3_lba_nalb_index_rw_pipe_data_unch.counts  = p3_lba_nalb_index_rw_pipe_data_odd.counts ;
    p3_lba_nalb_index_rw_pipe_data_unch.indexes = p3_lba_nalb_index_rw_pipe_data_odd.indexes ;
  end
  if ( p3_lba_ctrl_pipe_f_pcm ) begin
    p3_lba_nalb_index_rw_pipe_data_pcm.counts   = { p3_lba_nalb_index_rw_pipe_data_odd.counts
                                                  , p3_lba_nalb_index_rw_pipe_data_even.counts
                                                  } ;
    p3_lba_nalb_index_rw_pipe_data_pcm.indexes  = { p3_lba_nalb_index_rw_pipe_data_odd.indexes [ 7 : 0 ]
                                                  , p3_lba_nalb_index_rw_pipe_data_even.indexes
                                                  } ;
  end
  else begin
    p3_lba_nalb_index_rw_pipe_data_pcm.counts   = { 24'h0, p3_lba_nalb_index_rw_pipe_data_x.counts } ;
    p3_lba_nalb_index_rw_pipe_data_pcm.indexes  = { 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [ 23 : 21 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [ 20 : 18 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [ 17 : 15 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [ 14 : 12 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [ 11 :  9 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [  8 :  6 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [  5 :  3 ]
                                                  , 1'b0, p3_lba_nalb_index_rw_pipe_data_x.indexes [  2 :  0 ]
                                                  } ;
  end
end // always


hqm_AW_rf_mem_3pipe_core #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_CQ >> 1 )
        , .WIDTH                ( HQM_LSP_LB_ARBINDEX_MEM_WIDTH )
) i_cq_atm_pri_arbindex_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_atm_pri_arbindex_pipe_status )

        // Read pipe
        , .p0_v_nxt             ( p1_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rd_v_nxt          ( p0_lba_pop_cq [0] )
        , .p0_addr_nxt          ( p1_lba_ctrl_pipe_nxt_sch_pcq )
        , .p0_hold              ( p1_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p1_lba_atm_index_v_f_nc )
        , .p0_addr_f            ( p1_lba_atm_index_rw_pipe_addr_f_nc )

        , .p1_hold              ( p2_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p2_lba_atm_index_v_f_nc )
        , .p1_addr_f            ( p2_lba_atm_index_rw_pipe_addr_f_nc )

        , .p2_hold              ( p3_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p3_lba_atm_index_v_f_nc )
        , .p2_addr_f            ( p3_lba_atm_index_rw_pipe_addr_f_nc )
        , .p2_data_f            ( p3_lba_atm_index_rw_pipe_data_f )
        , .p2_data_nobyp_f      ( p3_lba_atm_index_rw_pipe_data_nobyp_f_nc )    // Unused
        , .p2_byp_v_nxt         ( 1'b0 )                                        // Unused
        , .p2_bypdata_nxt       ( { HQM_LSP_LB_ARBINDEX_MEM_WIDTH { 1'b0 } } )  // Unused

        // Write pipe
        , .pw_v_nxt             ( p4_lba_atm_sch_arb_update )
        , .pw_addr_nxt          ( p4_lba_ctrl_pipe_f_sch_pcq )
        , .pw_data_nxt          ( p4_lba_atm_index_rw_pipe_data_struct )
        , .pw_v_f               ( pw_lba_atm_index_v_f_nc )
        , .pw_addr_f            ( pw_lba_atm_index_rw_pipe_addr_f_nc )
        , .pw_data_f            ( pw_lba_atm_index_rw_pipe_data_f_nc )

        // mem intf
        , .mem_write            ( func_cq_atm_pri_arbindex_mem_we )
        , .mem_read             ( func_cq_atm_pri_arbindex_mem_re )
        , .mem_write_addr       ( func_cq_atm_pri_arbindex_mem_waddr )
        , .mem_read_addr        ( func_cq_atm_pri_arbindex_mem_raddr )
        , .mem_write_data       ( func_cq_atm_pri_arbindex_mem_wdata )
        , .mem_read_data        ( func_cq_atm_pri_arbindex_mem_rdata )
) ;

always_comb begin
  p3_lba_atm_index_rw_pipe_data_struct          = p3_lba_atm_index_rw_pipe_data_f ;
  p3_lba_atm_index_rw_pipe_data_odd.counts      = p3_lba_atm_index_rw_pipe_data_struct.counts_odd ;
  p3_lba_atm_index_rw_pipe_data_odd.indexes     = p3_lba_atm_index_rw_pipe_data_struct.indexes_odd ;
  p3_lba_atm_index_rw_pipe_data_even.counts     = p3_lba_atm_index_rw_pipe_data_struct.counts_even ;
  p3_lba_atm_index_rw_pipe_data_even.indexes    = p3_lba_atm_index_rw_pipe_data_struct.indexes_even ;

  if ( p3_lba_ctrl_pipe_f.sch_cq[0] ) begin
    p3_lba_atm_index_rw_pipe_data_x.counts      = p3_lba_atm_index_rw_pipe_data_odd.counts ;
    p3_lba_atm_index_rw_pipe_data_x.indexes     = p3_lba_atm_index_rw_pipe_data_odd.indexes ;
    p3_lba_atm_index_rw_pipe_data_unch.counts   = p3_lba_atm_index_rw_pipe_data_even.counts ;
    p3_lba_atm_index_rw_pipe_data_unch.indexes  = p3_lba_atm_index_rw_pipe_data_even.indexes ;
  end
  else begin
    p3_lba_atm_index_rw_pipe_data_x.counts      = p3_lba_atm_index_rw_pipe_data_even.counts ;
    p3_lba_atm_index_rw_pipe_data_x.indexes     = p3_lba_atm_index_rw_pipe_data_even.indexes ;
    p3_lba_atm_index_rw_pipe_data_unch.counts   = p3_lba_atm_index_rw_pipe_data_odd.counts ;
    p3_lba_atm_index_rw_pipe_data_unch.indexes  = p3_lba_atm_index_rw_pipe_data_odd.indexes ;
  end
  if ( p3_lba_ctrl_pipe_f_pcm ) begin
    p3_lba_atm_index_rw_pipe_data_pcm.counts    = { p3_lba_atm_index_rw_pipe_data_odd.counts
                                                  , p3_lba_atm_index_rw_pipe_data_even.counts
                                                  } ;
    p3_lba_atm_index_rw_pipe_data_pcm.indexes   = { p3_lba_atm_index_rw_pipe_data_odd.indexes [ 7 : 0 ]
                                                  , p3_lba_atm_index_rw_pipe_data_even.indexes
                                                  } ;
  end
  else begin
    p3_lba_atm_index_rw_pipe_data_pcm.counts    = { 24'h0, p3_lba_atm_index_rw_pipe_data_x.counts } ;
    p3_lba_atm_index_rw_pipe_data_pcm.indexes   = { 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [ 23 : 21 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [ 20 : 18 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [ 17 : 15 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [ 14 : 12 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [ 11 :  9 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [  8 :  6 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [  5 :  3 ]
                                                  , 1'b0, p3_lba_atm_index_rw_pipe_data_x.indexes [  2 :  0 ]
                                                  } ;
  end
end // always

//-------------------------------------------------------------------------------------------------
// cq_wu_cnt, cq_wu_lim
// Track if a CQ is overworked : sum(scheduled work) > limit

// Note: the FIFOs for qed_lsp_deq and aqed_lsp_deq are instantiated inside hqm_lsp_wu_pipe

hqm_lsp_wu_pipe # (
          .NUM_CQ                                       ( HQM_LSP_ARCH_NUM_LB_CQ )
        , .WU_CNT_WIDTH                                 ( HQM_LSP_LBWU_CQ_WU_CNT_WIDTH )
        , .DEPTH_QED_LSP_DEQ_FIFO                       ( 24 )
        , .DEPTH_AQED_LSP_DEQ_FIFO                      ( 24 )
) i_hqm_lsp_wu_pipe (
          .hqm_gated_clk                                ( hqm_gated_clk )
        , .hqm_gated_rst_n                              ( hqm_gated_rst_n )

        , .cfg_control_qed_lsp_deq_high_pri_wm          ( cfg_control_qed_lsp_deq_high_pri_wm )
        , .cfg_control_aqed_lsp_deq_high_pri_wm         ( cfg_control_aqed_lsp_deq_high_pri_wm )
        , .cfg_control_qe_wt_blk                        ( cfg_control_qe_wt_blk )
        , .cfg_control_qe_wt_frc_v                      ( cfg_control_qe_wt_frc_v )
        , .cfg_control_qe_wt_frc_val                    ( cfg_control_qe_wt_frc_val )
        , .cfg_control_disable_wu_res_chk               ( cfg_control_disable_wu_res_chk )
        , .cfg_qed_deq_pipeline_credit_limit_pnc        ( cfg_qed_deq_pipeline_credit_limit_pnc )
        , .cfg_aqed_deq_pipeline_credit_limit_pnc       ( cfg_aqed_deq_pipeline_credit_limit_pnc )

        , .cfg_mem_addr                                 ( cfg_mem_addr )
        , .cfgsc_cfg_mem_wdata                          ( cfgsc_cfg_mem_wdata )
        , .cfgsc_cfg_mem_wdata_par                      ( cfgsc_cfg_mem_wdata_par )
        , .cfgsc_cfg_mem_wdata_res                      ( cfgsc_cfg_mem_wdata_res )
        , .cfgsc_wu_cfg_data_f                          ( cfgsc_wu_cfg_data_f )

        , .cfgsc_cq_ldb_wu_count_mem_re                 ( cfgsc_cq_ldb_wu_count_mem_re )
        , .cfgsc_cq_ldb_wu_count_mem_we                 ( cfgsc_cq_ldb_wu_count_mem_we )
        , .cfgsc_cfg_cq_ldb_wu_limit_mem_re             ( cfgsc_cfg_cq_ldb_wu_limit_mem_re )
        , .cfgsc_cfg_cq_ldb_wu_limit_mem_we             ( cfgsc_cfg_cq_ldb_wu_limit_mem_we )

        , .cfgsc_wu_count_wr_ack                        ( cfgsc_wu_count_wr_ack )
        , .cfgsc_wu_count_rd_ack                        ( cfgsc_wu_count_rd_ack )
        , .cfgsc_wu_limit_wr_ack                        ( cfgsc_wu_limit_wr_ack )
        , .cfgsc_wu_limit_rd_ack                        ( cfgsc_wu_limit_rd_ack )

        , .qed_lsp_deq_v                                ( qed_lsp_deq_v )
        , .qed_lsp_deq_data_parity                      ( qed_lsp_deq_data.parity )
        , .qed_lsp_deq_data_cq                          ( qed_lsp_deq_data.cq )
        , .qed_lsp_deq_data_qe_wt                       ( qed_lsp_deq_data.qe_wt )

        , .qed_lsp_deq_fifo_of                          ( qed_lsp_deq_fifo_of )
        , .qed_lsp_deq_fifo_uf                          ( qed_lsp_deq_fifo_uf )
        , .qed_lsp_deq_fifo_empty                       ( qed_lsp_deq_fifo_empty)
        , .qed_deq_credit_empty                         ( qed_deq_credit_empty )
        , .qed_deq_credit_error                         ( qed_deq_credit_error )

        , .aqed_lsp_deq_v                               ( aqed_lsp_deq_v )
        , .aqed_lsp_deq_data_parity                     ( aqed_lsp_deq_data.parity )
        , .aqed_lsp_deq_data_cq                         ( aqed_lsp_deq_data.cq )
        , .aqed_lsp_deq_data_qe_wt                      ( aqed_lsp_deq_data.qe_wt )

        , .aqed_lsp_deq_fifo_of                         ( aqed_lsp_deq_fifo_of )
        , .aqed_lsp_deq_fifo_uf                         ( aqed_lsp_deq_fifo_uf )
        , .aqed_lsp_deq_fifo_empty                      ( aqed_lsp_deq_fifo_empty)
        , .aqed_deq_credit_empty                        ( aqed_deq_credit_empty )
        , .aqed_deq_credit_error                        ( aqed_deq_credit_error )

        , .p0_lba_nalb_credit_count_inc                 ( p0_lba_nalb_credit_count_inc )
        , .p4_lba_nalb_credit_count_dec_miss            ( p4_lba_nalb_credit_count_dec_miss )
        , .p4_lba_atm_credit_count_dec_miss             ( p4_lba_atm_credit_count_dec_miss )
        , .qed_deq_credit_afull                         ( qed_deq_credit_afull )
        , .aqed_deq_credit_afull                        ( aqed_deq_credit_afull )

        , .lbi_inp_cq_cmp_cq                            ( lbi_inp_cq_cmp_cq )
        , .lbi_inp_cq_cmp_qe_wt                         ( lbi_inp_cq_cmp_qe_wt )
        , .lbi_inp_cq_cmp_cq_wt_p                       ( lbi_inp_cq_cmp_cq_wt_p )
        , .lbi_cq_cmp_req_taken                         ( lbi_cq_cmp_req_taken )
        , .p0_lba_supress_cq_cmp                        ( p0_lba_supress_cq_cmp )

        , .p0_lba_sch_state_ready_for_work              ( p0_lba_sch_state_ready_for_work ) 

        , .p3_lbwu_cq_wu_cnt_upd_v_func                 ( p3_lbwu_cq_wu_cnt_upd_v_func )

        , .p4_lbwu_cq_wu_cnt_upd_v_f                    ( p4_lbwu_cq_wu_cnt_upd_v_f )
        , .p4_lbwu_cq_wu_cnt_upd_cq_f                   ( p4_lbwu_cq_wu_cnt_upd_cq_f )
        , .p4_lbwu_cq_wu_cnt_upd_gt_lim_f               ( p4_lbwu_cq_wu_cnt_upd_gt_lim_f )

        , .p1_lbwu_ctrl_pipe_v_f                        ( p1_lbwu_ctrl_pipe_v_f )
        , .p2_lbwu_ctrl_pipe_v_f                        ( p2_lbwu_ctrl_pipe_v_f )
        , .p3_lbwu_ctrl_pipe_v_f                        ( p3_lbwu_ctrl_pipe_v_f )
        , .p4_lbwu_ctrl_pipe_v_f                        ( p4_lbwu_ctrl_pipe_v_f )

        , .lbwu_cq_wu_cnt_rmw_pipe_status               ( lbwu_cq_wu_cnt_rmw_pipe_status )

        , .p3_lbwu_cq_wu_cnt_res_err_cond               ( p3_lbwu_cq_wu_cnt_res_err_cond )
        , .p3_lbwu_cq_wu_lim_par_err_cond               ( p3_lbwu_cq_wu_lim_par_err_cond )
        , .p3_lbwu_inp_par_err_cond                     ( p3_lbwu_inp_par_err_cond )

        , .smon_qed_lsp_deq_v                           ( smon_qed_lsp_deq_v )
        , .smon_qed_lsp_deq_data_parity                 ( smon_qed_lsp_deq_data_parity_nc )
        , .smon_qed_lsp_deq_data_cq                     ( smon_qed_lsp_deq_data_cq )
        , .smon_qed_lsp_deq_data_qe_wt                  ( smon_qed_lsp_deq_data_qe_wt_nc )

        , .smon_aqed_lsp_deq_v                          ( smon_aqed_lsp_deq_v )
        , .smon_aqed_lsp_deq_data_parity                ( smon_aqed_lsp_deq_data_parity_nc )
        , .smon_aqed_lsp_deq_data_cq                    ( smon_aqed_lsp_deq_data_cq )
        , .smon_aqed_lsp_deq_data_qe_wt                 ( smon_aqed_lsp_deq_data_qe_wt_nc )

        , .func_qed_lsp_deq_fifo_mem_re                 ( func_qed_lsp_deq_fifo_mem_re )
        , .func_qed_lsp_deq_fifo_mem_raddr              ( func_qed_lsp_deq_fifo_mem_raddr )
        , .func_qed_lsp_deq_fifo_mem_waddr              ( func_qed_lsp_deq_fifo_mem_waddr )
        , .func_qed_lsp_deq_fifo_mem_we                 ( func_qed_lsp_deq_fifo_mem_we )
        , .func_qed_lsp_deq_fifo_mem_wdata              ( func_qed_lsp_deq_fifo_mem_wdata )
        , .func_qed_lsp_deq_fifo_mem_rdata              ( func_qed_lsp_deq_fifo_mem_rdata ) 

        , .func_aqed_lsp_deq_fifo_mem_re                ( func_aqed_lsp_deq_fifo_mem_re )
        , .func_aqed_lsp_deq_fifo_mem_raddr             ( func_aqed_lsp_deq_fifo_mem_raddr )
        , .func_aqed_lsp_deq_fifo_mem_waddr             ( func_aqed_lsp_deq_fifo_mem_waddr )
        , .func_aqed_lsp_deq_fifo_mem_we                ( func_aqed_lsp_deq_fifo_mem_we )
        , .func_aqed_lsp_deq_fifo_mem_wdata             ( func_aqed_lsp_deq_fifo_mem_wdata )
        , .func_aqed_lsp_deq_fifo_mem_rdata             ( func_aqed_lsp_deq_fifo_mem_rdata ) 

        , .func_cq_ldb_wu_count_mem_re                  ( func_cq_ldb_wu_count_mem_re )
        , .func_cq_ldb_wu_count_mem_raddr               ( func_cq_ldb_wu_count_mem_raddr )
        , .func_cq_ldb_wu_count_mem_waddr               ( func_cq_ldb_wu_count_mem_waddr )
        , .func_cq_ldb_wu_count_mem_we                  ( func_cq_ldb_wu_count_mem_we )
        , .func_cq_ldb_wu_count_mem_wdata               ( func_cq_ldb_wu_count_mem_wdata )
        , .func_cq_ldb_wu_count_mem_rdata               ( func_cq_ldb_wu_count_mem_rdata )

        , .func_cfg_cq_ldb_wu_limit_mem_re              ( func_cfg_cq_ldb_wu_limit_mem_re )
        , .func_cfg_cq_ldb_wu_limit_mem_raddr           ( func_cfg_cq_ldb_wu_limit_mem_raddr )
        , .func_cfg_cq_ldb_wu_limit_mem_waddr           ( func_cfg_cq_ldb_wu_limit_mem_waddr )
        , .func_cfg_cq_ldb_wu_limit_mem_we              ( func_cfg_cq_ldb_wu_limit_mem_we )
        , .func_cfg_cq_ldb_wu_limit_mem_wdata           ( func_cfg_cq_ldb_wu_limit_mem_wdata )
        , .func_cfg_cq_ldb_wu_limit_mem_rdata           ( func_cfg_cq_ldb_wu_limit_mem_rdata )
) ;

//-------------------------------------------------------------------------------------------------
// Error reporting
//
// If there is a p5 calculation error (e.g. an if count overflow on a schedule request), don't block
// the request, don't want to hang or have timing issue or loop.  Just detect - will require at least
// a vas reset if not a pf_reset.

always_comb begin
  // Don't hold - 1-clock pulse to report
  p8_lba_qid_enq_cnt_uflow_err_nxt      = 1'b0 ;
  p8_lba_qid_enq_cnt_oflow_err_nxt      = 1'b0 ;
  p8_lba_qid_if_cnt_uflow_err_nxt       = 1'b0 ;
  p8_lba_qid_if_cnt_oflow_err_nxt       = 1'b0 ;
  p8_lba_cq_tok_cnt_oflow_err_nxt       = 1'b0 ;
  p8_lba_cq_tok_cnt_uflow_err_nxt       = 1'b0 ;
  p8_lba_cq_if_cnt_uflow_err_nxt        = 1'b0 ;
  p8_lba_cq_if_cnt_oflow_err_nxt        = 1'b0 ;
  p8_lba_tot_if_cnt_uflow_err_nxt       = 1'b0 ;
  p8_lba_tot_if_cnt_oflow_err_nxt       = 1'b0 ;

  p3_lba_inp_tok_cnt_res_err_nxt        = 1'b0 ;
  p8_lba_qid_enq_cnt_res_err_nxt        = 1'b0 ;
  p8_lba_qid_dpth_thrsh_par_err_nxt     = 1'b0 ;
  p8_lba_qid_if_cnt_res_err_nxt         = 1'b0 ;
  p8_lba_qid_if_lim_par_err_nxt         = 1'b0 ;
  p8_lba_cq_tok_cnt_res_err_nxt         = 1'b0 ;
  p8_lba_cq_tok_lim_par_err_nxt         = 1'b0 ;
  p8_lba_cq_if_cnt_res_err_nxt          = 1'b0 ;
  p8_lba_cq_if_lim_par_err_nxt          = 1'b0 ;
  p8_lba_inp_qid_par_err_nxt            = 1'b0 ;
  p8_lba_inp_cq_par_err_nxt             = 1'b0 ;
  p8_lba_tot_if_cnt_res_err_nxt         = 1'b0 ;

  p4_lba_cq2qid_priov_par_err_nxt       = 1'b0 ;
  p4_lba_cq2qid_qid0_par_err_nxt        = 1'b0 ;
  p4_lba_cq2qid_qid1_par_err_nxt        = 1'b0 ;

  if ( p2_lba_ctrl_pipe_v_f & ~ p3_lba_ctrl_pipe.hold ) begin
    p3_lba_inp_tok_cnt_res_err_nxt      = p2_lba_inp_tok_cnt_res_err_cond & ~ p2_lba_inp_tok_cq_disable ;
  end
  if ( p3_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold ) begin
    p4_lba_cq2qid_priov_par_err_nxt     = ( p3_lba_cq2qid_priov_par_err_cond | cfg_error_inject_f [ 5 ] ) & ~ p3_lba_cq2qid_cq_disable_x ;
    p4_lba_cq2qid_qid0_par_err_nxt      = p3_lba_cq2qid_qid0_par_err_cond & ~ p3_lba_cq2qid_cq_disable_x ;
    p4_lba_cq2qid_qid1_par_err_nxt      = p3_lba_cq2qid_qid1_par_err_cond & ~ p3_lba_cq2qid_cq_disable_x ;
  end
  if ( p7_lba_ctrl_pipe_v_f & ~ p8_lba_ctrl_pipe.hold ) begin
    p8_lba_qid_enq_cnt_uflow_err_nxt    = p7_lba_ctrl_pipe_f.sch_nalb_v & p7_lba_qid_enq_cnt_uflow_cond ;
    p8_lba_qid_enq_cnt_oflow_err_nxt    = p7_lba_ctrl_pipe_f.enq_v & ( p7_lba_qid_enq_cnt_oflow_cond ) ;
    p8_lba_qid_if_cnt_uflow_err_nxt     = ( p7_lba_ctrl_pipe_f.qid_cmp_v | p7_lba_ctrl_pipe_f.qid_if_dec_v ) & ( p7_lba_qid_if_cnt_uflow_cond ) ;
    p8_lba_qid_if_cnt_oflow_err_nxt     = p7_lba_ctrl_pipe_f.sch_nalb_v & p7_lba_qid_if_cnt_oflow_cond  ;
    p8_lba_cq_tok_cnt_uflow_err_nxt     = p7_lba_ctrl_pipe_f.tok_v & ( p7_lba_cq_tok_cnt_uflow_cond | cfg_error_inject_f [ 17 ] ) & ~ p7_lba_tok_cnt_cq_disable ;
    p8_lba_cq_tok_cnt_oflow_err_nxt     = ( p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.sch_atm_v ) & p7_lba_cq_tok_cnt_oflow_cond & ~ p7_lba_tok_cnt_cq_disable ;
    p8_lba_cq_if_cnt_uflow_err_nxt      = p7_lba_ctrl_pipe_f.cq_cmp_v & ( p7_lba_cq_if_cnt_uflow_cond | cfg_error_inject_f [ 1 ] ) & ~ p7_lba_if_cnt_cq_disable ;
    p8_lba_cq_if_cnt_oflow_err_nxt      = ( p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.sch_atm_v ) & p7_lba_cq_if_cnt_oflow_cond & ~ p7_lba_if_cnt_cq_disable ;
    p8_lba_tot_if_cnt_uflow_err_nxt     = p7_lba_ctrl_pipe_f.cq_cmp_v & p7_lba_tot_if_cnt_uflow_cond ;
    p8_lba_tot_if_cnt_oflow_err_nxt     = ( p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.sch_atm_v ) & p7_lba_tot_if_cnt_oflow_cond ;

    p8_lba_qid_enq_cnt_res_err_nxt      = p7_lba_qid_enq_cnt_res_err_cond ;
    p8_lba_qid_dpth_thrsh_par_err_nxt   = p7_lba_qid_dpth_thrsh_par_err_cond ;
    p8_lba_qid_if_cnt_res_err_nxt       = p7_lba_qid_if_cnt_res_err_cond ;
    p8_lba_qid_if_lim_par_err_nxt       = p7_lba_qid_if_lim_par_err_cond ;
    p8_lba_cq_tok_cnt_res_err_nxt       = p7_lba_cq_tok_cnt_res_err_cond & ~ p7_lba_tok_cnt_cq_disable ;
    p8_lba_cq_tok_lim_par_err_nxt       = p7_lba_cq_tok_lim_par_err_cond & ~ p7_lba_tok_cnt_cq_disable ;
    p8_lba_cq_if_cnt_res_err_nxt        = p7_lba_cq_if_cnt_res_err_cond & ~ p7_lba_if_cnt_cq_disable ;
    p8_lba_cq_if_lim_par_err_nxt        = ( p7_lba_cq_if_lim_par_err_cond | p7_lba_cq_if_thr_par_err_cond ) & ~ p7_lba_if_cnt_cq_disable ;
    p8_lba_inp_qid_par_err_nxt          = p7_lba_inp_qid_par_err_cond ;
    p8_lba_inp_cq_par_err_nxt           = p7_lba_inp_cq_par_err_cond ;
    p8_lba_tot_if_cnt_res_err_nxt       = p7_lba_tot_if_cnt_res_err_cond ;
  end

  p4_lbwu_inp_par_err_nxt               = 1'b0 ;
  p4_lbwu_cq_wu_cnt_res_err_nxt         = 1'b0 ;
  p4_lbwu_cq_wu_lim_par_err_nxt         = 1'b0 ;
  if ( p3_lbwu_cq_wu_cnt_upd_v_func ) begin     // Only do integrity checks on functional usage, not config reads
    p4_lbwu_inp_par_err_nxt             = p3_lbwu_inp_par_err_cond ;
    p4_lbwu_cq_wu_cnt_res_err_nxt       = p3_lbwu_cq_wu_cnt_res_err_cond ;
    p4_lbwu_cq_wu_lim_par_err_nxt       = p3_lbwu_cq_wu_lim_par_err_cond ;
  end

end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_lba_inp_tok_cnt_res_err_f        <= 1'b0 ;

    p8_lba_qid_enq_cnt_uflow_err_f      <= 1'b0 ;
    p8_lba_qid_enq_cnt_oflow_err_f      <= 1'b0 ;
    p8_lba_qid_if_cnt_uflow_err_f       <= 1'b0 ;
    p8_lba_qid_if_cnt_oflow_err_f       <= 1'b0 ;
    p8_lba_cq_tok_cnt_oflow_err_f       <= 1'b0 ;
    p8_lba_cq_tok_cnt_uflow_err_f       <= 1'b0 ;
    p8_lba_cq_if_cnt_uflow_err_f        <= 1'b0 ;
    p8_lba_cq_if_cnt_oflow_err_f        <= 1'b0 ;
    p8_lba_tot_if_cnt_uflow_err_f       <= 1'b0 ;
    p8_lba_tot_if_cnt_oflow_err_f       <= 1'b0 ;

    p8_lba_qid_enq_cnt_res_err_f        <= 1'b0 ;
    p8_lba_qid_dpth_thrsh_par_err_f     <= 1'b0 ;
    p8_lba_qid_if_cnt_res_err_f         <= 1'b0 ;
    p8_lba_qid_if_lim_par_err_f         <= 1'b0 ;
    p8_lba_cq_tok_cnt_res_err_f         <= 1'b0 ;
    p8_lba_cq_tok_lim_par_err_f         <= 1'b0 ;
    p8_lba_cq_if_cnt_res_err_f          <= 1'b0 ;
    p8_lba_cq_if_lim_par_err_f          <= 1'b0 ;
    p8_lba_inp_qid_par_err_f            <= 1'b0 ;
    p8_lba_inp_cq_par_err_f             <= 1'b0 ;
    p8_lba_tot_if_cnt_res_err_f         <= 1'b0 ;

    p9_lba_tot_enq_cnt_res_err_f        <= 1'b0 ;
    p9_lba_tot_sch_cnt_res_err_f        <= 1'b0 ;

    p4_lba_cq2qid_priov_par_err_f       <= 1'b0 ;
    p4_lba_cq2qid_qid0_par_err_f        <= 1'b0 ;
    p4_lba_cq2qid_qid1_par_err_f        <= 1'b0 ;

    p4_lbwu_inp_par_err_f               <= 1'b0 ;
    p4_lbwu_cq_wu_cnt_res_err_f         <= 1'b0 ;
    p4_lbwu_cq_wu_lim_par_err_f         <= 1'b0 ;
  end
  else begin
    p3_lba_inp_tok_cnt_res_err_f        <= p3_lba_inp_tok_cnt_res_err_nxt ;

    p8_lba_qid_enq_cnt_uflow_err_f      <= p8_lba_qid_enq_cnt_uflow_err_nxt ;
    p8_lba_qid_enq_cnt_oflow_err_f      <= p8_lba_qid_enq_cnt_oflow_err_nxt ;
    p8_lba_qid_if_cnt_uflow_err_f       <= p8_lba_qid_if_cnt_uflow_err_nxt ;
    p8_lba_qid_if_cnt_oflow_err_f       <= p8_lba_qid_if_cnt_oflow_err_nxt ;
    p8_lba_cq_tok_cnt_oflow_err_f       <= p8_lba_cq_tok_cnt_oflow_err_nxt ;
    p8_lba_cq_tok_cnt_uflow_err_f       <= p8_lba_cq_tok_cnt_uflow_err_nxt ;
    p8_lba_cq_if_cnt_uflow_err_f        <= p8_lba_cq_if_cnt_uflow_err_nxt ;
    p8_lba_cq_if_cnt_oflow_err_f        <= p8_lba_cq_if_cnt_oflow_err_nxt ;
    p8_lba_tot_if_cnt_uflow_err_f       <= p8_lba_tot_if_cnt_uflow_err_nxt ;
    p8_lba_tot_if_cnt_oflow_err_f       <= p8_lba_tot_if_cnt_oflow_err_nxt ;

    p8_lba_qid_enq_cnt_res_err_f        <= p8_lba_qid_enq_cnt_res_err_nxt ;
    p8_lba_qid_dpth_thrsh_par_err_f     <= p8_lba_qid_dpth_thrsh_par_err_nxt ;
    p8_lba_qid_if_cnt_res_err_f         <= p8_lba_qid_if_cnt_res_err_nxt ;
    p8_lba_qid_if_lim_par_err_f         <= p8_lba_qid_if_lim_par_err_nxt ;
    p8_lba_cq_tok_cnt_res_err_f         <= p8_lba_cq_tok_cnt_res_err_nxt ;
    p8_lba_cq_tok_lim_par_err_f         <= p8_lba_cq_tok_lim_par_err_nxt ;
    p8_lba_cq_if_cnt_res_err_f          <= p8_lba_cq_if_cnt_res_err_nxt ;
    p8_lba_cq_if_lim_par_err_f          <= p8_lba_cq_if_lim_par_err_nxt ;
    p8_lba_inp_qid_par_err_f            <= p8_lba_inp_qid_par_err_nxt ;
    p8_lba_inp_cq_par_err_f             <= p8_lba_inp_cq_par_err_nxt ;
    p8_lba_tot_if_cnt_res_err_f         <= p8_lba_tot_if_cnt_res_err_nxt ;

    p9_lba_tot_enq_cnt_res_err_f        <= p9_lba_tot_enq_cnt_res_err_nxt ;
    p9_lba_tot_sch_cnt_res_err_f        <= p9_lba_tot_sch_cnt_res_err_nxt ;

    p4_lba_cq2qid_priov_par_err_f       <= p4_lba_cq2qid_priov_par_err_nxt ;
    p4_lba_cq2qid_qid0_par_err_f        <= p4_lba_cq2qid_qid0_par_err_nxt ;
    p4_lba_cq2qid_qid1_par_err_f        <= p4_lba_cq2qid_qid1_par_err_nxt ;

    p4_lbwu_inp_par_err_f               <= p4_lbwu_inp_par_err_nxt ;
    p4_lbwu_cq_wu_cnt_res_err_f         <= p4_lbwu_cq_wu_cnt_res_err_nxt ;
    p4_lbwu_cq_wu_lim_par_err_f         <= p4_lbwu_cq_wu_lim_par_err_nxt ;
  end
end // always

assign p8_lba_cq_tok_cnt_uflow_err_rid  = { 1'b1 , 1'b0  , p8_lba_cq_tok_cnt_rmw_pipe_f_pnc.cq } ;      // is_ldb, spare, cq[5:0]
assign p8_lba_tot_if_cnt_uflow_err_rid  = { 1'b1 , 1'b0 , p8_lba_cq_if_cnt_rmw_pipe_f_pnc.cq } ;        // is_ldb, spare, cq[5:0]
assign p8_lba_cq_if_cnt_uflow_err_rid   = { 1'b1 , 1'b0 , p8_lba_cq_if_cnt_rmw_pipe_f_pnc.cq } ;        // is_ldb, spare, cq[5:0]
assign p8_lba_qid_if_cnt_uflow_err_rid  = { 1'b1 , p8_lba_qid_if_cnt_rmw_pipe_f_pnc.qid } ;             // is_ldb, qid[6:0]

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB ATM scheduling
//-----------------------------------------------------------------------------------------------------
// Add in cq p and qid p
assign p4_lba_ctrl_pipe_cmp_p                   = ^ ( { p4_lba_ctrl_pipe_f.cmp_p ,
                                                        p4_lba_ctrl_pipe_f.cmp_cq_p ,
                                                        p4_lba_ctrl_pipe_f.cmp_qid_atm_p } ) ;

hqm_AW_parity_gen #( .WIDTH( 1 + HQM_LSP_ARCH_NUM_LB_QIDB2 + 3 ) ) i_lba_lsp_ap_atm_sched_par_gen (
          .d            ( { p4_lba_ctrl_pipe_f.sch_cq_p ,
                            p4_lba_sch_arb_winner_qid ,                         // Add in qid
                            p4_lba_sch_arb_winner_qidix } )                     // Add in qidix
        , .odd          ( 1'b0 )                                                // Subtracting bits to existing parity so just want XOR
        , .p            ( p4_lsp_ap_atm_sched_p )
) ;

assign lsp_ap_atm_v             = p4_lba_ctrl_pipe_v_f & ~ p5_lba_ctrl_pipe.hold &
                                  ( p4_lba_sch_arb_atm | ( p4_lba_ctrl_pipe_f.cq_cmp_v & p4_lba_ctrl_pipe_f.cmp_atm ) ) ;

always_comb begin
  p4_lba_sch_atm_pri_scaled_pnc                                 = '0 ;
  p4_lba_sch_atm_pri_scaled_pnc [HQM_LSP_NUM_PRI_BINSB2-1:0]    = p4_lba_sch_atm_pri_f ;

  lsp_ap_atm_data.pcm = p4_lba_ctrl_pipe_f_pcm ; 
  if ( p4_lba_sch_arb_atm ) begin
    if ( p4_lba_sch_atm_rlist_f )
      lsp_ap_atm_data.cmd                       = LSP_AP_ATM_SCH_RLST ;
    else
      lsp_ap_atm_data.cmd                       = LSP_AP_ATM_SCH_SLST ;
    lsp_ap_atm_data.cq                          = p4_lba_ctrl_pipe_f_pcm ? { 2'h0 , p4_lba_ctrl_pipe_f.sch_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , p4_lba_sch_arb_winner_qidix_msb } : { 2'h0 , p4_lba_ctrl_pipe_f.sch_cq } ;
    lsp_ap_atm_data.qid                         = p4_lba_sch_arb_winner_qid ;
    lsp_ap_atm_data.qidix_msb                   = p4_lba_sch_arb_winner_qidix_msb ;
    lsp_ap_atm_data.qidix                       = p4_lba_sch_arb_winner_qidix ;
    lsp_ap_atm_data.qpri                        = ( p4_lba_sch_atm_pri_scaled_pnc << HQM_LSP_PRI_BIN_FACTOR ) ;
    lsp_ap_atm_data.parity                      = p4_lba_ctrl_pipe_f_pcm ? p4_lsp_ap_atm_sched_p ^ p4_lba_sch_arb_winner_qidix_msb ^ p4_lba_ctrl_pipe_f.sch_cq [ 0 ] : p4_lsp_ap_atm_sched_p ;
    lsp_ap_atm_data.fid                         = 12'h0 ;               // Unused
    lsp_ap_atm_data.fid_parity                  = 1'b1 ;                // Unused
    lsp_ap_atm_data.hid                         = 16'h0 ;               // Unused
    lsp_ap_atm_data.hid_parity                  = 1'b1 ;                // Unused
    lsp_ap_atm_data.hqm_core_flags.pad_ok                       = '0 ;
    lsp_ap_atm_data.hqm_core_flags.ignore_cq_depth              = p4_lba_sch_arb_winner_qidix_msb ;        // repurpose to carry qidix_msb 
    lsp_ap_atm_data.hqm_core_flags.cq_is_ldb                    = 1'b1 ;
    lsp_ap_atm_data.hqm_core_flags.write_buffer_optimization    = 2'h0 ;        // Not used for ldb
    lsp_ap_atm_data.hqm_core_flags.congestion_management        = p4_lba_sch_arb_winner_cm_code ;
    lsp_ap_atm_data.hqm_core_flags.parity                       = ~ ( ^ ( {             // Potential timing issue
                                                                            1'b1
                                                                          , p4_lba_sch_arb_winner_qidix_msb
                                                                          , p4_lba_sch_arb_winner_cm_code } ) ) ;
  end

  else begin
    lsp_ap_atm_data.cmd                         = LSP_AP_ATM_CMP ;
    lsp_ap_atm_data.cq                          = p4_lba_ctrl_pipe_f_pcm ? { 2'h0 , p4_lba_ctrl_pipe_f.cmp_cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , p4_lba_ctrl_pipe_f.cmp_qidix_msb } : { 2'h0 , p4_lba_ctrl_pipe_f.cmp_cq } ;
    lsp_ap_atm_data.qid                         = p4_lba_ctrl_pipe_f.cmp_qid_atm ;
    lsp_ap_atm_data.qidix_msb                   = p4_lba_ctrl_pipe_f.cmp_qidix_msb ;
    lsp_ap_atm_data.qidix                       = p4_lba_ctrl_pipe_f.cmp_qidix ;
    lsp_ap_atm_data.qpri                        = p4_lba_ctrl_pipe_f.cmp_qpri ;
    lsp_ap_atm_data.parity                      = p4_lba_ctrl_pipe_f_pcm ? p4_lba_ctrl_pipe_cmp_p ^ p4_lba_ctrl_pipe_f.cmp_qidix_msb ^ p4_lba_ctrl_pipe_f.cmp_cq [ 0 ] : p4_lba_ctrl_pipe_cmp_p ;              // Includes all of the above fields except cmd
    lsp_ap_atm_data.fid                         = p4_lba_ctrl_pipe_f.cmp_fid ;
    lsp_ap_atm_data.fid_parity                  = p4_lba_ctrl_pipe_f.cmp_fid_p ;
    lsp_ap_atm_data.hid                         = p4_lba_ctrl_pipe_f.cmp_hid ;
    lsp_ap_atm_data.hid_parity                  = p4_lba_ctrl_pipe_f.cmp_hid_p ;
    lsp_ap_atm_data.hqm_core_flags              = '0 ;                                  // Unused
    lsp_ap_atm_data.hqm_core_flags.parity       = 1'b1 ;
  end
end // always

assign p4_lba_atm_sch_hold      = lsp_ap_atm_v & ~ lsp_ap_atm_ready ;

//-------------------------------------------------------------------------------------------------
// Manage storage for per-qid cqidix map for blasting.  Since only needed for blasting only read
// when scheduling (both nalb and atm).
// p0/1/2/3 for the rw_pipe is pipe levels p5/p6/p7/p8
// Split into 16 memories to simplify config access.
// Only written by config.

always_comb begin
  if ( p4_lba_sch_arb_winner_v ) begin
    p5_lba_blast_qid2cqidix_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_READ ;                          // Don't do lookup unless necessary
  end
  else begin
    p5_lba_blast_qid2cqidix_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_NOOP ;
  end
  p5_lba_blast_qid2cqidix_rw_pipe_nxt.qid         = p4_lba_sch_arb_winner_qid ;
  p5_lba_blast_qid2cqidix_rw_pipe_nxt.data        = { $bits ( lsp_cfg_qid2cqidix_t ) { 1'b0 } } ; // Unused - cfg write done elsewhere
end // always

// Same as i_lba_qid2cqidix_pipe, replicated because of PD concerns about size/distance of blast logic and "spraying" logic
hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LB_QID2CQIDIX_MEM_WIDTH )
) i_lba_blast_qid2cqidix_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lba_blast_qid2cqidix_rmw_pipe_status_nc )                     // Unused - same as lba_cq_tok_cnt_rmw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p5_lba_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p5_lba_blast_qid2cqidix_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p5_lba_blast_qid2cqidix_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p5_lba_blast_qid2cqidix_rw_pipe_nxt.data )
        , .p0_hold              ( p5_lba_ctrl_pipe.hold )
        , .p0_v_f               ( p5_lba_blast_qid2cqidix_rw_pipe_v_f_nc )              // Unused - duplicate
        , .p0_rw_f              ( p5_lba_blast_qid2cqidix_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p5_lba_blast_qid2cqidix_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p5_lba_blast_qid2cqidix_rw_pipe_data_f_nc )

        , .p1_hold              ( p6_lba_ctrl_pipe.hold )
        , .p1_v_f               ( p6_lba_blast_qid2cqidix_rw_pipe_v_f_nc )              // Unused - duplicate
        , .p1_rw_f              ( p6_lba_blast_qid2cqidix_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p6_lba_blast_qid2cqidix_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p6_lba_blast_qid2cqidix_rw_pipe_data_f_nc )

        , .p2_hold              ( p7_lba_ctrl_pipe.hold )
        , .p2_v_f               ( p7_lba_blast_qid2cqidix_rw_pipe_v_f_nc )              // Unused - duplicate
        , .p2_rw_f              ( p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.rw_cmd )        // Used to distinguish parity check
        , .p2_addr_f            ( p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.qid )           // Unused
        , .p2_data_f            ( p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.data )

        , .p3_hold              ( p8_lba_ctrl_pipe.hold )
        , .p3_v_f               ( p8_lba_blast_qid2cqidix_rw_pipe_v_f_nc )              // Unused
        , .p3_rw_f              ( p8_lba_blast_qid2cqidix_rw_pipe_f_nc.rw_cmd )         // Unused
        , .p3_addr_f            ( p8_lba_blast_qid2cqidix_rw_pipe_f_nc.qid )            // Unused
        , .p3_data_f            ( p8_lba_blast_qid2cqidix_rw_pipe_f_nc.data )           // Unused


        // mem intf
        , .mem_write            ( func_cfg_qid_ldb_qid2cqidix2_mem_we )                 // Never used - cfg writes done elsewhere
        , .mem_read             ( func_cfg_qid_ldb_qid2cqidix2_mem_re )
        , .mem_addr             ( func_cfg_qid_ldb_qid2cqidix2_mem_addr )
        , .mem_write_data       ( func_cfg_qid_ldb_qid2cqidix2_mem_wdata )              // Never used - cfg writes done elsewhere
        , .mem_read_data        ( func_cfg_qid_ldb_qid2cqidix2_mem_rdata )
) ;

// "Spray" the scheduling status winning sch_atm qid to all cq/qidix pairs which also map to that qid.
assign p7_lba_blast_qid2cqidix_v        = p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.data.qidixv ;

assign p7_lba_blast_qid2cqidix_p        = p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.data.parity ;         // 16 bits

assign p7_lba_blast_nalb                = p7_lba_ctrl_pipe_v_1_f & ~ p8_lba_ctrl_pipe.hold & p7_lba_ctrl_pipe_f.sch_nalb_v ;
assign p7_lba_blast_slist               = p7_lba_ctrl_pipe_v_1_f & ~ p8_lba_ctrl_pipe.hold & p7_lba_ctrl_pipe_f.sch_atm_v & ~ p7_lba_ctrl_pipe_f.sch_atm_rlist ;
assign p7_lba_blast_rlist               = p7_lba_ctrl_pipe_v_1_f & ~ p8_lba_ctrl_pipe.hold & p7_lba_ctrl_pipe_f.sch_atm_v &   p7_lba_ctrl_pipe_f.sch_atm_rlist ;

// Include sw error case where ldb_sched_control was used to turn on a "haswork" but but the qid did not have work.  Avoids lba_sch_state machine hang
assign p7_lba_sched                     = p7_lba_ctrl_pipe_v_1_f & ~ p8_lba_ctrl_pipe.hold & p7_lba_ctrl_pipe_f.sch_v ;

assign p7_lba_set_cmpblast              = p7_lba_blast_slist & p8_lba_ctrl_pipe_nxt.sch_cmpblast_qidixv [ { p7_lba_ctrl_pipe_f.sch_qidix_msb , p7_lba_ctrl_pipe_f.sch_qidix } ] ;

assign p7_lba_blast_qid2cqidix_par_chk_en       = p7_lba_ctrl_pipe_v_f & ( p7_lba_blast_qid2cqidix_rw_pipe_f_pnc.rw_cmd == HQM_AW_RWPIPE_READ ) ;

generate
  for ( genvar gi = 0 ; gi < 16 ; gi = gi + 1 ) begin: gen_qid2cqidix2_par_chk
    hqm_AW_parity_check # ( .WIDTH ( 32 ) ) i_lba_qid2cqidix2_par_chk (
          .p                    ( p7_lba_blast_qid2cqidix_p [gi] )
        , .d                    ( p7_lba_blast_qid2cqidix_v [ ( gi * 32 ) +: 32 ] )
        , .e                    ( p7_lba_blast_qid2cqidix_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p7_lba_blast_qid2cqidix_par_err_cond [gi] )
    ) ;
  end
endgenerate

always_comb begin
  p8_lba_blast_qid2cqidix_v_nxt         = p8_lba_blast_qid2cqidix_v_f ;

  // Don't hold - 1-clock pulse to report
  p8_lba_blast_qid2cqidix_par_err_nxt   = 16'h0 ;

  if ( p8_lba_ctrl_pipe.en & p7_lba_ctrl_pipe_f.sch_nalb_v ) begin
    p8_lba_blast_qid2cqidix_v_nxt       = p7_lba_blast_qid2cqidix_v ;
    p8_lba_blast_qid2cqidix_par_err_nxt = p7_lba_blast_qid2cqidix_par_err_cond ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p8_lba_blast_qid2cqidix_v_f         <= 512'h0 ;
    p8_lba_blast_qid2cqidix_par_err_f   <= 16'h0 ;
  end
  else begin
    p8_lba_blast_qid2cqidix_v_f         <= p8_lba_blast_qid2cqidix_v_nxt ;
    p8_lba_blast_qid2cqidix_par_err_f   <= p8_lba_blast_qid2cqidix_par_err_nxt ;
  end
end // always

assign p8_lba_blast_qid2cqidix_par_err_any        = | p8_lba_blast_qid2cqidix_par_err_f ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB Update status vectors for next iteration
//-----------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// Per-CQ status - used for both nalb and atomic

assign p7_lba_cq_if_v_upd               = p7_lba_ctrl_pipe_f.sch_v | p7_lba_ctrl_pipe_f.cq_cmp_v ;
assign p7_lba_cq_tok_v_upd              = p7_lba_ctrl_pipe_f.sch_v | p7_lba_ctrl_pipe_f.tok_v ;

always_comb begin
  p8_lba_cq_tok_v_nxt           = p8_lba_cq_tok_v_f ;
  p8_lba_cq_if_v_nxt            = p8_lba_cq_if_v_f ;
  p8_lba_cq_thr_v_nxt           = p8_lba_cq_thr_v_f ;
  p8_lba_tot_if_v_nxt           = p8_lba_tot_if_v_f ;
  p8_lba_cq_tok_v_upd_nxt       = 1'b0 ;                                // No need to hold - unconditionally takes effect next clock
  p8_lba_cq_if_v_upd_nxt        = 1'b0 ;                                // No need to hold - unconditionally takes effect next clock
  p8_lba_cq_tok_cnt_v_nxt       = p8_lba_cq_tok_cnt_v_f ;
  p8_lba_cq_if_cnt_v_nxt        = p8_lba_cq_if_cnt_v_f ;

  // p8_lba_cq_if_v, p8_lba_cq_if_cnt_v and p8_lba_tot_if_v should be properly updated on a successful vas reset drain
  for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
    if ( p8_lba_ctrl_pipe.en ) begin
      if ( ( p7_lba_cq_tok_cnt_rmw_pipe_f.cq == i ) & p7_lba_cq_tok_v_upd ) begin
        p8_lba_cq_tok_v_nxt [i]         = p7_lba_cq_tok_cnt_upd_lt_lim_next ;
        p8_lba_cq_tok_cnt_v_nxt [i]     = p7_lba_cq_tok_cnt_upd_gt_0 ;
      end
      //--------
      if ( ( p7_lba_cq_if_cnt_rmw_pipe_f.cq == i ) & p7_lba_cq_if_v_upd ) begin
        p8_lba_cq_if_v_nxt [i]          = p7_lba_cq_if_cnt_upd_lt_lim ;
        p8_lba_cq_if_cnt_v_nxt [i]      = p7_lba_cq_if_cnt_upd_gt_0 ;

        // Note: Not possible to have a simultaneous set and clear, since one is on a sch and the other is on a cmp
        if ( p7_lba_ctrl_pipe_f.cq_cmp_v & p7_lba_cq_if_cnt_upd_le_thr ) begin
          p8_lba_cq_thr_v_nxt [i]       = 1'b1 ;
        end
        else if ( p7_lba_ctrl_pipe_f.sch_v & ( ~ p7_lba_cq_if_cnt_upd_lt_lim ) & cfg_control_enable_inflight_thresh ) begin
          p8_lba_cq_thr_v_nxt [i]       = 1'b0 ;
        end
      end
    end

    if ( cfgsc_cq_ldb_token_count_mem_we & ( cfg_mem_addr [HQM_NUM_LB_CQB2-1:0] == i ) ) begin          // Should only be done as part of vas reset or cq configuration
        p8_lba_cq_tok_v_nxt [i]         = 1'b1 ;
        p8_lba_cq_tok_cnt_v_nxt [i]     = 1'b0 ;
    end // if cfg wr
  end // for i

  if ( p8_lba_ctrl_pipe.en ) begin
    p8_lba_cq_tok_v_upd_nxt     = p7_lba_cq_tok_v_upd ;
    p8_lba_cq_if_v_upd_nxt      = p7_lba_cq_if_v_upd ;
  end // if en

  if ( p8_lba_ctrl_pipe.en & p7_lba_cq_if_v_upd ) begin
    p8_lba_tot_if_v_nxt         = p7_lba_tot_if_cnt_upd_lt_lim ;
  end
end // always_comb

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p8_lba_cq_tok_v_f           <= { HQM_NUM_LB_CQ { 1'b1 } } ;
    p8_lba_cq_if_v_f            <= { HQM_NUM_LB_CQ { 1'b1 } } ;
    p8_lba_cq_thr_v_f           <= { HQM_NUM_LB_CQ { 1'b1 } } ;
    p8_lba_tot_if_v_f           <= 1'b1 ;
    p8_lba_cq_tok_v_upd_f       <= 1'b0 ;
    p8_lba_cq_if_v_upd_f        <= 1'b0 ;
    p8_lba_cq_tok_cnt_v_f       <= { HQM_NUM_LB_CQ { 1'b0 } } ;
    p8_lba_cq_if_cnt_v_f        <= { HQM_NUM_LB_CQ { 1'b0 } } ;
  end
  else begin
    p8_lba_cq_tok_v_f           <= p8_lba_cq_tok_v_nxt ;
    p8_lba_cq_if_v_f            <= p8_lba_cq_if_v_nxt ;
    p8_lba_cq_thr_v_f           <= p8_lba_cq_thr_v_nxt ;
    p8_lba_tot_if_v_f           <= p8_lba_tot_if_v_nxt ;
    p8_lba_cq_tok_v_upd_f       <= p8_lba_cq_tok_v_upd_nxt ;
    p8_lba_cq_if_v_upd_f        <= p8_lba_cq_if_v_upd_nxt ;
    p8_lba_cq_tok_cnt_v_f       <= p8_lba_cq_tok_cnt_v_nxt ;
    p8_lba_cq_if_cnt_v_f        <= p8_lba_cq_if_cnt_v_nxt ;
  end
end // always

assign p8_lba_cq_has_space      = p8_lba_cq_tok_v_f &
                                  p8_lba_cq_thr_v_f & p8_lba_cq_if_v_f & { HQM_NUM_LB_CQ { p8_lba_tot_if_v_f } } ;      // Bitwise

assign cfg_cq_ldb_if_v_status   = p8_lba_cq_if_v_f ;
assign cfg_cq_ldb_thr_v_status  = p8_lba_cq_thr_v_f ;
assign cfg_cq_ldb_tok_v_status  = p8_lba_cq_tok_v_f ;

//-------------------------------------------------------------------------------------------------
// Per-qidix status - used only by nalb.  Atomic uses slist_v/rlist_v provided by AP for "has work",
// but does also track per-QID inflight.

// "Spray" the updated sch/if status for the winning qid to all cq/qidix pairs which also map to that qid.

// For completion (or RELEASE) need to update for all CQs (for that QID) even though completed for a particular CQ.
assign p7_lba_qidix_if_v_upd            = p7_lba_ctrl_pipe_f.sch_v      | p7_lba_ctrl_pipe_f.qid_cmp_v | p7_lba_ctrl_pipe_f.qid_if_dec_v ;      // Both LB and ATM sch
assign p7_lba_qidix_sch_v_upd           = p7_lba_ctrl_pipe_f.sch_nalb_v | p7_lba_ctrl_pipe_f.enq_v ;

always_comb begin
  // Should be correctly adjusted as part of a successful vas reset drain
  p8_lba_qidix_sch_v_nxt                = p8_lba_qidix_sch_v_f ;
  p8_lba_qidix_if_v_nxt                 = p8_lba_qidix_if_v_f ;
  p8_lba_qidix_sch_v_upd_nxt            = 1'b0 ;                        // No need to hold - unconditionally takes effect next clock
  p8_lba_qidix_if_v_upd_nxt             = 1'b0 ;                        // No need to hold - unconditionally takes effect next clock

  if ( p8_lba_ctrl_pipe.en ) begin
    p8_lba_qidix_sch_v_upd_nxt          = p7_lba_qidix_sch_v_upd ;
    p8_lba_qidix_if_v_upd_nxt           = p7_lba_qidix_if_v_upd ;
  end // if en
  if ( cfg_ldb_sched_control_inflight_ok_v ) begin
    p8_lba_qidix_if_v_upd_nxt          = 1'b1 ;
  end
  if ( cfg_ldb_sched_control_nalb_haswork_v ) begin
    p8_lba_qidix_sch_v_upd_nxt          = 1'b1 ;
  end

  for ( int i = 0 ; i < HQM_LSP_NUM_LB_CQQIDIX ; i = i + 1 ) begin
    if ( p8_lba_ctrl_pipe.en ) begin
      if ( p7_lba_qid2cqidix_v [i] & p7_lba_qidix_sch_v_upd ) begin
        p8_lba_qidix_sch_v_nxt [i]      = p7_lba_qid_enq_cnt_upd_gt0 ;
      end
      //--------
      if ( p7_lba_qid2cqidix_v [i] & p7_lba_qidix_if_v_upd ) begin
        p8_lba_qidix_if_v_nxt [i]       = p7_lba_qid_if_cnt_upd_lt_lim ;
      end
    end // if en
    if ( cfg_ldb_sched_control_inflight_ok_v & ( cfg_ldb_sched_control_cq_qidix == i ) ) begin
      p8_lba_qidix_if_v_nxt [i]         = cfg_ldb_sched_control_value ;
    end
    if ( cfg_ldb_sched_control_nalb_haswork_v & ( cfg_ldb_sched_control_cq_qidix == i ) ) begin
      p8_lba_qidix_sch_v_nxt [i]        = cfg_ldb_sched_control_value ;
    end
  end // for i
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p8_lba_qidix_if_v_f         <= { 512 { 1'b1 } } ;
    p8_lba_qidix_sch_v_f        <= { 512 { 1'b0 } } ;
    p8_lba_qidix_if_v_upd_f     <= 1'b0 ;
    p8_lba_qidix_sch_v_upd_f    <= 1'b0 ;
  end
  else begin
    p8_lba_qidix_if_v_f         <= p8_lba_qidix_if_v_nxt ;
    p8_lba_qidix_sch_v_f        <= p8_lba_qidix_sch_v_nxt ;
    p8_lba_qidix_if_v_upd_f     <= p8_lba_qidix_if_v_upd_nxt ;
    p8_lba_qidix_sch_v_upd_f    <= p8_lba_qidix_sch_v_upd_nxt ;
  end
end // always

assign p8_lba_qidix_has_work            = p8_lba_qidix_if_v_f & p8_lba_qidix_sch_v_f ;

assign cfg_qid_ldb_if_v_status          = p8_lba_qidix_if_v_f ;
assign cfg_qid_ldb_sch_v_status         = p8_lba_qidix_sch_v_f ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBARB Schedule output
//-----------------------------------------------------------------------------------------------------
// Need to include qid and slot/qidix parity in output, don't do in previous stage due to delay reasons
hqm_AW_parity_gen #( .WIDTH( HQM_LSP_ARCH_NUM_LB_QIDB2 + 3 + 1) ) i_lba_sch_par_gen (
          .d            ( { p8_lba_sch_pipe_f.parity ,                          // Just the cq parity in p8
                            p8_lba_sch_pipe_f.qid ,
                            p8_lba_sch_pipe_f.slot } )
        , .odd          ( 1'b0 )                // Adding bits to existing parity so just want XOR
        , .p            ( p8_lba_sch_pipe_gp )
) ;

assign p9_lba_nalb_sch_err_nxt                  = nalb_sel_nalb_fifo_credit_err_cond & ~ nalb_sel_nalb_fifo_cerr_reported_f ;

// sticky, only clearable by pf reset
assign nalb_sel_nalb_fifo_cerr_reported_nxt     = nalb_sel_nalb_fifo_cerr_reported_f | nalb_sel_nalb_fifo_credit_err_cond ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    nalb_sel_nalb_fifo_cerr_reported_f  <= 1'b0 ;
    p9_lba_nalb_sch_err_f               <= 1'b0 ;
  end
  else begin
    nalb_sel_nalb_fifo_cerr_reported_f  <= nalb_sel_nalb_fifo_cerr_reported_nxt ;
    p9_lba_nalb_sch_err_f               <= p9_lba_nalb_sch_err_nxt ;
  end
end // always

// Note: Pipe is not held; this condition should never occur if the FIFO wm and credit limit are properly configured.
// See comments in pipeline hold/en section.
assign nalb_sel_nalb_fifo_credit_err_cond       = p8_lba_ctrl_pipe_v_f & p8_lba_ctrl_pipe_f.sch_nalb_v & nalb_sel_nalb_fifo_afull ;

assign nalb_sel_nalb_fifo_push  = p8_lba_ctrl_pipe_v_f & p8_lba_ctrl_pipe_f.sch_nalb_v & ~ nalb_sel_nalb_fifo_afull ; // ~afull should be redundant if config OK

assign nalb_sel_nalb_fifo_push_data.cq          = p8_lba_ctrl_pipe_f_pcm ? { 2'h0 , p8_lba_sch_pipe_f.cq [ HQM_LSP_ARCH_NUM_LB_CQB2-1 : 1 ] , 1'b0  } : { 2'h0 , p8_lba_sch_pipe_f.cq } ;
assign nalb_sel_nalb_fifo_push_data.qid         = p8_lba_sch_pipe_f.qid ;
assign nalb_sel_nalb_fifo_push_data.qidix       = p8_lba_sch_pipe_f.slot ;
assign nalb_sel_nalb_fifo_push_data.parity      = p8_lba_sch_pipe_gp ^ cfg_error_inject_f [ 11 ] ^ ( p8_lba_ctrl_pipe_f_pcm & p8_lba_ctrl_pipe_f.sch_cq [ 0 ] ) ;
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.pad_ok                       = '0 ;
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.ignore_cq_depth              = p8_lba_ctrl_pipe_f.sch_qidix_msb ;        // repurpose to carry qidix_msb 
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.cq_is_ldb                    = 1'b1 ;
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.write_buffer_optimization    = 2'h0 ;        // Not used for ldb
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.congestion_management        = p8_lba_sch_pipe_f.cm_code ;
assign nalb_sel_nalb_fifo_push_data.hqm_core_flags.parity       = ~ ( ^ ( {             // Potential timing issue
                                                                              1'b1
                                                                            , p8_lba_ctrl_pipe_f.sch_qidix_msb
                                                                            , p8_lba_sch_pipe_f.cm_code
                                                                            , cfg_error_inject_f [ 12 ] } ) ) ;

//-------------------------------------------------------------------------------------------------

assign nalb_sel_nalb_fifo_hwm           = HQM_LSP_NALB_SEL_NALB_FIFO_DEPTH [HQM_LSP_NALB_SEL_NALB_FIFO_WMWIDTH-1:0] ;

hqm_AW_fifo_control #(
          .DEPTH                ( HQM_LSP_NALB_SEL_NALB_FIFO_DEPTH )
        , .DWIDTH               ( HQM_LSP_NALB_SEL_NALB_FIFO_DWIDTH )
) i_nalb_sel_nalb_if_fifo (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )

        , .push                 ( nalb_sel_nalb_fifo_push )
        , .push_data            ( nalb_sel_nalb_fifo_push_data )
        , .pop                  ( nalb_sel_nalb_fifo_pop )
        , .pop_data             ( nalb_sel_nalb_fifo_pop_data )

        , .cfg_high_wm          ( nalb_sel_nalb_fifo_hwm )

        , .mem_we               ( func_nalb_sel_nalb_fifo_mem_we )
        , .mem_waddr            ( func_nalb_sel_nalb_fifo_mem_waddr )
        , .mem_wdata            ( func_nalb_sel_nalb_fifo_mem_wdata )
        , .mem_re               ( func_nalb_sel_nalb_fifo_mem_re )
        , .mem_raddr            ( func_nalb_sel_nalb_fifo_mem_raddr )
        , .mem_rdata            ( func_nalb_sel_nalb_fifo_mem_rdata )

        , .fifo_status          ( nalb_sel_nalb_fifo_status_pnc )
        , .fifo_full            ( nalb_sel_nalb_fifo_full_nc )
        , .fifo_afull           ( nalb_sel_nalb_fifo_afull )
        , .fifo_empty           ( nalb_sel_nalb_fifo_empty )
) ;


assign nalb_sel_nalb_fifo_of                            = nalb_sel_nalb_fifo_status_pnc [1] ;
assign nalb_sel_nalb_fifo_uf                            = nalb_sel_nalb_fifo_status_pnc [0] ;

assign nalb_sel_nalb_fifo_pop_data_v       = ~ nalb_sel_nalb_fifo_empty ;
assign nalb_sel_nalb_fifo_pop              = nalb_sel_nalb_fifo_pop_data_v & lsp_nalb_sch_unoord_in_ready ;

// nalb_sel_nalb_fifo_pop_data goes to i_hqm_AW_tx_sync_lsp_nalb_sch_unoord

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: ATQ pipe - Detects initial atomic (ATQ) enqueue notifications and schedules to the NALB, and
// notifications from AQED that an ATQ has been sent out (pseudo-completion, actual completion occurs
// later but LSP doesn't need to wait that long since it is only protecting the AQED storage).
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: ATQ input pipe arbitration
//-----------------------------------------------------------------------------------------------------
// There are 3 functional inputs to the atq enqueue and aqed-active pipes: enqueue requests (E),
// aqed pseudo-completions (C) and schedule requests (S).  S ties up both pipes; C and E each tie up
// only their respective pipes.  In order to maximize efficiency, the logic only allows E and C requests
// to go if they are both present or if there are no S requests.  The algorithm is:
// S * E * C            : use arbiter; if S loses, allow both E and C to go (either way ties up both)
// S * ( ~E + ~C )      : Allow S to go (ties up both)
// ~S                   : Allow E or C (or both) to go if they are valid
assign atq_input_arb_new_both           = enq_atq_fifo_pop_data_vreq & send_atm_to_cq_fifo_pop_data_vreq ;
assign atq_input_arb_new_either         = enq_atq_fifo_pop_data_vreq | send_atm_to_cq_fifo_pop_data_vreq ;

assign atq_input_arb_reqs [0]           = atq_input_arb_new_either & ( atq_input_arb_new_both | ~ p4_atq_sch_v_f ) ;

assign atq_input_arb_reqs [1]           = p4_atq_sch_v_f ;

assign atq_input_arb_update             = p0_atq_ctrl_pipe.en ;

hqm_AW_rr_arb # ( .NUM_REQS ( 2 ) ) i_atq_input_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( atq_input_arb_reqs )
        , .update               ( atq_input_arb_update )
        , .winner_v             ( atq_input_arb_winner_pre_v )
        , .winner               ( atq_input_arb_winner )
) ;

assign atq_input_arb_winner_v   = atq_input_arb_winner_pre_v &
                                  ~ ( ( cfg_control_single_op_atq & ( ( ~ atq_upipe_idle_f ) | p0_atq_ctrl_pipe_v_f ) ) |
                                      ( cfg_control_half_bw_atq & p0_atq_ctrl_pipe_v_f ) ) ;

assign atq_input_arb_pre_enq    = atq_input_arb_winner_v & ~ atq_input_arb_winner & ~ p0_atq_ctrl_pipe.hold & enq_atq_fifo_pop_data_vreq ;
assign atq_input_arb_pre_cmp    = atq_input_arb_winner_v & ~ atq_input_arb_winner & ~ p0_atq_ctrl_pipe.hold & send_atm_to_cq_fifo_pop_data_vreq ;
assign atq_input_arb_sch        = atq_input_arb_winner_v &   atq_input_arb_winner & ~ p0_atq_ctrl_pipe.hold ;
assign atq_input_arb_sch_qid    = p4_atq_sch_qid_f ;

// Disable if arbiter has allowed multiple ops and disabled by config and toggle does not allow
assign atq_input_arb_enq        = atq_input_arb_pre_enq & ~ ( cfg_control_disable_multi_op_atq & atq_input_arb_pre_cmp & atq_input_arb_tog_f ) ;
assign atq_input_arb_cmp        = atq_input_arb_pre_cmp & ~ ( cfg_control_disable_multi_op_atq & atq_input_arb_pre_enq & ~ atq_input_arb_tog_f ) ;

always_comb begin
  atq_input_arb_tog_nxt         = atq_input_arb_tog_f ;
  if ( cfg_control_disable_multi_op_atq & atq_input_arb_pre_enq & atq_input_arb_pre_cmp )
    atq_input_arb_tog_nxt       = ~ atq_input_arb_tog_f ;
end // always

assign aqed_lsp_dec_fid_cnt_v_last_nxt  = aqed_lsp_dec_fid_cnt_v_f ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    atq_input_arb_tog_f                 <= 1'b0 ;
    aqed_lsp_dec_fid_cnt_v_f            <= 1'b0 ;
    aqed_lsp_dec_fid_cnt_v_last_f       <= 1'b0 ;
  end
  else begin
    atq_input_arb_tog_f                 <= atq_input_arb_tog_nxt ;
    aqed_lsp_dec_fid_cnt_v_f            <= aqed_lsp_dec_fid_cnt_v ;
    aqed_lsp_dec_fid_cnt_v_last_f       <= aqed_lsp_dec_fid_cnt_v_last_nxt ;
  end
end // always
assign aqed_lsp_dec_fid_cnt_v_idle      = ~ aqed_lsp_dec_fid_cnt_v_f & ~ aqed_lsp_dec_fid_cnt_v_last_f ;        // Need second stage to cover cfg_fid_inflight_count_f,
                                                                                                                // whose comparison feeds into atq arb_winner_v

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: ATQ enqueue count, aqed active count, aqed active limit pipe
//-----------------------------------------------------------------------------------------------------

assign atq_input_req_v          = atq_input_arb_enq | atq_input_arb_cmp | atq_input_arb_sch ;

// atq_input_req_v is effectively the "pipeline valid" for the atq inputs
assign p0_atq_ctrl_pipe.hold    = p0_atq_ctrl_pipe_v_f & p1_atq_ctrl_pipe.hold ;
assign p0_atq_ctrl_pipe.en      = atq_input_req_v & ~ p0_atq_ctrl_pipe.hold ;
assign p0_atq_ctrl_pipe_v_nxt   = atq_input_req_v | p0_atq_ctrl_pipe.hold ;
assign p0_atq_ctrl_pipe_v_nxt_gated     = p0_atq_ctrl_pipe_v_nxt & ~ p0_atq_ctrl_pipe.hold ;    // rmw can't handle p0_v_nxt & p0_hold

assign enq_atq_fifo_pop_data_qid_p              = enq_atq_fifo_pop_data.parity ^ ( ^ ( enq_atq_fifo_pop_data.qtype ) ) ;
assign send_atm_to_cq_fifo_pop_data_qid_p       = send_atm_to_cq_fifo_pop_data.parity ^
                                                  ( ^ ( { send_atm_to_cq_fifo_pop_data.cq , send_atm_to_cq_fifo_pop_data.qidix } ) ) ;

always_comb begin
  p0_atq_ctrl_pipe_nxt                  = p0_atq_ctrl_pipe_f ;
  if ( p0_atq_ctrl_pipe.en ) begin
    p0_atq_ctrl_pipe_nxt                = '0 ;                                  // Safety belt just in case any bits missed
    p0_atq_ctrl_pipe_nxt.sch_v          = atq_input_arb_sch ;
    p0_atq_ctrl_pipe_nxt.sch_qid_p      = atq_input_arb_sch_qid.qid_p ;
    p0_atq_ctrl_pipe_nxt.enq_v          = atq_input_arb_enq ;
    p0_atq_ctrl_pipe_nxt.enq_qid_p      = enq_atq_fifo_pop_data_qid_p ;         // arb_enq can only=1 if FIFO is valid
    p0_atq_ctrl_pipe_nxt.cmp_v          = atq_input_arb_cmp ;
    p0_atq_ctrl_pipe_nxt.cmp_qid_p      = send_atm_to_cq_fifo_pop_data_qid_p ;  // arb_cmp can only=1 if FIFO is valid
    p0_atq_ctrl_pipe_nxt.blast_enq      = atq_input_arb_enq &
                                          ( ( p4_atq_sch_v_f &   ( enq_atq_fifo_pop_data.qid == p4_atq_sch_qid_f.qid ) ) |
                                            ( p3_atq_sch_start & ( enq_atq_fifo_pop_data.qid == p3_atq_sch_start_qid ) ) ) ;
    p0_atq_ctrl_pipe_nxt.blast_cmp      = atq_input_arb_cmp &
                                          ( ( p4_atq_sch_v_f &   ( send_atm_to_cq_fifo_pop_data.qid == p4_atq_sch_qid_f.qid ) ) |
                                            ( p3_atq_sch_start & ( send_atm_to_cq_fifo_pop_data.qid == p3_atq_sch_start_qid ) ) ) ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p0_atq_ctrl_pipe_f            <= p0_atq_ctrl_pipe_nxt ;
  p1_atq_ctrl_pipe_f            <= p1_atq_ctrl_pipe_nxt ;
  p2_atq_ctrl_pipe_f            <= p2_atq_ctrl_pipe_nxt ;
end // always

assign p1_atq_ctrl_pipe.hold    = p1_atq_ctrl_pipe_v_f & p2_atq_ctrl_pipe.hold ;
assign p1_atq_ctrl_pipe.en      = p0_atq_ctrl_pipe_v_f & ~ p1_atq_ctrl_pipe.hold ;

assign p2_atq_ctrl_pipe.hold    = p2_atq_ctrl_pipe_v_f & p3_atq_ctrl_pipe.hold ;
assign p2_atq_ctrl_pipe.en      = p1_atq_ctrl_pipe_v_f & ~ p2_atq_ctrl_pipe.hold ;

assign p3_atq_ctrl_pipe.hold    = 1'b0 ;                                        // p3 qid status FFs always able to load
assign p3_atq_ctrl_pipe.en      = p2_atq_ctrl_pipe_v_f & ~ p3_atq_ctrl_pipe.hold ;

assign p4_atq_ctrl_pipe_en      = p3_atq_ctrl_pipe_v_f ;

always_comb begin
  p1_atq_ctrl_pipe_nxt          = p1_atq_ctrl_pipe_f ;
  p2_atq_ctrl_pipe_nxt          = p2_atq_ctrl_pipe_f ;

  if ( p1_atq_ctrl_pipe.en ) begin
    p1_atq_ctrl_pipe_nxt                = p0_atq_ctrl_pipe_f ;
    p1_atq_ctrl_pipe_nxt.blast_enq      = p0_atq_ctrl_pipe_f.blast_enq |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p0_atq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p0_atq_ctrl_pipe_f.enq_v ) ;
    p1_atq_ctrl_pipe_nxt.blast_cmp      = p0_atq_ctrl_pipe_f.blast_cmp |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p0_atq_aqed_act_cnt_rmw_pipe_f_pnc.qid ) &
                                            p0_atq_ctrl_pipe_f.cmp_v ) ;
  end
  else if ( p1_atq_ctrl_pipe.hold ) begin       // Need to blast writes which are holding
    p1_atq_ctrl_pipe_nxt.blast_enq      = p1_atq_ctrl_pipe_f.blast_enq |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p1_atq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_atq_ctrl_pipe_f.enq_v ) ;
    p1_atq_ctrl_pipe_nxt.blast_cmp      = p1_atq_ctrl_pipe_f.blast_cmp |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p1_atq_aqed_act_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_atq_ctrl_pipe_f.cmp_v ) ;
  end

  if ( p2_atq_ctrl_pipe.en ) begin
    p2_atq_ctrl_pipe_nxt                = p1_atq_ctrl_pipe_f ;
    p2_atq_ctrl_pipe_nxt.blast_enq      = p1_atq_ctrl_pipe_f.blast_enq |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p1_atq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_atq_ctrl_pipe_f.enq_v ) ;
    p2_atq_ctrl_pipe_nxt.blast_cmp      = p1_atq_ctrl_pipe_f.blast_cmp |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p1_atq_aqed_act_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_atq_ctrl_pipe_f.cmp_v ) ;
  end
  else if ( p2_atq_ctrl_pipe.hold ) begin       // Need to blast writes which are holding
    p2_atq_ctrl_pipe_nxt.blast_enq      = p2_atq_ctrl_pipe_f.blast_enq |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p2_atq_enq_cnt_rmw_pipe_f.qid ) &
                                            p2_atq_ctrl_pipe_f.enq_v ) ;
    p2_atq_ctrl_pipe_nxt.blast_cmp      = p2_atq_ctrl_pipe_f.blast_cmp |
                                          ( p3_atq_sch_start & ( p3_atq_sch_start_qid == p2_atq_aqed_act_cnt_rmw_pipe_f.qid ) &
                                            p2_atq_ctrl_pipe_f.cmp_v ) ;
  end
end // always

assign p2_atq_enq_cnt_upd_v             = ( p2_atq_enq_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_atq_ctrl_pipe.en ;
assign p2_atq_tot_enq_cnt_upd_v         = ( p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_atq_ctrl_pipe.en ;
assign p2_atq_aqed_act_cnt_upd_v        = ( p2_atq_aqed_act_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_atq_ctrl_pipe.en ;
assign p2_atq_atm_active_sum_v          = p2_atq_aqed_act_cnt_upd_v ;

always_comb begin
  if ( atq_input_arb_sch | atq_input_arb_enq ) begin
    p0_atq_enq_cnt_rmw_pipe_nxt.rw_cmd          = HQM_AW_RMWPIPE_RMW ;
  end
  else begin
    p0_atq_enq_cnt_rmw_pipe_nxt.rw_cmd          = HQM_AW_RMWPIPE_NOOP ;
  end
  if ( atq_input_arb_sch | atq_input_arb_cmp ) begin
    p0_atq_aqed_act_cnt_rmw_pipe_nxt.rw_cmd     = HQM_AW_RMWPIPE_RMW ;
    p0_atq_aqed_act_lim_rw_pipe_nxt.rw_cmd      = HQM_AW_RWPIPE_READ ;
    p0_atq_atm_active_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_READ ;         // Writes only occur via RMW bypsss
    p0_atq_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_READ ;
  end
  else begin
    p0_atq_aqed_act_cnt_rmw_pipe_nxt.rw_cmd     = HQM_AW_RMWPIPE_NOOP ;
    p0_atq_aqed_act_lim_rw_pipe_nxt.rw_cmd      = HQM_AW_RWPIPE_NOOP ;
    p0_atq_atm_active_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_NOOP ;
    p0_atq_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd    = HQM_AW_RWPIPE_NOOP ;
  end
  if ( atq_input_arb_enq )
    p0_atq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_RMW ;
  else
    p0_atq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd      = HQM_AW_RMWPIPE_NOOP ;
  if ( atq_input_arb_sch ) begin
    p0_atq_enq_cnt_rmw_pipe_nxt.qid             = atq_input_arb_sch_qid.qid ;
    p0_atq_aqed_act_cnt_rmw_pipe_nxt.qid        = atq_input_arb_sch_qid.qid ;
    p0_atq_aqed_act_lim_rw_pipe_nxt.qid         = atq_input_arb_sch_qid.qid ;
    p0_atq_atm_active_rmw_pipe_nxt.qid          = atq_input_arb_sch_qid.qid ;
    p0_atq_qid_dpth_thrsh_rw_pipe_nxt.qid       = atq_input_arb_sch_qid.qid ;
  end
  else begin
    p0_atq_enq_cnt_rmw_pipe_nxt.qid             = enq_atq_fifo_pop_data.qid ;           // enq
    p0_atq_aqed_act_cnt_rmw_pipe_nxt.qid        = send_atm_to_cq_fifo_pop_data.qid ;    // "cmp"
    p0_atq_aqed_act_lim_rw_pipe_nxt.qid         = send_atm_to_cq_fifo_pop_data.qid ;    // "cmp"
    p0_atq_atm_active_rmw_pipe_nxt.qid          = send_atm_to_cq_fifo_pop_data.qid ;    // "cmp"
    p0_atq_qid_dpth_thrsh_rw_pipe_nxt.qid       = send_atm_to_cq_fifo_pop_data.qid ;    // "cmp"
  end
  p0_atq_tot_enq_cnt_rmw_pipe_nxt.qid           = enq_atq_fifo_pop_data.qid ;
  p0_atq_enq_cnt_rmw_pipe_nxt.data              = { $bits ( lsp_atq_enq_cnt_t ) { 1'b0 } } ;            // Unused - cfg write done elsewhere
  p0_atq_atm_active_rmw_pipe_nxt.data           = { $bits ( lsp_atq_atm_active_t ) { 1'b0 } } ;         // Unused - cfg write done elsewhere
  p0_atq_qid_dpth_thrsh_rw_pipe_nxt.data        = { $bits ( lsp_atq_qid_dpth_thrsh_t ) { 1'b0 } } ;     // Unused - cfg write done elsewhere
  p0_atq_aqed_act_cnt_rmw_pipe_nxt.data         = { $bits ( lsp_atq_aqed_act_cnt_t ) { 1'b0 } } ;       // Unused - cfg write done elsewhere
  p0_atq_aqed_act_lim_rw_pipe_nxt.data          = { $bits ( lsp_atq_aqed_act_lim_t ) { 1'b0 } } ;       // Unused - cfg write done elsewhere
  p0_atq_tot_enq_cnt_rmw_pipe_nxt.data          = { $bits ( lsp_arch_cnt_t ) { 1'b0 } } ;               // Unused - cfg write done elsewhere
end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for atq enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ATQ_ENQ_CNT_MEM_WIDTH )
) i_atq_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_enq_cnt_rmw_pipe_status )

        // cmd input
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_atq_ctrl_pipe_v_f )
        , .p0_rw_f              ( p0_atq_enq_cnt_rmw_pipe_f_pnc.rw_cmd )        // Unused
        , .p0_addr_f            ( p0_atq_enq_cnt_rmw_pipe_f_pnc.qid )           // Used by blast logic
        , .p0_data_f            ( p0_atq_enq_cnt_rmw_pipe_f_pnc.data )          // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_ctrl_pipe_v_f )
        , .p1_rw_f              ( p1_atq_enq_cnt_rmw_pipe_f_pnc.rw_cmd )        // Unused
        , .p1_addr_f            ( p1_atq_enq_cnt_rmw_pipe_f_pnc.qid )           // Used by blast logic
        , .p1_data_f            ( p1_atq_enq_cnt_rmw_pipe_f_pnc.data )          // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_ctrl_pipe_v_f )
        , .p2_rw_f              ( p2_atq_enq_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_atq_enq_cnt_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_atq_enq_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_atq_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_atq_enq_cnt_upd )
        , .p3_v_f               ( p3_atq_ctrl_pipe_v_f )
        , .p3_rw_f              ( p3_atq_enq_cnt_rmw_pipe_f_nc.rw_cmd )         // Unused
        , .p3_addr_f            ( p3_atq_enq_cnt_rmw_pipe_f_nc.qid )            // Unused
        , .p3_data_f            ( p3_atq_enq_cnt_rmw_pipe_f_nc.data )           // Unused

        // mem intf
        , .mem_write            ( func_qid_atq_enqueue_count_mem_we )
        , .mem_read             ( func_qid_atq_enqueue_count_mem_re )
        , .mem_write_addr       ( func_qid_atq_enqueue_count_mem_waddr )
        , .mem_read_addr        ( func_qid_atq_enqueue_count_mem_raddr )
        , .mem_write_data       ( func_qid_atq_enqueue_count_mem_wdata )
        , .mem_read_data        ( func_qid_atq_enqueue_count_mem_rdata )
    ) ;

hqm_AW_residue_add i_atq_enq_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p2_atq_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_atq_enq_cnt_res_p1 )
) ;

hqm_AW_residue_sub i_atq_enq_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p2_atq_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_atq_enq_cnt_res_m1 )
) ;

assign { p2_atq_enq_cnt_p1_carry , p2_atq_enq_cnt_p1 }  = { 1'b0 , p2_atq_enq_cnt_rmw_pipe_f.data.cnt } + 15'h1 ;
assign { p2_atq_enq_cnt_m1_borrow , p2_atq_enq_cnt_m1 } = { 1'b0 , p2_atq_enq_cnt_rmw_pipe_f.data.cnt } - 15'h1 ;

always_comb begin
  p2_atq_enq_cnt_oflow_cond                     = 1'b0 ;
  p2_atq_enq_cnt_uflow_cond                     = 1'b0 ;
  if ( p2_atq_ctrl_pipe_f.sch_v ) begin
    if ( p2_atq_enq_cnt_m1_borrow ) begin
      p2_atq_enq_cnt_upd                        = p2_atq_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_atq_enq_cnt_uflow_cond                 = 1'b1 ;
    end
    else begin
      p2_atq_enq_cnt_upd.cnt                    = p2_atq_enq_cnt_m1 ;
      p2_atq_enq_cnt_upd.cnt_res                = p2_atq_enq_cnt_res_m1 ;
    end
  end
  else begin
    if ( p2_atq_enq_cnt_p1_carry ) begin
      p2_atq_enq_cnt_upd                        = p2_atq_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_atq_enq_cnt_oflow_cond                 = 1'b1 ;
    end
    else begin
      p2_atq_enq_cnt_upd.cnt                    = p2_atq_enq_cnt_p1 ;
      p2_atq_enq_cnt_upd.cnt_res                = p2_atq_enq_cnt_res_p1 ;
    end
  end
end // always

assign p2_atq_enq_cnt_upd_gt0                   = | ( p2_atq_enq_cnt_upd.cnt ) ;

assign p2_atq_enq_cnt_res_chk_en                = p2_atq_enq_cnt_upd_v ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ATQ_ENQ_CNT_WIDTH ) ) i_atq_enq_cnt_res_chk (
          .r                    ( p2_atq_enq_cnt_upd.cnt_res )
        , .d                    ( p2_atq_enq_cnt_upd.cnt )
        , .e                    ( p2_atq_enq_cnt_res_chk_en )
        , .err                  ( p2_atq_enq_cnt_res_err_cond )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for atm active count
// Only covers span of atq enqueue, but accessible when aqed_active is also being read.
// This count is added to the aqed_active count as an input to the count vs. depth calculation, effectively
// covering the lifespan of atq plus atm.
// Reads are in sync with aqed_act_cnt accesses, writes are accomplished via bypass input and occur when the
// atq_enq_cnt is being updated.  When an atq schedule occurs, atq_atm_active will have a read operation at p2
// due to the aqed_act_cnt increment, and a bypass write operation due to the atq_enq_cnt decrement.
// AW_rmw handles bypass r/w collisions, so regfile will be decremented.
// cm_code calculation is pipelined to avoid deep path: p2_atq_enq_cnt -> upd -> sum -> tot -> (calc_thresh_code) -> cm_code

assign p3_atq_atm_active_bypdata_sel_nxt        = p2_atq_enq_cnt_upd_v ;
assign p3_atq_atm_active_bypdata_nxt            = p2_atq_enq_cnt_upd ;
assign p3_atq_atm_active_bypaddr_sel_nxt        = p2_atq_enq_cnt_upd_v ;
assign p3_atq_atm_active_bypaddr_nxt            = p2_atq_enq_cnt_rmw_pipe_f.qid ;

hqm_AW_rmw_mem_4pipe_waddr #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ATQ_ATM_ACTIVE_MEM_WIDTH )
) i_atq_atm_active_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_atm_active_rmw_pipe_status_nc )         // Unused, same as aqed_act_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_atm_active_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_atm_active_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_atm_active_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_atq_atm_active_rmw_pipe_v_f_nc )         // Unused: same as aqed_act_cnt pipe
        , .p0_rw_f              ( p0_atq_atm_active_rmw_pipe_rw_f_nc )        // Unused
        , .p0_addr_f            ( p0_atq_atm_active_rmw_pipe_addr_f_nc )      // Unused
        , .p0_data_f            ( p0_atq_atm_active_rmw_pipe_data_f_nc )      // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_atm_active_rmw_pipe_v_f_nc )         // Unused: same as aqed_act_cnt pipe
        , .p1_rw_f              ( p1_atq_atm_active_rmw_pipe_rw_f_nc )        // Unused
        , .p1_addr_f            ( p1_atq_atm_active_rmw_pipe_addr_f_nc )      // Unused
        , .p1_data_f            ( p1_atq_atm_active_rmw_pipe_data_f_nc )      // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_atm_active_rmw_pipe_v_f_nc )         // Unused: same as aqed_act_cnt pipe
        , .p2_rw_f              ( p2_atq_atm_active_rmw_pipe_f_pnc.rw_cmd )   // Unused
        , .p2_addr_f            ( p2_atq_atm_active_rmw_pipe_f_pnc.qid )
        , .p2_data_f            ( p2_atq_atm_active_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_bypdata_sel_nxt   ( p3_atq_atm_active_bypdata_sel_nxt )
        , .p3_bypdata_nxt       ( p3_atq_atm_active_bypdata_nxt )
        , .p3_bypaddr_sel_nxt   ( p3_atq_atm_active_bypaddr_sel_nxt )
        , .p3_bypaddr_nxt       ( p3_atq_atm_active_bypaddr_nxt )

        , .p3_v_f               ( p3_atq_atm_active_rmw_pipe_v_f_nc )         // Unused: same as aqed_act_cnt pipe
        , .p3_rw_f              ( p3_atq_atm_active_rmw_pipe_f_nc.rw_cmd )    // Unused
        , .p3_addr_f            ( p3_atq_atm_active_rmw_pipe_f_nc.qid )       // Unused
        , .p3_data_f            ( p3_atq_atm_active_rmw_pipe_f_nc.data )      // Unused

        // mem intf
        , .mem_write            ( func_qid_atm_active_mem_we )
        , .mem_read             ( func_qid_atm_active_mem_re )
        , .mem_write_addr       ( func_qid_atm_active_mem_waddr )
        , .mem_read_addr        ( func_qid_atm_active_mem_raddr )
        , .mem_write_data       ( func_qid_atm_active_mem_wdata )
        , .mem_read_data        ( func_qid_atm_active_mem_rdata )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for atomic depth threshold
// Reads occur in sync with aqed_act_cnt updates since that's when it's needed for the cm_code calculation.

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ATQ_QID_DPTH_THRSH_MEM_WIDTH )
) i_atq_qid_dpth_thrsh_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_qid_dpth_thrsh_rw_pipe_status_nc )          // Unused: same as atq_aqed_act_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_qid_dpth_thrsh_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_qid_dpth_thrsh_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_qid_dpth_thrsh_rw_pipe_nxt.data )
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_atq_qid_dpth_thrsh_rw_pipe_v_f_nc )          // Unused: same as atq_enq_cnt pipe
        , .p0_rw_f              ( p0_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc )         // Unused
        , .p0_addr_f            ( p0_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc )       // Unused
        , .p0_data_f            ( p0_atq_qid_dpth_thrsh_rw_pipe_data_f_nc )       // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_qid_dpth_thrsh_rw_pipe_v_f_nc )          // Unused: same as atq_enq_cnt pipe
        , .p1_rw_f              ( p1_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc )         // Unused
        , .p1_addr_f            ( p1_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc )       // Unused
        , .p1_data_f            ( p1_atq_qid_dpth_thrsh_rw_pipe_data_f_nc )       // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_qid_dpth_thrsh_rw_pipe_v_f_nc )          // Unused: same as qid_enq_cnt_pipe
        , .p2_rw_f              ( p2_atq_qid_dpth_thrsh_rw_pipe_f_pnc.rw_cmd )    // Unused
        , .p2_addr_f            ( p2_atq_qid_dpth_thrsh_rw_pipe_f_pnc.qid )       // Unused
        , .p2_data_f            ( p2_atq_qid_dpth_thrsh_rw_pipe_f_pnc.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_v_f               ( p3_atq_qid_dpth_thrsh_rw_pipe_v_f_nc )          // Unused
        , .p3_rw_f              ( p3_atq_qid_dpth_thrsh_rw_pipe_rw_f_nc )         // Unused
        , .p3_addr_f            ( p3_atq_qid_dpth_thrsh_rw_pipe_addr_f_nc )       // Unused
        , .p3_data_f            ( p3_atq_qid_dpth_thrsh_rw_pipe_data_f_nc )       // Unused

        // mem intf
        , .mem_write            ( func_cfg_atm_qid_dpth_thrsh_mem_we )
        , .mem_read             ( func_cfg_atm_qid_dpth_thrsh_mem_re )
        , .mem_addr             ( func_cfg_atm_qid_dpth_thrsh_mem_addr )
        , .mem_write_data       ( func_cfg_atm_qid_dpth_thrsh_mem_wdata )
        , .mem_read_data        ( func_cfg_atm_qid_dpth_thrsh_mem_rdata )
    ) ;

always_comb begin
  if ( p2_atq_ctrl_pipe_f.sch_v ) begin
    p2_atq_atm_active_curr                      = p2_atq_enq_cnt_upd ;                          // SCH: ATQ count decremented for scheduled qe; aqed_act_cnt will already include +1
  end
  else begin
    p2_atq_atm_active_curr                      = p2_atq_atm_active_rmw_pipe_f_pnc.data ;       // CMP: Current ATQ value, not changed on completion
  end
end // always

always_comb begin
  p3_atq_atm_active_sum_v_nxt                   = 1'b0 ;
  p3_atq_aqed_act_cnt_upd_nxt                   = p3_atq_aqed_act_cnt_upd_f ;
  p3_atq_atm_active_curr_nxt                    = p3_atq_atm_active_curr_f ;
  p3_atq_qid_dpth_thrsh_nxt                     = p3_atq_qid_dpth_thrsh_f ;
  p3_atq_aqed_act_cnt_qid_nxt                   = p3_atq_aqed_act_cnt_qid_f ;
  if ( p2_atq_atm_active_sum_v ) begin
    p3_atq_atm_active_sum_v_nxt                 = 1'b1 ;
    p3_atq_aqed_act_cnt_upd_nxt                 = p2_atq_aqed_act_cnt_upd ;
    p3_atq_atm_active_curr_nxt                  = p2_atq_atm_active_curr ;
    p3_atq_qid_dpth_thrsh_nxt                   = p2_atq_qid_dpth_thrsh_rw_pipe_f_pnc.data ;
    p3_atq_aqed_act_cnt_qid_nxt                 = p2_atq_aqed_act_cnt_rmw_pipe_f.qid [HQM_NUM_LB_QIDB2-1:0] ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_atq_atm_active_sum_v_f                   <= 1'b0 ;
  end
  else begin
    p3_atq_atm_active_sum_v_f                   <= p3_atq_atm_active_sum_v_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p3_atq_aqed_act_cnt_upd_f                     <= p3_atq_aqed_act_cnt_upd_nxt ;
  p3_atq_atm_active_curr_f                      <= p3_atq_atm_active_curr_nxt ;
  p3_atq_qid_dpth_thrsh_f                       <= p3_atq_qid_dpth_thrsh_nxt ;
  p3_atq_aqed_act_cnt_qid_f                     <= p3_atq_aqed_act_cnt_qid_nxt ;
end // always

hqm_AW_residue_add i_atq_atm_active_res_add (
          .a                    ( p3_atq_aqed_act_cnt_upd_f.cnt_res )
        , .b                    ( p3_atq_atm_active_curr_f.cnt_res )
        , .r                    ( p3_atq_atm_active_sum.cnt_res )
) ;

always_comb begin
  { p3_atq_atm_active_sum_carry , p3_atq_atm_active_sum.cnt }   = { 1'b0 , 2'h0 , p3_atq_aqed_act_cnt_upd_f.cnt } + { 1'b0 , p3_atq_atm_active_curr_f.cnt } ;

  p3_atq_atm_active_oflow_cond                  = 1'b0 ;
  p3_atq_atm_active_tot                         = p3_atq_atm_active_curr_f ;
  if ( p3_atq_atm_active_sum_v_f ) begin
    if ( p3_atq_atm_active_sum_carry ) begin
      p3_atq_atm_active_tot                     = p3_atq_atm_active_curr_f ;    // Don't multiply errors
      p3_atq_atm_active_oflow_cond              = 1'b1 ;
    end
    else begin
      p3_atq_atm_active_tot                     = p3_atq_atm_active_sum ;
    end
  end
end // always

assign p3_atq_atm_active_res_chk_en             = p3_atq_atm_active_sum_v_f ;
assign p3_atq_qid_dpth_thrsh_par_chk_en         = p3_atq_atm_active_sum_v_f ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ATQ_ATM_ACTIVE_WIDTH ) ) i_atq_atm_active_res_chk (
          .r                    ( p3_atq_atm_active_tot.cnt_res )
        , .d                    ( p3_atq_atm_active_tot.cnt )
        , .e                    ( p3_atq_atm_active_res_chk_en )
        , .err                  ( p3_atq_atm_active_res_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH ) ) i_atq_qid_dpth_thrsh_par_chk (
          .p                    ( p3_atq_qid_dpth_thrsh_f.thrsh_p )
        , .d                    ( p3_atq_qid_dpth_thrsh_f.thrsh )
        , .e                    ( p3_atq_qid_dpth_thrsh_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p3_atq_qid_dpth_thrsh_par_err_cond )
) ;

assign p3_atq_qid_dpth_thrsh_cm_code    = hqm_lsp_calc_thresh_code (   p3_atq_atm_active_tot.cnt
                                                                     , p3_atq_qid_dpth_thrsh_f.thrsh ) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for atq aqed active count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ATQ_AQED_ACT_CNT_MEM_WIDTH )
) i_atq_aqed_act_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_aqed_act_cnt_rmw_pipe_status_nc )         // Unused, same as atq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_aqed_act_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_aqed_act_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_aqed_act_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_atq_aqed_act_cnt_rmw_pipe_v_f_nc )         // Unused: same as atq_enq_cnt pipe
        , .p0_rw_f              ( p0_atq_aqed_act_cnt_rmw_pipe_f_pnc.rw_cmd )   // Unused
        , .p0_addr_f            ( p0_atq_aqed_act_cnt_rmw_pipe_f_pnc.qid )      // Used by blast logic
        , .p0_data_f            ( p0_atq_aqed_act_cnt_rmw_pipe_f_pnc.data )     // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_aqed_act_cnt_rmw_pipe_v_f_nc )         // Unused: same as atq_enq_cnt pipe
        , .p1_rw_f              ( p1_atq_aqed_act_cnt_rmw_pipe_f_pnc.rw_cmd )   // Unused
        , .p1_addr_f            ( p1_atq_aqed_act_cnt_rmw_pipe_f_pnc.qid )      // Used by blast logic
        , .p1_data_f            ( p1_atq_aqed_act_cnt_rmw_pipe_f_pnc.data )     // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_aqed_act_cnt_rmw_pipe_v_f_nc )         // Unused: same as atq_enq_cnt pipe
        , .p2_rw_f              ( p2_atq_aqed_act_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_atq_aqed_act_cnt_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_atq_aqed_act_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_atq_aqed_act_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_atq_aqed_act_cnt_upd )
        , .p3_v_f               ( p3_atq_aqed_act_cnt_rmw_pipe_v_f_nc )         // Unused: same as atq_enq_cnt pipe
        , .p3_rw_f              ( p3_atq_aqed_act_cnt_rmw_pipe_f_nc.rw_cmd )    // Unused
        , .p3_addr_f            ( p3_atq_aqed_act_cnt_rmw_pipe_f_nc.qid )       // Unused
        , .p3_data_f            ( p3_atq_aqed_act_cnt_rmw_pipe_f_nc.data )      // Unused

        // mem intf
        , .mem_write            ( func_qid_aqed_active_count_mem_we )
        , .mem_read             ( func_qid_aqed_active_count_mem_re )
        , .mem_write_addr       ( func_qid_aqed_active_count_mem_waddr )
        , .mem_read_addr        ( func_qid_aqed_active_count_mem_raddr )
        , .mem_write_data       ( func_qid_aqed_active_count_mem_wdata )
        , .mem_read_data        ( func_qid_aqed_active_count_mem_rdata )
) ;

hqm_AW_residue_add i_atq_aqed_act_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p2_atq_aqed_act_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_atq_aqed_act_cnt_res_p1 )
) ;
hqm_AW_residue_sub i_atq_aqed_act_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p2_atq_aqed_act_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_atq_aqed_act_cnt_res_m1 )
) ;

assign { p2_atq_aqed_act_cnt_p1_carry , p2_atq_aqed_act_cnt_p1 }        = { 1'b0 , p2_atq_aqed_act_cnt_rmw_pipe_f.data.cnt } + 13'h1 ;
assign { p2_atq_aqed_act_cnt_m1_borrow , p2_atq_aqed_act_cnt_m1 }       = { 1'b0 , p2_atq_aqed_act_cnt_rmw_pipe_f.data.cnt } - 13'h1 ;

always_comb begin
  p2_atq_aqed_act_cnt_oflow_cond                        = 1'b0 ;
  p2_atq_aqed_act_cnt_uflow_cond                        = 1'b0 ;
  if ( p2_atq_ctrl_pipe_f.sch_v ) begin
    if ( p2_atq_aqed_act_cnt_p1_carry ) begin
      p2_atq_aqed_act_cnt_upd                           = p2_atq_aqed_act_cnt_rmw_pipe_f.data ;         // Saturate, no residue error
      p2_atq_aqed_act_cnt_oflow_cond                    = 1'b1 ;
    end
    else begin
      p2_atq_aqed_act_cnt_upd.cnt                       = p2_atq_aqed_act_cnt_p1 ;
      p2_atq_aqed_act_cnt_upd.cnt_res                   = p2_atq_aqed_act_cnt_res_p1 ;
    end
  end
  else begin
    if ( p2_atq_aqed_act_cnt_m1_borrow ) begin
      p2_atq_aqed_act_cnt_upd                           = p2_atq_aqed_act_cnt_rmw_pipe_f.data ;         // Saturate, no residue error
      p2_atq_aqed_act_cnt_uflow_cond                    = 1'b1 ;
    end
    else begin
      p2_atq_aqed_act_cnt_upd.cnt                       = p2_atq_aqed_act_cnt_m1 ;
      p2_atq_aqed_act_cnt_upd.cnt_res                   = p2_atq_aqed_act_cnt_res_m1 ;
    end
  end
end // always

assign p2_atq_aqed_act_cnt_upd_lt_lim           = ( p2_atq_aqed_act_cnt_upd.cnt < p2_atq_aqed_act_lim_rw_pipe_f_pnc.data.lim ) ;
assign p2_atq_aqed_act_cnt_upd_gt_0             = | p2_atq_aqed_act_cnt_upd.cnt ;
assign p2_atq_aqed_act_cnt_upd_eq_0             = ~ p2_atq_aqed_act_cnt_upd_gt_0 ;

//--------
// Increment occurs when schedule is generated from p3.
// Decrement occurs when cmp advances from p2 to p3
assign p3_atq_tot_act_cnt_upd_inc       = p3_atq_sch_req ;                      // Already includes hold/enable
assign p3_atq_tot_act_cnt_upd_dec       = p2_atq_ctrl_pipe_v_f & p2_atq_ctrl_pipe_f.cmp_v & ~ p3_atq_ctrl_pipe.hold ;
assign p3_atq_tot_act_cnt_upd_v         = p3_atq_tot_act_cnt_upd_inc | p3_atq_tot_act_cnt_upd_dec ;

hqm_AW_residue_add i_atq_tot_act_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p3_atq_tot_act_cnt_f.cnt_res )
        , .r                    ( p3_atq_tot_act_cnt_res_p1 )
) ;
hqm_AW_residue_sub i_atq_tot_act_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p3_atq_tot_act_cnt_f.cnt_res )
        , .r                    ( p3_atq_tot_act_cnt_res_m1 )
) ;

assign { p3_atq_tot_act_cnt_p1_carry , p3_atq_tot_act_cnt_p1 }          = { 1'b0 , p3_atq_tot_act_cnt_f.cnt } + {{HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH{1'b0}}, 1'b1} ;
assign { p3_atq_tot_act_cnt_m1_borrow , p3_atq_tot_act_cnt_m1 }         = { 1'b0 , p3_atq_tot_act_cnt_f.cnt } - {{HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH{1'b0}}, 1'b1} ;

always_comb begin
  p3_atq_tot_act_cnt_oflow_cond                         = 1'b0 ;
  p3_atq_tot_act_cnt_uflow_cond                         = 1'b0 ;
  p3_atq_tot_act_cnt_upd                                = p3_atq_tot_act_cnt_f ;

  // Simultaneous is possible
  case ( { p3_atq_tot_act_cnt_upd_inc , p3_atq_tot_act_cnt_upd_dec } )
    2'b01 : begin
      if ( p3_atq_tot_act_cnt_m1_borrow ) begin
        p3_atq_tot_act_cnt_upd                  = p3_atq_tot_act_cnt_f ;                        // Saturate, no residue error
        p3_atq_tot_act_cnt_uflow_cond           = 1'b1 ;
      end
      else begin
        p3_atq_tot_act_cnt_upd.cnt              = p3_atq_tot_act_cnt_m1 ;
        p3_atq_tot_act_cnt_upd.cnt_res          = p3_atq_tot_act_cnt_res_m1 ;
      end
    end // 01
    2'b10 : begin
      if ( p3_atq_tot_act_cnt_p1_carry ) begin
        p3_atq_tot_act_cnt_upd                  = p3_atq_tot_act_cnt_f ;                        // Saturate, no residue error
        p3_atq_tot_act_cnt_oflow_cond           = 1'b1 ;
      end
      else begin
        p3_atq_tot_act_cnt_upd.cnt              = p3_atq_tot_act_cnt_p1 ;
        p3_atq_tot_act_cnt_upd.cnt_res          = p3_atq_tot_act_cnt_res_p1 ;
      end
    end // 10
    default : begin                     // Same as default assigns above
        p3_atq_tot_act_cnt_oflow_cond           = 1'b0 ;
        p3_atq_tot_act_cnt_uflow_cond           = 1'b0 ;
        p3_atq_tot_act_cnt_upd                  = p3_atq_tot_act_cnt_f ;
    end
  endcase
end // always

assign p3_atq_tot_act_cnt_lt_lim                = ( p3_atq_tot_act_cnt_f.cnt <  cfg_aqed_tot_enqueue_limit_f ) ;
assign p3_atq_tot_act_cnt_eq_lim                = ( p3_atq_tot_act_cnt_f.cnt == cfg_aqed_tot_enqueue_limit_f ) ;
assign p3_atq_tot_act_cnt_gt_lim                = ( p3_atq_tot_act_cnt_f.cnt >  cfg_aqed_tot_enqueue_limit_f ) ;

// Should be correctly adjusted as part of a successful vas reset drain
always_comb begin
  cfg_aqed_tot_enqueue_count_nxt                = cfg_aqed_tot_enqueue_count_f ;
  if ( p3_atq_tot_act_cnt_upd_v ) begin
    cfg_aqed_tot_enqueue_count_nxt              = p3_atq_tot_act_cnt_upd ;
  end
end // always

assign p3_atq_tot_act_cnt_f                     = cfg_aqed_tot_enqueue_count_f ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH ) ) i_aqed_tot_enq_cnt_res_chk (
          .r                    ( cfg_aqed_tot_enqueue_count_f.cnt_res )
        , .d                    ( cfg_aqed_tot_enqueue_count_f.cnt )
        , .e                    ( p3_atq_tot_act_cnt_upd_v )
        , .err                  ( p3_atq_aqed_tot_enq_cnt_res_err_cond )
) ;

//--------
assign p3_atq_fid_inflight_cnt_upd_inc  = p3_atq_sch_req ;                      // Already includes hold/enable
assign p3_atq_fid_inflight_cnt_upd_dec  = aqed_lsp_dec_fid_cnt_v_f ;            // Pulse from aqed
assign p3_atq_fid_inflight_cnt_upd_v    = p3_atq_fid_inflight_cnt_upd_inc | p3_atq_fid_inflight_cnt_upd_dec ;

hqm_AW_residue_add i_atq_fid_inflight_count_res_add (
          .a                    ( 2'h1 )
        , .b                    ( cfg_fid_inflight_count_f.cnt_res )
        , .r                    ( p3_atq_fid_inflight_cnt_res_p1 )
) ;
hqm_AW_residue_sub i_atq_fid_inflight_count_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( cfg_fid_inflight_count_f.cnt_res )
        , .r                    ( p3_atq_fid_inflight_cnt_res_m1 )
) ;
assign { p3_atq_fid_inflight_cnt_p1_carry , p3_atq_fid_inflight_cnt_p1 }        = { 1'b0 , cfg_fid_inflight_count_f.cnt } + 13'h1 ;
assign { p3_atq_fid_inflight_cnt_m1_borrow , p3_atq_fid_inflight_cnt_m1 }       = { 1'b0 , cfg_fid_inflight_count_f.cnt } - 13'h1 ;


always_comb begin
  p3_atq_fid_inflight_cnt_oflow_cond            = 1'b0 ;
  p3_atq_fid_inflight_cnt_uflow_cond            = 1'b0 ;
  p3_atq_fid_inflight_cnt_upd                   = cfg_fid_inflight_count_f ;
  // Simultaneous is possible
  case ( { p3_atq_fid_inflight_cnt_upd_inc , p3_atq_fid_inflight_cnt_upd_dec } )
    2'b01 : begin
      if ( p3_atq_fid_inflight_cnt_m1_borrow ) begin
        p3_atq_fid_inflight_cnt_upd             = cfg_fid_inflight_count_f ;                    // Saturate, no residue error
        p3_atq_fid_inflight_cnt_uflow_cond      = 1'b1 ;
      end
      else begin
        p3_atq_fid_inflight_cnt_upd.cnt         = p3_atq_fid_inflight_cnt_m1 ;
        p3_atq_fid_inflight_cnt_upd.cnt_res     = p3_atq_fid_inflight_cnt_res_m1 ;
      end
    end // 01
    2'b10 : begin
      if ( p3_atq_fid_inflight_cnt_p1_carry ) begin
        p3_atq_fid_inflight_cnt_upd             = cfg_fid_inflight_count_f ;                    // Saturate, no residue error
        p3_atq_fid_inflight_cnt_oflow_cond      = 1'b1 ;
      end
      else begin
        p3_atq_fid_inflight_cnt_upd.cnt         = p3_atq_fid_inflight_cnt_p1 ;
        p3_atq_fid_inflight_cnt_upd.cnt_res     = p3_atq_fid_inflight_cnt_res_p1 ;
      end
    end // 10
    default : begin                     // Same as default assigns above
      p3_atq_fid_inflight_cnt_oflow_cond        = 1'b0 ;
      p3_atq_fid_inflight_cnt_uflow_cond        = 1'b0 ;
      p3_atq_fid_inflight_cnt_upd               = cfg_fid_inflight_count_f ;
    end
  endcase
end // always

assign p3_atq_fid_inflight_cnt_lt_lim           = ( cfg_fid_inflight_count_f.cnt <  cfg_fid_inflight_limit_f ) ;
assign p3_atq_fid_inflight_cnt_eq_lim           = ( cfg_fid_inflight_count_f.cnt == cfg_fid_inflight_limit_f ) ;
assign p3_atq_fid_inflight_cnt_gt_lim           = ( cfg_fid_inflight_count_f.cnt >  cfg_fid_inflight_limit_f ) ;

always_comb begin
  cfg_fid_inflight_count_nxt                    = cfg_fid_inflight_count_f ;
  if ( p3_atq_fid_inflight_cnt_upd_v )
    cfg_fid_inflight_count_nxt                  = p3_atq_fid_inflight_cnt_upd ;
end // always

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ATQ_FID_IF_CNT_WIDTH ) ) i_atq_fid_inflight_cnt_res_chk (
          .r                    ( cfg_fid_inflight_count_f.cnt_res )
        , .d                    ( cfg_fid_inflight_count_f.cnt )
        , .e                    ( p3_atq_fid_inflight_cnt_upd_v )
        , .err                  ( p3_atq_fid_inflight_cnt_res_err_cond )
) ;


//-------------------------------------------------------------------------------------------------
// Manage storage for atq aqed active limit
hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ATQ_AQED_ACT_LIM_MEM_WIDTH )
) i_atq_aqed_act_lim_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_aqed_act_lim_rw_pipe_status_nc )          // Unused: same as atq_aqed_act_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_aqed_act_lim_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_aqed_act_lim_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_aqed_act_lim_rw_pipe_nxt.data )
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_atq_aqed_act_lim_rw_pipe_v_f_nc )          // Unused: same as atq_enq_cnt pipe
        , .p0_rw_f              ( p0_atq_aqed_act_lim_rw_pipe_rw_f_nc )         // Unused
        , .p0_addr_f            ( p0_atq_aqed_act_lim_rw_pipe_addr_f_nc )       // Unused
        , .p0_data_f            ( p0_atq_aqed_act_lim_rw_pipe_data_f_nc )       // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_aqed_act_lim_rw_pipe_v_f_nc )          // Unused: same as atq_enq_cnt pipe
        , .p1_rw_f              ( p1_atq_aqed_act_lim_rw_pipe_rw_f_nc )         // Unused
        , .p1_addr_f            ( p1_atq_aqed_act_lim_rw_pipe_addr_f_nc )       // Unused
        , .p1_data_f            ( p1_atq_aqed_act_lim_rw_pipe_data_f_nc )       // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_aqed_act_lim_rw_pipe_v_f_nc )          // Unused: same as qid_enq_cnt_pipe
        , .p2_rw_f              ( p2_atq_aqed_act_lim_rw_pipe_f_pnc.rw_cmd )    // Unused
        , .p2_addr_f            ( p2_atq_aqed_act_lim_rw_pipe_f_pnc.qid )       // Unused
        , .p2_data_f            ( p2_atq_aqed_act_lim_rw_pipe_f_pnc.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_v_f               ( p3_atq_aqed_act_lim_rw_pipe_v_f_nc )          // Unused
        , .p3_rw_f              ( p3_atq_aqed_act_lim_rw_pipe_rw_f_nc )         // Unused
        , .p3_addr_f            ( p3_atq_aqed_act_lim_rw_pipe_addr_f_nc )       // Unused
        , .p3_data_f            ( p3_atq_aqed_act_lim_rw_pipe_data_f_nc )       // Unused

        // mem intf
        , .mem_write            ( func_cfg_qid_aqed_active_limit_mem_we )
        , .mem_read             ( func_cfg_qid_aqed_active_limit_mem_re )
        , .mem_addr             ( func_cfg_qid_aqed_active_limit_mem_addr )
        , .mem_write_data       ( func_cfg_qid_aqed_active_limit_mem_wdata )
        , .mem_read_data        ( func_cfg_qid_aqed_active_limit_mem_rdata )
    ) ;

assign p2_atq_aqed_act_cnt_res_chk_en              = p2_atq_aqed_act_cnt_upd_v ;
assign p2_atq_aqed_act_lim_par_chk_en              = p2_atq_aqed_act_cnt_res_chk_en ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH ) ) i_atq_aqed_act_cnt_res_chk (
          .r                    ( p2_atq_aqed_act_cnt_upd.cnt_res )
        , .d                    ( p2_atq_aqed_act_cnt_upd.cnt )
        , .e                    ( p2_atq_aqed_act_cnt_res_chk_en )
        , .err                  ( p2_atq_aqed_act_cnt_res_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ATQ_AQED_ACT_LIM_WIDTH ) ) i_atq_act_lim_par_chk (
          .p                    ( p2_atq_aqed_act_lim_rw_pipe_f_pnc.data.lim_p )
        , .d                    ( p2_atq_aqed_act_lim_rw_pipe_f_pnc.data.lim )
        , .e                    ( p2_atq_aqed_act_lim_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_atq_aqed_act_lim_par_err_cond )
) ;

assign p2_atq_inp_enq_qid_par_chk_en    = p2_atq_enq_cnt_upd_v ;
assign p2_atq_inp_cmp_qid_par_chk_en    = p2_atq_aqed_act_cnt_upd_v ;

always_comb begin
  if ( p2_atq_ctrl_pipe_f.sch_v ) begin
    p2_atq_inp_enq_qid_p                = p2_atq_ctrl_pipe_f.sch_qid_p ;
    p2_atq_inp_cmp_qid_p                = p2_atq_ctrl_pipe_f.sch_qid_p ;
  end
  else begin
    p2_atq_inp_enq_qid_p                = p2_atq_ctrl_pipe_f.enq_qid_p ;
    p2_atq_inp_cmp_qid_p                = p2_atq_ctrl_pipe_f.cmp_qid_p ;
  end
end // always

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_atq_inp_enq_qid_par_chk (
          .p                    ( p2_atq_inp_enq_qid_p )
        , .d                    ( p2_atq_enq_cnt_rmw_pipe_f.qid )
        , .e                    ( p2_atq_inp_enq_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_atq_inp_enq_qid_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_atq_inp_cmp_qid_par_chk (
          .p                    ( p2_atq_inp_cmp_qid_p )
        , .d                    ( p2_atq_aqed_act_cnt_rmw_pipe_f.qid )
        , .e                    ( p2_atq_inp_cmp_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_atq_inp_cmp_qid_par_err_cond )
) ;

assign p2_atq_inp_qid_par_err_cond      = p2_atq_inp_enq_qid_par_err_cond | p2_atq_inp_cmp_qid_par_err_cond ;


//-------------------------------------------------------------------------------------------------
// Manage storage for atq total enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_ARCH_CNT_MEM_WIDTH )
) i_atq_tot_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( atq_tot_enq_cnt_rmw_pipe_status_nc )          // Unused, same as atq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_atq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_atq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_atq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_atq_tot_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_atq_tot_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_atq_tot_enq_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p0_rw_f              ( p0_atq_tot_enq_cnt_rmw_pipe_rw_f_nc )         // Unused
        , .p0_addr_f            ( p0_atq_tot_enq_cnt_rmw_pipe_addr_f_nc )       // Unused
        , .p0_data_f            ( p0_atq_tot_enq_cnt_rmw_pipe_data_f_nc )       // Unused

        , .p1_hold              ( p1_atq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_atq_tot_enq_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p1_rw_f              ( p1_atq_tot_enq_cnt_rmw_pipe_rw_f_nc )         // Unused
        , .p1_addr_f            ( p1_atq_tot_enq_cnt_rmw_pipe_addr_f_nc )       // Unused
        , .p1_data_f            ( p1_atq_tot_enq_cnt_rmw_pipe_data_f_nc )       // Unused

        , .p2_hold              ( p2_atq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_atq_tot_enq_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p2_rw_f              ( p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd )    // Used for upd_v
        , .p2_addr_f            ( p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.qid )       // Unused
        , .p2_data_f            ( p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p3_atq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_atq_tot_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_atq_tot_enq_cnt_upd )
        , .p3_v_f               ( p3_atq_tot_enq_cnt_rmw_pipe_v_f_nc )          // Unused
        , .p3_rw_f              ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd )    // Used for res_chk_en
        , .p3_addr_f            ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.qid )       // Unused
        , .p3_data_f            ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.data )      // Used for res_chk

        // mem intf
        , .mem_write            ( cfgsc_func_qid_atm_tot_enq_cnt_mem_we )
        , .mem_read             ( func_qid_atm_tot_enq_cnt_mem_re )
        , .mem_write_addr       ( cfgsc_func_qid_atm_tot_enq_cnt_mem_waddr )
        , .mem_read_addr        ( func_qid_atm_tot_enq_cnt_mem_raddr )
        , .mem_write_data       ( cfgsc_func_qid_atm_tot_enq_cnt_mem_wdata )
        , .mem_read_data        ( func_qid_atm_tot_enq_cnt_mem_rdata )
    ) ;

hqm_AW_residue_add i_atq_tot_enq_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .r                    ( p2_atq_tot_enq_cnt_res_p1 )
) ;

assign p2_atq_tot_enq_cnt_p1            = p2_atq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt + 64'h1 ;          // wrap

assign p2_atq_tot_enq_cnt_upd.cnt       = p2_atq_tot_enq_cnt_p1 ;
assign p2_atq_tot_enq_cnt_upd.cnt_res   = p2_atq_tot_enq_cnt_res_p1 ;

assign p3_atq_tot_enq_cnt_res_chk_en    = p4_atq_ctrl_pipe_en & ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ARCH_CNT_WIDTH ) ) i_atq_tot_enq_cnt_res_chk (
          .r                    ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .d                    ( p3_atq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt )
        , .e                    ( p3_atq_tot_enq_cnt_res_chk_en )
        , .err                  ( p4_atq_tot_enq_cnt_res_err_nxt )
) ;

//-------------------------------------------------------------------------------------------------
// Underflow/overflow errors - some are impossible, some may be caused by software/config errors
//
always_comb begin
  // Don't hold - 1-clock pulse to report
  p3_atq_enq_cnt_uflow_err_nxt          = 1'b0 ;
  p3_atq_enq_cnt_oflow_err_nxt          = 1'b0 ;
  p3_atq_aqed_act_cnt_uflow_err_nxt     = 1'b0 ;
  p3_atq_aqed_act_cnt_oflow_err_nxt     = 1'b0 ;

  p4_atq_tot_act_cnt_uflow_err_nxt      = 1'b0 ;
  p4_atq_tot_act_cnt_oflow_err_nxt      = 1'b0 ;
  p4_atq_fid_inflight_cnt_uflow_err_nxt = 1'b0 ;
  p4_atq_fid_inflight_cnt_oflow_err_nxt = 1'b0 ;

  p3_atq_enq_cnt_res_err_nxt            = 1'b0 ;
  p3_atq_aqed_act_cnt_res_err_nxt       = 1'b0 ;
  p3_atq_aqed_act_lim_par_err_nxt       = 1'b0 ;
  p3_atq_inp_qid_par_err_nxt            = 1'b0 ;

  p4_atq_atm_active_oflow_err_nxt       = 1'b0 ;
  p4_atq_atm_active_res_err_nxt         = 1'b0 ;
  p4_atq_qid_dpth_thrsh_par_err_nxt     = 1'b0 ;

  p4_atq_aqed_tot_enq_cnt_res_err_nxt   = 1'b0 ;
  p4_atq_fid_inflight_cnt_res_err_nxt   = 1'b0 ;

  if ( p2_atq_ctrl_pipe_v_f & ~ p3_atq_ctrl_pipe.hold ) begin
    p3_atq_enq_cnt_uflow_err_nxt        = p2_atq_ctrl_pipe_f.sch_v & p2_atq_enq_cnt_uflow_cond ;
    p3_atq_enq_cnt_oflow_err_nxt        = p2_atq_ctrl_pipe_f.enq_v & p2_atq_enq_cnt_oflow_cond ;
    p3_atq_aqed_act_cnt_uflow_err_nxt   = p2_atq_ctrl_pipe_f.cmp_v & p2_atq_aqed_act_cnt_uflow_cond ;
    p3_atq_aqed_act_cnt_oflow_err_nxt   = p2_atq_ctrl_pipe_f.sch_v & p2_atq_aqed_act_cnt_oflow_cond ;

    p3_atq_enq_cnt_res_err_nxt          = p2_atq_enq_cnt_res_err_cond ;
    p3_atq_aqed_act_cnt_res_err_nxt     = p2_atq_aqed_act_cnt_res_err_cond ;
    p3_atq_aqed_act_lim_par_err_nxt     = p2_atq_aqed_act_lim_par_err_cond | cfg_error_inject_f [ 2 ] ;
    p3_atq_inp_qid_par_err_nxt          = p2_atq_inp_qid_par_err_cond ;
  end
  if ( p3_atq_atm_active_sum_v_f ) begin
    p4_atq_atm_active_oflow_err_nxt     = p3_atq_atm_active_oflow_cond ;
    p4_atq_atm_active_res_err_nxt       = p3_atq_atm_active_res_err_cond ;
    p4_atq_qid_dpth_thrsh_par_err_nxt   = p3_atq_qid_dpth_thrsh_par_err_cond ;
  end
  if ( p3_atq_fid_inflight_cnt_upd_v ) begin
    p4_atq_fid_inflight_cnt_oflow_err_nxt       = p3_atq_fid_inflight_cnt_oflow_cond ;
    p4_atq_fid_inflight_cnt_uflow_err_nxt       = p3_atq_fid_inflight_cnt_uflow_cond ;
    p4_atq_fid_inflight_cnt_res_err_nxt         = p3_atq_fid_inflight_cnt_res_err_cond ;
  end
  if ( p3_atq_tot_act_cnt_upd_v ) begin
    p4_atq_tot_act_cnt_uflow_err_nxt    = p3_atq_tot_act_cnt_uflow_cond ;
    p4_atq_tot_act_cnt_oflow_err_nxt    = p3_atq_tot_act_cnt_oflow_cond ;
    p4_atq_aqed_tot_enq_cnt_res_err_nxt = p3_atq_aqed_tot_enq_cnt_res_err_cond ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_atq_enq_cnt_uflow_err_f          <= 1'b0 ;
    p3_atq_enq_cnt_oflow_err_f          <= 1'b0 ;
    p3_atq_aqed_act_cnt_uflow_err_f     <= 1'b0 ;
    p3_atq_aqed_act_cnt_oflow_err_f     <= 1'b0 ;

    p4_atq_tot_act_cnt_uflow_err_f      <= 1'b0 ;
    p4_atq_tot_act_cnt_oflow_err_f      <= 1'b0 ;
    p4_atq_fid_inflight_cnt_uflow_err_f <= 1'b0 ;
    p4_atq_fid_inflight_cnt_oflow_err_f <= 1'b0 ;

    p3_atq_enq_cnt_res_err_f            <= 1'b0 ;
    p3_atq_aqed_act_cnt_res_err_f       <= 1'b0 ;
    p3_atq_aqed_act_lim_par_err_f       <= 1'b0 ;
    p3_atq_inp_qid_par_err_f            <= 1'b0 ;

    p4_atq_atm_active_oflow_err_f       <= 1'b0 ;
    p4_atq_atm_active_res_err_f         <= 1'b0 ;
    p4_atq_qid_dpth_thrsh_par_err_f     <= 1'b0 ;
    p4_atq_aqed_tot_enq_cnt_res_err_f   <= 1'b0 ;
    p4_atq_fid_inflight_cnt_res_err_f   <= 1'b0 ;
    p4_atq_tot_enq_cnt_res_err_f        <= 1'b0 ;
  end
  else begin
    p3_atq_enq_cnt_uflow_err_f          <= p3_atq_enq_cnt_uflow_err_nxt ;
    p3_atq_enq_cnt_oflow_err_f          <= p3_atq_enq_cnt_oflow_err_nxt ;
    p3_atq_aqed_act_cnt_uflow_err_f     <= p3_atq_aqed_act_cnt_uflow_err_nxt ;
    p3_atq_aqed_act_cnt_oflow_err_f     <= p3_atq_aqed_act_cnt_oflow_err_nxt ;

    p4_atq_tot_act_cnt_uflow_err_f      <= p4_atq_tot_act_cnt_uflow_err_nxt ;
    p4_atq_tot_act_cnt_oflow_err_f      <= p4_atq_tot_act_cnt_oflow_err_nxt ;
    p4_atq_fid_inflight_cnt_uflow_err_f <= p4_atq_fid_inflight_cnt_uflow_err_nxt ;
    p4_atq_fid_inflight_cnt_oflow_err_f <= p4_atq_fid_inflight_cnt_oflow_err_nxt ;

    p3_atq_enq_cnt_res_err_f            <= p3_atq_enq_cnt_res_err_nxt ;
    p3_atq_aqed_act_cnt_res_err_f       <= p3_atq_aqed_act_cnt_res_err_nxt ;
    p3_atq_aqed_act_lim_par_err_f       <= p3_atq_aqed_act_lim_par_err_nxt ;
    p3_atq_inp_qid_par_err_f            <= p3_atq_inp_qid_par_err_nxt ;

    p4_atq_atm_active_oflow_err_f       <= p4_atq_atm_active_oflow_err_nxt ;
    p4_atq_atm_active_res_err_f         <= p4_atq_atm_active_res_err_nxt ;
    p4_atq_qid_dpth_thrsh_par_err_f     <= p4_atq_qid_dpth_thrsh_par_err_nxt ;
    p4_atq_aqed_tot_enq_cnt_res_err_f   <= p4_atq_aqed_tot_enq_cnt_res_err_nxt ;
    p4_atq_fid_inflight_cnt_res_err_f   <= p4_atq_fid_inflight_cnt_res_err_nxt ;
    p4_atq_tot_enq_cnt_res_err_f        <= p4_atq_tot_enq_cnt_res_err_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: ATQ p3 qid_v, aqed_nfull and aqed_empty status vectors
//-----------------------------------------------------------------------------------------------------
// See comments under DIRENQ regarding scheduling terminology

assign atq_fid_cnt_upd_v_nxt            = aqed_lsp_fid_cnt_upd_v ;
assign atq_fid_cnt_upd_val_nxt          = aqed_lsp_fid_cnt_upd_val ;
assign atq_fid_cnt_upd_qid_nxt          = aqed_lsp_fid_cnt_upd_qid ;
assign atq_fid_cnt_upd_last_v_nxt       = atq_fid_cnt_upd_v_f ;
assign atq_fid_cnt_upd_idle             = ~ atq_fid_cnt_upd_v_f & ~ atq_fid_cnt_upd_last_v_f ;  // Need second stage to cover p3_atq_qid_en_f which feeds into atq arb_winner_v

assign atq_stop_atqatm_nxt              = aqed_lsp_stop_atqatm ;
assign atq_stop_atqatm_last_nxt         = atq_stop_atqatm_f ;
assign atq_stop_atqatm_change           = atq_stop_atqatm_f ^ atq_stop_atqatm_last_f ;
assign atq_stop_atqatm_idle             = ~ atq_stop_atqatm_change ;                            // Only need single stage, feeds into atq arb_winner_v

hqm_AW_bindec #( .WIDTH( HQM_NUM_LB_QIDB2 ) ) i_p3_atq_sch_start_qid_bindec (
          .a                            ( p3_atq_sch_start_qid [HQM_NUM_LB_QIDB2-1:0] )
        , .enable                       ( p3_atq_sch_start )
        , .dec                          ( p3_atq_sch_hit )
) ;

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
    // Bypass update from sch takes precedence over update from p2; sch update will cause subsequent write
    // of latest/correct value of counts caused by this scheduling.
    // enq/cmp updates from upper pipe must be supressed from "enabling" if they were blasted by newer scheduling.
    p3_atq_p2_enq_hit[i]                = p3_atq_ctrl_pipe.en & ( p2_atq_ctrl_pipe_f.enq_v | p2_atq_ctrl_pipe_f.sch_v ) &
                                          ( p2_atq_enq_cnt_rmw_pipe_f.qid == i ) & ~ p2_atq_ctrl_pipe_f.blast_enq ;
    p3_atq_p2_cmp_hit[i]                = p3_atq_ctrl_pipe.en & ( p2_atq_ctrl_pipe_f.cmp_v | p2_atq_ctrl_pipe_f.sch_v ) &
                                          ( p2_atq_aqed_act_cnt_rmw_pipe_f.qid == i ) & ~ p2_atq_ctrl_pipe_f.blast_cmp ;
  end // for
end // always

// For each atq qid maintain state for "qid has data" (qid_v), "aqed not full" (aqed_nfull) and "aqed empty".
// Update (set to 0 or 1) when enq count or aqed avail count is updated, reset when that qid is selected to be scheduled.
// All should be cleared as part of a successful vas reset drain
always_comb begin
  p3_atq_qid_v_nxt                              = p3_atq_qid_v_f ;
  if ( p3_atq_sch_start | p3_atq_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      if ( p3_atq_sch_hit [i] ) begin
        p3_atq_qid_v_nxt [i]                    = 1'b0 ;
      end
      else if ( p3_atq_p2_enq_hit [i] ) begin
        p3_atq_qid_v_nxt [i]                    = p2_atq_enq_cnt_upd_gt0 ;
      end
    end // for i
  end // if

  p4_atq_cm_code_nxt                            = p4_atq_cm_code_f ;
  if ( cfgsc_cfg_atm_qid_dpth_thrsh_mem_we | p3_atq_atm_active_sum_v_f ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      if ( cfgsc_cfg_atm_qid_dpth_thrsh_mem_we & ( cfg_mem_addr [HQM_NUM_LB_QIDB2-1:0] == i ) ) begin
        p4_atq_cm_code_nxt [i]                  = 2'h0 ;
      end
      else if ( p3_atq_atm_active_sum_v_f & ( p3_atq_aqed_act_cnt_qid_f == i ) ) begin   // sch_v or cmp_v
        p4_atq_cm_code_nxt [i]                  = p3_atq_qid_dpth_thrsh_cm_code ;
      end
    end // for i
  end // if

  p3_atq_aqed_nfull_nxt                         = p3_atq_aqed_nfull_f ;
  p3_atq_aqed_empty_nxt                         = p3_atq_aqed_empty_f ;
  p3_atq_aqed_act_v_nxt                         = p3_atq_aqed_act_v_f ;
  if ( p3_atq_sch_start | p3_atq_ctrl_pipe.en | cfg_ldb_sched_control_aqed_nfull_v ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      if ( p3_atq_sch_hit [i] ) begin
        p3_atq_aqed_nfull_nxt [i]               = 1'b0 ;
        p3_atq_aqed_empty_nxt [i]               = 1'b0 ;
        p3_atq_aqed_act_v_nxt [i]               = 1'b1 ;
      end
      else if ( p3_atq_p2_cmp_hit[i] ) begin
        p3_atq_aqed_nfull_nxt [i]               = p2_atq_aqed_act_cnt_upd_lt_lim ;
        p3_atq_aqed_empty_nxt [i]               = p2_atq_aqed_act_cnt_upd_eq_0 ;
        p3_atq_aqed_act_v_nxt [i]               = p2_atq_aqed_act_cnt_upd_gt_0 ;
      end
      if ( cfg_ldb_sched_control_aqed_nfull_v & ( cfg_ldb_sched_control_qid == i ) ) begin
        p3_atq_aqed_nfull_nxt [i]               = cfg_ldb_sched_control_value ;
      end
    end // for i
  end // if

  p3_atq_qid_en_nxt                             = p3_atq_qid_en_f ;
  if ( atq_fid_cnt_upd_v_f ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      if ( atq_fid_cnt_upd_v_f & ( atq_fid_cnt_upd_qid_f == i ) ) begin
        p3_atq_qid_en_nxt [i]                   = atq_fid_cnt_upd_val_f ;
      end
    end // for i
  end // if
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_atq_aqed_nfull_f                         <= { HQM_NUM_LB_QID { 1'b1 } } ;
    p3_atq_aqed_empty_f                         <= { HQM_NUM_LB_QID { 1'b1 } } ;
    p3_atq_qid_v_f                              <= { HQM_NUM_LB_QID { 1'b0 } } ;

    atq_fid_cnt_upd_v_f                         <= 1'b0 ;
    atq_fid_cnt_upd_val_f                       <= 1'b0 ;
    atq_fid_cnt_upd_qid_f                       <= { HQM_LSP_ARCH_NUM_LB_QIDB2 { 1'b0 } } ;
    atq_fid_cnt_upd_last_v_f                    <= 1'b0 ;
    atq_stop_atqatm_f                           <= 1'b0 ;
    atq_stop_atqatm_last_f                      <= 1'b0 ;
    p3_atq_qid_en_f                             <= { HQM_NUM_LB_QID { 1'b1 } } ;
    p3_atq_aqed_act_v_f                         <= { HQM_NUM_LB_QID { 1'b0 } } ;

    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      p4_atq_cm_code_f [i]                      <= 2'h0 ;
    end
  end
  else begin
    p3_atq_aqed_nfull_f                         <= p3_atq_aqed_nfull_nxt ;
    p3_atq_aqed_empty_f                         <= p3_atq_aqed_empty_nxt ;
    p3_atq_qid_v_f                              <= p3_atq_qid_v_nxt ;

    atq_fid_cnt_upd_v_f                         <= atq_fid_cnt_upd_v_nxt ;
    atq_fid_cnt_upd_val_f                       <= atq_fid_cnt_upd_val_nxt ;
    atq_fid_cnt_upd_qid_f                       <= atq_fid_cnt_upd_qid_nxt ;
    atq_fid_cnt_upd_last_v_f                    <= atq_fid_cnt_upd_last_v_nxt ;
    atq_stop_atqatm_f                           <= atq_stop_atqatm_nxt ;
    atq_stop_atqatm_last_f                      <= atq_stop_atqatm_last_nxt ;
    p3_atq_qid_en_f                             <= p3_atq_qid_en_nxt ;
    p3_atq_aqed_act_v_f                         <= p3_atq_aqed_act_v_nxt ;

    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      p4_atq_cm_code_f [i]                      <= p4_atq_cm_code_nxt [i] ;
    end
  end // else rst_n

end // always

assign p3_atq_qid_avail                 = p3_atq_qid_en_f ;

always_comb begin
  p3_atq_nfull_arb_reqs                 = p3_atq_qid_v_f & p3_atq_aqed_nfull_f & p3_atq_qid_avail ;
  p3_atq_empty_arb_reqs                 = p3_atq_qid_v_f & p3_atq_aqed_empty_f & p3_atq_qid_avail ;

  cfg_qid_atq_sch_v_status              = p3_atq_qid_v_f ;
  cfg_qid_atq_aqed_avail_status         = p3_atq_aqed_nfull_f ;
  // Note: per-qid aqed_empty status can be determined from config-readable "aqed active".  AND readable in diag status 0
end // always

// Use external index to keep the two arbiters in sync
hqm_AW_rr_arb_windex # ( .NUM_REQS ( HQM_NUM_LB_QID ) ) i_atq_nfull_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p3_atq_nfull_arb_reqs )
        , .index_f              ( p3_atq_arb_index_0_f )
        , .winner_v             ( p3_atq_nfull_arb_winner_v )
        , .winner               ( p3_atq_nfull_arb_winner )
) ;

hqm_AW_rr_arb_windex # ( .NUM_REQS ( HQM_NUM_LB_QID ) ) i_atq_empty_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p3_atq_empty_arb_reqs )
        , .index_f              ( p3_atq_arb_index_1_f )
        , .winner_v             ( p3_atq_empty_arb_winner_pre_v )
        , .winner               ( p3_atq_empty_arb_winner )
) ;
assign p3_atq_empty_arb_winner_v        = p3_atq_empty_arb_winner_pre_v & ~ cfg_control_disable_atq_empty_arb ;

// Give priority to empty aqed to put reasonable max bounds on how long it will take a given atq qid to be
// "scheduled" (moved from atq to atm) when space becomes available.
always_comb begin
  if ( p3_atq_empty_arb_winner_v ) begin
    p3_atq_arb_winner_pre_v     = 1'b1 ;
    p3_atq_arb_winner           = p3_atq_empty_arb_winner ;
  end
  else begin
    p3_atq_arb_winner_pre_v     = p3_atq_nfull_arb_winner_v ;
    p3_atq_arb_winner           = p3_atq_nfull_arb_winner ;
  end
  p3_atq_arb_winner_p1          = p3_atq_arb_winner + { { ( HQM_NUM_LB_QIDB2-1) { 1'b0 } } , 1'b1 } ;
end // always

assign p3_atq_arb_winner_v      = p3_atq_arb_winner_pre_v   & p3_atq_fid_inflight_cnt_lt_lim & p3_atq_tot_act_cnt_lt_lim &
                                  ~ atq_stop_atqatm_f & ~ cause_pipe_idle ;

// No need to include redundant (for purposes of idle) "empty arb" logic or transient config access
assign cfg_atq_arb_winner_v_nxt = p3_atq_nfull_arb_winner_v & p3_atq_fid_inflight_cnt_lt_lim & p3_atq_tot_act_cnt_lt_lim &
                                  ~ atq_stop_atqatm_f ;


hqm_AW_parity_gen #( .WIDTH( HQM_NUM_LB_QIDB2 ) ) i_atq_qid_par_gen (
          .d            ( p3_atq_arb_winner )
        , .odd          ( 1'b1 )
        , .p            ( p3_atq_arb_winner_gp )
) ;

assign p3_atq_sch_req                   = p3_atq_arb_winner_v & ~ atq_sel_ap_fifo_hold & ~ p4_atq_sch_hold ;
assign p3_atq_sch_stall_smon            = p3_atq_arb_winner_v &   atq_sel_ap_fifo_hold & ~ p4_atq_sch_hold ;    // For smon only

always_comb begin
  p3_atq_sch_req_qid.qid                        = { HQM_LSP_ARCH_NUM_LB_QIDB2 { 1'b0 } } ;
  p3_atq_sch_req_qid.qid [HQM_NUM_LB_QIDB2-1:0] = p3_atq_arb_winner ;
  p3_atq_sch_req_qid.qid_p                      = p3_atq_arb_winner_gp ;
end // always

assign p3_atq_arb_update                = p3_atq_sch_req ;

assign p3_atq_sch_start                 = p3_atq_sch_req ;
assign p3_atq_sch_start_qid             = p3_atq_sch_req_qid.qid ;

assign p4_atq_sch_hold                  = p4_atq_sch_v_f & ~ atq_input_arb_sch ;
assign p4_atq_sch_v_nxt                 = p3_atq_sch_req | p4_atq_sch_hold ;

always_comb begin
  p3_atq_arb_index_0_nxt                = p3_atq_arb_index_0_f ;        // Duplicated for drive
  p3_atq_arb_index_1_nxt                = p3_atq_arb_index_1_f ;        // Duplicated for drive
  p4_atq_sch_qid_nxt                    = p4_atq_sch_qid_f ;

  if ( p3_atq_arb_update ) begin
    p3_atq_arb_index_0_nxt              = p3_atq_arb_winner_p1 ;
    p3_atq_arb_index_1_nxt              = p3_atq_arb_winner_p1 ;
  end 

  if ( p3_atq_sch_req & ~ p4_atq_sch_hold ) begin
    p4_atq_sch_qid_nxt                  = p3_atq_sch_req_qid ;
  end
end //always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_atq_arb_index_0_f                <= { HQM_NUM_LB_QIDB2 { 1'b0 } } ;
    p3_atq_arb_index_1_f                <= { HQM_NUM_LB_QIDB2 { 1'b0 } } ;
    p4_atq_sch_v_f                      <= 1'b0 ;
  end
  else begin
    p3_atq_arb_index_0_f                <= p3_atq_arb_index_0_nxt ;
    p3_atq_arb_index_1_f                <= p3_atq_arb_index_1_nxt ;
    p4_atq_sch_v_f                      <= p4_atq_sch_v_nxt ;
  end
end // always
always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p4_atq_sch_qid_f                    <= '0 ;
  end
  else begin
    p4_atq_sch_qid_f                    <= p4_atq_sch_qid_nxt ;
  end
end
//-------------------------------------------------------------------------------------------------
// Output FIFO (DB) - for static timing isolation
assign atq_sel_ap_fifo_push             = p3_atq_sch_req ;                      // sch_req already has afull in equation
assign atq_sel_ap_fifo_push_data.qid    = p3_atq_sch_req_qid.qid ;
assign atq_sel_ap_fifo_push_data.parity = p3_atq_sch_req_qid.qid_p ^ cfg_error_inject_f [ 13 ] ;

assign atq_sel_ap_db_in_valid           = atq_sel_ap_fifo_push ;
assign atq_sel_ap_db_in_data            = atq_sel_ap_fifo_push_data ;
assign atq_sel_ap_fifo_afull            = ~ atq_sel_ap_db_in_ready ;
assign atq_sel_ap_fifo_empty            = atq_sel_ap_tx_sync_idle ;
assign atq_sel_ap_fifo_hold             = atq_sel_ap_fifo_afull | ( cfg_control_single_out_atq & ~ atq_sel_ap_fifo_empty ) ;

// atq_sel_ap_db_in_data goes to i_hqm_AW_tx_sync_atq_sel_ap

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: DIRENQ pipe - Detects Directed enqueue notifications and schedules to the Dir Pipe unit
//*****************************************************************************************************
//*****************************************************************************************************

// SUBSECTION: DIRENQ input pipe arbitration
// Besides config, there are 3 inputs to the direnq enqueue and token pipes: enqueue requests (E),
// token returns (T) and schedule requests (S).  S ties up both pipes; T and E each tie up only their
// respective pipes.  In order to maximize efficiency, the logic only allows E and T requests to go
// if they are both present or if there are no S requests.  The algorithm is:
// S * E * T            : use arbiter; if S loses, allow both E and T to go (either way ties up both)
// S * ( ~E + ~T )      : Allow S to go (ties up both)
// ~S                   : Allow E or T (or both) to go if they are valid


assign dp_lsp_enq_dir_fifo_pop_data_v           = core_dp_lsp_enq_dir_v ;
assign dp_lsp_enq_dir_fifo_pop_data_vreq        = dp_lsp_enq_dir_fifo_pop_data_v & ~ cause_pipe_idle ;
assign dp_lsp_enq_dir_fifo_pop_data             = core_dp_lsp_enq_dir_data ;

assign core_dp_lsp_enq_dir_ready                = dp_lsp_enq_dir_fifo_pop ;
assign dp_lsp_enq_dir_fifo_pop                  = direnq_input_arb_enq ;


assign direnq_input_arb_new_both        = dp_lsp_enq_dir_fifo_pop_data_vreq & dir_tokrtn_fifo_pop_data_vreq ;
assign direnq_input_arb_new_either      = dp_lsp_enq_dir_fifo_pop_data_vreq | dir_tokrtn_fifo_pop_data_vreq ;
assign direnq_input_arb_reqs [0]        = direnq_input_arb_new_either & ( direnq_input_arb_new_both | ~ p4_direnq_sch_v_f ) ;

assign direnq_input_arb_reqs [1]        = p4_direnq_sch_v_f ;

assign direnq_input_arb_update          = p0_direnq_ctrl_pipe.en ;

// Note: rr used (instead of 50/50 wrand) because with wrand if extremely biased sch can go out of LSP but be stuck in p4 so long that
// corresponding token returns, wins the wrand arb and decrements (underflows) the token count.
hqm_AW_rr_arb # ( .NUM_REQS ( 2 ) ) i_direnq_input_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( direnq_input_arb_reqs )
        , .update               ( direnq_input_arb_update )
        , .winner_v             ( direnq_input_arb_winner_pre_v )
        , .winner               ( direnq_input_arb_winner )
) ;

assign direnq_input_arb_winner_v        = direnq_input_arb_winner_pre_v &
                                          ~ ( ( cfg_control_single_op_direnq & ( ( ~ direnq_upipe_idle_f ) | p0_direnq_ctrl_pipe_v_f ) ) |
                                              ( cfg_control_half_bw_direnq & p0_direnq_ctrl_pipe_v_f ) ) ;

assign direnq_input_arb_pre_enq = direnq_input_arb_winner_v & ~ direnq_input_arb_winner & ~ p0_direnq_ctrl_pipe.hold & dp_lsp_enq_dir_fifo_pop_data_vreq ;
assign direnq_input_arb_pre_tok = direnq_input_arb_winner_v & ~ direnq_input_arb_winner & ~ p0_direnq_ctrl_pipe.hold & dir_tokrtn_fifo_pop_data_vreq ;
assign direnq_input_arb_sch     = direnq_input_arb_winner_v &   direnq_input_arb_winner & ~ p0_direnq_ctrl_pipe.hold ;
assign direnq_input_arb_sch_qid = p4_direnq_sch_qid_f ;
assign direnq_input_arb_sch_beats       = { 1'b0 , p4_direnq_calc_rem_beats } + 3'h1 ;          // Total beats including this one (1..4)

// Disable if arbiter has allowed multiple ops and disabled by config and toggle does not allow
assign direnq_input_arb_enq     = direnq_input_arb_pre_enq & ~ ( cfg_control_disable_multi_op_direnq & direnq_input_arb_pre_tok & direnq_input_arb_tog_f ) ;
assign direnq_input_arb_tok     = direnq_input_arb_pre_tok & ~ ( cfg_control_disable_multi_op_direnq & direnq_input_arb_pre_enq & ~ direnq_input_arb_tog_f ) ;

always_comb begin
  direnq_input_arb_tog_nxt      = direnq_input_arb_tog_f ;
  if ( cfg_control_disable_multi_op_direnq & direnq_input_arb_pre_enq & direnq_input_arb_pre_tok )
    direnq_input_arb_tog_nxt    = ~ direnq_input_arb_tog_f ;
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    direnq_input_arb_tog_f      <= 1'b0 ;
  end
  else begin
    direnq_input_arb_tog_f      <= direnq_input_arb_tog_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: DIRENQ enqueue count, token count and token limit pipe
//-----------------------------------------------------------------------------------------------------
// The p3 status FFs are always able to be updated by the direnq_enq and direnq_tok pipes from p2.

assign direnq_input_req_v               = direnq_input_arb_enq | direnq_input_arb_tok | direnq_input_arb_sch ;

// direnq_input_req_v is effectively the "pipeline valid" for the direnq inputs
assign p0_direnq_ctrl_pipe.hold         = p0_direnq_ctrl_pipe_v_f & p1_direnq_ctrl_pipe.hold ;
assign p0_direnq_ctrl_pipe.en           = direnq_input_req_v & ~ p0_direnq_ctrl_pipe.hold ;
assign p0_direnq_ctrl_pipe_v_nxt        = direnq_input_req_v | p0_direnq_ctrl_pipe.hold ;
assign p0_direnq_ctrl_pipe_v_nxt_gated  = p0_direnq_ctrl_pipe_v_nxt & ~ p0_direnq_ctrl_pipe.hold ;

assign dir_tokrtn_fifo_pop_data_cq_p    = dir_tokrtn_fifo_pop_data.parity ^ dir_tokrtn_fifo_pop_data.is_ldb ;

always_comb begin
  p0_direnq_ctrl_pipe_nxt                       = p0_direnq_ctrl_pipe_f ;
  dir_tokrtn_fifo_pop_data_count_ms_nc          = dir_tokrtn_fifo_pop_data.count[12:11] ;       // Unused ms token count bits
  if ( p0_direnq_ctrl_pipe.en ) begin
    p0_direnq_ctrl_pipe_nxt                     = '0 ;                                  // Safety belt just in case any bits missed
    p0_direnq_ctrl_pipe_nxt.sch_v               = direnq_input_arb_sch ;
    p0_direnq_ctrl_pipe_nxt.sch_qid_p           = direnq_input_arb_sch_qid.qid_p ;
    p0_direnq_ctrl_pipe_nxt.sch_beats           = direnq_input_arb_sch_beats ;
    p0_direnq_ctrl_pipe_nxt.enq_v               = direnq_input_arb_enq ;
    p0_direnq_ctrl_pipe_nxt.enq_qid_p           = dp_lsp_enq_dir_fifo_pop_data.parity ; // arb_enq can only=1 if FIFO is valid
    p0_direnq_ctrl_pipe_nxt.tok_v               = direnq_input_arb_tok ;
    p0_direnq_ctrl_pipe_nxt.tok_cq_p            = dir_tokrtn_fifo_pop_data_cq_p ;       // arb_tok can only=1 if FIFO is valid
    p0_direnq_ctrl_pipe_nxt.tok_delta.cnt       = dir_tokrtn_fifo_pop_data.count[HQM_LSP_DIR_TOK_DELTA_WIDTH-1:0] ;
    p0_direnq_ctrl_pipe_nxt.tok_delta.cnt_res   = dir_tokrtn_fifo_pop_data.count_residue ;
    p0_direnq_ctrl_pipe_nxt.blast_enq           = direnq_input_arb_enq &
                                                  ( ( p4_direnq_sch_v_f &   ( dp_lsp_enq_dir_fifo_pop_data.qid == p4_direnq_sch_qid_f.qid ) ) |
                                                    ( p3_direnq_sch_start & ( dp_lsp_enq_dir_fifo_pop_data.qid == p3_direnq_sch_start_qid ) ) ) ;
    p0_direnq_ctrl_pipe_nxt.blast_tok           = direnq_input_arb_tok &
                                                  ( ( p4_direnq_sch_v_f &   ( dir_tokrtn_fifo_pop_data_cq == p4_direnq_sch_qid_f.qid ) ) |      // For DIR, CQ = QID
                                                    ( p3_direnq_sch_start & ( dir_tokrtn_fifo_pop_data_cq == p3_direnq_sch_start_qid ) ) ) ;    // For DIR, CQ = QID
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p0_direnq_ctrl_pipe_f                 <= p0_direnq_ctrl_pipe_nxt ;
  p1_direnq_ctrl_pipe_f                 <= p1_direnq_ctrl_pipe_nxt ;
  p2_direnq_ctrl_pipe_f                 <= p2_direnq_ctrl_pipe_nxt ;
end // always

assign p1_direnq_ctrl_pipe.hold         = p1_direnq_ctrl_pipe_v_f & p2_direnq_ctrl_pipe.hold ;
assign p1_direnq_ctrl_pipe.en           = p0_direnq_ctrl_pipe_v_f & ~ p1_direnq_ctrl_pipe.hold ;

assign p2_direnq_ctrl_pipe.hold         = p2_direnq_ctrl_pipe_v_f & p3_direnq_ctrl_pipe.hold ;
assign p2_direnq_ctrl_pipe.en           = p1_direnq_ctrl_pipe_v_f & ~ p2_direnq_ctrl_pipe.hold ;

assign p3_direnq_ctrl_pipe.hold         = 1'b0 ;                                        // p3 qid status FFs always able to load
assign p3_direnq_ctrl_pipe.en           = p2_direnq_ctrl_pipe_v_f & ~ p3_direnq_ctrl_pipe.hold ;

assign p4_direnq_ctrl_pipe_en           = p3_direnq_ctrl_pipe_v_f ;

always_comb begin
  p1_direnq_ctrl_pipe_nxt               = p1_direnq_ctrl_pipe_f ;
  p2_direnq_ctrl_pipe_nxt               = p2_direnq_ctrl_pipe_f ;

  if ( p1_direnq_ctrl_pipe.en ) begin   // Only blast when sch request gets in to p4 (for fill arbiter, only 1st clock of 4)
    p1_direnq_ctrl_pipe_nxt             = p0_direnq_ctrl_pipe_f ;
    p1_direnq_ctrl_pipe_nxt.blast_enq   = p0_direnq_ctrl_pipe_f.blast_enq |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p0_direnq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p0_direnq_ctrl_pipe_f.enq_v ) ;
    p1_direnq_ctrl_pipe_nxt.blast_tok   = p0_direnq_ctrl_pipe_f.blast_tok |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p0_direnq_tok_cnt_rmw_pipe_f_pnc.cq ) &
                                            p0_direnq_ctrl_pipe_f.tok_v ) ;
  end
  else if ( p1_direnq_ctrl_pipe.hold ) begin    // Need to blast writes which are holding
    p1_direnq_ctrl_pipe_nxt.blast_enq   = p1_direnq_ctrl_pipe_f.blast_enq |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p1_direnq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_direnq_ctrl_pipe_f.enq_v ) ;
    p1_direnq_ctrl_pipe_nxt.blast_tok   = p1_direnq_ctrl_pipe_f.blast_tok |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p1_direnq_tok_cnt_rmw_pipe_f_pnc.cq )  &
                                            p1_direnq_ctrl_pipe_f.tok_v ) ;
  end

  if ( p2_direnq_ctrl_pipe.en ) begin
    p2_direnq_ctrl_pipe_nxt             = p1_direnq_ctrl_pipe_f ;
    p2_direnq_ctrl_pipe_nxt.blast_enq   = p1_direnq_ctrl_pipe_f.blast_enq |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p1_direnq_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_direnq_ctrl_pipe_f.enq_v ) ;
    p2_direnq_ctrl_pipe_nxt.blast_tok   = p1_direnq_ctrl_pipe_f.blast_tok |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p1_direnq_tok_cnt_rmw_pipe_f_pnc.cq ) &
                                            p1_direnq_ctrl_pipe_f.tok_v ) ;
  end
  else if ( p2_direnq_ctrl_pipe.hold ) begin    // Need to blast writes which are holding
    p2_direnq_ctrl_pipe_nxt.blast_enq   = p2_direnq_ctrl_pipe_f.blast_enq |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p2_direnq_enq_cnt_rmw_pipe_f.qid ) &
                                            p2_direnq_ctrl_pipe_f.enq_v ) ;
    p2_direnq_ctrl_pipe_nxt.blast_tok   = p2_direnq_ctrl_pipe_f.blast_tok |
                                          ( p3_direnq_sch_start & ( p3_direnq_sch_start_qid == p2_direnq_tok_cnt_rmw_pipe_f.cq ) &
                                            p2_direnq_ctrl_pipe_f.tok_v ) ;
  end
end // always

assign p2_direnq_enq_cnt_upd_v          = ( p2_direnq_enq_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_direnq_ctrl_pipe.en ;
assign p2_direnq_tok_cnt_upd_v          = ( p2_direnq_tok_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_direnq_ctrl_pipe.en ;
assign p2_direnq_tot_enq_cnt_upd_v      = ( p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_direnq_ctrl_pipe.en ;
assign p2_direnq_tot_sch_cnt_upd_v      = ( p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_direnq_ctrl_pipe.en ;
assign p2_direnq_max_enq_depth_upd_v    = ( p2_direnq_max_enq_depth_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_READ ) & p3_direnq_ctrl_pipe.en & p2_direnq_enq_cnt_gt_max_depth ;

always_comb begin
  if ( direnq_input_arb_sch | direnq_input_arb_enq ) begin
    p0_direnq_enq_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_RMW ;
    p0_direnq_dpth_thrsh_rw_pipe_nxt.rw_cmd     = HQM_AW_RWPIPE_READ ;
    p0_direnq_max_enq_depth_rmw_pipe_nxt.rw_cmd = HQM_AW_RMWPIPE_READ ;         // Also check on sch (decrement) in case RW/C (sets to 0) is followed by sch and depth is > 0
                                                                                // Update occurs via bypass at going into p3 if curr upd depth > curr max
  end
  else begin
    p0_direnq_enq_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_NOOP ;
    p0_direnq_dpth_thrsh_rw_pipe_nxt.rw_cmd     = HQM_AW_RWPIPE_NOOP ;
    p0_direnq_max_enq_depth_rmw_pipe_nxt.rw_cmd = HQM_AW_RMWPIPE_NOOP ;
  end
  if ( direnq_input_arb_sch | direnq_input_arb_tok ) begin
    p0_direnq_tok_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_RMW ;
    p0_direnq_tok_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_READ ;
  end
  else begin
    p0_direnq_tok_cnt_rmw_pipe_nxt.rw_cmd       = HQM_AW_RMWPIPE_NOOP ;
    p0_direnq_tok_lim_rw_pipe_nxt.rw_cmd        = HQM_AW_RWPIPE_NOOP ;
  end
  if ( direnq_input_arb_enq )
    p0_direnq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd   = HQM_AW_RMWPIPE_RMW ;
  else
    p0_direnq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd   = HQM_AW_RMWPIPE_NOOP ;
  if ( direnq_input_arb_sch )
    p0_direnq_tot_sch_cnt_rmw_pipe_nxt.rw_cmd   = HQM_AW_RMWPIPE_RMW ;
  else
    p0_direnq_tot_sch_cnt_rmw_pipe_nxt.rw_cmd   = HQM_AW_RMWPIPE_NOOP ;
  //--------------------------------------------------------------------------
  if ( direnq_input_arb_sch ) begin
    p0_direnq_enq_cnt_rmw_pipe_nxt.qid          = direnq_input_arb_sch_qid.qid ;
    p0_direnq_dpth_thrsh_rw_pipe_nxt.qid        = direnq_input_arb_sch_qid.qid ;
    p0_direnq_tok_cnt_rmw_pipe_nxt.cq           = direnq_input_arb_sch_qid.qid ;        // direct mapping of qid to cq
    p0_direnq_tok_lim_rw_pipe_nxt.cq            = direnq_input_arb_sch_qid.qid ;        // direct mapping of qid to cq
    p0_direnq_max_enq_depth_rmw_pipe_nxt.qid    = direnq_input_arb_sch_qid.qid ;
  end
  else begin
    p0_direnq_enq_cnt_rmw_pipe_nxt.qid          = dp_lsp_enq_dir_fifo_pop_data.qid ;
    p0_direnq_dpth_thrsh_rw_pipe_nxt.qid        = dp_lsp_enq_dir_fifo_pop_data.qid ;
    p0_direnq_tok_cnt_rmw_pipe_nxt.cq           = dir_tokrtn_fifo_pop_data_cq ;
    p0_direnq_tok_lim_rw_pipe_nxt.cq            = dir_tokrtn_fifo_pop_data_cq ;
    p0_direnq_max_enq_depth_rmw_pipe_nxt.qid    = dp_lsp_enq_dir_fifo_pop_data.qid ;
  end
  p0_direnq_tot_enq_cnt_rmw_pipe_nxt.qid        = dp_lsp_enq_dir_fifo_pop_data.qid ;
  p0_direnq_tot_sch_cnt_rmw_pipe_nxt.cq         = direnq_input_arb_sch_qid.qid ;        // direct mapping of qid to cq
  //--------------------------------------------------------------------------
  p0_direnq_enq_cnt_rmw_pipe_nxt.data           = { $bits ( lsp_direnq_enq_cnt_t ) { 1'b0 } } ;         // Unused - cfg write done elsewhere
  p0_direnq_dpth_thrsh_rw_pipe_nxt.data         = { $bits ( lsp_direnq_dpth_thrsh_t ) { 1'b0 } } ;      // Unused - cfg write done elsewhere
  p0_direnq_tok_cnt_rmw_pipe_nxt.data           = { $bits ( lsp_direnq_tok_cnt_t ) { 1'b0 } } ;         // Unused - cfg write done elsewhere
  p0_direnq_tok_lim_rw_pipe_nxt.data            = { $bits ( lsp_direnq_tok_lim_t ) { 1'b0 } } ;         // Unused - cfg write done elsewhere
  p0_direnq_tot_enq_cnt_rmw_pipe_nxt.data       = { $bits ( lsp_arch_cnt_t ) { 1'b0 } } ;               // Unused - cfg write done elsewhere
  p0_direnq_tot_sch_cnt_rmw_pipe_nxt.data       = { $bits ( lsp_arch_cnt_t ) { 1'b0 } } ;               // Unused - cfg write done elsewhere
  p0_direnq_max_enq_depth_rmw_pipe_nxt.data     = { HQM_LSP_DIRENQ_ENQ_CNT_WIDTH { 1'b0 } } ;           // Unused - cfg write done elsewhere
end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq enq count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_QID )
        , .WIDTH                ( HQM_LSP_DIRENQ_ENQ_CNT_MEM_WIDTH )
) i_direnq_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_enq_cnt_rmw_pipe_status )

        // cmd input
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_direnq_enq_cnt_rmw_pipe_nxt.data )
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_direnq_ctrl_pipe_v_f )
        , .p0_rw_f              ( p0_direnq_enq_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p0_addr_f            ( p0_direnq_enq_cnt_rmw_pipe_f_pnc.qid )                // Used by blast logic
        , .p0_data_f            ( p0_direnq_enq_cnt_rmw_pipe_f_pnc.data )               // Unused

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_ctrl_pipe_v_f ) 
        , .p1_rw_f              ( p1_direnq_enq_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p1_addr_f            ( p1_direnq_enq_cnt_rmw_pipe_f_pnc.qid )                // Used by blast logic
        , .p1_data_f            ( p1_direnq_enq_cnt_rmw_pipe_f_pnc.data )               // Unused

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_ctrl_pipe_v_f ) 
        , .p2_rw_f              ( p2_direnq_enq_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_direnq_enq_cnt_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_direnq_enq_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_direnq_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_direnq_enq_cnt_upd )
        , .p3_v_f               ( p3_direnq_ctrl_pipe_v_f ) 
        , .p3_rw_f              ( p3_direnq_enq_cnt_rmw_pipe_f_nc.rw_cmd )              // Unused
        , .p3_addr_f            ( p3_direnq_enq_cnt_rmw_pipe_f_nc.qid )                 // Unused
        , .p3_data_f            ( p3_direnq_enq_cnt_rmw_pipe_f_nc.data )                // Unused


        // mem intf
        , .mem_write            ( func_dir_enq_cnt_mem_we )
        , .mem_read             ( func_dir_enq_cnt_mem_re )
        , .mem_write_addr       ( func_dir_enq_cnt_mem_waddr )
        , .mem_read_addr        ( func_dir_enq_cnt_mem_raddr )
        , .mem_write_data       ( func_dir_enq_cnt_mem_wdata )
        , .mem_read_data        ( func_dir_enq_cnt_mem_rdata )
) ;

always_comb begin
  p2_direnq_ctrl_pipe_enq_delta                 = { HQM_LSP_DIRENQ_ENQ_CNT_WIDTH { 1'b0 } } ;
  p2_direnq_ctrl_pipe_enq_delta [2:0]           = p2_direnq_ctrl_pipe_f.sch_beats ;
  p2_direnq_ctrl_pipe_sch_delta                 = { HQM_LSP_DIRENQ_TOK_CNT_WIDTH { 1'b0 } } ;
  p2_direnq_ctrl_pipe_sch_delta [2:0]           = p2_direnq_ctrl_pipe_f.sch_beats ;
  case ( p2_direnq_ctrl_pipe_f.sch_beats )
    3'h3 : p2_direnq_ctrl_pipe_sch_delta_res            = 2'h0 ;
    3'h4 : p2_direnq_ctrl_pipe_sch_delta_res            = 2'h1 ;
    default : p2_direnq_ctrl_pipe_sch_delta_res         = p2_direnq_ctrl_pipe_f.sch_beats [1:0] ;
  endcase
end // always

hqm_AW_residue_add i_direnq_enq_cnt_res_inc (
          .a                    ( 2'h1 )
        , .b                    ( p2_direnq_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_direnq_enq_cnt_res_p1 )
) ;

hqm_AW_residue_sub i_direnq_enq_cnt_res_dec (
          .a                    ( p2_direnq_ctrl_pipe_sch_delta_res )
        , .b                    ( p2_direnq_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_direnq_enq_cnt_res_mn )
) ;

assign { p2_direnq_enq_cnt_p1_carry , p2_direnq_enq_cnt_p1 }    = { 1'b0 , p2_direnq_enq_cnt_rmw_pipe_f.data.cnt } + { 1'b0 , { (HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-1) { 1'b0 } } , 1'b1 };
assign { p2_direnq_enq_cnt_mn_borrow , p2_direnq_enq_cnt_mn }   = { 1'b0 , p2_direnq_enq_cnt_rmw_pipe_f.data.cnt } - { 1'b0 , p2_direnq_ctrl_pipe_enq_delta } ;

always_comb begin
  p2_direnq_enq_cnt_oflow_cond                  = 1'b0 ;
  p2_direnq_enq_cnt_uflow_cond                  = 1'b0 ;
  if ( p2_direnq_ctrl_pipe_f.sch_v ) begin
    if ( p2_direnq_enq_cnt_mn_borrow ) begin
      p2_direnq_enq_cnt_upd                     = p2_direnq_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_direnq_enq_cnt_uflow_cond              = 1'b1 ;
    end
    else begin
      p2_direnq_enq_cnt_upd.cnt                 = p2_direnq_enq_cnt_mn ;
      p2_direnq_enq_cnt_upd.cnt_res             = p2_direnq_enq_cnt_res_mn ;
    end
  end
  else begin
    if ( p2_direnq_enq_cnt_p1_carry ) begin
      p2_direnq_enq_cnt_upd                     = p2_direnq_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_direnq_enq_cnt_oflow_cond              = 1'b1 ;
    end
    else begin
      p2_direnq_enq_cnt_upd.cnt                 = p2_direnq_enq_cnt_p1 ;
      p2_direnq_enq_cnt_upd.cnt_res             = p2_direnq_enq_cnt_res_p1 ;
    end
  end
end // always

assign p2_direnq_enq_cnt_upd_ge4        = ( p2_direnq_enq_cnt_upd.cnt >= { { { (HQM_LSP_DIRENQ_ENQ_CNT_WIDTH-3) { 1'b0 } } , 3'h4 } } ) ;

assign p2_direnq_dpth_thrsh_cm_code     = hqm_lsp_calc_thresh_code (   p2_direnq_enq_cnt_rmw_pipe_f.data.cnt
                                                                     , p2_direnq_dpth_thrsh_rw_pipe_f_pnc.data.thrsh ) ;

assign p2_direnq_enq_cnt_res_chk_en     = p2_direnq_enq_cnt_upd_v ;
assign p2_direnq_dpth_thrsh_par_chk_en  = p2_direnq_enq_cnt_res_chk_en ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_DIRENQ_ENQ_CNT_WIDTH ) ) i_direnq_enq_cnt_res_chk (
          .r                    ( p2_direnq_enq_cnt_upd.cnt_res )
        , .d                    ( p2_direnq_enq_cnt_upd.cnt )
        , .e                    ( p2_direnq_enq_cnt_res_chk_en )
        , .err                  ( p2_direnq_enq_cnt_res_err_cond )
) ;

assign p2_direnq_inp_enq_qid_par_chk_en = p2_direnq_enq_cnt_upd_v ;
assign p2_direnq_inp_tok_cq_par_chk_en  = p2_direnq_tok_cnt_upd_v ;

always_comb begin
  if ( p2_direnq_ctrl_pipe_f.sch_v ) begin
    p2_direnq_inp_enq_qid_p             = p2_direnq_ctrl_pipe_f.sch_qid_p ;
    p2_direnq_inp_tok_cq_p              = p2_direnq_ctrl_pipe_f.sch_qid_p ;
  end
  else begin
    p2_direnq_inp_enq_qid_p             = p2_direnq_ctrl_pipe_f.enq_qid_p ;
    p2_direnq_inp_tok_cq_p              = p2_direnq_ctrl_pipe_f.tok_cq_p ;
  end
end // always

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_DIR_QIDB2 ) ) i_direnq_inp_enq_qid_par_chk (
          .p                    ( p2_direnq_inp_enq_qid_p )
        , .d                    ( p2_direnq_enq_cnt_rmw_pipe_f.qid )
        , .e                    ( p2_direnq_inp_enq_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_direnq_inp_enq_qid_par_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_DIR_CQB2 ) ) i_direnq_inp_tok_cq_par_chk (
          .p                    ( p2_direnq_inp_tok_cq_p )
        , .d                    ( p2_direnq_tok_cnt_rmw_pipe_f.cq )
        , .e                    ( p2_direnq_inp_tok_cq_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_direnq_inp_tok_cq_par_err_cond )
) ;

assign p2_direnq_inp_qid_cq_par_err_cond   = p2_direnq_inp_enq_qid_par_err_cond | p2_direnq_inp_tok_cq_par_err_cond | cfg_error_inject_f [ 6 ] ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq per-qid dpth_thrsh

hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_CQ )
        , .WIDTH                ( HQM_LSP_DIRENQ_DPTH_THRSH_MEM_WIDTH )
) i_direnq_dpth_thrsh_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_dpth_thrsh_rw_pipe_status_nc )         // Unused: same as direnq_tok_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_dpth_thrsh_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_dpth_thrsh_rw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_direnq_dpth_thrsh_rw_pipe_nxt.data )
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_direnq_dpth_thrsh_rw_pipe_v_f_nc )         // Unused: same as enq_cnt_pipe
        , .p0_rw_f              ( p0_direnq_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p0_direnq_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p0_direnq_dpth_thrsh_rw_pipe_data_f_nc )

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_dpth_thrsh_rw_pipe_v_f_nc )         // Unused: same as enq_cnt_pipe
        , .p1_rw_f              ( p1_direnq_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p1_direnq_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p1_direnq_dpth_thrsh_rw_pipe_data_f_nc )

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_dpth_thrsh_rw_pipe_v_f_nc )         // Unused: same as enq_cnt_pipe
        , .p2_rw_f              ( p2_direnq_dpth_thrsh_rw_pipe_f_pnc.rw_cmd )   // Unused
        , .p2_addr_f            ( p2_direnq_dpth_thrsh_rw_pipe_f_pnc.qid )      // Unused
        , .p2_data_f            ( p2_direnq_dpth_thrsh_rw_pipe_f_pnc.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_v_f               ( p3_direnq_dpth_thrsh_rw_pipe_v_f_nc )         // Unused: same as enq_cnt_pipe
        , .p3_rw_f              ( p3_direnq_dpth_thrsh_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p3_direnq_dpth_thrsh_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p3_direnq_dpth_thrsh_rw_pipe_data_f_nc )


        // mem intf
        , .mem_write            ( func_cfg_dir_qid_dpth_thrsh_mem_we )
        , .mem_read             ( func_cfg_dir_qid_dpth_thrsh_mem_re )
        , .mem_addr             ( func_cfg_dir_qid_dpth_thrsh_mem_addr )
        , .mem_write_data       ( func_cfg_dir_qid_dpth_thrsh_mem_wdata )
        , .mem_read_data        ( func_cfg_dir_qid_dpth_thrsh_mem_rdata )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH ) ) i_direnq_dpth_thrsh_par_chk (
          .p                    ( p2_direnq_dpth_thrsh_rw_pipe_f_pnc.data.thrsh_p )
        , .d                    ( p2_direnq_dpth_thrsh_rw_pipe_f_pnc.data.thrsh )
        , .e                    ( p2_direnq_dpth_thrsh_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_direnq_dpth_thrsh_par_err_cond )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq token count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_CQ )
        , .WIDTH                ( HQM_LSP_DIRENQ_TOK_CNT_MEM_WIDTH )
) i_direnq_tok_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_tok_cnt_rmw_pipe_status_nc )                   // Unused, same as direnq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_tok_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_tok_cnt_rmw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p0_direnq_tok_cnt_rmw_pipe_nxt.data )
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_direnq_tok_cnt_rmw_pipe_v_f_nc )                   // Unused: same as enq_cnt_pipe
        , .p0_rw_f              ( p0_direnq_tok_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p0_addr_f            ( p0_direnq_tok_cnt_rmw_pipe_f_pnc.cq )                 // Used by blast logic and cq disable
        , .p0_data_f            ( p0_direnq_tok_cnt_rmw_pipe_f_pnc.data )               // Unused

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_tok_cnt_rmw_pipe_v_f_nc )                   // Unused: same as enq_cnt_pipe
        , .p1_rw_f              ( p1_direnq_tok_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p1_addr_f            ( p1_direnq_tok_cnt_rmw_pipe_f_pnc.cq )                 // Used for input error rid and blast
        , .p1_data_f            ( p1_direnq_tok_cnt_rmw_pipe_f_pnc.data )               // Unused

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_tok_cnt_rmw_pipe_v_f_nc )                   // Unused: same as enq_cnt_pipe
        , .p2_rw_f              ( p2_direnq_tok_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_direnq_tok_cnt_rmw_pipe_f.cq )
        , .p2_data_f            ( p2_direnq_tok_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_direnq_tok_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_direnq_tok_cnt_upd )
        , .p3_v_f               ( p3_direnq_tok_cnt_rmw_pipe_v_f_nc )                   // Unused: same as enq_cnt_pipe
        , .p3_rw_f              ( p3_direnq_tok_cnt_rmw_pipe_f_pnc.rw_cmd )             // Unused
        , .p3_addr_f            ( p3_direnq_tok_cnt_rmw_pipe_f_pnc.cq )                 // Used for error rid
        , .p3_data_f            ( p3_direnq_tok_cnt_rmw_pipe_f_pnc.data )               // Unused


        // mem intf
        , .mem_write            ( func_dir_tok_cnt_mem_we )
        , .mem_read             ( func_dir_tok_cnt_mem_re )
        , .mem_write_addr       ( func_dir_tok_cnt_mem_waddr )
        , .mem_read_addr        ( func_dir_tok_cnt_mem_raddr )
        , .mem_write_data       ( func_dir_tok_cnt_mem_wdata )
        , .mem_read_data        ( func_dir_tok_cnt_mem_rdata )
) ;

hqm_AW_residue_add i_direnq_tok_cnt_res_add (
          .a                    ( p2_direnq_ctrl_pipe_sch_delta_res )
        , .b                    ( p2_direnq_tok_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_direnq_tok_cnt_res_pn )
) ;

hqm_AW_residue_sub i_direnq_tok_cnt_res_sub (
          .a                    ( p2_direnq_ctrl_pipe_f.tok_delta.cnt_res )
        , .b                    ( p2_direnq_tok_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_direnq_tok_cnt_res_mn )
) ;
assign { p2_direnq_tok_cnt_pn_carry , p2_direnq_tok_cnt_pn }    = { 1'b0 , p2_direnq_tok_cnt_rmw_pipe_f.data.cnt } + { 1'b0 , p2_direnq_ctrl_pipe_sch_delta } ;
assign { p2_direnq_tok_cnt_mn_borrow , p2_direnq_tok_cnt_mn }   = { 1'b0 , p2_direnq_tok_cnt_rmw_pipe_f.data.cnt } -
                                                                  { 1'b0 , p2_direnq_ctrl_pipe_f.tok_delta.cnt } ;

always_comb begin
  p2_direnq_tok_cnt_oflow_cond                  = 1'b0 ;
  p2_direnq_tok_cnt_uflow_cond                  = 1'b0 ;
  if ( p2_direnq_ctrl_pipe_f.sch_v ) begin
    if ( p2_direnq_tok_cnt_pn_carry ) begin
      p2_direnq_tok_cnt_upd                     = p2_direnq_tok_cnt_rmw_pipe_f.data ;         // Saturate, no residue error
      p2_direnq_tok_cnt_oflow_cond              = 1'b1 ;
    end
    else begin
      p2_direnq_tok_cnt_upd.cnt                 = p2_direnq_tok_cnt_pn ;
      p2_direnq_tok_cnt_upd.cnt_res             = p2_direnq_tok_cnt_res_pn ;
    end
  end
  else begin
    if ( p2_direnq_tok_cnt_mn_borrow ) begin    // Decrement to 0, no residue error
      p2_direnq_tok_cnt_upd.cnt                 = { HQM_LSP_DIRENQ_TOK_CNT_WIDTH { 1'b0 } } ;
      p2_direnq_tok_cnt_upd.cnt_res             = 2'h0 ;
      p2_direnq_tok_cnt_uflow_cond              = 1'b1 ;
    end
    else begin
      p2_direnq_tok_cnt_upd.cnt                 = p2_direnq_tok_cnt_mn ;
      p2_direnq_tok_cnt_upd.cnt_res             = p2_direnq_tok_cnt_res_mn ;
    end
  end
end // always

always_comb begin
  case ( p2_direnq_tok_lim_rw_pipe_f_pnc.data.lim_sel )
    4'h0 : p2_direnq_tok_limit     = 11'h004 ;
    4'h1 : p2_direnq_tok_limit     = 11'h008 ;
    4'h2 : p2_direnq_tok_limit     = 11'h010 ;
    4'h3 : p2_direnq_tok_limit     = 11'h020 ;
    4'h4 : p2_direnq_tok_limit     = 11'h040 ;
    4'h5 : p2_direnq_tok_limit     = 11'h080 ;
    4'h6 : p2_direnq_tok_limit     = 11'h100 ;
    4'h7 : p2_direnq_tok_limit     = 11'h200 ;
    4'h8 : p2_direnq_tok_limit     = 11'h400 ;
    default :  p2_direnq_tok_limit = 11'h000 ;
  endcase
end // always

assign p2_direnq_tok_cnt_upd_space_sub  = { 1'b0 , p2_direnq_tok_limit } - { 1'b0 , p2_direnq_tok_cnt_upd.cnt } ;
assign p2_direnq_tok_cnt_upd_space      = ( p2_direnq_tok_cnt_upd_space_sub [HQM_LSP_DIRENQ_TOK_CNT_WIDTH] )    // borrow, should be impossible
                                            ? { HQM_LSP_DIRENQ_TOK_CNT_WIDTH { 1'b0 } }
                                            : p2_direnq_tok_cnt_upd_space_sub [HQM_LSP_DIRENQ_TOK_CNT_WIDTH-1:0] ;
assign p2_direnq_tok_cnt_upd_space_ge4  = ( p2_direnq_tok_cnt_upd_space >= { { (HQM_LSP_DIRENQ_TOK_CNT_WIDTH-3) { 1'b0 } } , 3'h4 } ) ;
assign p2_direnq_tok_cnt_upd_gt_0       = | p2_direnq_tok_cnt_upd.cnt ;


assign p0_direnq_inp_tok_cnt_res_chk_en = p0_direnq_ctrl_pipe_v_f & p1_direnq_ctrl_pipe.en & p0_direnq_ctrl_pipe_f.tok_v ;
assign p2_direnq_tok_cnt_res_chk_en     = p2_direnq_tok_cnt_upd_v ;
assign p2_direnq_tok_lim_par_chk_en     = p2_direnq_tok_cnt_res_chk_en ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_DIR_TOK_DELTA_WIDTH ) ) i_direnq_inp_tok_cnt_res_chk (
          .r                    ( p0_direnq_ctrl_pipe_f.tok_delta.cnt_res )
        , .d                    ( p0_direnq_ctrl_pipe_f.tok_delta.cnt )
        , .e                    ( p0_direnq_inp_tok_cnt_res_chk_en )
        , .err                  ( p0_direnq_inp_tok_cnt_res_err_cond )
) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_DIRENQ_TOK_CNT_WIDTH ) ) i_direnq_tok_cnt_res_chk (
          .r                    ( p2_direnq_tok_cnt_upd.cnt_res )
        , .d                    ( p2_direnq_tok_cnt_upd.cnt )
        , .e                    ( p2_direnq_tok_cnt_res_chk_en )
        , .err                  ( p2_direnq_tok_cnt_res_err_cond )
) ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_DIRENQ_TOK_LIM_SEL_WIDTH + 1 ) ) i_direnq_tok_lim_par_chk (
          .p                    ( p2_direnq_tok_lim_rw_pipe_f_pnc.data.lim_p )
        , .d                    ( {   p2_direnq_tok_lim_rw_pipe_f_pnc.data.disab_opt
                                    , p2_direnq_tok_lim_rw_pipe_f_pnc.data.lim_sel } )
        , .e                    ( p2_direnq_tok_lim_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_direnq_tok_lim_par_err_cond )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq per-cq limit
hqm_AW_rw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_CQ )
        , .WIDTH                ( HQM_LSP_DIRENQ_TOK_LIM_MEM_WIDTH )
) i_direnq_tok_lim_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_tok_lim_rw_pipe_status_nc )            // Unused: same as direnq_tok_cnt_rw_pipe_status

        // cmd input
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_tok_lim_rw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_tok_lim_rw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p0_direnq_tok_lim_rw_pipe_nxt.data )
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_f               ( p0_direnq_tok_lim_rw_pipe_v_f_nc )            // Unused: same as enq_cnt_pipe
        , .p0_rw_f              ( p0_direnq_tok_lim_rw_pipe_rw_f_nc )
        , .p0_addr_f            ( p0_direnq_tok_lim_rw_pipe_addr_f_nc )
        , .p0_data_f            ( p0_direnq_tok_lim_rw_pipe_data_f_nc )

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_tok_lim_rw_pipe_v_f_nc )            // Unused: same as enq_cnt_pipe
        , .p1_rw_f              ( p1_direnq_tok_lim_rw_pipe_rw_f_nc )
        , .p1_addr_f            ( p1_direnq_tok_lim_rw_pipe_addr_f_nc )
        , .p1_data_f            ( p1_direnq_tok_lim_rw_pipe_data_f_nc )

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_tok_lim_rw_pipe_v_f_nc )            // Unused: same as enq_cnt_pipe
        , .p2_rw_f              ( p2_direnq_tok_lim_rw_pipe_f_pnc.rw_cmd )      // Unused
        , .p2_addr_f            ( p2_direnq_tok_lim_rw_pipe_f_pnc.cq )          // Unused
        , .p2_data_f            ( p2_direnq_tok_lim_rw_pipe_f_pnc.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_v_f               ( p3_direnq_tok_lim_rw_pipe_v_f_nc )            // Unused: same as enq_cnt_pipe
        , .p3_rw_f              ( p3_direnq_tok_lim_rw_pipe_rw_f_nc )
        , .p3_addr_f            ( p3_direnq_tok_lim_rw_pipe_addr_f_nc )
        , .p3_data_f            ( p3_direnq_tok_lim_rw_pipe_data_f_nc )


        // mem intf
        , .mem_write            ( func_dir_tok_lim_mem_we )
        , .mem_read             ( func_dir_tok_lim_mem_re )
        , .mem_addr             ( func_dir_tok_lim_mem_addr )
        , .mem_write_data       ( func_dir_tok_lim_mem_wdata )
        , .mem_read_data        ( func_dir_tok_lim_mem_rdata )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq total enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_QID )
        , .WIDTH                ( HQM_LSP_ARCH_CNT_MEM_WIDTH )
) i_direnq_tot_enq_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_tot_enq_cnt_rmw_pipe_status_nc )               // Unused, same as direnq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_tot_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_tot_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_direnq_tot_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_direnq_tot_enq_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p0_rw_f              ( p0_direnq_tot_enq_cnt_rmw_pipe_rw_f_nc )      // Unused
        , .p0_addr_f            ( p0_direnq_tot_enq_cnt_rmw_pipe_addr_f_nc )    // Unused
        , .p0_data_f            ( p0_direnq_tot_enq_cnt_rmw_pipe_data_f_nc )    // Unused

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_tot_enq_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p1_rw_f              ( p1_direnq_tot_enq_cnt_rmw_pipe_rw_f_nc )      // Unused
        , .p1_addr_f            ( p1_direnq_tot_enq_cnt_rmw_pipe_addr_f_nc )    // Unused
        , .p1_data_f            ( p1_direnq_tot_enq_cnt_rmw_pipe_data_f_nc )    // Unused

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_tot_enq_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p2_rw_f              ( p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd ) // Used to determine upd_v
        , .p2_addr_f            ( p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.qid )    // Unused
        , .p2_data_f            ( p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_direnq_tot_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_direnq_tot_enq_cnt_upd )
        , .p3_v_f               ( p3_direnq_tot_enq_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p3_rw_f              ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd ) // Used for res_chk_en
        , .p3_addr_f            ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.qid )    // Unused
        , .p3_data_f            ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data )   // Used for res_chk

        // mem intf
        , .mem_write            ( cfgsc_func_qid_dir_tot_enq_cnt_mem_we )
        , .mem_read             ( func_qid_dir_tot_enq_cnt_mem_re )
        , .mem_write_addr       ( cfgsc_func_qid_dir_tot_enq_cnt_mem_waddr )
        , .mem_read_addr        ( func_qid_dir_tot_enq_cnt_mem_raddr )
        , .mem_write_data       ( cfgsc_func_qid_dir_tot_enq_cnt_mem_wdata )
        , .mem_read_data        ( func_qid_dir_tot_enq_cnt_mem_rdata )
) ;

hqm_AW_residue_add i_direnq_tot_enq_cnt_res_add (
          .a                    ( 2'h1 )
        , .b                    ( p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .r                    ( p2_direnq_tot_enq_cnt_res_p1 )
) ;

assign p2_direnq_tot_enq_cnt_p1                 = p2_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt + 64'h1 ;               // wrap

assign p2_direnq_tot_enq_cnt_upd.cnt            = p2_direnq_tot_enq_cnt_p1 ;
assign p2_direnq_tot_enq_cnt_upd.cnt_res        = p2_direnq_tot_enq_cnt_res_p1 ;

assign p3_direnq_tot_enq_cnt_res_chk_en         = p4_direnq_ctrl_pipe_en & ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ARCH_CNT_WIDTH ) ) i_direnq_tot_enq_cnt_res_chk (
          .r                    ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .d                    ( p3_direnq_tot_enq_cnt_rmw_pipe_f_pnc.data.cnt )
        , .e                    ( p3_direnq_tot_enq_cnt_res_chk_en )
        , .err                  ( p4_direnq_tot_enq_cnt_res_err_nxt )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq total schedule count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_CQ )
        , .WIDTH                ( HQM_LSP_ARCH_CNT_MEM_WIDTH )
) i_direnq_tot_sch_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_tot_sch_cnt_rmw_pipe_status_nc )               // Unused, direnq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_tot_sch_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_tot_sch_cnt_rmw_pipe_nxt.cq )
        , .p0_write_data_nxt    ( p0_direnq_tot_sch_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_direnq_tot_sch_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p0_rw_f              ( p0_direnq_tot_sch_cnt_rmw_pipe_rw_f_nc )      // Unused
        , .p0_addr_f            ( p0_direnq_tot_sch_cnt_rmw_pipe_addr_f_nc )    // Unused
        , .p0_data_f            ( p0_direnq_tot_sch_cnt_rmw_pipe_data_f_nc )    // Unused

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_tot_sch_cnt_rmw_pipe_v_f_nc )       // Unused
        , .p1_rw_f              ( p1_direnq_tot_sch_cnt_rmw_pipe_rw_f_nc )      // Unused
        , .p1_addr_f            ( p1_direnq_tot_sch_cnt_rmw_pipe_addr_f_nc )    // Unused
        , .p1_data_f            ( p1_direnq_tot_sch_cnt_rmw_pipe_data_f_nc )    // Unused

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_tot_sch_cnt_rmw_pipe_v_f_nc )
        , .p2_rw_f              ( p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd ) // Used to determine upd_v
        , .p2_addr_f            ( p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.cq )     // Unused
        , .p2_data_f            ( p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_direnq_tot_sch_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_direnq_tot_sch_cnt_upd )
        , .p3_v_f               ( p3_direnq_tot_sch_cnt_rmw_pipe_v_f_nc )
        , .p3_rw_f              ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd ) // Used for res_chk_en
        , .p3_addr_f            ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.cq )     // Unused
        , .p3_data_f            ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data )   // Used for res_chk

        // mem intf
        , .mem_write            ( cfgsc_func_cq_dir_tot_sch_cnt_mem_we )
        , .mem_read             ( func_cq_dir_tot_sch_cnt_mem_re )
        , .mem_write_addr       ( cfgsc_func_cq_dir_tot_sch_cnt_mem_waddr )
        , .mem_read_addr        ( func_cq_dir_tot_sch_cnt_mem_raddr )
        , .mem_write_data       ( cfgsc_func_cq_dir_tot_sch_cnt_mem_wdata )
        , .mem_read_data        ( func_cq_dir_tot_sch_cnt_mem_rdata )
    ) ;

hqm_AW_residue_add i_direnq_tot_sch_cnt_res_add (
          .a                    ( p2_direnq_ctrl_pipe_sch_delta_res )
        , .b                    ( p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .r                    ( p2_direnq_tot_sch_cnt_res_pn )
) ;

assign p2_direnq_tot_sch_cnt_pn                 = p2_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt + { { ( 64 - HQM_LSP_DIRENQ_TOK_CNT_WIDTH ) { 1'b0 } } , p2_direnq_ctrl_pipe_sch_delta } ;      // wrap

assign p2_direnq_tot_sch_cnt_upd.cnt            = p2_direnq_tot_sch_cnt_pn ;
assign p2_direnq_tot_sch_cnt_upd.cnt_res        = p2_direnq_tot_sch_cnt_res_pn ;

assign p3_direnq_tot_sch_cnt_res_chk_en         = p4_direnq_ctrl_pipe_en & ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.rw_cmd == HQM_AW_RMWPIPE_RMW ) ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_ARCH_CNT_WIDTH ) ) i_direnq_tot_sch_cnt_res_chk (
          .r                    ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt_res )
        , .d                    ( p3_direnq_tot_sch_cnt_rmw_pipe_f_pnc.data.cnt )
        , .e                    ( p3_direnq_tot_sch_cnt_res_chk_en )
        , .err                  ( p4_direnq_tot_sch_cnt_res_err_nxt )
) ;

//-------------------------------------------------------------------------------------------------
// Manage storage for direnq total enqueue count
hqm_AW_rmw_mem_4pipe_waddr #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_DIR_QID )
        , .WIDTH                ( HQM_LSP_DIRENQ_ENQ_CNT_WIDTH )
) i_direnq_max_enq_depth_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( direnq_max_enq_depth_rmw_pipe_status_nc )     // Unused, direnq_enq_cnt_rmw_pipe_status

        // cmd input
        , .p0_hold              ( p0_direnq_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_direnq_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_direnq_max_enq_depth_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_direnq_max_enq_depth_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_direnq_max_enq_depth_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_direnq_max_enq_depth_rmw_pipe_v_f_nc )     // Unused
        , .p0_rw_f              ( p0_direnq_max_enq_depth_rmw_pipe_rw_f_nc )    // Unused
        , .p0_addr_f            ( p0_direnq_max_enq_depth_rmw_pipe_addr_f_nc )  // Unused
        , .p0_data_f            ( p0_direnq_max_enq_depth_rmw_pipe_data_f_nc )  // Unused

        , .p1_hold              ( p1_direnq_ctrl_pipe.hold )
        , .p1_v_f               ( p1_direnq_max_enq_depth_rmw_pipe_v_f_nc )     // Unused
        , .p1_rw_f              ( p1_direnq_max_enq_depth_rmw_pipe_rw_f_nc )    // Unused
        , .p1_addr_f            ( p1_direnq_max_enq_depth_rmw_pipe_addr_f_nc )  // Unused
        , .p1_data_f            ( p1_direnq_max_enq_depth_rmw_pipe_data_f_nc )  // Unused

        , .p2_hold              ( p2_direnq_ctrl_pipe.hold )
        , .p2_v_f               ( p2_direnq_max_enq_depth_rmw_pipe_v_f_nc )
        , .p2_rw_f              ( p2_direnq_max_enq_depth_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_direnq_max_enq_depth_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_direnq_max_enq_depth_rmw_pipe_f.data )

        , .p3_hold              ( p3_direnq_ctrl_pipe.hold )
        , .p3_bypdata_sel_nxt   ( p2_direnq_max_enq_depth_upd_v )
        , .p3_bypdata_nxt       ( p2_direnq_max_enq_depth_upd )
        , .p3_bypaddr_sel_nxt   ( p2_direnq_max_enq_depth_upd_v )
        , .p3_bypaddr_nxt       ( p2_direnq_max_enq_depth_rmw_pipe_f.qid )
        , .p3_v_f               ( p3_direnq_max_enq_depth_rmw_pipe_v_f_nc )
        , .p3_rw_f              ( p3_direnq_max_enq_depth_rmw_pipe_f_nc.rw_cmd )        // Unused
        , .p3_addr_f            ( p3_direnq_max_enq_depth_rmw_pipe_f_nc.qid )           // Unused
        , .p3_data_f            ( p3_direnq_max_enq_depth_rmw_pipe_f_nc.data )          // Unused

        // mem intf
        , .mem_write            ( func_qid_dir_max_depth_mem_we )
        , .mem_read             ( func_qid_dir_max_depth_mem_re )
        , .mem_write_addr       ( func_qid_dir_max_depth_mem_waddr )
        , .mem_read_addr        ( func_qid_dir_max_depth_mem_raddr )
        , .mem_write_data       ( func_qid_dir_max_depth_mem_wdata )
        , .mem_read_data        ( func_qid_dir_max_depth_mem_rdata )
) ;

assign p2_direnq_enq_cnt_gt_max_depth           = ( p2_direnq_enq_cnt_upd.cnt > p2_direnq_max_enq_depth_rmw_pipe_f.data ) ;
assign p2_direnq_max_enq_depth_upd              = p2_direnq_enq_cnt_upd.cnt ;

//-------------------------------------------------------------------------------------------------
// Underflow/overflow errors - some are impossible, some may be caused by software/config errors
//

always_comb begin
  // Don't hold - 1-clock pulse to report
  p3_direnq_enq_cnt_uflow_err_nxt       = 1'b0 ;
  p3_direnq_enq_cnt_oflow_err_nxt       = 1'b0 ;
  p3_direnq_tok_cnt_uflow_err_nxt       = 1'b0 ;
  p3_direnq_tok_cnt_oflow_err_nxt       = 1'b0 ;

  p1_direnq_inp_tok_cnt_res_err_nxt     = 1'b0 ;
  p3_direnq_enq_cnt_res_err_nxt         = 1'b0 ;
  p3_direnq_dpth_thrsh_par_err_nxt      = 1'b0 ;
  p3_direnq_tok_cnt_res_err_nxt         = 1'b0 ;
  p3_direnq_tok_lim_par_err_nxt         = 1'b0 ;
  p3_direnq_inp_qid_cq_par_err_nxt      = 1'b0 ;

  if ( p0_direnq_ctrl_pipe_v_f & ~ p1_direnq_ctrl_pipe.hold ) begin
    p1_direnq_inp_tok_cnt_res_err_nxt   = p0_direnq_inp_tok_cnt_res_err_cond & ~ p0_direnq_inp_tok_cq_disable ;
  end

  if ( p2_direnq_ctrl_pipe_v_f & ~ p3_direnq_ctrl_pipe.hold ) begin
    p3_direnq_enq_cnt_uflow_err_nxt     = p2_direnq_ctrl_pipe_f.sch_v & p2_direnq_enq_cnt_uflow_cond & ~ p2_direnq_enq_cnt_cq_disable ;
    p3_direnq_enq_cnt_oflow_err_nxt     = p2_direnq_ctrl_pipe_f.enq_v & p2_direnq_enq_cnt_oflow_cond & ~ p2_direnq_enq_cnt_cq_disable ;
    p3_direnq_tok_cnt_uflow_err_nxt     = p2_direnq_ctrl_pipe_f.tok_v & ( p2_direnq_tok_cnt_uflow_cond | cfg_error_inject_f [ 16 ] ) & ~ p2_direnq_tok_cnt_cq_disable ;
    p3_direnq_tok_cnt_oflow_err_nxt     = p2_direnq_ctrl_pipe_f.sch_v & p2_direnq_tok_cnt_oflow_cond & ~ p2_direnq_tok_cnt_cq_disable ;

    p3_direnq_enq_cnt_res_err_nxt       = p2_direnq_enq_cnt_res_err_cond & ~ p2_direnq_enq_cnt_cq_disable ;
    p3_direnq_dpth_thrsh_par_err_nxt    = p2_direnq_dpth_thrsh_par_err_cond & ~ p2_direnq_enq_cnt_cq_disable ;
    p3_direnq_tok_cnt_res_err_nxt       = p2_direnq_tok_cnt_res_err_cond & ~ p2_direnq_tok_cnt_cq_disable ;
    p3_direnq_tok_lim_par_err_nxt       = ( p2_direnq_tok_lim_par_err_cond | cfg_error_inject_f [ 3 ] ) & ~ p2_direnq_tok_cnt_cq_disable ;
    p3_direnq_inp_qid_cq_par_err_nxt    = p2_direnq_inp_qid_cq_par_err_cond ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_direnq_enq_cnt_uflow_err_f       <= 1'b0 ;
    p3_direnq_enq_cnt_oflow_err_f       <= 1'b0 ;
    p3_direnq_tok_cnt_uflow_err_f       <= 1'b0 ;
    p3_direnq_tok_cnt_oflow_err_f       <= 1'b0 ;

    p1_direnq_inp_tok_cnt_res_err_f     <= 1'b0 ;
    p3_direnq_enq_cnt_res_err_f         <= 1'b0 ;
    p3_direnq_dpth_thrsh_par_err_f      <= 1'b0 ;
    p3_direnq_tok_cnt_res_err_f         <= 1'b0 ;
    p3_direnq_tok_lim_par_err_f         <= 1'b0 ;
    p3_direnq_inp_qid_cq_par_err_f      <= 1'b0 ;

    p4_direnq_tot_enq_cnt_res_err_f     <= 1'b0 ;
    p4_direnq_tot_sch_cnt_res_err_f     <= 1'b0 ;
  end
  else begin
    p3_direnq_enq_cnt_uflow_err_f       <= p3_direnq_enq_cnt_uflow_err_nxt ;
    p3_direnq_enq_cnt_oflow_err_f       <= p3_direnq_enq_cnt_oflow_err_nxt ;
    p3_direnq_tok_cnt_uflow_err_f       <= p3_direnq_tok_cnt_uflow_err_nxt ;
    p3_direnq_tok_cnt_oflow_err_f       <= p3_direnq_tok_cnt_oflow_err_nxt ;

    p1_direnq_inp_tok_cnt_res_err_f     <= p1_direnq_inp_tok_cnt_res_err_nxt ;
    p3_direnq_enq_cnt_res_err_f         <= p3_direnq_enq_cnt_res_err_nxt ;
    p3_direnq_dpth_thrsh_par_err_f      <= p3_direnq_dpth_thrsh_par_err_nxt ;
    p3_direnq_tok_cnt_res_err_f         <= p3_direnq_tok_cnt_res_err_nxt ;
    p3_direnq_tok_lim_par_err_f         <= p3_direnq_tok_lim_par_err_nxt ;
    p3_direnq_inp_qid_cq_par_err_f      <= p3_direnq_inp_qid_cq_par_err_nxt ;

    p4_direnq_tot_enq_cnt_res_err_f     <= p4_direnq_tot_enq_cnt_res_err_nxt ;
    p4_direnq_tot_sch_cnt_res_err_f     <= p4_direnq_tot_sch_cnt_res_err_nxt ;
  end
end // always

assign p3_direnq_tok_cnt_uflow_err_rid  = { 1'b0 , p3_direnq_tok_cnt_rmw_pipe_f_pnc.cq } ;              // is_ldb, cq[6:0]

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: DIRENQ status bits, arbiter and output buffering
//-----------------------------------------------------------------------------------------------------
// In general, for all of the non-load-balanced pipes, when the arbiter determines that there is a schedule
// ready to go, it is only allowed to go if the destination(s) are ready to accept it.
// - all schedules go to the output FIFO, so the output FIFO afull must = 0
// - If the schedule request goes through a FIFO/DB/register level before feeding into the input arbiter,
//   that FIFO/DB/register must be available.  If the request feeds directly into the input arbiter, the
//   schedule is only allowed to go if it wins the arbitration.  Currently the requests all feed back
//   into a staging register.
// If the schedule is allowed to go, several actions must be taken:
// - a request must go through the input arbiter in order to update the counts via the RMW pipe(s)
// - the p3 status bits must be updated to temporarily prevent a schedule from being (possibly incorrectly)
//   initiated on the subsequent clock(s), until the correct count update occurs.
// - the upper pipeline stages must have any pending updates for this same qid "blasted", meaning that
//   they must not be allowed to update the p3 status bits once they reach p3 (they must still update the
//   the regfile count(s).
// - the output FIFO must be pushed to actually cause the schedule to occur
//
// In the case of the ATQ and two RPL pipelines, one schedule arbitration causes each of these actions to
// occur once.  In the case of the DIRENQ pipeline, one scheduled arbitration causes 1 to 4 pushes to the
// output FIFO on consecutive clocks (when there is space) but only a single occurence of the other three.
// The signal naming for each of these events is consistent across all 4 non-lb pipes:
// - <pipe>_sch_req - arbiter determines sch ready to go and destination(s) can accept it.  In the case
//   where there is no FIFO/DB/register for this update request, the sch still might not be allowed to go
//   if the input arbiter does not select it
// - <pipe>_input_arb_reqs[i] - sch request to the input arbiter (to get into p0)
// - <pipe>_input_arb_sch - input arbiter picks sch as winner and it is not held up by pipeline
// - <pipe>_sch_start - sch request meets all requirements and may be initiated.  In the case of DIRENQ fill
//   sequences, this is just the first of the 1..4 clocks.
// - <pipe_sch_out> - sch request is generating an output schedule.  Except for DIRENQ schedules, this
//   is the same as <pipe>_sch_start.  For DIRENQ schedules, this is asserted for all 1..4 output clocks.
// e.g.:
// p3_direnq_sch_req
// direnq_input_arb_reqs[1]
// direnq_input_arb_sch
// p3_direnq_sch_start
// p3_direnq_sch_out

//-------------------------------------------------------------------------------------------------
function automatic [1:0] hqm_lsp_dir_rem_beats ;
// Calculate max number of beats to perform after the current one, based on the availabilty of
// data, CQ space, and space on the current cache line (max 4 beats per line).
  input logic [2:0] qid_v ;     // 0..4
  input logic [2:0] cq_avail ;  // 0..4
  input logic [1:0] wp ;        // 0..3
  logic [2:0] num_beats ;       // Number of beats including this one, not accounting for wp (1..4)
  logic [1:0] rem_beats ;       // 0..3
  begin
    if ( ( qid_v == 3'h4 ) & ( cq_avail == 3'h4 ) )
      num_beats = 3'h4 ;
    else if ( ( qid_v >= 3'h3 ) & ( cq_avail >= 3'h3 ) )
      num_beats = 3'h3 ;
    else if ( ( qid_v >= 3'h2 ) & ( cq_avail >= 3'h2 ) )
      num_beats = 3'h2 ;
    else
      num_beats = 3'h1 ;

    if ( ( num_beats == 3'h4 ) & ( wp == 2'h0 ) )
      rem_beats = 2'h3 ;
    else if ( ( num_beats >= 3'h3 ) & ( wp <= 2'h1 ) )
      rem_beats = 2'h2 ;
    else if ( ( num_beats >= 3'h2 ) & ( wp <= 2'h2 ) )
      rem_beats = 2'h1 ;
    else
      rem_beats = 2'h0 ;
  end
  return rem_beats ;
endfunction // hqm_lsp_dir_rem_beats

//-------------------------------------------------------------------------------------------------

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
    // Bypass update from sch takes precedence over update from p2; sch update will cause subsequent write
    // of latest/correct value of counts caused by this scheduling.  If entering a fill sequence, do the full inc/dec by 4
    // on the first clock, set fill_count to force the subsequent 3 writes for the same qid/cq, do not update status on
    // final 3 clocks.
    // Do not let enq or tok writes which have been blasted update the arbiter status vector; the subsequent sch update which caused
    // the blast will update with the correct status when it reaches p2.
 
    p3_direnq_sch_hit[i]                        = p3_direnq_sch_start & ( p3_direnq_sch_start_qid == i ) ;

    p3_direnq_p2_enq_hit[i]                     = p3_direnq_ctrl_pipe.en & ( p2_direnq_ctrl_pipe_f.enq_v | p2_direnq_ctrl_pipe_f.sch_v ) &
                                                  ( p2_direnq_enq_cnt_rmw_pipe_f.qid == i ) & ~ p2_direnq_ctrl_pipe_f.blast_enq ;

    p3_direnq_p2_tok_hit[i]                     = p3_direnq_ctrl_pipe.en & ( p2_direnq_ctrl_pipe_f.tok_v | p2_direnq_ctrl_pipe_f.sch_v ) &
                                                  ( p2_direnq_tok_cnt_rmw_pipe_f.cq == i )  & ~ p2_direnq_ctrl_pipe_f.blast_tok ;

    // Any output to this CQ.  Update must be correct before sch gets back down to p2 and re-enables scheduling.
    // Do on clock after schedule start for delay reasons, on clock where calc is done.
    p3_direnq_wp_en [i]                         = p4_direnq_sch_first_clock_f & ( p4_direnq_sch_qid_f.qid[HQM_NUM_DIR_QIDB2-1:0] == i ) ;
  end // for
end // always

// For each Directed qid and its corresponding cq, maintain state required for each arbiter.
// Update (potentially set) when enq count or token count is updated, reset when that qid/cq is selected to be scheduled.
always_comb begin
  p3_direnq_arb_stat_nxt                        = p3_direnq_arb_stat_f ;
  p3_direnq_tok_cnt_v_nxt                       = p3_direnq_tok_cnt_v_f ;
  if ( p3_direnq_sch_start | p3_direnq_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
      // Should be cleared to 0 on a successful vas reset drain
      if ( p3_direnq_sch_hit [i] ) begin
        p3_direnq_arb_stat_nxt[i].qid_v         = 3'h0 ;
      end
      else if ( p3_direnq_p2_enq_hit[i] ) begin
        if ( p2_direnq_enq_cnt_upd_ge4 ) begin
          p3_direnq_arb_stat_nxt[i].qid_v       = 3'h4 ;
        end
        else begin
          p3_direnq_arb_stat_nxt[i].qid_v       = { 1'b0 , p2_direnq_enq_cnt_upd.cnt [1:0] } ;
        end
      end
    end // for i
  end // if
  if ( cfgsc_dir_tok_cnt_mem_we | p3_direnq_sch_start | p3_direnq_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_CQ ; i = i + 1 ) begin
      if ( cfgsc_dir_tok_cnt_mem_we & ( cfg_mem_addr [HQM_NUM_DIR_CQB2-1:0] == i ) ) begin      // Should only be done as part of vas reset
        p3_direnq_arb_stat_nxt[i].cq_avail      = 3'h1 ;                        // Don't yet know actual configured depth, just enable it
        p3_direnq_tok_cnt_v_nxt [i]             = 1'b0 ;
      end
      else if ( p3_direnq_sch_hit [i] ) begin
        p3_direnq_arb_stat_nxt[i].cq_avail      = 3'h0 ;
        p3_direnq_tok_cnt_v_nxt [i]             = 1'b1 ;
      end
      else if ( p3_direnq_p2_tok_hit [i] ) begin
        if ( p2_direnq_tok_cnt_upd_space_ge4 ) begin
          p3_direnq_arb_stat_nxt[i].cq_avail    = 3'h4 ;
        end
        else begin
          p3_direnq_arb_stat_nxt[i].cq_avail    = { 1'b0 , p2_direnq_tok_cnt_upd_space [1:0] } ;
        end
        p3_direnq_tok_cnt_v_nxt [i]             = p2_direnq_tok_cnt_upd_gt_0 ;
      end
    end // for i
  end // if

  // Update latest enq count vs. cfg threshold status
  p3_direnq_cm_code_nxt                         = p3_direnq_cm_code_f ;
  if ( cfgsc_dir_tok_cnt_mem_we | cfgsc_cfg_dir_qid_dpth_thrsh_mem_we | p3_direnq_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
      if ( cfgsc_dir_tok_cnt_mem_we & ( cfg_mem_addr [HQM_NUM_DIR_QIDB2-1:0] == i ) ) begin     // DIR CQ = QID so ok.  Should only be done as part of vas reset
        p3_direnq_cm_code_nxt [i]               = 2'h0 ;
      end
      else if ( cfgsc_cfg_dir_qid_dpth_thrsh_mem_we & ( cfg_mem_addr [HQM_NUM_DIR_QIDB2-1:0] == i ) ) begin
        p3_direnq_cm_code_nxt [i]               = 2'h0 ;
      end
      else if ( p3_direnq_p2_enq_hit[i] ) begin         // enq or re-inserted sch, same conditions which functionally update the enq_cnt
        p3_direnq_cm_code_nxt [i]               = p2_direnq_dpth_thrsh_cm_code ;
      end
    end // for i
  end // if

  // Increment wp for cq being scheduled
  p3_direnq_wp_nxt                              = p3_direnq_wp_f ;
  if ( cfgsc_dir_tok_cnt_mem_we | p4_direnq_sch_first_clock_f ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_CQ ; i = i + 1 ) begin
      if ( cfgsc_dir_tok_cnt_mem_we & ( cfg_mem_addr [HQM_NUM_DIR_CQB2-1:0] == i ) ) begin                      // Should only be done as part of vas reset
        p3_direnq_wp_nxt [i]                    = 2'h0 ;
      end
      else if ( p3_direnq_wp_en [i] ) begin
        p3_direnq_wp_nxt [i]                    = p4_direnq_sch_wp_f + p4_direnq_calc_rem_beats + 2'h1 ;        // mod 4
      end
    end // for i
  end // if

  cfg_dir_tok_lim_disab_opt_nxt                    = cfg_dir_tok_lim_disab_opt_f ;
  if ( cfgsc_dir_tok_lim_mem_we ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_CQ ; i = i + 1 ) begin
      if ( cfgsc_dir_tok_lim_mem_we & ( cfg_mem_addr [HQM_NUM_DIR_CQB2-1:0] == i ) ) begin
        cfg_dir_tok_lim_disab_opt_nxt [i]          = cfgsc_dir_tok_lim_mem_wdata_struct.disab_opt ;
      end
    end // for
  end // if
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
      p3_direnq_arb_stat_f[i].cq_avail          <= 3'h1 ;
      p3_direnq_arb_stat_f[i].qid_v             <= 3'h0 ;
      p3_direnq_cm_code_f [i]                   <= 2'h0 ;
      p3_direnq_wp_f[i]                         <= 2'h0 ;
    end
    p3_direnq_tok_cnt_v_f                       <= { HQM_NUM_DIR_CQ { 1'b0 } } ;
  end
  else begin
    for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
      p3_direnq_arb_stat_f[i]                   <= p3_direnq_arb_stat_nxt[i] ;
      p3_direnq_cm_code_f [i]                   <= p3_direnq_cm_code_nxt [i] ;
      p3_direnq_wp_f[i]                         <= p3_direnq_wp_nxt[i] ;
    end // for i
    p3_direnq_tok_cnt_v_f                       <= p3_direnq_tok_cnt_v_nxt ;
  end // else rst_n
end // always

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_DIR_QID ; i = i + 1 ) begin
    p3_qid_dir_sch_v_status [i]         = ( | p3_direnq_arb_stat_f[i].qid_v ) ;
    p3_cq_dir_tok_v_status [i]          = ( | p3_direnq_arb_stat_f[i].cq_avail ) ;      // num DIR cq will always = num DIR qid so OK in this loop
  end // for i
end // always
assign p3_direnq_arb_reqs               = p3_qid_dir_sch_v_status & p3_cq_dir_tok_v_status & ( ~ cfg_cq_dir_disable_f ) ;

hqm_AW_rr_arb # ( .NUM_REQS ( HQM_NUM_DIR_QID ) ) i_direnq_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p3_direnq_arb_reqs )
        , .update               ( p3_direnq_arb_update )
        , .winner_v             ( p3_direnq_arb_winner_pre_v )
        , .winner               ( p3_direnq_arb_winner )
) ;


assign p3_direnq_arb_winner_v   = p3_direnq_arb_winner_pre_v & ~ cause_pipe_idle ;

always_comb begin
  p3_direnq_arb_winner_qid.qid                          = { HQM_LSP_ARCH_NUM_DIR_QIDB2 { 1'b0 } } ;
  p3_direnq_arb_winner_qid.qid [HQM_NUM_DIR_QIDB2-1:0]  = p3_direnq_arb_winner ;
end // always

hqm_AW_parity_gen #( .WIDTH ( HQM_LSP_ARCH_NUM_DIR_QIDB2 ) ) i_direnq_arb_winner_qid_par_gen (
          .d            ( p3_direnq_arb_winner_qid.qid )
        , .odd          ( 1'b1 )
        , .p            ( p3_direnq_arb_winner_qid.qid_p )
) ;

assign p3_direnq_sch_req                = p3_direnq_arb_winner_v & ~ p3_direnq_fill_in_progress & ~ dir_sel_dp_fifo_hold & ~ p4_direnq_sch_hold ;
assign p3_direnq_sch_req_qid            = p3_direnq_arb_winner_qid.qid ;

// Timing might be tight, 64:1 arbiter -> 64:1 mux
assign p3_direnq_arb_winner_qid_v       = p3_direnq_arb_stat_f[ p3_direnq_arb_winner ].qid_v ;
assign p3_direnq_arb_winner_cq_avail    = p3_direnq_arb_stat_f[ p3_direnq_arb_winner ].cq_avail ;
assign p3_direnq_arb_winner_cm_code     = p3_direnq_cm_code_f[ p3_direnq_arb_winner ] ;
assign p3_direnq_arb_winner_wp          = p3_direnq_wp_f[ p3_direnq_arb_winner ] ;
assign p3_direnq_arb_winner_disab_opt   = cfg_dir_tok_lim_disab_opt_f [ p3_direnq_arb_winner ] ;

assign p4_direnq_calc_rem_beats_enab    = hqm_lsp_dir_rem_beats ( p4_direnq_sch_qid_v_f , p4_direnq_sch_cq_avail_f , p4_direnq_sch_wp_f ) ;
assign p4_direnq_calc_rem_beats         = ( p4_direnq_sch_disab_opt_f ) ? 2'h0 : p4_direnq_calc_rem_beats_enab ;
assign p3_direnq_rem_beats              = ( p4_direnq_sch_first_beat_f ) ? p4_direnq_calc_rem_beats : p4_direnq_sch_rem_beats_f ;
assign p3_direnq_fill_in_progress       = | p3_direnq_rem_beats ;
assign p3_direnq_rem_beats_m1           = ( p3_direnq_rem_beats - 2'h1 ) ;              // In "underflow" case will be ignored, fill not in progress
assign p4_direnq_sch_rem_beats_m1       = ( p4_direnq_sch_rem_beats_f - 2'h1 ) ;        // In "underflow" case will be ignored, fill not in progress

assign p3_direnq_sch_start              = p3_direnq_sch_req ;
assign p3_direnq_sch_start_qid          = p3_direnq_sch_req_qid ;
assign p3_direnq_arb_update             = p3_direnq_sch_start ;

always_comb begin
  if ( p3_direnq_fill_in_progress ) begin       // Use the saved qid during fill sequence, sched whenever no bp - no p4 hold consideration
    p3_direnq_sch_out_qid               = p4_direnq_sch_qid_f.qid [HQM_NUM_DIR_QIDB2-1:0] ;
    p3_direnq_sch_out_cm_code           = p4_direnq_sch_cm_code_f ;
    p3_direnq_sch_out                   = ~ dir_sel_dp_fifo_hold ;
  end
  else begin
    p3_direnq_sch_out_qid               = p3_direnq_arb_winner_qid.qid [HQM_NUM_DIR_QIDB2-1:0] ;
    p3_direnq_sch_out_cm_code           = p3_direnq_arb_winner_cm_code ;
    p3_direnq_sch_out                   = p3_direnq_sch_start & ~ dir_sel_dp_fifo_hold ;
  end

  p4_direnq_sch_rem_beats_nxt           = p4_direnq_sch_rem_beats_f ;
  p4_direnq_sch_qid_v_nxt               = p4_direnq_sch_qid_v_f ;
  p4_direnq_sch_cq_avail_nxt            = p4_direnq_sch_cq_avail_f ;
  p4_direnq_sch_wp_nxt                  = p4_direnq_sch_wp_f ;
  p4_direnq_sch_qid_nxt                 = p4_direnq_sch_qid_f ;
  p4_direnq_sch_cm_code_nxt             = p4_direnq_sch_cm_code_f ;
  p4_direnq_sch_disab_opt_nxt           = p4_direnq_sch_disab_opt_f ;
  p4_direnq_sch_first_beat_nxt          = p4_direnq_sch_first_beat_f ;
  p4_direnq_sch_first_clock_nxt         = p4_direnq_sch_first_clock_f ;

  if ( p3_direnq_sch_start ) begin      // Capture new winner and all related info
    p4_direnq_sch_rem_beats_nxt         = 2'h0 ;                // Should be a don't care since calculated on the fly for first beat, but clean it up
    p4_direnq_sch_qid_v_nxt             = p3_direnq_arb_winner_qid_v ;
    p4_direnq_sch_cq_avail_nxt          = p3_direnq_arb_winner_cq_avail ;
    p4_direnq_sch_wp_nxt                = p3_direnq_arb_winner_wp ;
    p4_direnq_sch_qid_nxt               = p3_direnq_arb_winner_qid ;
    p4_direnq_sch_disab_opt_nxt         = p3_direnq_arb_winner_disab_opt ;
    p4_direnq_sch_cm_code_nxt           = p3_direnq_arb_winner_cm_code ;
    p4_direnq_sch_first_beat_nxt        = 1'b1 ;
    p4_direnq_sch_first_clock_nxt       = 1'b1 ;
  end
  else begin
    if ( p3_direnq_sch_out & p3_direnq_fill_in_progress ) begin
      p4_direnq_sch_first_beat_nxt      = 1'b0 ;
      if ( p4_direnq_sch_first_beat_f ) begin
        p4_direnq_sch_rem_beats_nxt     = p3_direnq_rem_beats_m1 ;      // Save the on-the-fly calculated value for the next iter (if any)
      end
      else begin
        p4_direnq_sch_rem_beats_nxt     = p4_direnq_sch_rem_beats_m1 ;  // Underflow wrap OK, in that case fill will be done
      end
    end
    p4_direnq_sch_first_clock_nxt       = 1'b0 ;                        // No hold; just update p3 wp on first clock of sched
  end
end // always

assign p4_direnq_sch_hold               = p4_direnq_sch_v_f & ~ direnq_input_arb_sch ;
assign p4_direnq_sch_v_nxt              = p3_direnq_sch_req | p4_direnq_sch_hold ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p4_direnq_sch_v_f                   <= 1'b0 ;
    p4_direnq_sch_qid_f.qid_p           <= 1'b1 ;
    p4_direnq_sch_qid_f.qid             <= { HQM_LSP_ARCH_NUM_DIR_QIDB2 { 1'b0 } } ;
    p4_direnq_sch_cm_code_f             <= 2'h0 ;
    p4_direnq_sch_rem_beats_f           <= 2'h0 ;
    p4_direnq_sch_qid_v_f               <= 3'h0 ;
    p4_direnq_sch_cq_avail_f            <= 3'h0 ;
    p4_direnq_sch_wp_f                  <= 2'h0 ;
    p4_direnq_sch_disab_opt_f           <= 1'b0 ;
    p4_direnq_sch_first_beat_f          <= 1'b0 ;
    p4_direnq_sch_first_clock_f         <= 1'b0 ;
  end
  else begin
    p4_direnq_sch_v_f                   <= p4_direnq_sch_v_nxt ;
    p4_direnq_sch_qid_f                 <= p4_direnq_sch_qid_nxt ;
    p4_direnq_sch_cm_code_f             <= p4_direnq_sch_cm_code_nxt ;
    p4_direnq_sch_rem_beats_f           <= p4_direnq_sch_rem_beats_nxt ;
    p4_direnq_sch_qid_v_f               <= p4_direnq_sch_qid_v_nxt ;
    p4_direnq_sch_cq_avail_f            <= p4_direnq_sch_cq_avail_nxt ;
    p4_direnq_sch_wp_f                  <= p4_direnq_sch_wp_nxt ;
    p4_direnq_sch_disab_opt_f           <= p4_direnq_sch_disab_opt_nxt ;
    p4_direnq_sch_first_beat_f          <= p4_direnq_sch_first_beat_nxt ;
    p4_direnq_sch_first_clock_f         <= p4_direnq_sch_first_clock_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
assign dir_sel_dp_fifo_push             = p3_direnq_sch_out ;             // Includes ~afull

always_comb begin
  dir_sel_dp_fifo_push_data.cq                                  = '0 ;
  dir_sel_dp_fifo_push_data.cq [HQM_NUM_DIR_CQB2-1:0]           = p3_direnq_sch_out_qid ;
  dir_sel_dp_fifo_push_data.qid                                 = '0 ;
  dir_sel_dp_fifo_push_data.qid [HQM_NUM_DIR_QIDB2-1:0]         = p3_direnq_sch_out_qid ;
  dir_sel_dp_fifo_push_data.qidix                               = 3'h0 ;                        // Unused by Directed
  dir_sel_dp_fifo_push_data.parity                              = 1'b1 ^ cfg_error_inject_f [ 9 ] ;     // qid & qid
  dir_sel_dp_fifo_push_data.hqm_core_flags.pad_ok                       = '0 ;
  dir_sel_dp_fifo_push_data.hqm_core_flags.ignore_cq_depth              = 1'b0 ;        // repurpose to carry qidix_msb
  dir_sel_dp_fifo_push_data.hqm_core_flags.cq_is_ldb                    = 1'b0 ;        // Directed, not lb
  dir_sel_dp_fifo_push_data.hqm_core_flags.write_buffer_optimization    = p3_direnq_rem_beats_m1 ;      // Conditionally overridden on output if not fill_in_progress
  dir_sel_dp_fifo_push_data.hqm_core_flags.congestion_management        = p3_direnq_sch_out_cm_code ;
  dir_sel_dp_fifo_push_data.hqm_core_flags.parity                       = 1'b0 ;        // Totally calculated on output; DB contents not protected by parity
  dir_sel_dp_fifo_push_data.fill_in_progress                    = p3_direnq_fill_in_progress ;
  dir_sel_dp_fifo_push_data.qid_v                               = p3_direnq_arb_winner_qid_v ;
  dir_sel_dp_fifo_push_data.cq_avail                            = p3_direnq_arb_winner_cq_avail ;
  dir_sel_dp_fifo_push_data.wp                                  = p3_direnq_arb_winner_wp ;
  dir_sel_dp_fifo_push_data.disab_opt                           = p3_direnq_arb_winner_disab_opt ;
end // always

assign dir_sel_dp_db_in_valid           = dir_sel_dp_fifo_push ;
assign dir_sel_dp_db_in_data            = dir_sel_dp_fifo_push_data ;
assign dir_sel_dp_fifo_afull            = ~ dir_sel_dp_db_in_ready ;
assign dir_sel_dp_fifo_empty            = lsp_dp_sch_dir_tx_sync_idle ;
assign dir_sel_dp_fifo_hold             = dir_sel_dp_fifo_afull | ( cfg_control_single_out_direnq & ~ dir_sel_dp_fifo_empty ) ;

// dir_sel_dp_db_in_data goes to i_hqm_AW_tx_sync_lsp_dp_sch_dir

assign lsp_dp_sch_dir_data_write_buffer_optimization       = ( lsp_dp_sch_dir_pre_data.fill_in_progress )
                                                               ? lsp_dp_sch_dir_pre_data.hqm_core_flags.write_buffer_optimization       // calc already OK for non-first iter
                                                               : ( lsp_dp_sch_dir_pre_data.disab_opt )
                                                                  ? 2'h0
                                                                  : hqm_lsp_dir_rem_beats (   lsp_dp_sch_dir_pre_data.qid_v             // calc on the fly for first iter
                                                                                            , lsp_dp_sch_dir_pre_data.cq_avail
                                                                                            , lsp_dp_sch_dir_pre_data.wp ) ;

assign lsp_dp_sch_dir_data.cq                              = lsp_dp_sch_dir_pre_data.cq ;
assign lsp_dp_sch_dir_data.qid                             = lsp_dp_sch_dir_pre_data.qid ;
assign lsp_dp_sch_dir_data.qidix                           = lsp_dp_sch_dir_pre_data.qidix ;
assign lsp_dp_sch_dir_data.parity                          = lsp_dp_sch_dir_pre_data.parity ;
assign lsp_dp_sch_dir_data.hqm_core_flags.pad_ok                        = lsp_dp_sch_dir_pre_data.hqm_core_flags.pad_ok ;
assign lsp_dp_sch_dir_data.hqm_core_flags.ignore_cq_depth               = 1'b0 ;    // repurpose to carry qidix_msb
assign lsp_dp_sch_dir_data.hqm_core_flags.cq_is_ldb                     = lsp_dp_sch_dir_pre_data.hqm_core_flags.cq_is_ldb ;
assign lsp_dp_sch_dir_data.hqm_core_flags.write_buffer_optimization     = lsp_dp_sch_dir_data_write_buffer_optimization ;
assign lsp_dp_sch_dir_data.hqm_core_flags.congestion_management         = lsp_dp_sch_dir_pre_data.hqm_core_flags.congestion_management ;

hqm_AW_parity_gen #( .WIDTH ( 4 ) ) i_dp_sch_dir_flag_par_gen (                         // Potential timing issue
          .d            ( {                                                                     // pad_ok always 0
                                                                                                // repurpose to carry qidix_msb, always 0 for dir 
                                                                                                // cq_is_ldb is always 0 (DIR)
                              lsp_dp_sch_dir_data_write_buffer_optimization                     // Modified on FIFO output, need to get
                            , lsp_dp_sch_dir_pre_data.hqm_core_flags.congestion_management } )  // No modification, straight from FIFO
        , .odd          ( 1'b1 )
        , .p            ( lsp_dp_sch_dir_data.hqm_core_flags.parity )
) ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: LBRPL pipe - Detects LB "reorder complete" notifications and adds the frag count
// to the specified qid's count, then schedules out replay requests one at a time.
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBRPL input pipe arbitration
//-----------------------------------------------------------------------------------------------------
// There are 2 functional inputs to the LBRPL pipe: fragment "enqueue" requests and replay "schedule"
// requests.  A simple 50/50 weighted random arbiter is used.
assign lbrpl_input_arb_reqs [0]        = nalbrpl_fifo_pop_data_vreq ;
assign lbrpl_input_arb_reqs [1]        = p4_lbrpl_sch_v_f ;

hqm_AW_wrand_arb # ( .NUM_REQS ( 2 ) , .SEED ( 1 ) ) i_lbrpl_input_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( lbrpl_input_arb_reqs )
        , .cfg_weight           ( { HQM_LSP_LBRPL_INPUT_ARB_WEIGHT_REQ1 ,               // Equal weights = random
                                    HQM_LSP_LBRPL_INPUT_ARB_WEIGHT_REQ0 } )
        , .winner_v             ( lbrpl_input_arb_winner_pre_v )
        , .winner               ( lbrpl_input_arb_winner )
) ;

assign lbrpl_input_arb_winner_v = lbrpl_input_arb_winner_pre_v &
                                  ~ ( ( cfg_control_single_op_lbrpl & ( ( ~ lbrpl_upipe_idle_f ) | p0_lbrpl_ctrl_pipe_v_f ) ) |
                                      ( cfg_control_half_bw_lbrpl & p0_lbrpl_ctrl_pipe_v_f ) ) ;

assign lbrpl_input_arb_sch      = lbrpl_input_arb_winner_v &   lbrpl_input_arb_winner & ~ p0_lbrpl_ctrl_pipe.hold ;
assign lbrpl_input_arb_enq      = lbrpl_input_arb_winner_v & ~ lbrpl_input_arb_winner & ~ p0_lbrpl_ctrl_pipe.hold ;
assign lbrpl_input_arb_sch_qid  = p4_lbrpl_sch_qid_f ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBRPL enqueue count pipe
//-----------------------------------------------------------------------------------------------------

assign lbrpl_input_req_v                = lbrpl_input_arb_enq | lbrpl_input_arb_sch ;

// lbrpl_input_req_v is effectively the "pipeline valid" for the lbrpl inputs
assign p0_lbrpl_ctrl_pipe.hold          = p0_lbrpl_ctrl_pipe_v_f & p1_lbrpl_ctrl_pipe.hold ;
assign p0_lbrpl_ctrl_pipe.en            = lbrpl_input_req_v & ~ p0_lbrpl_ctrl_pipe.hold ;
assign p0_lbrpl_ctrl_pipe_v_nxt         = lbrpl_input_req_v | p0_lbrpl_ctrl_pipe.hold ;
assign p0_lbrpl_ctrl_pipe_v_nxt_gated   = p0_lbrpl_ctrl_pipe_v_nxt & ~ p0_lbrpl_ctrl_pipe.hold ;


always_comb begin
  p0_lbrpl_ctrl_pipe_nxt                        = p0_lbrpl_ctrl_pipe_f ;
  if ( p0_lbrpl_ctrl_pipe.en ) begin
    p0_lbrpl_ctrl_pipe_nxt                      = '0 ;                                  // Safety belt just in case any bits missed
    p0_lbrpl_ctrl_pipe_nxt.enq_v                = lbrpl_input_arb_enq ;
    if ( lbrpl_input_arb_sch )
      p0_lbrpl_ctrl_pipe_nxt.qid_p              = lbrpl_input_arb_sch_qid.qid_p ;
    else
      p0_lbrpl_ctrl_pipe_nxt.qid_p              = nalbrpl_fifo_pop_data.parity ^ ( ^ nalbrpl_fifo_pop_data.qtype ) ;    // subtract out qtype parity
    p0_lbrpl_ctrl_pipe_nxt.frag_cnt             = nalbrpl_fifo_pop_data.frag_cnt ;
    p0_lbrpl_ctrl_pipe_nxt.frag_cnt_res         = nalbrpl_fifo_pop_data.frag_residue ;
    p0_lbrpl_ctrl_pipe_nxt.sch_v                = lbrpl_input_arb_sch ;
    p0_lbrpl_ctrl_pipe_nxt.blast_enq            = lbrpl_input_arb_enq &
                                                  ( ( p4_lbrpl_sch_v_f &   ( nalbrpl_fifo_pop_data.qid == p4_lbrpl_sch_qid_f.qid ) ) |
                                                    ( p3_lbrpl_sch_start & ( nalbrpl_fifo_pop_data.qid == p3_lbrpl_sch_start_qid ) ) ) ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p0_lbrpl_ctrl_pipe_f                  <= p0_lbrpl_ctrl_pipe_nxt ;
  p1_lbrpl_ctrl_pipe_f                  <= p1_lbrpl_ctrl_pipe_nxt ;
  p2_lbrpl_ctrl_pipe_f                  <= p2_lbrpl_ctrl_pipe_nxt ;
end // always

assign p1_lbrpl_ctrl_pipe.hold          = p1_lbrpl_ctrl_pipe_v_f & p2_lbrpl_ctrl_pipe.hold ;
assign p1_lbrpl_ctrl_pipe.en            = p0_lbrpl_ctrl_pipe_v_f & ~ p1_lbrpl_ctrl_pipe.hold ;

assign p2_lbrpl_ctrl_pipe.hold          = p2_lbrpl_ctrl_pipe_v_f & p3_lbrpl_ctrl_pipe.hold ;
assign p2_lbrpl_ctrl_pipe.en            = p1_lbrpl_ctrl_pipe_v_f & ~ p2_lbrpl_ctrl_pipe.hold ;

assign p3_lbrpl_ctrl_pipe.hold          = 1'b0 ;                                        // p3 qid status FFs always able to load
assign p3_lbrpl_ctrl_pipe.en            = p2_lbrpl_ctrl_pipe_v_f & ~ p3_lbrpl_ctrl_pipe.hold ;

always_comb begin
  p1_lbrpl_ctrl_pipe_nxt                = p1_lbrpl_ctrl_pipe_f ;
  p2_lbrpl_ctrl_pipe_nxt                = p2_lbrpl_ctrl_pipe_f ;

  if ( p1_lbrpl_ctrl_pipe.en ) begin
    p1_lbrpl_ctrl_pipe_nxt              = p0_lbrpl_ctrl_pipe_f ;
    p1_lbrpl_ctrl_pipe_nxt.blast_enq    = p0_lbrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_lbrpl_sch_start & ( p3_lbrpl_sch_start_qid == p0_lbrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p0_lbrpl_ctrl_pipe_f.enq_v ) ;
  end
  else if ( p1_lbrpl_ctrl_pipe.hold ) begin     // Need to blast writes which are holding
    p1_lbrpl_ctrl_pipe_nxt.blast_enq    = p1_lbrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_lbrpl_sch_start & ( p3_lbrpl_sch_start_qid == p1_lbrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_lbrpl_ctrl_pipe_f.enq_v ) ;
  end

  if ( p2_lbrpl_ctrl_pipe.en ) begin
    p2_lbrpl_ctrl_pipe_nxt              = p1_lbrpl_ctrl_pipe_f ;
    p2_lbrpl_ctrl_pipe_nxt.blast_enq    = p1_lbrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_lbrpl_sch_start & ( p3_lbrpl_sch_start_qid == p1_lbrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_lbrpl_ctrl_pipe_f.enq_v ) ;
  end
  else if ( p2_lbrpl_ctrl_pipe.hold ) begin     // Need to blast writes which are holding
    p2_lbrpl_ctrl_pipe_nxt.blast_enq    = p2_lbrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_lbrpl_sch_start & ( p3_lbrpl_sch_start_qid == p2_lbrpl_enq_cnt_rmw_pipe_f.qid ) &
                                            p2_lbrpl_ctrl_pipe_f.enq_v ) ;
  end
end // always

assign p2_lbrpl_enq_cnt_upd_v           = ( p2_lbrpl_enq_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_lbrpl_ctrl_pipe.en ;

always_comb begin
  p0_lbrpl_enq_cnt_rmw_pipe_nxt.rw_cmd          = HQM_AW_RMWPIPE_RMW ;
  if ( lbrpl_input_arb_sch ) begin
    p0_lbrpl_enq_cnt_rmw_pipe_nxt.qid           = lbrpl_input_arb_sch_qid.qid ;
  end
  else begin
    p0_lbrpl_enq_cnt_rmw_pipe_nxt.qid           = nalbrpl_fifo_pop_data.qid ;
  end
  p0_lbrpl_enq_cnt_rmw_pipe_nxt.data            = { $bits ( lsp_lbrpl_enq_cnt_t ) { 1'b0 } } ;          // Unused - cfg write done elsewhere
end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for lbrpl enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )
        , .WIDTH                ( HQM_LSP_LBRPL_ENQ_CNT_MEM_WIDTH )
) i_lb_replay_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( lbrpl_enq_cnt_rmw_pipe_status )

        // cmd input
        , .p0_hold              ( p0_lbrpl_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_lbrpl_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_lbrpl_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_lbrpl_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_lbrpl_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_lbrpl_ctrl_pipe_v_f )
        , .p0_rw_f              ( p0_lbrpl_enq_cnt_rmw_pipe_f_pnc.rw_cmd )      // Unused
        , .p0_addr_f            ( p0_lbrpl_enq_cnt_rmw_pipe_f_pnc.qid )         // Used by blast logic
        , .p0_data_f            ( p0_lbrpl_enq_cnt_rmw_pipe_f_pnc.data )        // Unused

        , .p1_hold              ( p1_lbrpl_ctrl_pipe.hold )
        , .p1_v_f               ( p1_lbrpl_ctrl_pipe_v_f )
        , .p1_rw_f              ( p1_lbrpl_enq_cnt_rmw_pipe_f_pnc.rw_cmd )      // Unused
        , .p1_addr_f            ( p1_lbrpl_enq_cnt_rmw_pipe_f_pnc.qid )         // Used by blast logic and input error rid
        , .p1_data_f            ( p1_lbrpl_enq_cnt_rmw_pipe_f_pnc.data )        // Unused

        , .p2_hold              ( p2_lbrpl_ctrl_pipe.hold )
        , .p2_v_f               ( p2_lbrpl_ctrl_pipe_v_f )
        , .p2_rw_f              ( p2_lbrpl_enq_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_lbrpl_enq_cnt_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_lbrpl_enq_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_lbrpl_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_lbrpl_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_lbrpl_enq_cnt_upd )
        , .p3_v_f               ( p3_lbrpl_ctrl_pipe_v_f )
        , .p3_rw_f              ( p3_lbrpl_enq_cnt_rmw_pipe_f_nc.rw_cmd )       // Unused
        , .p3_addr_f            ( p3_lbrpl_enq_cnt_rmw_pipe_f_nc.qid )          // Unused
        , .p3_data_f            ( p3_lbrpl_enq_cnt_rmw_pipe_f_nc.data )         // Unused

        // mem intf
        , .mem_write            ( func_qid_ldb_replay_count_mem_we )
        , .mem_read             ( func_qid_ldb_replay_count_mem_re )
        , .mem_write_addr       ( func_qid_ldb_replay_count_mem_waddr )
        , .mem_read_addr        ( func_qid_ldb_replay_count_mem_raddr )
        , .mem_write_data       ( func_qid_ldb_replay_count_mem_wdata )
        , .mem_read_data        ( func_qid_ldb_replay_count_mem_rdata )
    ) ;

hqm_AW_residue_add i_lbrpl_enq_cnt_res_add (
          .a                    ( p2_lbrpl_ctrl_pipe_f.frag_cnt_res )
        , .b                    ( p2_lbrpl_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_lbrpl_enq_cnt_res_pn )
) ;

hqm_AW_residue_sub i_lbrpl_enq_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p2_lbrpl_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_lbrpl_enq_cnt_res_m1 )
) ;

// Interface supports 15-bit frag_cnt, max possible total count is 14 bits (8K LDB credits), count memory supports 16 bits (2 spares)
assign { p2_lbrpl_enq_cnt_pn_carry , p2_lbrpl_enq_cnt_pn }      = { 1'b0 , p2_lbrpl_enq_cnt_rmw_pipe_f.data.cnt } + { 2'h0 , p2_lbrpl_ctrl_pipe_f.frag_cnt } ;
assign { p2_lbrpl_enq_cnt_m1_borrow , p2_lbrpl_enq_cnt_m1 }     = { 1'b0 , p2_lbrpl_enq_cnt_rmw_pipe_f.data.cnt } - {{HQM_LSP_LBRPL_ENQ_CNT_WIDTH{1'b0}}, 1'b1} ;

always_comb begin
  p2_lbrpl_enq_cnt_oflow_cond                   = 1'b0 ;
  p2_lbrpl_enq_cnt_uflow_cond                   = 1'b0 ;
  if ( p2_lbrpl_ctrl_pipe_f.sch_v ) begin
    if ( p2_lbrpl_enq_cnt_m1_borrow ) begin
      p2_lbrpl_enq_cnt_upd                      = p2_lbrpl_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_lbrpl_enq_cnt_uflow_cond               = 1'b1 ;
    end
    else begin
      p2_lbrpl_enq_cnt_upd.cnt                  = p2_lbrpl_enq_cnt_m1 ;
      p2_lbrpl_enq_cnt_upd.cnt_res              = p2_lbrpl_enq_cnt_res_m1 ;
    end
  end
  else begin
    if ( p2_lbrpl_enq_cnt_pn_carry ) begin
      p2_lbrpl_enq_cnt_upd                      = p2_lbrpl_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_lbrpl_enq_cnt_oflow_cond               = 1'b1 ;
    end
    else begin
      p2_lbrpl_enq_cnt_upd.cnt                  = p2_lbrpl_enq_cnt_pn ;
      p2_lbrpl_enq_cnt_upd.cnt_res              = p2_lbrpl_enq_cnt_res_pn ;
    end
  end
end // always

assign p2_lbrpl_enq_cnt_upd_gt0                 = | ( p2_lbrpl_enq_cnt_upd.cnt ) ;



assign p0_lbrpl_inp_frag_cnt_res_chk_en         = p0_lbrpl_ctrl_pipe_f.enq_v ;

hqm_AW_residue_check #( .WIDTH ( 15 ) ) i_lbrpl_inp_frag_cnt_res_chk (
          .r                    ( p0_lbrpl_ctrl_pipe_f.frag_cnt_res )
        , .d                    ( p0_lbrpl_ctrl_pipe_f.frag_cnt )
        , .e                    ( p0_lbrpl_inp_frag_cnt_res_chk_en )
        , .err                  ( p0_lbrpl_inp_frag_cnt_res_err_cond )
) ;



assign p2_lbrpl_enq_cnt_res_chk_en              = p2_lbrpl_enq_cnt_upd_v ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_LBRPL_ENQ_CNT_WIDTH ) ) i_lbrpl_enq_cnt_res_chk (
          .r                    ( p3_lbrpl_enq_cnt_f.cnt_res )
        , .d                    ( p3_lbrpl_enq_cnt_f.cnt )
        , .e                    ( p3_lbrpl_enq_cnt_res_chk_en_f )
        , .err                  ( p3_lbrpl_enq_cnt_res_err )
) ;

assign p2_lbrpl_inp_qid_par_chk_en = p2_lbrpl_enq_cnt_upd_v ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_lbrpl_inp_qid_par_chk (
          .p                    ( p2_lbrpl_ctrl_pipe_f.qid_p )
        , .d                    ( p2_lbrpl_enq_cnt_rmw_pipe_f.qid )
        , .e                    ( p2_lbrpl_inp_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_lbrpl_inp_qid_par_err_cond )
) ;

//-------------------------------------------------------------------------------------------------
// Underflow/overflow errors - some are impossible, some may be caused by software/config errors
//

always_comb begin
  // Don't hold error flops - 1-clock pulse to report
  p3_lbrpl_enq_cnt_uflow_err_nxt        = 1'b0 ;
  p3_lbrpl_enq_cnt_oflow_err_nxt        = 1'b0 ;

  p1_lbrpl_inp_frag_cnt_res_err_nxt     = 1'b0 ;
  p3_lbrpl_inp_qid_par_err_nxt          = 1'b0 ;

  p3_lbrpl_enq_cnt_res_chk_en_nxt       = 1'b0 ;
  p3_lbrpl_enq_cnt_nxt                  = p3_lbrpl_enq_cnt_f ;

  if ( p0_lbrpl_ctrl_pipe_v_f & ~ p1_lbrpl_ctrl_pipe.hold ) begin
    p1_lbrpl_inp_frag_cnt_res_err_nxt   = p0_lbrpl_inp_frag_cnt_res_err_cond ;
  end

  if ( p2_lbrpl_ctrl_pipe_v_f & ~ p3_lbrpl_ctrl_pipe.hold ) begin
    p3_lbrpl_enq_cnt_uflow_err_nxt      = p2_lbrpl_ctrl_pipe_f.sch_v & p2_lbrpl_enq_cnt_uflow_cond ;
    p3_lbrpl_enq_cnt_oflow_err_nxt      = p2_lbrpl_ctrl_pipe_f.enq_v & p2_lbrpl_enq_cnt_oflow_cond ;

    p3_lbrpl_inp_qid_par_err_nxt        = p2_lbrpl_inp_qid_par_err_cond ;

    p3_lbrpl_enq_cnt_res_chk_en_nxt     = p2_lbrpl_enq_cnt_res_chk_en ;
    p3_lbrpl_enq_cnt_nxt                = p2_lbrpl_enq_cnt_upd ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_lbrpl_enq_cnt_uflow_err_f        <= 1'b0 ;
    p3_lbrpl_enq_cnt_oflow_err_f        <= 1'b0 ;

    p1_lbrpl_inp_frag_cnt_res_err_f     <= 1'b0 ;
    p3_lbrpl_inp_qid_par_err_f          <= 1'b0 ;

    p3_lbrpl_enq_cnt_res_chk_en_f       <= 1'b0 ;
  end
  else begin
    p3_lbrpl_enq_cnt_uflow_err_f        <= p3_lbrpl_enq_cnt_uflow_err_nxt ;
    p3_lbrpl_enq_cnt_oflow_err_f        <= p3_lbrpl_enq_cnt_oflow_err_nxt ;

    p1_lbrpl_inp_frag_cnt_res_err_f     <= p1_lbrpl_inp_frag_cnt_res_err_nxt ;
    p3_lbrpl_inp_qid_par_err_f          <= p3_lbrpl_inp_qid_par_err_nxt ;

    p3_lbrpl_enq_cnt_res_chk_en_f       <= p3_lbrpl_enq_cnt_res_chk_en_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p3_lbrpl_enq_cnt_f                    <= p3_lbrpl_enq_cnt_nxt ;
end // always

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: LBRPL p3 qid_v status vector
//-----------------------------------------------------------------------------------------------------
// See comments under DIRENQ regarding scheduling terminology

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
    // Bypass update from sch takes precedence over update from p2; sch update will cause subsequent write
    // of latest/correct value of count caused by this scheduling.
    // enq updates from upper pipe must be supressed from "enabling" if they were blasted by newer scheduling.
    p3_lbrpl_sch_hit[i]                 = p3_lbrpl_sch_start & ( p3_lbrpl_sch_start_qid == i ) ;
    p3_lbrpl_p2_enq_hit[i]              = p3_lbrpl_ctrl_pipe.en & ( p2_lbrpl_ctrl_pipe_f.enq_v | p2_lbrpl_ctrl_pipe_f.sch_v ) &
                                           ( p2_lbrpl_enq_cnt_rmw_pipe_f.qid == i ) & ~ p2_lbrpl_ctrl_pipe_f.blast_enq ;
  end // for
end // always

// For each lbrpl qid maintain state for "qid has data" (qid_v)
// Update (set to 0 or 1) when enq count is updated, reset when that qid is selected to be scheduled.
// Should be cleared as part of a successful vas reset drain
always_comb begin
  p3_lbrpl_arb_stat_nxt                 = p3_lbrpl_arb_stat_f ;
  if ( p3_lbrpl_sch_start | p3_lbrpl_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      if ( p3_lbrpl_sch_hit[i] )
        p3_lbrpl_arb_stat_nxt[i].qid_v          = 1'b0 ;
      else if ( p3_lbrpl_p2_enq_hit[i] )
        p3_lbrpl_arb_stat_nxt[i].qid_v          = p2_lbrpl_enq_cnt_upd_gt0 ;
    end // for i
  end // if
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      p3_lbrpl_arb_stat_f[i].qid_v      <= 1'b0 ;
    end
  end
  else begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
      p3_lbrpl_arb_stat_f[i]            <= p3_lbrpl_arb_stat_nxt[i] ;
    end // for i
  end // else rst_n

end // always

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
    p3_lbrpl_arb_reqs [i]               = p3_lbrpl_arb_stat_f[i].qid_v ;
    cfg_qid_ldb_replay_v_status [i]     = p3_lbrpl_arb_stat_f[i].qid_v ;
  end // for i
end // always

hqm_AW_rr_arb # ( .NUM_REQS ( HQM_NUM_LB_QID ) ) i_lbrpl_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p3_lbrpl_arb_reqs )
        , .update               ( p3_lbrpl_arb_update )
        , .winner_v             ( p3_lbrpl_arb_winner_pre_v )
        , .winner               ( p3_lbrpl_arb_winner )
) ;
assign p3_lbrpl_arb_winner_v            = p3_lbrpl_arb_winner_pre_v & ~ cause_pipe_idle ;

hqm_AW_parity_gen #( .WIDTH( HQM_NUM_LB_QIDB2 ) ) i_lbrpl_sch_qid_par_gen (
          .d            ( p3_lbrpl_arb_winner )
        , .odd          ( 1'b1 )
        , .p            ( p3_lbrpl_arb_winner_gp )
) ;

always_comb begin
  p3_lbrpl_sch_req                                      = p3_lbrpl_arb_winner_v & ~ rpl_ldb_nalb_fifo_hold & ~ p4_lbrpl_sch_hold ;
  p3_lbrpl_sch_stall_smon                               = p3_lbrpl_arb_winner_v &   rpl_ldb_nalb_fifo_hold & ~ p4_lbrpl_sch_hold ;      // For smon only
  p3_lbrpl_sch_req_qid.qid                              = { HQM_LSP_ARCH_NUM_LB_QIDB2 { 1'b0 } } ;
  p3_lbrpl_sch_req_qid.qid [HQM_NUM_LB_QIDB2-1:0]       = p3_lbrpl_arb_winner ;
  p3_lbrpl_sch_req_qid.qid_p                            = p3_lbrpl_arb_winner_gp ;
end // always

assign p3_lbrpl_arb_update              = p3_lbrpl_sch_req ;

assign p3_lbrpl_sch_start               = p3_lbrpl_sch_req ;
assign p3_lbrpl_sch_start_qid           = p3_lbrpl_sch_req_qid.qid ;

assign p4_lbrpl_sch_hold                = p4_lbrpl_sch_v_f & ~ lbrpl_input_arb_sch ;
assign p4_lbrpl_sch_v_nxt               = p3_lbrpl_sch_req | p4_lbrpl_sch_hold ;

always_comb begin
  p4_lbrpl_sch_qid_nxt                  = p4_lbrpl_sch_qid_f ;
  if ( p3_lbrpl_sch_req & ~ p4_lbrpl_sch_hold )
    p4_lbrpl_sch_qid_nxt                = p3_lbrpl_sch_req_qid ;
end //always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p4_lbrpl_sch_v_f                    <= 1'b0 ;
  end
  else begin
    p4_lbrpl_sch_v_f                    <= p4_lbrpl_sch_v_nxt ;
  end
end // always
always_ff @ ( posedge hqm_gated_clk ) begin
  p4_lbrpl_sch_qid_f                    <= p4_lbrpl_sch_qid_nxt ;
end // always

//-------------------------------------------------------------------------------------------------
// Output FIFO (DB) - for static timing isolation
assign rpl_ldb_nalb_fifo_push                   = p3_lbrpl_sch_req ;            // sch_req already has afull in equation
assign rpl_ldb_nalb_fifo_push_data.parity       = p3_lbrpl_sch_req_qid.qid_p ^ cfg_error_inject_f [ 14 ] ;
assign rpl_ldb_nalb_fifo_push_data.qid          = p3_lbrpl_sch_req_qid.qid ;

assign rpl_ldb_nalb_db_in_valid                 = rpl_ldb_nalb_fifo_push ;
assign rpl_ldb_nalb_db_in_data                  = rpl_ldb_nalb_fifo_push_data ;
assign rpl_ldb_nalb_fifo_afull                  = ~ rpl_ldb_nalb_db_in_ready ;
assign rpl_ldb_nalb_fifo_empty                  = rpl_ldb_nalb_tx_sync_idle ;
assign rpl_ldb_nalb_fifo_hold                   = rpl_ldb_nalb_fifo_afull | ( cfg_control_single_out_lbrpl & ~ rpl_ldb_nalb_fifo_empty ) ;

// rpl_ldb_nalb_db_in_data goes to i_hqm_AW_tx_sync_rpl_ldb_nalb

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: DIRRPL pipe - Detects directed "reorder complete" notifications and adds the frag count
// to the specified qid's count, then schedules out replay requests one at a time.  Note that qid is
// the originating (ORD) qid (load-balanced), so structures are scaled by LB QID.
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: DIRRPL input pipe arbitration
//-----------------------------------------------------------------------------------------------------
// There are 2 functional inputs to the DIRRPL pipe: fragment "enqueue" requests and replay "schedule"
// requests.  A simple 50/50 weighted random arbiter is used.
assign dirrpl_input_arb_reqs [0]        = dirrpl_fifo_pop_data_vreq ;
assign dirrpl_input_arb_reqs [1]        = p4_dirrpl_sch_v_f ;

hqm_AW_wrand_arb # ( .NUM_REQS ( 2 ) , .SEED ( 1 ) ) i_dirrpl_input_arb (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( dirrpl_input_arb_reqs )
        , .cfg_weight           ( { HQM_LSP_DIRRPL_INPUT_ARB_WEIGHT_REQ1 ,              // Equal weights = random
                                    HQM_LSP_DIRRPL_INPUT_ARB_WEIGHT_REQ0 } )
        , .winner_v             ( dirrpl_input_arb_winner_pre_v )
        , .winner               ( dirrpl_input_arb_winner )
) ;

assign dirrpl_input_arb_winner_v        = dirrpl_input_arb_winner_pre_v &
                                          ~ ( ( cfg_control_single_op_dirrpl & ( ( ~ dirrpl_upipe_idle_f ) | p0_dirrpl_ctrl_pipe_v_f ) ) |
                                              ( cfg_control_half_bw_dirrpl & p0_dirrpl_ctrl_pipe_v_f ) ) ;

assign dirrpl_input_arb_sch     = dirrpl_input_arb_winner_v &   dirrpl_input_arb_winner & ~ p0_dirrpl_ctrl_pipe.hold ;
assign dirrpl_input_arb_enq     = dirrpl_input_arb_winner_v & ~ dirrpl_input_arb_winner & ~ p0_dirrpl_ctrl_pipe.hold ;
assign dirrpl_input_arb_sch_qid = p4_dirrpl_sch_qid_f ;

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: DIRRPL enqueue count pipe
//-----------------------------------------------------------------------------------------------------

assign dirrpl_input_req_v               = dirrpl_input_arb_enq | dirrpl_input_arb_sch ;

// dirrpl_input_req_v is effectively the "pipeline valid" for the dirrpl inputs
assign p0_dirrpl_ctrl_pipe.hold         = p0_dirrpl_ctrl_pipe_v_f & p1_dirrpl_ctrl_pipe.hold ;
assign p0_dirrpl_ctrl_pipe.en           = dirrpl_input_req_v & ~ p0_dirrpl_ctrl_pipe.hold ;
assign p0_dirrpl_ctrl_pipe_v_nxt        = dirrpl_input_req_v | p0_dirrpl_ctrl_pipe.hold ;
assign p0_dirrpl_ctrl_pipe_v_nxt_gated  = p0_dirrpl_ctrl_pipe_v_nxt & ~ p0_dirrpl_ctrl_pipe.hold ;

always_comb begin
  p0_dirrpl_ctrl_pipe_nxt                       = p0_dirrpl_ctrl_pipe_f ;
  if ( p0_dirrpl_ctrl_pipe.en ) begin
    p0_dirrpl_ctrl_pipe_nxt                     = '0 ;                                  // Safety belt just in case any bits missed
    p0_dirrpl_ctrl_pipe_nxt.enq_v               = dirrpl_input_arb_enq ;
    if ( dirrpl_input_arb_sch )
      p0_dirrpl_ctrl_pipe_nxt.qid_p             = dirrpl_input_arb_sch_qid.qid_p ;
    else
      p0_dirrpl_ctrl_pipe_nxt.qid_p             = dirrpl_fifo_pop_data.parity ;
    p0_dirrpl_ctrl_pipe_nxt.frag_cnt            = dirrpl_fifo_pop_data.frag_cnt ;
    p0_dirrpl_ctrl_pipe_nxt.frag_cnt_res        = dirrpl_fifo_pop_data.frag_residue ;
    p0_dirrpl_ctrl_pipe_nxt.sch_v               = dirrpl_input_arb_sch ;
    p0_dirrpl_ctrl_pipe_nxt.blast_enq           = dirrpl_input_arb_enq &
                                                  ( ( p4_dirrpl_sch_v_f &   ( dirrpl_fifo_pop_data.qid == p4_dirrpl_sch_qid_f.qid ) ) |
                                                    ( p3_dirrpl_sch_start & ( dirrpl_fifo_pop_data.qid == p3_dirrpl_sch_start_qid ) ) ) ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p0_dirrpl_ctrl_pipe_f                 <= p0_dirrpl_ctrl_pipe_nxt ;
  p1_dirrpl_ctrl_pipe_f                 <= p1_dirrpl_ctrl_pipe_nxt ;
  p2_dirrpl_ctrl_pipe_f                 <= p2_dirrpl_ctrl_pipe_nxt ;
end // always

assign p1_dirrpl_ctrl_pipe.hold         = p1_dirrpl_ctrl_pipe_v_f & p2_dirrpl_ctrl_pipe.hold ;
assign p1_dirrpl_ctrl_pipe.en           = p0_dirrpl_ctrl_pipe_v_f & ~ p1_dirrpl_ctrl_pipe.hold ;

assign p2_dirrpl_ctrl_pipe.hold         = p2_dirrpl_ctrl_pipe_v_f & p3_dirrpl_ctrl_pipe.hold ;
assign p2_dirrpl_ctrl_pipe.en           = p1_dirrpl_ctrl_pipe_v_f & ~ p2_dirrpl_ctrl_pipe.hold ;

assign p3_dirrpl_ctrl_pipe.hold         = 1'b0 ;                                        // p3 qid status FFs always able to load
assign p3_dirrpl_ctrl_pipe.en           = p2_dirrpl_ctrl_pipe_v_f & ~ p3_dirrpl_ctrl_pipe.hold ;

always_comb begin
  p1_dirrpl_ctrl_pipe_nxt               = p1_dirrpl_ctrl_pipe_f ;
  p2_dirrpl_ctrl_pipe_nxt               = p2_dirrpl_ctrl_pipe_f ;

  if ( p1_dirrpl_ctrl_pipe.en ) begin
    p1_dirrpl_ctrl_pipe_nxt             = p0_dirrpl_ctrl_pipe_f ;
    p1_dirrpl_ctrl_pipe_nxt.blast_enq   = p0_dirrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_dirrpl_sch_start & ( p3_dirrpl_sch_start_qid == p0_dirrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p0_dirrpl_ctrl_pipe_f.enq_v ) ;
  end
  else if ( p1_dirrpl_ctrl_pipe.hold ) begin    // Need to blast writes which are holding
    p1_dirrpl_ctrl_pipe_nxt.blast_enq   = p1_dirrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_dirrpl_sch_start & ( p3_dirrpl_sch_start_qid == p1_dirrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_dirrpl_ctrl_pipe_f.enq_v ) ;
  end

  if ( p2_dirrpl_ctrl_pipe.en ) begin
    p2_dirrpl_ctrl_pipe_nxt             = p1_dirrpl_ctrl_pipe_f ;
    p2_dirrpl_ctrl_pipe_nxt.blast_enq   = p1_dirrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_dirrpl_sch_start & ( p3_dirrpl_sch_start_qid == p1_dirrpl_enq_cnt_rmw_pipe_f_pnc.qid ) &
                                            p1_dirrpl_ctrl_pipe_f.enq_v ) ;
  end
  else if ( p2_dirrpl_ctrl_pipe.hold ) begin    // Need to blast writes which are holding
    p2_dirrpl_ctrl_pipe_nxt.blast_enq   = p2_dirrpl_ctrl_pipe_f.blast_enq |
                                          ( p3_dirrpl_sch_start & ( p3_dirrpl_sch_start_qid == p2_dirrpl_enq_cnt_rmw_pipe_f.qid ) &
                                            p2_dirrpl_ctrl_pipe_f.enq_v ) ;
  end
end // always

assign p2_dirrpl_enq_cnt_upd_v          = ( p2_dirrpl_enq_cnt_rmw_pipe_f.rw_cmd == HQM_AW_RMWPIPE_RMW ) & p3_dirrpl_ctrl_pipe.en ;

always_comb begin
  p0_dirrpl_enq_cnt_rmw_pipe_nxt.rw_cmd         = HQM_AW_RMWPIPE_RMW ;
  if ( dirrpl_input_arb_sch ) begin
    p0_dirrpl_enq_cnt_rmw_pipe_nxt.qid          = dirrpl_input_arb_sch_qid.qid ;
  end
  else begin
    p0_dirrpl_enq_cnt_rmw_pipe_nxt.qid          = dirrpl_fifo_pop_data.qid ;
  end
  p0_dirrpl_enq_cnt_rmw_pipe_nxt.data           = { $bits ( lsp_dirrpl_enq_cnt_t ) { 1'b0 } } ;       // Unused - cfg write done elsewhere
end // always

//-------------------------------------------------------------------------------------------------
// Manage storage for dirrpl enqueue count
hqm_AW_rmw_mem_4pipe #(
          .DEPTH                ( HQM_LSP_ARCH_NUM_LB_QID )                     // Orig ORD qid
        , .WIDTH                ( HQM_LSP_DIRRPL_ENQ_CNT_MEM_WIDTH )
) i_dir_replay_cnt_pipe (
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .status               ( dirrpl_enq_cnt_rmw_pipe_status )

        // cmd input
        , .p0_hold              ( p0_dirrpl_ctrl_pipe.hold )
        , .p0_v_nxt             ( p0_dirrpl_ctrl_pipe_v_nxt_gated )
        , .p0_rw_nxt            ( p0_dirrpl_enq_cnt_rmw_pipe_nxt.rw_cmd )
        , .p0_addr_nxt          ( p0_dirrpl_enq_cnt_rmw_pipe_nxt.qid )
        , .p0_write_data_nxt    ( p0_dirrpl_enq_cnt_rmw_pipe_nxt.data )
        , .p0_v_f               ( p0_dirrpl_ctrl_pipe_v_f )
        , .p0_rw_f              ( p0_dirrpl_enq_cnt_rmw_pipe_f_pnc.rw_cmd )     // Unused
        , .p0_addr_f            ( p0_dirrpl_enq_cnt_rmw_pipe_f_pnc.qid )        // Used by blast logic
        , .p0_data_f            ( p0_dirrpl_enq_cnt_rmw_pipe_f_pnc.data )       // Unused

        , .p1_hold              ( p1_dirrpl_ctrl_pipe.hold )
        , .p1_v_f               ( p1_dirrpl_ctrl_pipe_v_f )
        , .p1_rw_f              ( p1_dirrpl_enq_cnt_rmw_pipe_f_pnc.rw_cmd )     // Unused
        , .p1_addr_f            ( p1_dirrpl_enq_cnt_rmw_pipe_f_pnc.qid )        // Used by blast logic and input error rid
        , .p1_data_f            ( p1_dirrpl_enq_cnt_rmw_pipe_f_pnc.data )       // Unused

        , .p2_hold              ( p2_dirrpl_ctrl_pipe.hold )
        , .p2_v_f               ( p2_dirrpl_ctrl_pipe_v_f )
        , .p2_rw_f              ( p2_dirrpl_enq_cnt_rmw_pipe_f.rw_cmd )
        , .p2_addr_f            ( p2_dirrpl_enq_cnt_rmw_pipe_f.qid )
        , .p2_data_f            ( p2_dirrpl_enq_cnt_rmw_pipe_f.data )

        , .p3_hold              ( p3_dirrpl_ctrl_pipe.hold )
        , .p3_bypsel_nxt        ( p2_dirrpl_enq_cnt_upd_v )
        , .p3_bypdata_nxt       ( p2_dirrpl_enq_cnt_upd )
        , .p3_v_f               ( p3_dirrpl_ctrl_pipe_v_f )
        , .p3_rw_f              ( p3_dirrpl_enq_cnt_rmw_pipe_f_nc.rw_cmd )      // Unused
        , .p3_addr_f            ( p3_dirrpl_enq_cnt_rmw_pipe_f_nc.qid )         // Unused
        , .p3_data_f            ( p3_dirrpl_enq_cnt_rmw_pipe_f_nc.data )        // Unused

        // mem intf
        , .mem_write            ( func_qid_dir_replay_count_mem_we )
        , .mem_read             ( func_qid_dir_replay_count_mem_re )
        , .mem_write_addr       ( func_qid_dir_replay_count_mem_waddr )
        , .mem_read_addr        ( func_qid_dir_replay_count_mem_raddr )
        , .mem_write_data       ( func_qid_dir_replay_count_mem_wdata )
        , .mem_read_data        ( func_qid_dir_replay_count_mem_rdata )
    ) ;

hqm_AW_residue_add i_dirrpl_enq_cnt_res_add (
          .a                    ( p2_dirrpl_ctrl_pipe_f.frag_cnt_res )
        , .b                    ( p2_dirrpl_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_dirrpl_enq_cnt_res_pn )
) ;

hqm_AW_residue_sub i_dirrpl_enq_cnt_res_sub (
          .a                    ( 2'h1 )
        , .b                    ( p2_dirrpl_enq_cnt_rmw_pipe_f.data.cnt_res )
        , .r                    ( p2_dirrpl_enq_cnt_res_m1 )
) ;

// Interface supports 13-bit frag_cnt, max possible total count is 13 bits (4K DIR credits), count memory supports 14 bits (1 spare)
assign { p2_dirrpl_enq_cnt_pn_carry , p2_dirrpl_enq_cnt_pn }  = { 1'b0 , p2_dirrpl_enq_cnt_rmw_pipe_f.data.cnt } + { 2'h0 , p2_dirrpl_ctrl_pipe_f.frag_cnt } ;
assign { p2_dirrpl_enq_cnt_m1_borrow , p2_dirrpl_enq_cnt_m1 } = { 1'b0 , p2_dirrpl_enq_cnt_rmw_pipe_f.data.cnt } - 15'h0001 ;

always_comb begin
  p2_dirrpl_enq_cnt_oflow_cond                  = 1'b0 ;
  p2_dirrpl_enq_cnt_uflow_cond                  = 1'b0 ;
  if ( p2_dirrpl_ctrl_pipe_f.sch_v ) begin
    if ( p2_dirrpl_enq_cnt_m1_borrow ) begin
      p2_dirrpl_enq_cnt_upd                     = p2_dirrpl_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_dirrpl_enq_cnt_uflow_cond              = 1'b1 ;
    end
    else begin
      p2_dirrpl_enq_cnt_upd.cnt                 = p2_dirrpl_enq_cnt_m1 ;
      p2_dirrpl_enq_cnt_upd.cnt_res             = p2_dirrpl_enq_cnt_res_m1 ;
    end
  end
  else begin
    if ( p2_dirrpl_enq_cnt_pn_carry ) begin
      p2_dirrpl_enq_cnt_upd                     = p2_dirrpl_enq_cnt_rmw_pipe_f.data ;      // Saturate, no residue error
      p2_dirrpl_enq_cnt_oflow_cond              = 1'b1 ;
    end
    else begin
      p2_dirrpl_enq_cnt_upd.cnt                 = p2_dirrpl_enq_cnt_pn ;
      p2_dirrpl_enq_cnt_upd.cnt_res             = p2_dirrpl_enq_cnt_res_pn ;
    end
  end
end // always

assign p2_dirrpl_enq_cnt_upd_gt0                = | ( p2_dirrpl_enq_cnt_upd.cnt ) ;

assign p0_dirrpl_inp_frag_cnt_res_chk_en        = p0_dirrpl_ctrl_pipe_f.enq_v ;

hqm_AW_residue_check #( .WIDTH ( 13 ) ) i_dirrpl_inp_frag_cnt_res_chk (
          .r                    ( p0_dirrpl_ctrl_pipe_f.frag_cnt_res )
        , .d                    ( p0_dirrpl_ctrl_pipe_f.frag_cnt )
        , .e                    ( p0_dirrpl_inp_frag_cnt_res_chk_en )
        , .err                  ( p0_dirrpl_inp_frag_cnt_res_err_cond )
) ;

assign p2_dirrpl_enq_cnt_res_chk_en             = p2_dirrpl_enq_cnt_upd_v ;

hqm_AW_residue_check #( .WIDTH ( HQM_LSP_DIRRPL_ENQ_CNT_WIDTH ) ) i_dirrpl_enq_cnt_res_chk (
          .r                    ( p3_dirrpl_enq_cnt_f.cnt_res )
        , .d                    ( p3_dirrpl_enq_cnt_f.cnt )
        , .e                    ( p3_dirrpl_enq_cnt_res_chk_en_f )
        , .err                  ( p3_dirrpl_enq_cnt_res_err )
) ;

assign p2_dirrpl_inp_qid_par_chk_en     = p2_dirrpl_enq_cnt_upd_v ;

hqm_AW_parity_check # ( .WIDTH ( HQM_LSP_ARCH_NUM_LB_QIDB2 ) ) i_dirrpl_inp_qid_par_chk (       // Orig ORD qid
          .p                    ( p2_dirrpl_ctrl_pipe_f.qid_p )
        , .d                    ( p2_dirrpl_enq_cnt_rmw_pipe_f.qid )
        , .e                    ( p2_dirrpl_inp_qid_par_chk_en )
        , .odd                  ( 1'b1 )
        , .err                  ( p2_dirrpl_inp_qid_par_err_cond )
) ;

//-------------------------------------------------------------------------------------------------
// Underflow/overflow errors - some are impossible, some may be caused by software/config errors
//

always_comb begin
  // Don't hold error flops - 1-clock pulse to report
  p3_dirrpl_enq_cnt_uflow_err_nxt       = 1'b0 ;
  p3_dirrpl_enq_cnt_oflow_err_nxt       = 1'b0 ;

  p1_dirrpl_inp_frag_cnt_res_err_nxt    = 1'b0 ;
  p3_dirrpl_inp_qid_par_err_nxt         = 1'b0 ;

  p3_dirrpl_enq_cnt_res_chk_en_nxt      = 1'b0 ;
  p3_dirrpl_enq_cnt_nxt                 = p3_dirrpl_enq_cnt_f ;

  if ( p0_dirrpl_ctrl_pipe_v_f & ~ p1_dirrpl_ctrl_pipe.hold ) begin
    p1_dirrpl_inp_frag_cnt_res_err_nxt  = p0_dirrpl_inp_frag_cnt_res_err_cond ;
  end

  if ( p2_dirrpl_ctrl_pipe_v_f & ~ p3_dirrpl_ctrl_pipe.hold ) begin
    p3_dirrpl_enq_cnt_uflow_err_nxt     = p2_dirrpl_ctrl_pipe_f.sch_v & p2_dirrpl_enq_cnt_uflow_cond ;
    p3_dirrpl_enq_cnt_oflow_err_nxt     = p2_dirrpl_ctrl_pipe_f.enq_v & p2_dirrpl_enq_cnt_oflow_cond ;

    p3_dirrpl_inp_qid_par_err_nxt       = p2_dirrpl_inp_qid_par_err_cond ;

    p3_dirrpl_enq_cnt_res_chk_en_nxt    = p2_dirrpl_enq_cnt_res_chk_en ;
    p3_dirrpl_enq_cnt_nxt               = p2_dirrpl_enq_cnt_upd ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p3_dirrpl_enq_cnt_uflow_err_f       <= 1'b0 ;
    p3_dirrpl_enq_cnt_oflow_err_f       <= 1'b0 ;

    p1_dirrpl_inp_frag_cnt_res_err_f    <= 1'b0 ;
    p3_dirrpl_inp_qid_par_err_f         <= 1'b0 ;

    p3_dirrpl_enq_cnt_res_chk_en_f      <= 1'b0 ;
  end
  else begin
    p3_dirrpl_enq_cnt_uflow_err_f       <= p3_dirrpl_enq_cnt_uflow_err_nxt ;
    p3_dirrpl_enq_cnt_oflow_err_f       <= p3_dirrpl_enq_cnt_oflow_err_nxt ;

    p1_dirrpl_inp_frag_cnt_res_err_f    <= p1_dirrpl_inp_frag_cnt_res_err_nxt ;
    p3_dirrpl_inp_qid_par_err_f         <= p3_dirrpl_inp_qid_par_err_nxt ;

    p3_dirrpl_enq_cnt_res_chk_en_f      <= p3_dirrpl_enq_cnt_res_chk_en_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  p3_dirrpl_enq_cnt_f                   <= p3_dirrpl_enq_cnt_nxt ;
end // always

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: DIRRPL p3 qid_v status vector
//-----------------------------------------------------------------------------------------------------
// See comments under DIRENQ regarding scheduling terminology

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin      // Orig ORD qid
    // Bypass update from sch takes precedence over update from p2; sch update will cause subsequent write
    // of latest/correct value of count caused by this scheduling.
    // enq updates from upper pipe must be supressed from "enabling" if they were blasted by newer scheduling.
    p3_dirrpl_sch_hit[i]                = p3_dirrpl_sch_start & ( p3_dirrpl_sch_start_qid == i ) ;
    p3_dirrpl_p2_enq_hit[i]             = p3_dirrpl_ctrl_pipe.en & ( p2_dirrpl_ctrl_pipe_f.enq_v | p2_dirrpl_ctrl_pipe_f.sch_v ) &
                                          ( p2_dirrpl_enq_cnt_rmw_pipe_f.qid == i ) & ~ p2_dirrpl_ctrl_pipe_f.blast_enq ;
  end // for
end // always

// For each dirrpl qid maintain state for "qid has data" (qid_v)
// Update (set to 0 or 1) when enq count is updated, reset when that qid is selected to be scheduled.
// Should be cleared as part of a successful vas reset drain
always_comb begin
  p3_dirrpl_arb_stat_nxt                = p3_dirrpl_arb_stat_f ;
  if ( p3_dirrpl_sch_start | p3_dirrpl_ctrl_pipe.en ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin    // Orig ORD qid
      if ( p3_dirrpl_sch_hit [i] ) begin
        p3_dirrpl_arb_stat_nxt[i].qid_v         = 1'b0 ;
      end
      else if ( p3_dirrpl_p2_enq_hit [i] ) begin
        p3_dirrpl_arb_stat_nxt[i].qid_v         = p2_dirrpl_enq_cnt_upd_gt0 ;
      end
    end // for i
  end // if
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin    // Orig ORD qid
      p3_dirrpl_arb_stat_f[i].qid_v     <= 1'b0 ;
    end
  end
  else begin
    for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin    // Orig ORD qid
      p3_dirrpl_arb_stat_f[i]           <= p3_dirrpl_arb_stat_nxt[i] ;
    end // for i
  end // else rst_n

end // always

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_QID ; i = i + 1 ) begin
    p3_dirrpl_arb_reqs [i]              = p3_dirrpl_arb_stat_f[i].qid_v ;
    cfg_qid_dir_replay_v_status [i]     = p3_dirrpl_arb_stat_f[i].qid_v ;
  end // for i
end // always

hqm_AW_rr_arb # ( .NUM_REQS ( HQM_NUM_LB_QID ) ) i_dirrpl_arb (         // Orig ORD qid
          .clk                  ( hqm_gated_clk )
        , .rst_n                ( hqm_gated_rst_n )
        , .reqs                 ( p3_dirrpl_arb_reqs )
        , .update               ( p3_dirrpl_arb_update )
        , .winner_v             ( p3_dirrpl_arb_winner_pre_v )
        , .winner               ( p3_dirrpl_arb_winner )
) ;
assign p3_dirrpl_arb_winner_v           = p3_dirrpl_arb_winner_pre_v & ~ cause_pipe_idle ;

hqm_AW_parity_gen #( .WIDTH( HQM_NUM_LB_QIDB2 ) ) i_dirrpl_sch_qid_par_gen (    // Orig ORD qid
          .d            ( p3_dirrpl_arb_winner )
        , .odd          ( 1'b1 )
        , .p            ( p3_dirrpl_arb_winner_gp )
) ;

always_comb begin
  p3_dirrpl_sch_req                                     = p3_dirrpl_arb_winner_v & ~ rpl_dir_dp_fifo_hold & ~ p4_dirrpl_sch_hold ;
  p3_dirrpl_sch_stall_smon                              = p3_dirrpl_arb_winner_v &   rpl_dir_dp_fifo_hold & ~ p4_dirrpl_sch_hold ;      // For smon only
  p3_dirrpl_sch_req_qid.qid                             = { HQM_LSP_ARCH_NUM_LB_QIDB2 { 1'b0 } } ;
  p3_dirrpl_sch_req_qid.qid [HQM_NUM_LB_QIDB2-1:0]      = p3_dirrpl_arb_winner ;
  p3_dirrpl_sch_req_qid.qid_p                           = p3_dirrpl_arb_winner_gp ;
end // always

assign p3_dirrpl_arb_update             = p3_dirrpl_sch_req ;

assign p3_dirrpl_sch_start              = p3_dirrpl_sch_req ;
assign p3_dirrpl_sch_start_qid          = p3_dirrpl_sch_req_qid.qid ;

assign p4_dirrpl_sch_hold               = p4_dirrpl_sch_v_f & ~ dirrpl_input_arb_sch ;
assign p4_dirrpl_sch_v_nxt              = p3_dirrpl_sch_req | p4_dirrpl_sch_hold ;

always_comb begin
  p4_dirrpl_sch_qid_nxt                 = p4_dirrpl_sch_qid_f ;
  if ( p3_dirrpl_sch_req & ~ p4_dirrpl_sch_hold )
    p4_dirrpl_sch_qid_nxt               = p3_dirrpl_sch_req_qid ;
end //always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    p4_dirrpl_sch_v_f                   <= 1'b0 ;
  end
  else begin
    p4_dirrpl_sch_v_f                   <= p4_dirrpl_sch_v_nxt ;
  end
end // always
always_ff @ ( posedge hqm_gated_clk ) begin
  p4_dirrpl_sch_qid_f                   <= p4_dirrpl_sch_qid_nxt ;
end // always

//-------------------------------------------------------------------------------------------------
// Output FIFO (DB) - for static timing isolation
assign rpl_dir_dp_fifo_push             = p3_dirrpl_sch_req ;                   // sch_req already has afull in equation
assign rpl_dir_dp_fifo_push_data.parity = p3_dirrpl_sch_req_qid.qid_p ^ cfg_error_inject_f [ 15 ] ;
assign rpl_dir_dp_fifo_push_data.qid    = p3_dirrpl_sch_req_qid.qid ;

assign rpl_dir_dp_db_in_valid           = rpl_dir_dp_fifo_push ;
assign rpl_dir_dp_db_in_data            = rpl_dir_dp_fifo_push_data ;
assign rpl_dir_dp_fifo_afull            = ~ rpl_dir_dp_db_in_ready ;
assign rpl_dir_dp_fifo_empty            = rpl_dir_dp_tx_sync_idle ;
assign rpl_dir_dp_fifo_hold             = rpl_dir_dp_fifo_afull | ( cfg_control_single_out_dirrpl & ~ rpl_dir_dp_fifo_empty ) ;

// rpl_dir_dp_db_in_data goes to i_hqm_AW_tx_sync_rpl_dir_dp

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: Sidecar logic
//*****************************************************************************************************
//*****************************************************************************************************

//-------------------------------------------------------------------------------------------------

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
    p0_lba_slist_cq_v [i]       = | ( p0_lba_slist_v_f [ ( i * HQM_QID_PER_CQ ) +: HQM_QID_PER_CQ ] ) ;
    p0_lba_rlist_cq_v [i]       = | ( p0_lba_rlist_v_f [ ( i * HQM_QID_PER_CQ ) +: HQM_QID_PER_CQ ] ) ;
  end // for i
end // always

assign cfg_qid_atq_sch_v_nxt            = | cfg_qid_atq_sch_v_status ;
assign cfg_qid_dir_replay_v_nxt         = | cfg_qid_dir_replay_v_status ;
assign cfg_qid_ldb_replay_v_nxt         = | cfg_qid_ldb_replay_v_status ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_qid_atq_sch_v_f                 <= 1'b0 ;
    cfg_qid_dir_replay_v_f              <= 1'b0 ;
    cfg_qid_ldb_replay_v_f              <= 1'b0 ;
    cfg_lba_cq_arb_reqs_f               <= 1'b0 ;
    cfg_direnq_arb_reqs_f               <= 1'b0 ;
    cfg_atq_arb_winner_v_f              <= 1'b0 ;
  end
  else begin
    cfg_qid_atq_sch_v_f                 <= cfg_qid_atq_sch_v_nxt ;
    cfg_qid_dir_replay_v_f              <= cfg_qid_dir_replay_v_nxt ;
    cfg_qid_ldb_replay_v_f              <= cfg_qid_ldb_replay_v_nxt ;
    cfg_lba_cq_arb_reqs_f               <= cfg_lba_cq_arb_reqs_nxt ;
    cfg_direnq_arb_reqs_f               <= cfg_direnq_arb_reqs_nxt ;
    cfg_atq_arb_winner_v_f              <= cfg_atq_arb_winner_v_nxt ;
  end
end // always


always_comb begin
  cfg_unit_idle_nxt             = cfg_unit_idle_f ;
  lsp_unit_pipeidle             = cfg_unit_idle_f.pipe_idle ;
  lsp_reset_done                = ~ ( hqm_gated_rst_n_active ) ;


reset_pf_counter_nxt = reset_pf_counter_f ;
reset_pf_active_nxt = reset_pf_active_f ;
reset_pf_done_nxt = reset_pf_done_f ;
hw_init_done_nxt = hw_init_done_f ;





  pf_dir_enq_cnt_mem_we                                 = 1'b0 ;
  pf_dir_enq_cnt_mem_waddr                              = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
  pf_dir_enq_cnt_mem_wdata                              = '0 ;
  pf_dir_enq_cnt_mem_re                                 = 1'b0 ;                                        // Unused
  pf_dir_enq_cnt_mem_raddr                              = '0 ;                                          // Unused
  pf_dir_enq_cnt_mem_rdata_nc                           = pf_dir_enq_cnt_mem_rdata ;                    // Unused

  pf_dir_tok_cnt_mem_we                                 = 1'b0 ;
  pf_dir_tok_cnt_mem_waddr                              = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0] ;
  pf_dir_tok_cnt_mem_wdata_struct.cnt_res               = 2'h0 ;
  pf_dir_tok_cnt_mem_wdata_struct.cnt                   = '0 ;
  pf_dir_tok_cnt_mem_wdata                              = pf_dir_tok_cnt_mem_wdata_struct ;
  pf_dir_tok_cnt_mem_re                                 = 1'b0 ;                                        // Unused
  pf_dir_tok_cnt_mem_raddr                              = '0 ;                                          // Unused
  pf_dir_tok_cnt_mem_rdata_nc                           = pf_dir_tok_cnt_mem_rdata ;                    // Unused

  pf_dir_tok_lim_mem_we                                 = 1'b0 ;
  pf_dir_tok_lim_mem_addr                               = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0] ;
  pf_dir_tok_lim_mem_wdata_struct.lim_p                 = 1'b1 ;
  pf_dir_tok_lim_mem_wdata_struct.spare                 = 2'h0 ;
  pf_dir_tok_lim_mem_wdata_struct.disab_opt             = 1'b0 ;
  pf_dir_tok_lim_mem_wdata_struct.lim_sel               = 4'h0 ;
  pf_dir_tok_lim_mem_wdata                              = pf_dir_tok_lim_mem_wdata_struct ;
  pf_dir_tok_lim_mem_re                                 = 1'b0 ;                                        // Unused
  pf_dir_tok_lim_mem_rdata_nc                           = pf_dir_tok_lim_mem_rdata ;                    // Unused

  pf_enq_nalb_fifo_mem_we                               = 1'b0 ;                                        // Unused
  pf_enq_nalb_fifo_mem_waddr                            = '0 ;                                          // Unused
  pf_enq_nalb_fifo_mem_wdata                            = '0 ;                                          // Unused
  pf_enq_nalb_fifo_mem_re                               = 1'b0 ;                                        // Unused
  pf_enq_nalb_fifo_mem_raddr                            = '0 ;                                          // Unused
  pf_enq_nalb_fifo_mem_rdata_nc                         = pf_enq_nalb_fifo_mem_rdata ;                  // Unused

  pf_uno_atm_cmp_fifo_mem_we                            = 1'b0 ;                                        // Unused
  pf_uno_atm_cmp_fifo_mem_waddr                         = '0 ;                                          // Unused
  pf_uno_atm_cmp_fifo_mem_wdata                         = '0 ;                                          // Unused
  pf_uno_atm_cmp_fifo_mem_re                            = 1'b0 ;                                        // Unused
  pf_uno_atm_cmp_fifo_mem_raddr                         = '0 ;                                          // Unused
  pf_uno_atm_cmp_fifo_mem_rdata_nc                      = pf_uno_atm_cmp_fifo_mem_rdata ;               // Unused

  pf_nalb_cmp_fifo_mem_we                               = 1'b0 ;                                        // Unused
  pf_nalb_cmp_fifo_mem_waddr                            = '0 ;                                          // Unused
  pf_nalb_cmp_fifo_mem_wdata                            = '0 ;                                          // Unused
  pf_nalb_cmp_fifo_mem_re                               = 1'b0 ;                                        // Unused
  pf_nalb_cmp_fifo_mem_raddr                            = '0 ;                                          // Unused
  pf_nalb_cmp_fifo_mem_rdata_nc                         = pf_nalb_cmp_fifo_mem_rdata ;                  // Unused

  pf_atm_cmp_fifo_mem_we                                = 1'b0 ;                                        // Unused
  pf_atm_cmp_fifo_mem_waddr                             = '0 ;                                          // Unused
  pf_atm_cmp_fifo_mem_wdata                             = '0 ;                                          // Unused
  pf_atm_cmp_fifo_mem_re                                = 1'b0 ;                                        // Unused
  pf_atm_cmp_fifo_mem_raddr                             = '0 ;                                          // Unused
  pf_atm_cmp_fifo_mem_rdata_nc                          = pf_atm_cmp_fifo_mem_rdata ;                   // Unused

  pf_ldb_token_rtn_fifo_mem_we                          = 1'b0 ;                                        // Unused
  pf_ldb_token_rtn_fifo_mem_waddr                       = '0 ;                                          // Unused
  pf_ldb_token_rtn_fifo_mem_wdata                       = '0 ;                                          // Unused
  pf_ldb_token_rtn_fifo_mem_re                          = 1'b0 ;                                        // Unused
  pf_ldb_token_rtn_fifo_mem_raddr                       = '0 ;                                          // Unused
  pf_ldb_token_rtn_fifo_mem_rdata_nc                    = pf_ldb_token_rtn_fifo_mem_rdata ;             // Unused

  pf_nalb_sel_nalb_fifo_mem_we                          = 1'b0 ;                                        // Unused
  pf_nalb_sel_nalb_fifo_mem_waddr                       = '0 ;                                          // Unused
  pf_nalb_sel_nalb_fifo_mem_wdata                       = '0 ;                                          // Unused
  pf_nalb_sel_nalb_fifo_mem_re                          = 1'b0 ;                                        // Unused
  pf_nalb_sel_nalb_fifo_mem_raddr                       = '0 ;                                          // Unused
  pf_nalb_sel_nalb_fifo_mem_rdata_nc                    = pf_nalb_sel_nalb_fifo_mem_rdata ;             // Unused

  pf_cfg_cq2priov_odd_mem_we                            = 1'b0 ;
  pf_cfg_cq2priov_odd_mem_addr                          = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2priov_odd_mem_wdata                         = 33'h100000000 ;                       // Must match initial values in RDL and pf reset
  pf_cfg_cq2priov_odd_mem_re                            = 1'b0 ;                                // Unused
  pf_cfg_cq2priov_odd_mem_rdata_nc                      = pf_cfg_cq2priov_odd_mem_rdata ;       // Unused

  pf_cfg_cq2priov_mem_we                                = 1'b0 ;
  pf_cfg_cq2priov_mem_addr                              = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2priov_mem_wdata                             = 33'h100000000 ;                       // Must match initial values in RDL and pf reset
  pf_cfg_cq2priov_mem_re                                = 1'b0 ;                                // Unused
  pf_cfg_cq2priov_mem_rdata_nc                          = pf_cfg_cq2priov_mem_rdata ;           // Unused

  pf_cfg_cq2qid_0_odd_mem_we                            = 1'b0 ;
  pf_cfg_cq2qid_0_odd_mem_addr                          = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2qid_0_odd_mem_wdata                         = 29'h10000000 ;                        // Must match initial values in RDL and pf reset
  pf_cfg_cq2qid_0_odd_mem_re                            = 1'b0 ;                                // Unused
  pf_cfg_cq2qid_0_odd_mem_rdata_nc                      = pf_cfg_cq2qid_0_odd_mem_rdata ;       // Unused

  pf_cfg_cq2qid_0_mem_we                                = 1'b0 ;
  pf_cfg_cq2qid_0_mem_addr                              = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2qid_0_mem_wdata                             = 29'h10000000 ;                        // Must match initial values in RDL and pf reset
  pf_cfg_cq2qid_0_mem_re                                = 1'b0 ;                                // Unused
  pf_cfg_cq2qid_0_mem_rdata_nc                          = pf_cfg_cq2qid_0_mem_rdata ;           // Unused

  pf_cfg_cq2qid_1_odd_mem_we                            = 1'b0 ;
  pf_cfg_cq2qid_1_odd_mem_addr                          = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2qid_1_odd_mem_wdata                         = 29'h10000000 ;                        // Must match initial values in RDL and pf reset
  pf_cfg_cq2qid_1_odd_mem_re                            = 1'b0 ;                                // Unused
  pf_cfg_cq2qid_1_odd_mem_rdata_nc                      = pf_cfg_cq2qid_1_odd_mem_rdata ;       // Unused

  pf_cfg_cq2qid_1_mem_we                                = 1'b0 ;
  pf_cfg_cq2qid_1_mem_addr                              = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_PCQB2-1:0] ;
  pf_cfg_cq2qid_1_mem_wdata                             = 29'h10000000 ;                        // Must match initial values in RDL and pf reset
  pf_cfg_cq2qid_1_mem_re                                = 1'b0 ;                                // Unused
  pf_cfg_cq2qid_1_mem_rdata_nc                          = pf_cfg_cq2qid_1_mem_rdata ;           // Unused

  pf_qid_ldb_enqueue_count_mem_we                       = 1'b0 ;
  pf_qid_ldb_enqueue_count_mem_waddr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_ldb_enqueue_count_mem_wdata                    = '0 ;
  pf_qid_ldb_enqueue_count_mem_re                       = 1'b0 ;                                // Unused
  pf_qid_ldb_enqueue_count_mem_raddr                    = '0 ;                                  // Unused
  pf_qid_ldb_enqueue_count_mem_rdata_nc                 = pf_qid_ldb_enqueue_count_mem_rdata ;  // Unused

  pf_qid_ldb_inflight_count_mem_we                      = 1'b0 ;
  pf_qid_ldb_inflight_count_mem_waddr                   = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_ldb_inflight_count_mem_wdata_struct.cnt_res    = 2'h0 ;
  pf_qid_ldb_inflight_count_mem_wdata_struct.cnt        = '0 ;
  pf_qid_ldb_inflight_count_mem_wdata                   = pf_qid_ldb_inflight_count_mem_wdata_struct ;
  pf_qid_ldb_inflight_count_mem_re                      = 1'b0 ;                                        // Unused
  pf_qid_ldb_inflight_count_mem_raddr                   = '0 ;                                          // Unused
  pf_qid_ldb_inflight_count_mem_rdata_nc                = pf_qid_ldb_inflight_count_mem_rdata ;         // Unused

  pf_cfg_qid_ldb_inflight_limit_mem_we                  = 1'b0 ;
  pf_cfg_qid_ldb_inflight_limit_mem_addr                = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_qid_ldb_inflight_limit_mem_wdata_struct.lim_p  = 1'b1 ;
  pf_cfg_qid_ldb_inflight_limit_mem_wdata_struct.lim    = '0 ;
  pf_cfg_qid_ldb_inflight_limit_mem_wdata               = pf_cfg_qid_ldb_inflight_limit_mem_wdata_struct ;
  pf_cfg_qid_ldb_inflight_limit_mem_re                  = 1'b0 ;                                         // Unused
  pf_cfg_qid_ldb_inflight_limit_mem_rdata_nc            = pf_cfg_qid_ldb_inflight_limit_mem_rdata ;      // Unused

  pf_cfg_qid_ldb_qid2cqidix_mem_we                      = 1'b0 ;
  pf_cfg_qid_ldb_qid2cqidix_mem_addr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_qid_ldb_qid2cqidix_mem_wdata                   = { 16'hffff , 512'h0 } ;
  pf_cfg_qid_ldb_qid2cqidix_mem_re                      = 1'b0 ;                                        // Unused
  pf_cfg_qid_ldb_qid2cqidix_mem_rdata_nc                = pf_cfg_qid_ldb_qid2cqidix_mem_rdata ;         // Unused

  pf_cfg_qid_ldb_qid2cqidix2_mem_we                     = 1'b0 ;
  pf_cfg_qid_ldb_qid2cqidix2_mem_addr                   = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_qid_ldb_qid2cqidix2_mem_wdata                  = { 16'hffff , 512'h0 } ;
  pf_cfg_qid_ldb_qid2cqidix2_mem_re                     = 1'b0 ;                                        // Unused
  pf_cfg_qid_ldb_qid2cqidix2_mem_rdata_nc               = pf_cfg_qid_ldb_qid2cqidix2_mem_rdata ;        // Unused

  pf_cq_ldb_token_count_mem_we                          = 1'b0 ;
  pf_cq_ldb_token_count_mem_waddr                       = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cq_ldb_token_count_mem_wdata                       = '0 ;
  pf_cq_ldb_token_count_mem_re                          = 1'b0 ;                                        // Unused
  pf_cq_ldb_token_count_mem_raddr                       = '0 ;                                          // Unused
  pf_cq_ldb_token_count_mem_rdata_nc                    = pf_cq_ldb_token_count_mem_rdata ;             // Unused

  pf_cfg_cq_ldb_token_depth_select_mem_we               = 1'b0 ;
  pf_cfg_cq_ldb_token_depth_select_mem_addr             = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cfg_cq_ldb_token_depth_select_mem_wdata_struct.lim_p      = 1'b1 ;
  pf_cfg_cq_ldb_token_depth_select_mem_wdata_struct.lim_sel    = 4'h0 ;                 // most restrictive, must be configured
  pf_cfg_cq_ldb_token_depth_select_mem_wdata            = pf_cfg_cq_ldb_token_depth_select_mem_wdata_struct ;
  pf_cfg_cq_ldb_token_depth_select_mem_re               = 1'b0 ;                                        // Unused
  pf_cfg_cq_ldb_token_depth_select_mem_rdata_nc         = pf_cfg_cq_ldb_token_depth_select_mem_rdata ;  // Unused

  pf_cq_ldb_inflight_count_mem_we                       = 1'b0 ;
  pf_cq_ldb_inflight_count_mem_waddr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cq_ldb_inflight_count_mem_wdata_struct.cnt_res     = 2'h0 ;
  pf_cq_ldb_inflight_count_mem_wdata_struct.cnt         = '0 ;
  pf_cq_ldb_inflight_count_mem_wdata                    = pf_cq_ldb_inflight_count_mem_wdata_struct ;
  pf_cq_ldb_inflight_count_mem_re                       = 1'b0 ;                                        // Unused
  pf_cq_ldb_inflight_count_mem_raddr                    = '0 ;                                          // Unused
  pf_cq_ldb_inflight_count_mem_rdata_nc                 = pf_cq_ldb_inflight_count_mem_rdata ;          // Unused

  pf_cfg_cq_ldb_inflight_limit_mem_we                   = 1'b0 ;
  pf_cfg_cq_ldb_inflight_limit_mem_addr                 = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cfg_cq_ldb_inflight_limit_mem_wdata_struct.lim_p   = 1'b1 ;
  pf_cfg_cq_ldb_inflight_limit_mem_wdata_struct.lim     = '0 ;
  pf_cfg_cq_ldb_inflight_limit_mem_wdata                = pf_cfg_cq_ldb_inflight_limit_mem_wdata_struct ;
  pf_cfg_cq_ldb_inflight_limit_mem_re                   = 1'b0 ;                                        // Unused
  pf_cfg_cq_ldb_inflight_limit_mem_rdata_nc             = pf_cfg_cq_ldb_inflight_limit_mem_rdata ;      // Unused

  pf_cfg_cq_ldb_inflight_threshold_mem_we                       = 1'b0 ;
  pf_cfg_cq_ldb_inflight_threshold_mem_addr                     = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cfg_cq_ldb_inflight_threshold_mem_wdata_struct.thr_p       = 1'b1 ;
  pf_cfg_cq_ldb_inflight_threshold_mem_wdata_struct.thr         = '0 ;
  pf_cfg_cq_ldb_inflight_threshold_mem_wdata                    = pf_cfg_cq_ldb_inflight_threshold_mem_wdata_struct ;
  pf_cfg_cq_ldb_inflight_threshold_mem_re                       = 1'b0 ;                                        // Unused
  pf_cfg_cq_ldb_inflight_threshold_mem_rdata_nc                 = pf_cfg_cq_ldb_inflight_threshold_mem_rdata ;  // Unused

  pf_cq_nalb_pri_arbindex_mem_we                        = 1'b0 ;
  pf_cq_nalb_pri_arbindex_mem_waddr                     = reset_pf_counter_f [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0] ;
  pf_cq_nalb_pri_arbindex_mem_wdata_struct.counts_odd   = { 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3 } ;          // If the config default changes this should be changed too
  pf_cq_nalb_pri_arbindex_mem_wdata_struct.indexes_odd  = '0 ;
  pf_cq_nalb_pri_arbindex_mem_wdata_struct.counts_even  = { 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3 } ;          // If the config default changes this should be changed too
  pf_cq_nalb_pri_arbindex_mem_wdata_struct.indexes_even = '0 ;
  pf_cq_nalb_pri_arbindex_mem_wdata                     = pf_cq_nalb_pri_arbindex_mem_wdata_struct ;
  pf_cq_nalb_pri_arbindex_mem_re                        = 1'b0 ;                                        // Unused
  pf_cq_nalb_pri_arbindex_mem_raddr                     = '0 ;                                          // Unused
  pf_cq_nalb_pri_arbindex_mem_rdata_nc                  = pf_cq_nalb_pri_arbindex_mem_rdata ;           // Unused

  pf_cq_atm_pri_arbindex_mem_we                         = 1'b0 ;
  pf_cq_atm_pri_arbindex_mem_waddr                      = reset_pf_counter_f [(HQM_LSP_ARCH_NUM_LB_CQB2-1)-1:0] ;
  pf_cq_atm_pri_arbindex_mem_wdata_struct.counts_odd    = { 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3 } ;          // If the config default changes this should be changed too
  pf_cq_atm_pri_arbindex_mem_wdata_struct.indexes_odd   = '0 ;
  pf_cq_atm_pri_arbindex_mem_wdata_struct.counts_even   = { 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3, 3'h3 } ;          // If the config default changes this should be changed too
  pf_cq_atm_pri_arbindex_mem_wdata_struct.indexes_even  = '0 ;
  pf_cq_atm_pri_arbindex_mem_wdata                      = pf_cq_atm_pri_arbindex_mem_wdata_struct ;
  pf_cq_atm_pri_arbindex_mem_re                         = 1'b0 ;                                        // Unused
  pf_cq_atm_pri_arbindex_mem_raddr                      = '0 ;                                          // Unused
  pf_cq_atm_pri_arbindex_mem_rdata_nc                   = pf_cq_atm_pri_arbindex_mem_rdata ;            // Unused

  pf_qid_atq_enqueue_count_mem_we                       = 1'b0 ;
  pf_qid_atq_enqueue_count_mem_waddr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_atq_enqueue_count_mem_wdata                    = '0 ;
  pf_qid_atq_enqueue_count_mem_re                       = 1'b0 ;                                        // Unused
  pf_qid_atq_enqueue_count_mem_raddr                    = '0 ;                                          // Unused
  pf_qid_atq_enqueue_count_mem_rdata_nc                 = pf_qid_atq_enqueue_count_mem_rdata ;          // Unused

  pf_qid_aqed_active_count_mem_we                       = 1'b0 ;
  pf_qid_aqed_active_count_mem_waddr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_aqed_active_count_mem_wdata                    = '0 ;
  pf_qid_aqed_active_count_mem_re                       = 1'b0 ;                                        // Unused
  pf_qid_aqed_active_count_mem_raddr                    = '0 ;                                          // Unused
  pf_qid_aqed_active_count_mem_rdata_nc                 = pf_qid_aqed_active_count_mem_rdata ;          // Unused

  pf_cfg_qid_aqed_active_limit_mem_we                   = 1'b0 ;
  pf_cfg_qid_aqed_active_limit_mem_addr                 = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_qid_aqed_active_limit_mem_wdata_struct.lim_p   = 1'b1 ;
  pf_cfg_qid_aqed_active_limit_mem_wdata_struct.lim     = '0 ;
  pf_cfg_qid_aqed_active_limit_mem_wdata                = pf_cfg_qid_aqed_active_limit_mem_wdata_struct ;
  pf_cfg_qid_aqed_active_limit_mem_re                   = 1'b0 ;                                        // Unused
  pf_cfg_qid_aqed_active_limit_mem_rdata_nc             = pf_cfg_qid_aqed_active_limit_mem_rdata ;      // Unused

  pf_qid_ldb_replay_count_mem_we                        = 1'b0 ;
  pf_qid_ldb_replay_count_mem_waddr                     = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_ldb_replay_count_mem_wdata                     = '0 ;      
  pf_qid_ldb_replay_count_mem_re                        = 1'b0 ;                                        // Unused
  pf_qid_ldb_replay_count_mem_raddr                     = '0 ;                                          // Unused
  pf_qid_ldb_replay_count_mem_rdata_nc                  = pf_qid_ldb_replay_count_mem_rdata ;           // Unused

  pf_qid_dir_replay_count_mem_we                        = 1'b0 ;
  pf_qid_dir_replay_count_mem_waddr                     = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_dir_replay_count_mem_wdata                     = '0 ;
  pf_qid_dir_replay_count_mem_re                        = 1'b0 ;                                        // Unused
  pf_qid_dir_replay_count_mem_raddr                     = '0 ;                                          // Unused
  pf_qid_dir_replay_count_mem_rdata_nc                  = pf_qid_dir_replay_count_mem_rdata ;           // Unused

  pf_qid_naldb_tot_enq_cnt_mem_we                       = 1'b0 ;
  pf_qid_naldb_tot_enq_cnt_mem_waddr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_naldb_tot_enq_cnt_mem_wdata                    = '0 ;          // Includes residue
  pf_qid_naldb_tot_enq_cnt_mem_re                       = 1'b0 ;                                        // Unused
  pf_qid_naldb_tot_enq_cnt_mem_raddr                    = '0 ;                                          // Unused
  pf_qid_naldb_tot_enq_cnt_mem_rdata_nc                 = pf_qid_naldb_tot_enq_cnt_mem_rdata ;          // Unused

  pf_qid_atm_tot_enq_cnt_mem_we                         = 1'b0 ;
  pf_qid_atm_tot_enq_cnt_mem_waddr                      = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_atm_tot_enq_cnt_mem_wdata                      = '0 ;          // Includes residue
  pf_qid_atm_tot_enq_cnt_mem_re                         = 1'b0 ;                                        // Unused
  pf_qid_atm_tot_enq_cnt_mem_raddr                      = '0 ;                                          // Unused
  pf_qid_atm_tot_enq_cnt_mem_rdata_nc                   = pf_qid_atm_tot_enq_cnt_mem_rdata ;            // Unused

  pf_cq_ldb_tot_sch_cnt_mem_we                          = 1'b0 ;
  pf_cq_ldb_tot_sch_cnt_mem_waddr                       = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cq_ldb_tot_sch_cnt_mem_wdata                       = '0 ;          // Includes residue
  pf_cq_ldb_tot_sch_cnt_mem_re                          = 1'b0 ;                                        // Unused
  pf_cq_ldb_tot_sch_cnt_mem_raddr                       = '0 ;                                          // Unused
  pf_cq_ldb_tot_sch_cnt_mem_rdata_nc                    = pf_cq_ldb_tot_sch_cnt_mem_rdata ;             // Unused

  pf_qid_dir_tot_enq_cnt_mem_we                         = 1'b0 ;
  pf_qid_dir_tot_enq_cnt_mem_waddr                      = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
  pf_qid_dir_tot_enq_cnt_mem_wdata                      = '0 ;          // Includes residue
  pf_qid_dir_tot_enq_cnt_mem_re                         = 1'b0 ;                                        // Unused
  pf_qid_dir_tot_enq_cnt_mem_raddr                      = '0 ;                                          // Unused
  pf_qid_dir_tot_enq_cnt_mem_rdata_nc                   = pf_qid_dir_tot_enq_cnt_mem_rdata ;            // Unused

  pf_cq_dir_tot_sch_cnt_mem_we                          = 1'b0 ;
  pf_cq_dir_tot_sch_cnt_mem_waddr                       = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_CQB2-1:0] ;
  pf_cq_dir_tot_sch_cnt_mem_wdata                       = '0 ;          // Includes residue
  pf_cq_dir_tot_sch_cnt_mem_re                          = 1'b0 ;                                        // Unused
  pf_cq_dir_tot_sch_cnt_mem_raddr                       = '0 ;                                          // Unused
  pf_cq_dir_tot_sch_cnt_mem_rdata_nc                    = pf_cq_dir_tot_sch_cnt_mem_rdata ;             // Unused

  pf_qid_naldb_max_depth_mem_we                         = 1'b0 ;
  pf_qid_naldb_max_depth_mem_waddr                      = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_naldb_max_depth_mem_wdata                      = '0 ;
  pf_qid_naldb_max_depth_mem_re                         = 1'b0 ;                                        // Unused
  pf_qid_naldb_max_depth_mem_raddr                      = '0 ;                                          // Unused
  pf_qid_naldb_max_depth_mem_rdata_nc                   = pf_qid_naldb_max_depth_mem_rdata ;            // Unused

  pf_qid_dir_max_depth_mem_we                           = 1'b0;
  pf_qid_dir_max_depth_mem_waddr                        = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
  pf_qid_dir_max_depth_mem_wdata                        = '0 ;
  pf_qid_dir_max_depth_mem_re                           = 1'b0 ;                                        // Unused
  pf_qid_dir_max_depth_mem_raddr                        = '0 ;                                          // Unused
  pf_qid_dir_max_depth_mem_rdata_nc                     = pf_qid_dir_max_depth_mem_rdata ;              // Unused

  pf_chp_lsp_token_rx_sync_fifo_mem_we                  = 1'b0 ;                                        // Unused
  pf_chp_lsp_token_rx_sync_fifo_mem_waddr               = '0 ;                                          // Unused
  pf_chp_lsp_token_rx_sync_fifo_mem_wdata               = '0 ;                                          // Unused
  pf_chp_lsp_token_rx_sync_fifo_mem_re                  = 1'b0 ;                                        // Unused
  pf_chp_lsp_token_rx_sync_fifo_mem_raddr               = '0 ;                                          // Unused
  pf_chp_lsp_token_rx_sync_fifo_mem_rdata_nc            = pf_chp_lsp_token_rx_sync_fifo_mem_rdata ;     // Unused

  pf_chp_lsp_cmp_rx_sync_fifo_mem_we                    = 1'b0 ;                                        // Unused
  pf_chp_lsp_cmp_rx_sync_fifo_mem_waddr                 = '0 ;                                          // Unused
  pf_chp_lsp_cmp_rx_sync_fifo_mem_wdata                 = '0 ;                                          // Unused
  pf_chp_lsp_cmp_rx_sync_fifo_mem_re                    = 1'b0 ;                                        // Unused
  pf_chp_lsp_cmp_rx_sync_fifo_mem_raddr                 = '0 ;                                          // Unused
  pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata_nc              = pf_chp_lsp_cmp_rx_sync_fifo_mem_rdata ;       // Unused

  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_we             = 1'b0 ;                                        // Unused
  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr          = '0 ;                                          // Unused
  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata          = '0 ;                                          // Unused
  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_re             = 1'b0 ;                                        // Unused
  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr          = '0 ;                                          // Unused
  pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata_nc       = pf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata ;        // Unused

  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we                = 1'b0 ;                                        // Unused
  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr             = '0 ;                                          // Unused
  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata             = '0 ;                                          // Unused
  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re                = 1'b0 ;                                        // Unused
  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr             = '0 ;                                          // Unused
  pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata_nc          = pf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata ;   // Unused

  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_we                 = 1'b0 ;                                        // Unused
  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr              = '0 ;                                          // Unused
  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata              = '0 ;                                          // Unused
  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_re                 = 1'b0 ;                                        // Unused
  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr              = '0 ;                                          // Unused
  pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata_nc           = pf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata ;    // Unused

  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we              = 1'b0 ;                                        // Unused
  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr           = '0 ;                                          // Unused
  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata           = '0 ;                                          // Unused
  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re              = 1'b0 ;                                        // Unused
  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr           = '0 ;                                          // Unused
  pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata_nc        = pf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata ;         // Unused

  pf_send_atm_to_cq_rx_sync_fifo_mem_we                 = 1'b0 ;                                        // Unused
  pf_send_atm_to_cq_rx_sync_fifo_mem_waddr              = '0 ;                                          // Unused
  pf_send_atm_to_cq_rx_sync_fifo_mem_wdata              = '0 ;                                          // Unused
  pf_send_atm_to_cq_rx_sync_fifo_mem_re                 = 1'b0 ;                                        // Unused
  pf_send_atm_to_cq_rx_sync_fifo_mem_raddr              = '0 ;                                          // Unused
  pf_send_atm_to_cq_rx_sync_fifo_mem_rdata_nc           = pf_send_atm_to_cq_rx_sync_fifo_mem_rdata ;    // Unused

  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we            = 1'b0 ;                                        // Unused
  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr         = '0 ;                                          // Unused
  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata         = '0 ;                                          // Unused
  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re            = 1'b0 ;                                        // Unused
  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr         = '0 ;                                          // Unused
  pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata_nc      = pf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata ;       // Unused

  pf_cfg_atm_qid_dpth_thrsh_mem_we                      = 1'b0 ;
  pf_cfg_atm_qid_dpth_thrsh_mem_addr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_atm_qid_dpth_thrsh_mem_wdata                   = { 1'b1 , { HQM_LSP_ATQ_QID_DPTH_THRSH_WIDTH { 1'b0 } } } ;    // Zero with good parity
  pf_cfg_atm_qid_dpth_thrsh_mem_re                      = 1'b0 ;                                        // Unused
  pf_cfg_atm_qid_dpth_thrsh_mem_rdata_nc                = pf_cfg_atm_qid_dpth_thrsh_mem_rdata ;         // Unused

  pf_cfg_nalb_qid_dpth_thrsh_mem_we                     = 1'b0 ;
  pf_cfg_nalb_qid_dpth_thrsh_mem_addr                   = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_cfg_nalb_qid_dpth_thrsh_mem_wdata                  = { 1'b1 , { HQM_LSP_LB_QID_DPTH_THRSH_WIDTH { 1'b0 } } } ;     // Zero with good parity
  pf_cfg_nalb_qid_dpth_thrsh_mem_re                     = 1'b0 ;                                        // Unused
  pf_cfg_nalb_qid_dpth_thrsh_mem_rdata_nc               = pf_cfg_nalb_qid_dpth_thrsh_mem_rdata ;        // Unused

  pf_cfg_dir_qid_dpth_thrsh_mem_we                      = 1'b0 ;
  pf_cfg_dir_qid_dpth_thrsh_mem_addr                    = reset_pf_counter_f [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
  pf_cfg_dir_qid_dpth_thrsh_mem_wdata                   = { 1'b1 , { HQM_LSP_DIRENQ_DPTH_THRSH_WIDTH { 1'b0 } } } ;     // Zero with good parity
  pf_cfg_dir_qid_dpth_thrsh_mem_re                      = 1'b0 ;                                        // Unused
  pf_cfg_dir_qid_dpth_thrsh_mem_rdata_nc                = pf_cfg_dir_qid_dpth_thrsh_mem_rdata ;         // Unused

  pf_qid_atm_active_mem_we                              = 1'b0 ;
  pf_qid_atm_active_mem_waddr                           = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
  pf_qid_atm_active_mem_wdata                           = '0 ;                                                          // Zero with good residue
  pf_qid_atm_active_mem_re                              = 1'b0 ;                                        // Unused
  pf_qid_atm_active_mem_raddr                           = '0 ;                                          // Unused
  pf_qid_atm_active_mem_rdata_nc                        = pf_qid_atm_active_mem_rdata ;                 // Unused

  pf_cq_ldb_wu_count_mem_we                             = 1'b0 ;
  pf_cq_ldb_wu_count_mem_waddr                          = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cq_ldb_wu_count_mem_wdata                          = { (2+HQM_LSP_LBWU_CQ_WU_CNT_WIDTH) { 1'b0 } } ;               // Will get linra warning if struct width changes
  pf_cq_ldb_wu_count_mem_re                             = 1'b0 ;                                        // Unused
  pf_cq_ldb_wu_count_mem_raddr                          = '0 ;                                          // Unused
  pf_cq_ldb_wu_count_mem_rdata_nc                       = pf_cq_ldb_wu_count_mem_rdata ;                // Unused

  pf_cfg_cq_ldb_wu_limit_mem_we                         = 1'b0 ;
  pf_cfg_cq_ldb_wu_limit_mem_waddr                      = reset_pf_counter_f [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
  pf_cfg_cq_ldb_wu_limit_mem_wdata                      = { 1'b1 , { (1+HQM_LSP_LBWU_CQ_WU_LIM_WIDTH) { 1'b0 } } } ;    // Will get linra warning if struct width changes
  pf_cfg_cq_ldb_wu_limit_mem_re                         = 1'b0 ;                                        // Unused
  pf_cfg_cq_ldb_wu_limit_mem_raddr                      = '0 ;                                          // Unused
  pf_cfg_cq_ldb_wu_limit_mem_rdata_nc                   = pf_cfg_cq_ldb_wu_limit_mem_rdata ;            // Unused

  pf_qed_lsp_deq_fifo_mem_we                    = 1'b0 ;                                        // Unused
  pf_qed_lsp_deq_fifo_mem_waddr                 = '0 ;                                          // Unused
  pf_qed_lsp_deq_fifo_mem_wdata                 = '0 ;                                          // Unused
  pf_qed_lsp_deq_fifo_mem_re                    = 1'b0 ;                                        // Unused
  pf_qed_lsp_deq_fifo_mem_raddr                 = '0 ;                                          // Unused
  pf_qed_lsp_deq_fifo_mem_rdata_nc              = pf_qed_lsp_deq_fifo_mem_rdata ;               // Unused

  pf_aqed_lsp_deq_fifo_mem_we                   = 1'b0 ;                                        // Unused
  pf_aqed_lsp_deq_fifo_mem_waddr                = '0 ;                                          // Unused
  pf_aqed_lsp_deq_fifo_mem_wdata                = '0 ;                                          // Unused
  pf_aqed_lsp_deq_fifo_mem_re                   = 1'b0 ;                                        // Unused
  pf_aqed_lsp_deq_fifo_mem_raddr                = '0 ;                                          // Unused
  pf_aqed_lsp_deq_fifo_mem_rdata_nc             = pf_aqed_lsp_deq_fifo_mem_rdata ;              // Unused


  cfg_lba_cq_arb_reqs_nxt       = | p0_lba_cq_arb_reqs ;
  cfg_direnq_arb_reqs_nxt       = | p3_direnq_arb_reqs ;

  cfg_lbwu_pipe_idle            = ~ ( | { p1_lbwu_ctrl_pipe_v_f , p2_lbwu_ctrl_pipe_v_f , p3_lbwu_ctrl_pipe_v_f , p4_lbwu_ctrl_pipe_v_f } ) ;

  cfg_unit_idle_nxt.pipe_idle   =       ~ ( | { cfg_pipe_health_valid_1_nxt , cfg_pipe_health_valid_0_nxt } ) ;
  cfg_unit_idle_nxt.unit_idle   =       ( cfg_unit_idle_nxt.pipe_idle
                                        //-------------------------------------------------------
                                        & cfg_lbwu_pipe_idle                            // Can't be in pipe_idle since lbwu pipe is not idled during cfg access
                                        // Input FIFOs/DBs
                                        & dir_tokrtn_fifo_empty                         // dir_tokrtn_db_status_pnc
                                        & ldb_token_rtn_fifo_empty
                                        & uno_atm_cmp_fifo_empty
                                        & nalb_cmp_fifo_empty
                                        & atm_cmp_fifo_empty
                                        & enq_nalb_fifo_empty
                                        & ( enq_atq_db_status_pnc [1:0] == 2'h0 )
                                        & qed_lsp_deq_fifo_empty
                                        & aqed_lsp_deq_fifo_empty
// The following Input rx_sync FIFO idle conditions are included in lsp_unit_idle signal calculated by hqm_AW_module_clock_control,
// so do not need to be included here.
// chp_lsp_token_rx_sync_idle
// chp_lsp_cmp_rx_sync_idle
// rop_lsp_reordercmp_rx_sync_idle
// nalb_lsp_enq_lb_rx_sync_idle
// nalb_lsp_enq_rorply_rx_sync_idle
// dp_lsp_enq_dir_rx_sync_idle
// dp_lsp_enq_rorply_rx_sync_idle
// send_atm_to_cq_rx_sync_idle

// The following interrupt serializer idle conditions are included in lsp_unit_idle signal calculated by hqm_AW_module_clock_control,
// so do not need to be included here.
// ( int_serializer_status_up [1:0] == 2'h0 )
// ( int_serializer_status_down [1:0] == 2'h0 )
                                        //-------------------------------------------------------
                                        // Output FIFOs/DBs
                                        & lsp_dp_sch_dir_tx_sync_idle                   // dir_sel_dp_db_status_nc
                                        & lsp_nalb_sch_unoord_tx_sync_idle              // lsp_nalb_sch_unoord_status_pnc
                                        & atq_sel_ap_tx_sync_idle                       // atq_sel_ap_db_status_pnc
                                        & rpl_ldb_nalb_tx_sync_idle                     // rpl_ldb_nalb_db_status_pnc
                                        & rpl_dir_dp_tx_sync_idle                       // rpl_dir_dp_db_status_pnc

                                        & nalb_sel_nalb_fifo_empty
                                        //-------------------------------------------------------
                                        // Pending scheduling work to do (enqueues), all types of QEs
                                        & ~ cfg_lba_cq_arb_reqs_f                                       // LB work to do (nalb, slist, rlist), not blocked by external dependencies
                                        & ~ cfg_direnq_arb_reqs_f                                       // DIR work to do, not blocked by external dependencies
                                        & ~ cfg_atq_arb_winner_v_f                                      // ATQ work to do, not blocked by external dependencies
                                        & ~ cfg_qid_dir_replay_v_f                                      // ORD REPLAY: "enqueue" DIR, not blocked by external dependencies
                                        & ~ cfg_qid_ldb_replay_v_f                                      // ORD REPLAY: "enqueue" LB, not blocked by external dependencies
                                        & ~ cfg_lba_atm_haswork                                         // LB: atomic - 1-clock gap on input
                                        //-------------------------------------------------------
                                        // Inputs from AQED which can not be backpressured, are not supressed by cause_pipe_idle, and must keep the clocks on
                                        & aqed_intf_idle
                                        //-------------------------------------------------------
                                        // Safety term - if credit count is > 0, something is valid in LSP (or AP - same clock domain so OK)
                                        & p0_lba_atm_credit_count_eq_0
                                        & p0_lba_nalb_credit_count_eq_0
                                        //-------------------------------------------------------
                                        & qed_deq_credit_empty                                          // Must be ready for qed_lsp_deq : no backpressure
                                        & aqed_deq_credit_empty                                         // Must be ready for aqed_lsp_deq : no backpressure
                                        //-------------------------------------------------------
                                        // Pending tokens, all types of QEs.
                                        & ( ~ cfg_control_include_tok_unit_idle |
                                            (
                                                ~ cfg_diag_status_0_f [ HQM_LSP_CFG_DIAG_0_DIR_TOK_V ]          // DIR: token
                                              & ~ cfg_diag_status_0_f [ HQM_LSP_CFG_DIAG_0_LB_TOK_V ]           // LB: token
                                            )
                                          )
                                        //-------------------------------------------------------
                                        // Pending completions.
                                        & ( ~ cfg_control_include_cmp_unit_idle |
                                            ~ cfg_diag_status_0_f [ HQM_LSP_CFG_DIAG_0_LB_CMP_V ]               // LB: completion
                                          )
                                        ) ;

  lsp_unit_idle_local           = ~ ( hqm_gated_rst_n_active ) & cfg_unit_idle_nxt.unit_idle ;

  lsp_unit_idle = ( wire_lsp_unit_idle 
                  & aqed_unit_idle
                  & ap_unit_idle                                  // Strictly speaking not necessary to include since LSP "covers" AP
                  ) ;

  //----------------------------------------------------------------------------------------------
  // PF reset
  reset_pf_count_lt_num_dir_qid         = ( reset_pf_counter_f < HQM_NUM_DIR_QID ) ;
  reset_pf_count_lt_num_dir_cq          = ( reset_pf_counter_f < HQM_NUM_DIR_CQ ) ;
  reset_pf_count_lt_num_lb_qid          = ( reset_pf_counter_f < HQM_NUM_LB_QID ) ;
  reset_pf_count_lt_num_lb_cq           = ( reset_pf_counter_f < HQM_NUM_LB_CQ ) ;
  reset_pf_count_lt_num_lb_pcq          = ( reset_pf_counter_f < HQM_NUM_LB_PCQ ) ;
  if ( hqm_gated_rst_n_start & reset_pf_active_f & ~ hw_init_done_f ) begin
    reset_pf_counter_nxt                = reset_pf_counter_f + 32'h1 ;

    if ( reset_pf_counter_f < HQM_LSP_CFG_RST_PFMAX ) begin
      pf_cfg_cq2priov_odd_mem_we                        = reset_pf_count_lt_num_lb_pcq ;
      pf_cfg_cq2priov_mem_we                            = reset_pf_count_lt_num_lb_pcq ;
      pf_cfg_cq2qid_0_odd_mem_we                        = reset_pf_count_lt_num_lb_pcq ;
      pf_cfg_cq2qid_0_mem_we                            = reset_pf_count_lt_num_lb_pcq ;
      pf_cfg_cq2qid_1_odd_mem_we                        = reset_pf_count_lt_num_lb_pcq ;
      pf_cfg_cq2qid_1_mem_we                            = reset_pf_count_lt_num_lb_pcq ;
      pf_cq_ldb_inflight_count_mem_we                   = reset_pf_count_lt_num_lb_cq ;
      pf_cfg_cq_ldb_inflight_limit_mem_we               = reset_pf_count_lt_num_lb_cq ;
      pf_cfg_cq_ldb_inflight_threshold_mem_we           = reset_pf_count_lt_num_lb_cq ;
      pf_cq_nalb_pri_arbindex_mem_we                    = reset_pf_count_lt_num_lb_pcq ;        // Not config accessible, but need to be initialized by pf reset
      pf_cq_atm_pri_arbindex_mem_we                     = reset_pf_count_lt_num_lb_pcq ;        // Not config accessible, but need to be initialized by pf reset
      pf_cq_ldb_token_count_mem_we                      = reset_pf_count_lt_num_lb_cq ;
      pf_cfg_cq_ldb_token_depth_select_mem_we           = reset_pf_count_lt_num_lb_cq ;
      pf_cq_ldb_tot_sch_cnt_mem_we                      = reset_pf_count_lt_num_lb_cq ;
      pf_cq_ldb_wu_count_mem_we                         = reset_pf_count_lt_num_lb_cq ;
      pf_cfg_cq_ldb_wu_limit_mem_we                     = reset_pf_count_lt_num_lb_cq ;

      pf_dir_tok_cnt_mem_we                             = reset_pf_count_lt_num_dir_cq ;
      pf_cq_dir_tot_sch_cnt_mem_we                      = reset_pf_count_lt_num_dir_cq ;
      pf_dir_tok_lim_mem_we                             = reset_pf_count_lt_num_dir_cq ;

      pf_cfg_qid_ldb_qid2cqidix_mem_we                  = reset_pf_count_lt_num_lb_qid ;
      pf_cfg_qid_ldb_qid2cqidix2_mem_we                 = reset_pf_count_lt_num_lb_qid ;
      pf_qid_ldb_replay_count_mem_we                    = reset_pf_count_lt_num_lb_qid ;
      pf_qid_ldb_enqueue_count_mem_we                   = reset_pf_count_lt_num_lb_qid ;
      pf_qid_aqed_active_count_mem_we                   = reset_pf_count_lt_num_lb_qid ;
      pf_cfg_qid_aqed_active_limit_mem_we               = reset_pf_count_lt_num_lb_qid ;
      pf_qid_ldb_inflight_count_mem_we                  = reset_pf_count_lt_num_lb_qid ;
      pf_cfg_qid_ldb_inflight_limit_mem_we              = reset_pf_count_lt_num_lb_qid ;
      pf_qid_atq_enqueue_count_mem_we                   = reset_pf_count_lt_num_lb_qid ;
      pf_qid_naldb_max_depth_mem_we                     = reset_pf_count_lt_num_lb_qid ;
      pf_qid_atm_tot_enq_cnt_mem_we                     = reset_pf_count_lt_num_lb_qid ;
      pf_qid_naldb_tot_enq_cnt_mem_we                   = reset_pf_count_lt_num_lb_qid ;
      pf_qid_dir_replay_count_mem_we                    = reset_pf_count_lt_num_lb_qid ;        // address = original ORD qid
      pf_cfg_atm_qid_dpth_thrsh_mem_we                  = reset_pf_count_lt_num_lb_qid ;
      pf_cfg_nalb_qid_dpth_thrsh_mem_we                 = reset_pf_count_lt_num_lb_qid ;
      pf_qid_atm_active_mem_we                          = reset_pf_count_lt_num_lb_qid ;

      pf_dir_enq_cnt_mem_we                             = reset_pf_count_lt_num_dir_qid ;
      pf_qid_dir_max_depth_mem_we                       = reset_pf_count_lt_num_dir_qid ;
      pf_qid_dir_tot_enq_cnt_mem_we                     = reset_pf_count_lt_num_dir_qid ;
      pf_cfg_dir_qid_dpth_thrsh_mem_we                  = reset_pf_count_lt_num_dir_qid ;

    end
    else begin
      reset_pf_counter_nxt              = reset_pf_counter_f;
      hw_init_done_nxt                  = 1'b1 ;
    end
  end

   // reset_active is set on reset.
   // reset_active is cleared when hw_init_done_f is set

   if ( reset_pf_active_f ) begin
       if ( hw_init_done_f ) begin
         reset_pf_counter_nxt = 32'd0 ;
         reset_pf_active_nxt = 1'b0 ;
         reset_pf_done_nxt = 1'b1 ;
         hw_init_done_nxt = 1'b0 ;
       end
   end


  // cfg_ignore_pipe_busy is handled by sidecar
  cfg_unit_idle_nxt.cfg_ready                   = ( ( ~ ( | { cfg_pipe_health_valid_1_nxt , cfg_pipe_health_valid_0_nxt } ) ) ) ;

end // always

assign cfg_req_ready            = cfg_unit_idle_f.cfg_ready ;

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: Memories
//*****************************************************************************************************
//*****************************************************************************************************

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: Config / Shared logic
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// Controlled by sidecar logic


//-----------------------------------------------------------------------------------------------------

//----
assign hqm_lsp_target_cfg_unit_idle_reg_nxt                     = cfg_unit_idle_nxt ;
assign cfg_unit_idle_f                                          = hqm_lsp_target_cfg_unit_idle_reg_f ;
//----

// Previously replicated to reduce transitive fanout, may need to do that again.
assign cfg_unit_idle_1_f_pnc                            = cfg_unit_idle_f ;
assign cfg_unit_idle_2_f_pnc                            = cfg_unit_idle_f ;

assign cause_pipe_idle          = cfg_req_idlepipe |
                                  ap_lsp_freeze ;       // Strictly speaking only requirement is to idle lba pipe, but not attempting to optimize

//-----------------------------------------------------------------------------------------------------
// Register for possible future use, currently nothing to connect
assign hqm_lsp_target_cfg_patch_control_reg_v           = 1'b0 ;
assign hqm_lsp_target_cfg_patch_control_reg_nxt         = hqm_lsp_target_cfg_patch_control_reg_f ;

//-----------------------------------------------------------------------------------------------------

//----
assign hqm_lsp_target_cfg_error_inject_reg_v            = 1'b0 ;
assign hqm_lsp_target_cfg_error_inject_reg_nxt          = cfg_error_inject_nxt ;
assign cfg_error_inject_f                               = hqm_lsp_target_cfg_error_inject_reg_f ;
//----

assign cfg_error_inject_nxt                     = cfg_error_inject_f ;

//-----------------------------------------------------------------------------------------------------
// Performance counters
// The intention of performance counters 0, 1, 2, 3 and 5 is that on each clock while the interval counter
// is active exactly one will count.  Count #3 aggregates multiple situations where scheduling can not be considered.
// If a CQ is busy, the has_space and ow vectors must be ignored.
// The accounting is as follows:
// If LSP is not in the "ready_for_work" state, or cause_pipe_idle or pipe holds prevent it from considering scheduling, count #3 (pipe friction)
// else if no CQs have work to do, count #0 (no work)
// else if all CQs with work to do are masked by blasting, count #3 (pipe friction)
// else if all CQs with post-blast work to do are disabled by config, count #0 (no work)
// else if any CQ is cfg enabled, has post-blast work to do, has space and is not busy, count #2 (sched)
// else if any CQ is cfg enabled, has post-blast work, is not busy and does not have space, count #1 (no space)
// else if any CQ is cfg enabled, has post-blast work, is not busy, has space but is overworked, count #7 (overworked)
// else (all cfg enabled CQs with post-blast work are busy), count #5 (pipe friction, will be merged with count #3)
// 
// The accounting assumes there is no agitation active, either in hardware or forced by simulation.

//---------------------------------------
// count #0
assign cfg_ldb_sched_perf_cq_disabled           = p0_lba_sch_state_ready_for_work & ~ cause_pipe_idle &
                                                  ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                  ( | p0_lba_cq_arb_any_has_work ) & ~ ( | ( p0_lba_cq_arb_any_has_work & ~ cfg_cq_ldb_disable_f ) ) ;

assign cfg_ldb_sched_perf_no_work               = p0_lba_sch_state_ready_for_work & ~ cause_pipe_idle &
                                                  ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                  ( ( ~ ( | { p0_lba_slist_v_f , p0_lba_rlist_v_f , p0_lba_nalb_v_f } ) ) | cfg_ldb_sched_perf_cq_disabled ) ;

//---------------------------------------
// count #1
assign cfg_ldb_sched_perf_no_space              = p0_lba_sch_state_ready_for_work & ~ cause_pipe_idle &
                                                  ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                  ( | ( p0_lba_cq_arb_any_has_work & ~ cfg_cq_ldb_disable_f & ~ p0_lba_cq_busy_sch_f & ~ p0_lba_cq_has_space_f ) ) &
                                                  ~ p0_lba_cq_arb_winner_pre_v [0] ;

//---------------------------------------
// count #2
assign cfg_ldb_sched_perf_sched                 = p0_lba_pop_cq [0] ;

//---------------------------------------
// count #3
assign cfg_ldb_sched_perf_pipe_frict_not_wait_work      = ~ p0_lba_sch_state_ready_for_work ;
assign cfg_ldb_sched_perf_pipe_frict_wait_work_hold     = p0_lba_sch_state_ready_for_work &
                                                          ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) ;
assign cfg_ldb_sched_perf_wait_blast                    = p0_lba_sch_state_ready_for_work &
                                                          ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                          ( | { p0_lba_slist_v_f , p0_lba_rlist_v_f , p0_lba_nalb_v_f } ) & ~ ( | p0_lba_cq_arb_any_has_work ) ;
assign cfg_ldb_sched_perf_pipe_frict_cause_pipe_idle    = cause_pipe_idle ;

assign cfg_ldb_sched_perf_3_inc                         =   cfg_ldb_sched_perf_pipe_frict_not_wait_work
                                                          | cfg_ldb_sched_perf_pipe_frict_wait_work_hold
                                                          | cfg_ldb_sched_perf_pipe_frict_cause_pipe_idle
                                                          | cfg_ldb_sched_perf_wait_blast ;

//---------------------------------------
// count #4
assign cfg_ldb_sched_perf_wait_tot_inflight     = ~ p8_lba_tot_if_v_f ;

//---------------------------------------
// count #5
assign cfg_ldb_sched_perf_wait_cq_busy          = p0_lba_sch_state_ready_for_work & ~ cause_pipe_idle &
                                                  ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                  ( | ( p0_lba_cq_arb_any_has_work & ~ cfg_cq_ldb_disable_f & p0_lba_cq_busy_sch_f ) ) &
                                                  ~ p0_lba_cq_arb_winner_pre_v [0] & ~ cfg_ldb_sched_perf_no_space & ~ cfg_ldb_sched_perf_overworked ;

//---------------------------------------
// count #6
assign cfg_ldb_sched_perf_wait_atq_fid_unavail  = p3_atq_fid_inflight_cnt_eq_lim | p3_atq_fid_inflight_cnt_gt_lim ;

//---------------------------------------
// count #7
assign cfg_ldb_sched_perf_overworked            = p0_lba_sch_state_ready_for_work & ~ cause_pipe_idle &
                                                  ~ ( p1_lba_ctrl_pipe.hold | p0_lba_ctrl_pipe_sch_hold_cond ) &
                                                  ( | ( p0_lba_cq_arb_any_has_work & ~ cfg_cq_ldb_disable_f & ~ p0_lba_cq_busy_sch_f & p0_lba_cq_has_space_f & p0_lba_cq_ow_f ) ) &
                                                  ~ p0_lba_cq_arb_winner_pre_v [0] ;


//----
assign hqm_lsp_target_cfg_ldb_sched_perf_control_reg_v          = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_control_reg_nxt        = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f ;


assign hqm_lsp_target_cfg_ldb_sched_perf_7_inc                  = cfg_ldb_sched_perf_overworked ;
assign hqm_lsp_target_cfg_ldb_sched_perf_7_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_7_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_7_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_7_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_7_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_6_inc                  = cfg_ldb_sched_perf_wait_atq_fid_unavail ;
assign hqm_lsp_target_cfg_ldb_sched_perf_6_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_6_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_6_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_6_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_6_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_5_inc                  = cfg_ldb_sched_perf_wait_cq_busy ;
assign hqm_lsp_target_cfg_ldb_sched_perf_5_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_5_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_5_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_5_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_5_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_4_inc                  = cfg_ldb_sched_perf_wait_tot_inflight ;
assign hqm_lsp_target_cfg_ldb_sched_perf_4_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_4_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_4_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_4_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_4_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_3_inc                  = cfg_ldb_sched_perf_3_inc ;
assign hqm_lsp_target_cfg_ldb_sched_perf_3_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_3_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_3_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_3_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_3_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_2_inc                  = cfg_ldb_sched_perf_sched ;
assign hqm_lsp_target_cfg_ldb_sched_perf_2_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_2_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_2_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_2_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_2_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_1_inc                  = cfg_ldb_sched_perf_no_space ;
assign hqm_lsp_target_cfg_ldb_sched_perf_1_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_1_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_1_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_1_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_1_count ;

assign hqm_lsp_target_cfg_ldb_sched_perf_0_inc                  = cfg_ldb_sched_perf_no_work ;
assign hqm_lsp_target_cfg_ldb_sched_perf_0_en                   = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 0 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_0_clr                  = hqm_lsp_target_cfg_ldb_sched_perf_control_reg_f [ 1 ] ;
assign hqm_lsp_target_cfg_ldb_sched_perf_0_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_ldb_sched_perf_0_count_nc             = hqm_lsp_target_cfg_ldb_sched_perf_0_count ;

//-----------------------------------------------------------------------------------------------------
// Global scheduling count across all CQs.

always_comb begin
  hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_nxt           = hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_f ;
  hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_nxt           = hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_f ;
  if ( p2_direnq_tot_sch_cnt_upd_v ) begin      // Whenever one of the per-CQ sched counts is incremented (by n), also increment the total count (by n)
    { hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_nxt , hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_nxt } =
    { hqm_lsp_target_cfg_lsp_perf_dir_sch_count_h_reg_f ,   hqm_lsp_target_cfg_lsp_perf_dir_sch_count_l_reg_f } + { {(64 - HQM_LSP_DIRENQ_TOK_CNT_WIDTH){1'b0}}, p2_direnq_ctrl_pipe_sch_delta } ;   // Wrap
  end
end // always

//----

assign hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_inc            = p7_lba_perf_sch_count_upd_v ;
assign hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_en             = 1'b1 ;
assign hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clr            = 1'b0 ;
assign hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_clrv           = 1'b0 ;
assign hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count_nc       = hqm_lsp_target_cfg_lsp_perf_ldb_sch_count_count ;

//-----------------------------------------------------------------------------------------------------
// Previously explicitly registered

assign hqm_lsp_target_cfg_interface_status_reg_f_nc     = hqm_lsp_target_cfg_interface_status_reg_f ;

assign hqm_lsp_target_cfg_interface_status_reg_nxt      = {   ~ lsp_ap_atm_ready                                                // 31  Internal intf.
                                                            ,   lsp_ap_atm_v                                                    // 30  Internal intf.
                                                            , ~ lsp_nalb_sch_unoord_ready                                       // 29
                                                            ,   lsp_nalb_sch_unoord_v                                           // 28
                                                            , ~ lsp_nalb_sch_atq_ready                                          // 27
                                                            ,   lsp_nalb_sch_atq_v                                              // 26
                                                            , ~ lsp_dp_sch_dir_ready                                            // 25
                                                            ,   lsp_dp_sch_dir_v                                                // 24
                                                            , ~ lsp_nalb_sch_rorply_ready                                       // 23
                                                            ,   lsp_nalb_sch_rorply_v                                           // 22
                                                            , ~ lsp_dp_sch_rorply_ready                                         // 21
                                                            ,   lsp_dp_sch_rorply_v                                             // 20
                                                            , 1'h0                                                              // 19
                                                            , ~ atm_clk_idle                                                    // 18
                                                            , ~ aqed_clk_idle                                                   // 17
                                                            , ~ int_idle                                                        // 16
                                                            , ~ core_chp_lsp_token_ready                                        // 15
                                                            , ~ chp_lsp_token_rx_sync_idle                                      // 14
                                                            , ~ core_chp_lsp_cmp_ready                                          // 13
                                                            , ~ chp_lsp_cmp_rx_sync_idle                                        // 12
                                                            , ( core_rop_lsp_reordercmp_v & ~ core_rop_lsp_reordercmp_ready )   // 11
                                                            , ~ rop_lsp_reordercmp_rx_sync_idle                                 // 10
                                                            , ~ core_nalb_lsp_enq_lb_ready                                      //  9  Not a "pop" signal so OK to not gate w/ v
                                                            , ~ nalb_lsp_enq_lb_rx_sync_idle                                    //  8
                                                            , ( core_nalb_lsp_enq_rorply_v & ~ core_nalb_lsp_enq_rorply_ready ) //  7
                                                            , ~ nalb_lsp_enq_rorply_rx_sync_idle                                //  6
                                                            , ( core_dp_lsp_enq_dir_v & ~ core_dp_lsp_enq_dir_ready )           //  5
                                                            , ~ dp_lsp_enq_dir_rx_sync_idle                                     //  4
                                                            , ( core_dp_lsp_enq_rorply_v & ~ core_dp_lsp_enq_rorply_ready )     //  3
                                                            , ~ dp_lsp_enq_rorply_rx_sync_idle                                  //  2
                                                            , ( send_atm_to_cq_v & ~ send_atm_to_cq_ready )                     //  1
                                                            , ~ send_atm_to_cq_rx_sync_idle                                     //  0
                                                          } ;

//-----------------------------------------------------------------------------------------------------
assign cfg_pipe_health_hold_0_nxt       = {       4'h0
                                                , p4_lba_atm_sch_hold
                                                , p4_from_p5_hold
                                                , p0_lba_atm_credit_hold_cond
                                                , p0_lba_nalb_credit_hold_cond
                                                , 14'h0
                                                , p9_lba_ctrl_pipe.hold
                                                , p8_lba_ctrl_pipe.hold
                                                , p7_lba_ctrl_pipe.hold
                                                , p6_lba_ctrl_pipe.hold
                                                , p5_lba_ctrl_pipe.hold
                                                , p4_lba_ctrl_pipe.hold
                                                , p3_lba_ctrl_pipe.hold
                                                , p2_lba_ctrl_pipe.hold
                                                , p1_lba_ctrl_pipe.hold
                                                , 1'b0
                                          } ;

assign cfg_pipe_health_hold_1_nxt       = {       3'h0
                                                , p4_lbrpl_sch_hold
                                                , p3_lbrpl_ctrl_pipe.hold
                                                , p2_lbrpl_ctrl_pipe.hold
                                                , p1_lbrpl_ctrl_pipe.hold
                                                , p0_lbrpl_ctrl_pipe.hold
                                                , 3'h0
                                                , p4_dirrpl_sch_hold
                                                , p3_dirrpl_ctrl_pipe.hold
                                                , p2_dirrpl_ctrl_pipe.hold
                                                , p1_dirrpl_ctrl_pipe.hold
                                                , p0_dirrpl_ctrl_pipe.hold
                                                , 3'h0
                                                , p4_atq_sch_hold
                                                , p3_atq_ctrl_pipe.hold
                                                , p2_atq_ctrl_pipe.hold
                                                , p1_atq_ctrl_pipe.hold
                                                , p0_atq_ctrl_pipe.hold
                                                , 3'h0
                                                , p4_direnq_sch_hold
                                                , p3_direnq_ctrl_pipe.hold
                                                , p2_direnq_ctrl_pipe.hold
                                                , p1_direnq_ctrl_pipe.hold
                                                , p0_direnq_ctrl_pipe.hold
                                          } ;

//----
// Previously registered
assign hqm_lsp_target_cfg_pipe_health_hold_01_status            = cfg_pipe_health_hold_1_nxt ;
assign hqm_lsp_target_cfg_pipe_health_hold_00_status            = cfg_pipe_health_hold_0_nxt ;
//----

//-----------------------------------------------------------------------------------------------------
assign cfg_pipe_health_valid_0_nxt      = {       23'h0
                                                , p8_lba_ctrl_pipe_v_f
                                                , p7_lba_ctrl_pipe_v_f
                                                , p6_lba_ctrl_pipe_v_f
                                                , p5_lba_ctrl_pipe_v_f
                                                , p4_lba_ctrl_pipe_v_f
                                                , p3_lba_ctrl_pipe_v_f
                                                , p2_lba_ctrl_pipe_v_f
                                                , p1_lba_ctrl_pipe_v_f
                                                , 1'b0
                                          } ;

assign cfg_pipe_health_valid_1_nxt      = {       3'h0
                                                , p4_lbrpl_sch_v_f
                                                , p3_lbrpl_ctrl_pipe_v_f
                                                , p2_lbrpl_ctrl_pipe_v_f
                                                , p1_lbrpl_ctrl_pipe_v_f
                                                , p0_lbrpl_ctrl_pipe_v_f
                                                , 3'h0
                                                , p4_dirrpl_sch_v_f
                                                , p3_dirrpl_ctrl_pipe_v_f
                                                , p2_dirrpl_ctrl_pipe_v_f
                                                , p1_dirrpl_ctrl_pipe_v_f
                                                , p0_dirrpl_ctrl_pipe_v_f
                                                , 3'h0
                                                , p4_atq_sch_v_f
                                                , p3_atq_ctrl_pipe_v_f
                                                , p2_atq_ctrl_pipe_v_f
                                                , p1_atq_ctrl_pipe_v_f
                                                , p0_atq_ctrl_pipe_v_f
                                                , 3'h0
                                                , p4_direnq_sch_v_f
                                                , p3_direnq_ctrl_pipe_v_f
                                                , p2_direnq_ctrl_pipe_v_f
                                                , p1_direnq_ctrl_pipe_v_f
                                                , p0_direnq_ctrl_pipe_v_f
                                          } ;

//----
assign hqm_lsp_target_cfg_pipe_health_valid_01_status           = cfg_pipe_health_valid_1_nxt ;
assign hqm_lsp_target_cfg_pipe_health_valid_00_status           = cfg_pipe_health_valid_0_nxt ;
//----

//-----------------------------------------------------------------------------------------------------
// Loaded when interrupt reported to serializer

//----
assign hqm_lsp_target_cfg_syndrome_hw_capture_v         = cfg_syndrome0_capture_v ;
assign hqm_lsp_target_cfg_syndrome_hw_capture_data      = cfg_syndrome0_capture_data ;
assign hqm_lsp_target_cfg_syndrome_hw_syndrome_data_nc  = hqm_lsp_target_cfg_syndrome_hw_syndrome_data ;
//----

//-----------------------------------------------------------------------------------------------------
// Loaded when interrupt reported to serializer

//----
assign hqm_lsp_target_cfg_syndrome_sw_capture_v         = cfg_syndrome1_capture_v ;
assign hqm_lsp_target_cfg_syndrome_sw_capture_data      = cfg_syndrome1_capture_data ;
assign hqm_lsp_target_cfg_syndrome_sw_syndrome_data_nc  = hqm_lsp_target_cfg_syndrome_sw_syndrome_data ;
//----

//-----------------------------------------------------------------------------------------------------
assign hqm_lsp_target_cfg_diagnostic_aw_status_status   = {   4'h0                                                      // 31:28        spare
                                                            ,   ~ int_serializer_status_up   [2]                        // 27
                                                            , ( | int_serializer_status_up   [1:0] )                    // 26
                                                            ,   ~ int_serializer_status_down [2]                        // 25
                                                            , ( | int_serializer_status_down [1:0] )                    // 24
                                                            , 4'h0                                                      // 23:20        spare
                                                            , ( dir_tokrtn_db_out_valid & ~ dir_tokrtn_fifo_pop )       // 19
                                                            , ( | dir_tokrtn_db_status_pnc [1:0] )                      // 18
                                                            , ( enq_atq_db_out_valid & ~ enq_atq_db_out_ready )         // 17
                                                            , ( | enq_atq_db_status_pnc [1:0] )                         // 16
                                                            , 4'h0                                                      // 15:12        spare
                                                            ,   ldb_token_rtn_fifo_afull                                // 11
                                                            , ~ ldb_token_rtn_fifo_empty                                // 10
                                                            ,   uno_atm_cmp_fifo_afull                                  //  9
                                                            , ~ uno_atm_cmp_fifo_empty                                  //  8
                                                            ,   nalb_cmp_fifo_afull                                     //  7
                                                            , ~ nalb_cmp_fifo_empty                                     //  6
                                                            ,   enq_nalb_fifo_afull                                     //  5
                                                            , ~ enq_nalb_fifo_empty                                     //  4
                                                            ,   atm_cmp_fifo_afull                                      //  3
                                                            , ~ atm_cmp_fifo_empty                                      //  2
                                                            ,   nalb_sel_nalb_fifo_afull                                //  1
                                                            , ~ nalb_sel_nalb_fifo_empty                                //  0
                                                          } ;

//-----------------------------------------------------------------------------------------------------
assign cfg_lba_rlist_v                  = | ( p0_lba_rlist_cq_v & ~ cfg_cq_ldb_disable_f & ~ core_chp_lsp_ldb_cq_off_f ) ;       // 64-bit OR
assign cfg_lba_rlist_blast              = | p0_lba_rlist_blast_f ;      // 512-bit OR - timing might be tight
assign cfg_lba_slist_v                  = | ( p0_lba_slist_cq_v & ~ cfg_cq_ldb_disable_f & ~ core_chp_lsp_ldb_cq_off_f ) ;       // 64-bit OR
assign cfg_lba_slist_blast              = | p0_lba_slist_blast_f ;      // 512-bit OR - timing might be tight
assign cfg_lba_nalb_v                   = | p0_lba_nalb_v_f ;           // 512-bit OR - timing might be tight
assign cfg_lba_nalb_blast               = | p0_lba_nalb_blast_f ;       // 512-bit OR - timing might be tight
assign cfg_lba_cmpblast_chkv            = | p0_lba_cmpblast_chkv_f ;    // 512-bit OR - timing might be tight
assign cfg_lba_cmpblast                 = | p0_lba_cmpblast_f ;         // 512-bit OR - timing might be tight
assign cfg_atq_qid_dis                  = | ( ~p3_atq_qid_en_f ) ;      // 128-bit OR
assign cfg_lba_cq_busy                  = | p0_lba_cq_busy_sch_f ;      // 64-bit OR
assign cfg_lba_cq_no_space              = | ( ~p0_lba_cq_has_space_f ); // 64-bit OR
assign cfg_direnq_tok_cnt_v             = | p3_direnq_tok_cnt_v_f ;     // 128-bit OR
assign cfg_atq_aqed_act_v               = | p3_atq_aqed_act_v_f ;       // 128-bit OR
assign cfg_lba_atm_haswork              = ( ap_lsp_haswork_rlst_v & ap_lsp_haswork_rlst_func ) |        // Cover gap where not in AP
                                          ( ap_lsp_haswork_slst_v & ap_lsp_haswork_slst_func ) ;
assign cfg_lba_cq_tok_cnt_v             = | p8_lba_cq_tok_cnt_v_f ;     // 64-bit OR
assign cfg_lba_cq_if_cnt_v              = | p8_lba_cq_if_cnt_v_f ;      // 64-bit OR
assign cfg_qid_atq_aqed_empty           = & p3_atq_aqed_empty_f ;       // 128-bit AND
assign cfg_lba_atm_if_v                 = & p0_lba_atm_if_v_f ;         // 512-bit AND - timing might be tight
assign cfg_lba_ow_any                   = | ( p0_lba_cq_ow_f ) ;        // 64-bit OR

always_comb begin
  cfg_diag_status_0_nxt                                         = 32'h0 ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_SLIST_V ]          = cfg_lba_slist_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_SLIST_BLAST ]      = cfg_lba_slist_blast ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_RLIST_V ]          = cfg_lba_rlist_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_RLIST_BLAST ]      = cfg_lba_rlist_blast ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_NALB_V ]           = cfg_lba_nalb_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_NALB_BLAST ]       = cfg_lba_nalb_blast ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_CMPBLAST_CHKV ]    = cfg_lba_cmpblast_chkv ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_CMPBLAST ]         = cfg_lba_cmpblast ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_ATQ_QID_DIS ]      = cfg_atq_qid_dis ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_CQ_BUSY ]          = cfg_lba_cq_busy ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_CQ_NO_SPACE ]      = cfg_lba_cq_no_space ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_DIR_TOK_V ]        = cfg_direnq_tok_cnt_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_ATQ_ACT_V ]        = cfg_atq_aqed_act_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_ATM_HASWORK_V ]    = cfg_lba_atm_haswork ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_TOK_V ]         = cfg_lba_cq_tok_cnt_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_CMP_V ]         = cfg_lba_cq_if_cnt_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT0 ]   = p0_lba_cq_arb_status [0] ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT1 ]   = p0_lba_cq_arb_status [1] ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT2 ]   = p0_lba_cq_arb_status [2] ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LB_CQARB_STAT3 ]   = p0_lba_cq_arb_status [3] ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_STOP_ATQATM ]      = atq_stop_atqatm_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_QED_CRED_AFULL ]   = qed_deq_credit_afull ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_AQED_CRED_AFULL ]  = aqed_deq_credit_afull ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LBA_OW_ANY ]       = cfg_lba_ow_any ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_NSN_FCERR_RPTD ]   = nalb_sel_nalb_fifo_cerr_reported_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_AQED_EMPTY ]       = cfg_qid_atq_aqed_empty ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_ATM_IF_V ]         = cfg_lba_atm_if_v ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_TOT_IF_V ]         = p8_lba_tot_if_v_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LBWU_P1_V ]        = p1_lbwu_ctrl_pipe_v_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LBWU_P2_V ]        = p2_lbwu_ctrl_pipe_v_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LBWU_P3_V ]        = p3_lbwu_ctrl_pipe_v_f ;
  cfg_diag_status_0_nxt [ HQM_LSP_CFG_DIAG_0_LBWU_P4_V ]        = p4_lbwu_ctrl_pipe_v_f ;
end

// Register bits are used functionally, concerned about timing
always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_diag_status_0_f         <= 32'h0 ;
  end
  else begin
    cfg_diag_status_0_f         <= cfg_diag_status_0_nxt ;
  end
end // always

//----
assign hqm_lsp_target_cfg_diagnostic_status_0_status            = cfg_diag_status_0_f ;
//----

//-----------------------------------------------------------------------------------------------------
// cfg_diag_status_2 is for non-synth checking code only and will be optimized out, no static timing or power concerns.
// Change from v1 functionality, only capture first error.  Also no cfg clear.

assign p3_lba_cq2qid_v_err              = p3_lba_cq2qid_v_err_cond & ~ p3_lba_cq2qid_cq_disable_x & p3_lba_ctrl_pipe_v_f & ~ p4_lba_ctrl_pipe.hold ;
assign p7_lba_qid2cqidix_sch_v_err      = p7_lba_qid2cqidix_sch_v_err_cond & p7_lba_ctrl_pipe_v_f & ~ p8_lba_ctrl_pipe.hold ;
assign p7_lba_qid2cqidix_enq_v_err      = p7_lba_qid2cqidix_enq_v_err_cond & p7_lba_ctrl_pipe_v_f & ~ p8_lba_ctrl_pipe.hold ;

always_comb begin
  cfg_diag_status_2_allow_load          = | cfg_diag_status_2_f [7:0] ;

  cfg_diag_status_2_nxt                 = cfg_diag_status_2_f ;
  if ( cfg_diag_status_2_allow_load ) begin
    cfg_diag_status_2_nxt               = '0 ;                                  // Clear out unused/spare bits
    cfg_diag_status_2_nxt [7:0]         = {   5'h0                              // 7:3 spare
                                            , p7_lba_qid2cqidix_enq_v_err       // 2
                                            , p7_lba_qid2cqidix_sch_v_err       // 1
                                            , p3_lba_cq2qid_v_err               // 0
                                          } ;
    cfg_diag_status_2_nxt [  8 +: HQM_LSP_ARCH_NUM_LB_CQB2 ]    = p3_lba_ctrl_pipe_f.sch_cq ;           // Should match { p3_lba_cq2qid_rw_pipe_f_pnc.pcq << 1 }
    cfg_diag_status_2_nxt [ 16 +: HQM_LSP_ARCH_NUM_LB_QIDB2 ]   = p7_lba_qid2cqidix_rw_pipe_f.qid ;
    cfg_diag_status_2_nxt [ 24 +: HQM_LSP_ARCH_NUM_LB_QIDB2 ]   = p7_lba_qid2cqidix_rw_pipe_f.qid ;
  end
end

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_diag_status_2_f         <= 32'h0 ;
  end
  else begin
    cfg_diag_status_2_f         <= cfg_diag_status_2_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// cfg_diag_status_4 is for non-synth checking code only and will be optimized out, no static timing or power concerns.

always_comb begin
  // In general, "1" means "unexpected"
  cfg_diag_status_4_nxt         = 32'h0 ;
  cfg_diag_status_4_nxt [00]    = ~ ( & p3_cq_dir_tok_v_status ) ;              // DIR CQ has space w.r.t. token limit          Expect all 1
  cfg_diag_status_4_nxt [01]    = | p3_qid_dir_sch_v_status ;                   // DIR QID has work to do                       Expect all 0
  cfg_diag_status_4_nxt [02]    = ~ ( & cfg_qid_atq_aqed_avail_status ) ;       // ATQ QID has space w.r.t. aqed active limit   Expect all 1
  cfg_diag_status_4_nxt [03]    = cfg_qid_atq_sch_v_f ;                         // ATQ QID has work to do                       Expect all 0
  cfg_diag_status_4_nxt [04]    = ~ ( & cfg_qid_ldb_if_v_status ) ;             // LB QID has space w.r.t. qid if limit         Expect all 1
  cfg_diag_status_4_nxt [05]    = ~ ( & cfg_cq_ldb_if_v_status ) ;              // LB CQ has space w.r.t. cq if limit           Expect all 1
  cfg_diag_status_4_nxt [06]    = ~ ( & cfg_cq_ldb_tok_v_status ) ;             // LB CQ has space w.r.t. token limit           Expect all 1
  cfg_diag_status_4_nxt [07]    = | cfg_qid_ldb_sch_v_status ;                  // NALB qid has work to do                      Expect all 0
  cfg_diag_status_4_nxt [08]    = cfg_qid_dir_replay_v_f ;                      // ORD QID has DIR frag work to do              Expect all 0
  cfg_diag_status_4_nxt [09]    = cfg_qid_ldb_replay_v_f ;                      // ORD QID has LB frag work to do               Expect all 0
  cfg_diag_status_4_nxt [10]    = ~ ( & cfg_cq_ldb_thr_v_status ) ;             // LB CQ has space w.r.t. cq if threshold       Expect all 1
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_diag_status_4_f_nc      <= 32'h0 ;
  end
  else begin
    cfg_diag_status_4_f_nc      <= cfg_diag_status_4_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// Residue bits are not accessible by config.  Read returns 0.  Register is read-only.

//----
// Zero the residue bits going into the config reg; append the residue bits for functional use
always_comb begin
  hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_nxt                                          = 32'h0 ;
  hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_nxt [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]         = cfg_cq_ldb_tot_inflight_count_nxt [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0] ;

  cfg_cq_ldb_tot_inflight_count_f [HQM_LSP_LB_CQ_IF_CNT_WIDTH +: 2]     = cfg_cq_ldb_tot_inflight_count_res_f ;
  cfg_cq_ldb_tot_inflight_count_f [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]      = hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_f [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0] ;
end // always
//----

assign cfg_cq_ldb_tot_inflight_count_f_nc               = hqm_lsp_target_cfg_cq_ldb_tot_inflight_count_reg_f [31:HQM_LSP_LB_CQ_IF_CNT_WIDTH] ;
assign cfg_cq_ldb_tot_inflight_count_res_nxt            = cfg_cq_ldb_tot_inflight_count_nxt [HQM_LSP_LB_CQ_IF_CNT_WIDTH +: 2] ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_cq_ldb_tot_inflight_count_res_f <= 2'h0 ;
  end
  else begin
    cfg_cq_ldb_tot_inflight_count_res_f <= cfg_cq_ldb_tot_inflight_count_res_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// Only written by config
assign cfg_cq_ldb_tot_inflight_limit_nxt        = cfg_cq_ldb_tot_inflight_limit_f ;

//----
always_comb begin
  hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_nxt                                          = 32'h0 ;
  hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_nxt [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0]         = cfg_cq_ldb_tot_inflight_limit_nxt [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0] ;
  cfg_cq_ldb_tot_inflight_limit_f       = hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_f [HQM_LSP_LB_CQ_IF_CNT_WIDTH-1:0] ;
  cfg_cq_ldb_tot_inflight_limit_f_nc    = hqm_lsp_target_cfg_cq_ldb_tot_inflight_limit_reg_f [31:HQM_LSP_LB_CQ_IF_CNT_WIDTH] ;
end // always
//----

//-----------------------------------------------------------------------------------------------------
// Residue bits are not accessible by config.  Read returns 0.  Register is read-only.
// Note: vf reset updates total to subtract any inflight for the qid being reset

//----
// Zero the residue bits going into the config reg; append the residue bits for functional use
always_comb begin
  hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_nxt                                             = 32'h0 ;
  hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_nxt [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]        = cfg_aqed_tot_enqueue_count_nxt [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0] ;

  cfg_aqed_tot_enqueue_count_f [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH +: 2]    = cfg_aqed_tot_enqueue_count_res_f ;
  cfg_aqed_tot_enqueue_count_f [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]     = hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_f [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0] ;
end // always
//----

assign cfg_aqed_tot_enqueue_count_f_nc                  = hqm_lsp_target_cfg_aqed_tot_enqueue_count_reg_f [31:HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH] ;
assign cfg_aqed_tot_enqueue_count_res_nxt               = cfg_aqed_tot_enqueue_count_nxt [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH +: 2] ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_aqed_tot_enqueue_count_res_f    <= 2'h0 ;
  end
  else begin
    cfg_aqed_tot_enqueue_count_res_f    <= cfg_aqed_tot_enqueue_count_res_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// Only written by config
assign cfg_aqed_tot_enqueue_limit_nxt           = cfg_aqed_tot_enqueue_limit_f ;

//----
always_comb begin
  hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_nxt                                             = 32'h0 ;
  hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_nxt [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0]        = cfg_aqed_tot_enqueue_limit_nxt [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0] ;
  cfg_aqed_tot_enqueue_limit_f          = hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_f [HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH-1:0] ;
  cfg_aqed_tot_enqueue_limit_f_nc       = hqm_lsp_target_cfg_aqed_tot_enqueue_limit_reg_f [31:HQM_LSP_ATQ_AQED_ACT_CNT_WIDTH] ;
end // always
//----

//-----------------------------------------------------------------------------------------------------
// Residue bits are not accessible by config.  Read returns 0.  Register is read-only.
// Note: vf reset does NOT adjust total; sw algorithm is intended to guarantee that the BCAM will be empty for this VAS.

//----
// Zero the residue bits going into the config reg; append the residue bits for functional use
always_comb begin
  hqm_lsp_target_cfg_fid_inflight_count_reg_nxt                                         = 32'h0 ;
  hqm_lsp_target_cfg_fid_inflight_count_reg_nxt [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0]      = cfg_fid_inflight_count_nxt.cnt ;

  cfg_fid_inflight_count_f.cnt_res                                = cfg_fid_inflight_count_res_f ;
  cfg_fid_inflight_count_f.cnt                                    = hqm_lsp_target_cfg_fid_inflight_count_reg_f [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0] ;
end // always
//----

assign cfg_fid_inflight_count_f_nc                      = hqm_lsp_target_cfg_fid_inflight_count_reg_f [31:HQM_LSP_ATQ_FID_IF_CNT_WIDTH] ;
assign cfg_fid_inflight_count_res_nxt                   = cfg_fid_inflight_count_nxt.cnt_res ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_fid_inflight_count_res_f        <= 2'h0 ;
  end
  else begin
    cfg_fid_inflight_count_res_f        <= cfg_fid_inflight_count_res_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// Only written by config
assign cfg_fid_inflight_limit_nxt           = cfg_fid_inflight_limit_f ;

//----
always_comb begin
  hqm_lsp_target_cfg_fid_inflight_limit_reg_nxt                                         = 32'h0 ;
  hqm_lsp_target_cfg_fid_inflight_limit_reg_nxt [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0]      = cfg_fid_inflight_limit_nxt [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0] ;
  cfg_fid_inflight_limit_f              = hqm_lsp_target_cfg_fid_inflight_limit_reg_f [HQM_LSP_ATQ_FID_IF_CNT_WIDTH-1:0] ;
  cfg_fid_inflight_limit_f_nc           = hqm_lsp_target_cfg_fid_inflight_limit_reg_f [31:HQM_LSP_ATQ_FID_IF_CNT_WIDTH] ;
end // always
//----

//-----------------------------------------------------------------------------------------------------

//----
assign hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_v                  = 1'b0 ;
assign hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_nxt                = cfg_arb_weight_ldb_issue_0_nxt ;
assign cfg_arb_weight_ldb_issue_0_f                                     = hqm_lsp_target_cfg_arb_weight_ldb_issue_0_reg_f ;
//----

assign cfg_arb_weight_ldb_issue_0_nxt           = cfg_arb_weight_ldb_issue_0_f ;
assign cfg_lbi_cq_cmp_arb_weight_atm            = cfg_arb_weight_ldb_issue_0_f [7:0] ;
assign cfg_lbi_cq_cmp_arb_weight_nalb           = cfg_arb_weight_ldb_issue_0_f [15:8] ;
assign cfg_lbi_qid_cmp_arb_weight_ord           = cfg_arb_weight_ldb_issue_0_f [23:16] ;
assign cfg_lbi_qid_cmp_arb_weight_uno_atm       = cfg_arb_weight_ldb_issue_0_f [31:24] ;

//-----------------------------------------------------------------------------------------------------
// HQM_LSP_TARGET_CFG_ARB_WEIGHT_DIR_QID - used in arb wtcfg

//-----------------------------------------------------------------------------------------------------
// Note: cfg_arb_weight_ldb_qid_0_f is no longer needed and could be removed
assign cfg_arb_weight_ldb_qid_0_nxt             = cfg_arb_weight_ldb_qid_0_f ;
// Note: cfg_arb_weight_ldb_qid_1_f is no longer needed and could be removed
assign cfg_arb_weight_ldb_qid_1_nxt             = cfg_arb_weight_ldb_qid_1_f ;

// Requestor 0 is priority 0 (highest priority), and so on.  8-bit weights, one for each priority bin.
// Assign the default weights to give requestor 0 highest priority, etc.  Effective weight (chance of
// winning) is delta from next lower requestor, e.g. req 1 has (8'hc0 - 8'h80)/255 chance of winning.

//----
assign hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_v            = 1'b0 ;
assign hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_nxt          = cfg_arb_weight_ldb_qid_0_nxt ;
assign cfg_arb_weight_ldb_qid_0_f                               = hqm_lsp_target_cfg_arb_weight_ldb_qid_0_reg_f ;

assign hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_v            = 1'b0 ;
assign hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_nxt          = cfg_arb_weight_ldb_qid_1_nxt ;
assign cfg_arb_weight_ldb_qid_1_f                               = hqm_lsp_target_cfg_arb_weight_ldb_qid_1_reg_f ;
//----

//-----------------------------------------------------------------------------------------------------
assign cfg_arb_weight_atm_nalb_qid_0_nxt        = cfg_arb_weight_atm_nalb_qid_0_f ;
assign cfg_arb_weight_atm_nalb_qid_1_nxt        = cfg_arb_weight_atm_nalb_qid_1_f ;

// Requestor 0 is priority 0 (highest priority), and so on.  8-bit weights, one for each priority bin.
// Assign the default weights to give requestor 0 highest priority, etc.  Effective weight (chance of
// winning) is delta from next lower requestor, e.g. req 1 has (8'hc0 - 8'h80)/255 chance of winning.

//----
assign hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_v               = 1'b0 ;
assign hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_nxt             = cfg_arb_weight_atm_nalb_qid_0_nxt ;
assign cfg_arb_weight_atm_nalb_qid_0_f                                  = hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_0_reg_f ;

assign hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_v               = 1'b0 ;
assign hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_nxt             = cfg_arb_weight_atm_nalb_qid_1_nxt ;
assign cfg_arb_weight_atm_nalb_qid_1_f                                  = hqm_lsp_target_cfg_arb_weight_atm_nalb_qid_1_reg_f ;
//----

//-----------------------------------------------------------------------------------------------------
assign cfg_control_general_0_nxt                = cfg_control_general_0_f ;
assign cfg_control_disable_atq_empty_arb        = cfg_control_general_0_f [00] ;
assign cfg_control_include_tok_unit_idle        = cfg_control_general_0_f [01] ;
assign cfg_control_disable_rlist_pri            = cfg_control_general_0_f [02] ;
assign cfg_control_include_cmp_unit_idle        = cfg_control_general_0_f [03] ;
assign cfg_control_enable_inflight_thresh       = cfg_control_general_0_f [04] ;
// 5 - spare
assign cfg_control_single_op_direnq             = cfg_control_general_0_f [06] ;
assign cfg_control_half_bw_direnq               = cfg_control_general_0_f [07] ;
assign cfg_control_single_out_direnq            = cfg_control_general_0_f [08] ;
assign cfg_control_disable_multi_op_direnq      = cfg_control_general_0_f [09] ;
assign cfg_control_single_op_atq                = cfg_control_general_0_f [10] ;
assign cfg_control_half_bw_atq                  = cfg_control_general_0_f [11] ;
assign cfg_control_single_out_atq               = cfg_control_general_0_f [12] ;
assign cfg_control_disable_multi_op_atq         = cfg_control_general_0_f [13] ;
assign cfg_control_single_op_dirrpl             = cfg_control_general_0_f [14] ;
assign cfg_control_half_bw_dirrpl               = cfg_control_general_0_f [15] ;
assign cfg_control_single_out_dirrpl            = cfg_control_general_0_f [16] ;
assign cfg_control_single_op_lbrpl              = cfg_control_general_0_f [17] ;
assign cfg_control_half_bw_lbrpl                = cfg_control_general_0_f [18] ;
assign cfg_control_single_out_lbrpl             = cfg_control_general_0_f [19] ;
assign cfg_control_single_op_lba                = cfg_control_general_0_f [20] ;
assign cfg_control_half_bw_lba                  = cfg_control_general_0_f [21] ;
assign cfg_control_disable_multi_op_lba         = cfg_control_general_0_f [22] ;
assign cfg_control_single_op_atm_sched          = cfg_control_general_0_f [23] ;
assign cfg_control_single_op_atm_cmp            = cfg_control_general_0_f [24] ;
assign cfg_control_ldb_ce_tog_arb               = cfg_control_general_0_f [25] ;
// 26 - spare
assign cfg_smon0_v_sel                          = cfg_control_general_0_f [28:27] ;
assign cfg_smon0_value_sel                      = cfg_control_general_0_f [29] ;
assign cfg_smon0_comp_sel                       = cfg_control_general_0_f [31:30] ;
//----
assign hqm_lsp_target_cfg_control_general_0_reg_v               = 1'b0 ;
assign hqm_lsp_target_cfg_control_general_0_reg_nxt             = cfg_control_general_0_nxt ;
assign cfg_control_general_0_f                                  = hqm_lsp_target_cfg_control_general_0_reg_f ;
//-----------------------------------------------------------------------------------------------------
assign cfg_control_general_1_nxt                = cfg_control_general_1_f ;

assign cfg_control_qe_wt_frc_val                = cfg_control_general_1_f [01:00] ;
assign cfg_control_qe_wt_frc_v                  = cfg_control_general_1_f [02] ;
assign cfg_control_qe_wt_blk                    = cfg_control_general_1_f [03] ;
assign cfg_control_qed_lsp_deq_high_pri_wm      = cfg_control_general_1_f [08:04] ;
assign cfg_control_disable_wu_res_chk           = cfg_control_general_1_f [09] ;
// 11:10 - spare
assign cfg_control_aqed_lsp_deq_high_pri_wm     = cfg_control_general_1_f [16:12] ;
// 31:17 - spare

//----
assign hqm_lsp_target_cfg_control_general_1_reg_v               = 1'b0 ;
assign hqm_lsp_target_cfg_control_general_1_reg_nxt             = cfg_control_general_1_nxt ;
assign cfg_control_general_1_f                                  = hqm_lsp_target_cfg_control_general_1_reg_f ;
//----

// Upper pipe levels - those feeding into the status vectors, the internal end of the pipe.
assign direnq_upipe_idle_nxt    = ~ ( p0_direnq_ctrl_pipe_v_f | p1_direnq_ctrl_pipe_v_f | p2_direnq_ctrl_pipe_v_f ) ;
assign atq_upipe_idle_nxt       = ~ ( p0_atq_ctrl_pipe_v_f    | p1_atq_ctrl_pipe_v_f    | p2_atq_ctrl_pipe_v_f ) ;
assign dirrpl_upipe_idle_nxt    = ~ ( p0_dirrpl_ctrl_pipe_v_f | p1_dirrpl_ctrl_pipe_v_f | p2_dirrpl_ctrl_pipe_v_f ) ;
assign lbrpl_upipe_idle_nxt     = ~ ( p0_lbrpl_ctrl_pipe_v_f  | p1_lbrpl_ctrl_pipe_v_f  | p2_lbrpl_ctrl_pipe_v_f ) ;

// Do not include p0 since that is the arbiter level
assign lba_pipe_idle_nxt        = ~ ( p1_lba_ctrl_pipe_v_f    | p2_lba_ctrl_pipe_v_f    | p3_lba_ctrl_pipe_v_f |
                                      p4_lba_ctrl_pipe_v_f    | p5_lba_ctrl_pipe_v_f    | p6_lba_ctrl_pipe_v_f |
                                      p7_lba_ctrl_pipe_v_f    | p8_lba_ctrl_pipe_v_f                           ) ;

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    direnq_upipe_idle_f                 <= 1'b1 ;
    atq_upipe_idle_f                    <= 1'b1 ;
    dirrpl_upipe_idle_f                 <= 1'b1 ;
    lbrpl_upipe_idle_f                  <= 1'b1 ;
    lba_pipe_idle_f                     <= 1'b1 ;
  end
  else begin
    direnq_upipe_idle_f                 <= direnq_upipe_idle_nxt ;
    atq_upipe_idle_f                    <= atq_upipe_idle_nxt ;
    dirrpl_upipe_idle_f                 <= dirrpl_upipe_idle_nxt ;
    lbrpl_upipe_idle_f                  <= lbrpl_upipe_idle_nxt ;
    lba_pipe_idle_f                     <= lba_pipe_idle_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
assign cfg_lsp_csr_control_nxt                          = cfg_lsp_csr_control_f ;

// 1:0 reserved for int_cor, 3:2 reserved for int_unc
assign cfg_control_disable_qid_if_uflow_interrupt       = cfg_lsp_csr_control_f [4] ;
assign cfg_control_disable_qid_if_uflow_synd_load       = cfg_lsp_csr_control_f [5] ;
assign cfg_control_disable_cq_if_uflow_interrupt        = cfg_lsp_csr_control_f [6] ;
assign cfg_control_disable_cq_if_uflow_synd_load        = cfg_lsp_csr_control_f [7] ;
assign cfg_control_disable_tok_uflow_interrupt          = cfg_lsp_csr_control_f [8] ;
assign cfg_control_disable_tok_uflow_synd_load          = cfg_lsp_csr_control_f [9] ;
assign cfg_control_disable_hwerr_interrupt              = cfg_lsp_csr_control_f [10] ;
assign cfg_control_disable_hwerr_synd_load              = cfg_lsp_csr_control_f [11] ;
assign cfg_control_disable_non_mc_interrupt             = cfg_lsp_csr_control_f [12] ;
assign cfg_control_disable_non_mc_synd_load             = cfg_lsp_csr_control_f [13] ;

assign cfg_control_ldb_wrr_count_base                   = cfg_lsp_csr_control_f [30:28] ;
assign cfg_control_atm_cq_qid_priority_prot             = cfg_lsp_csr_control_f [31] ;

//----
assign hqm_lsp_target_cfg_lsp_csr_control_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_lsp_csr_control_reg_nxt       = cfg_lsp_csr_control_nxt ;
assign cfg_lsp_csr_control_f                            = hqm_lsp_target_cfg_lsp_csr_control_reg_f ;
//----

//-----------------------------------------------------------------------------------------------------
always_comb begin
  cfg_ldb_sched_control_nxt                     = cfg_ldb_sched_control_f_pnc ;
  cfg_ldb_sched_control_nxt [16:12]             = 5'h0 ;                        // Self-clearing
end // always

assign cfg_ldb_sched_control_cq                 = cfg_ldb_sched_control_f_pnc [5:0] ;
assign cfg_ldb_sched_control_qidix              = cfg_ldb_sched_control_f_pnc [10:8] ;
assign cfg_ldb_sched_control_value              = cfg_ldb_sched_control_f_pnc [11] ;
assign cfg_ldb_sched_control_nalb_haswork_v     = cfg_ldb_sched_control_f_pnc [12] ;    // Self-clearing
assign cfg_ldb_sched_control_rlist_haswork_v    = cfg_ldb_sched_control_f_pnc [13] ;    // Self-clearing
assign cfg_ldb_sched_control_slist_haswork_v    = cfg_ldb_sched_control_f_pnc [14] ;    // Self-clearing
assign cfg_ldb_sched_control_inflight_ok_v      = cfg_ldb_sched_control_f_pnc [15] ;    // Self-clearing
assign cfg_ldb_sched_control_aqed_nfull_v       = cfg_ldb_sched_control_f_pnc [16] ;    // Self-clearing

assign cfg_ldb_sched_control_cq_qidix           = { cfg_ldb_sched_control_cq , cfg_ldb_sched_control_qidix } ;
assign cfg_ldb_sched_control_qid                = cfg_ldb_sched_control_cq_qidix [6:0] ;

//----
assign hqm_lsp_target_cfg_ldb_sched_control_reg_nxt             = cfg_ldb_sched_control_nxt ;
assign cfg_ldb_sched_control_f_pnc                              = hqm_lsp_target_cfg_ldb_sched_control_reg_f ;
//----

//-----------------------------------------------------------------------------------------------------
assign cfg_control_pipeline_credits_nxt         = cfg_control_pipeline_credits_f ;
assign cfg_lba_pipeline_credit_limit            = cfg_control_pipeline_credits_f [7:0] ;
assign cfg_atm_pipeline_credit_limit            = cfg_control_pipeline_credits_f [15:8] ;
assign cfg_qed_deq_pipeline_credit_limit_pnc    = cfg_control_pipeline_credits_f [23:16] ;
assign cfg_aqed_deq_pipeline_credit_limit_pnc   = cfg_control_pipeline_credits_f [31:24] ;

//----
assign hqm_lsp_target_cfg_control_pipeline_credits_reg_v                = 1'b0 ;
assign hqm_lsp_target_cfg_control_pipeline_credits_reg_nxt              = cfg_control_pipeline_credits_nxt ;
assign cfg_control_pipeline_credits_f                                   = hqm_lsp_target_cfg_control_pipeline_credits_reg_f ;
//----

//-----------------------------------------------------------------------------------------------------
// New V2 registers

assign hqm_lsp_target_cfg_cos_ctrl_reg_v        = 1'b0 ;
assign hqm_lsp_target_cfg_cos_ctrl_reg_nxt      = hqm_lsp_target_cfg_cos_ctrl_reg_f ;

// Only changed by shdw load
always_comb begin
  cfg_range_cos0_reg_nxt                        = cfg_range_cos0_reg_f ;
  cfg_range_cos1_reg_nxt                        = cfg_range_cos1_reg_f ;
  cfg_range_cos2_reg_nxt                        = cfg_range_cos2_reg_f ;
  cfg_range_cos3_reg_nxt                        = cfg_range_cos3_reg_f ;

  if ( cfg_shdw_ctrl_load ) begin
    cfg_range_cos0_reg_nxt                      = hqm_lsp_target_cfg_shdw_range_cos0_reg_f ;
    cfg_range_cos1_reg_nxt                      = hqm_lsp_target_cfg_shdw_range_cos1_reg_f ;
    cfg_range_cos2_reg_nxt                      = hqm_lsp_target_cfg_shdw_range_cos2_reg_f ;
    cfg_range_cos3_reg_nxt                      = hqm_lsp_target_cfg_shdw_range_cos3_reg_f ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_range_cos0_reg_f                <= { 23'h0 , HQM_LSP_CFG_RANGE_COS0_DEFAULT } ;
    cfg_range_cos1_reg_f                <= { 23'h0 , HQM_LSP_CFG_RANGE_COS1_DEFAULT } ;
    cfg_range_cos2_reg_f                <= { 23'h0 , HQM_LSP_CFG_RANGE_COS2_DEFAULT } ;
    cfg_range_cos3_reg_f                <= { 23'h0 , HQM_LSP_CFG_RANGE_COS3_DEFAULT } ;
  end
  else begin
    cfg_range_cos0_reg_f                <= cfg_range_cos0_reg_nxt ;
    cfg_range_cos1_reg_f                <= cfg_range_cos1_reg_nxt ;
    cfg_range_cos2_reg_f                <= cfg_range_cos2_reg_nxt ;
    cfg_range_cos3_reg_f                <= cfg_range_cos3_reg_nxt ;
  end
end // always

assign cfg_range_cos0_f                 = cfg_range_cos0_reg_f [8:0] ;
assign cfg_range_cos1_f                 = cfg_range_cos1_reg_f [8:0] ;
assign cfg_range_cos2_f                 = cfg_range_cos2_reg_f [8:0] ;
assign cfg_range_cos3_f                 = cfg_range_cos3_reg_f [8:0] ;
assign cfg_no_extra_credit0_f           = cfg_range_cos0_reg_f [31] ;
assign cfg_no_extra_credit1_f           = cfg_range_cos1_reg_f [31] ;
assign cfg_no_extra_credit2_f           = cfg_range_cos2_reg_f [31] ;
assign cfg_no_extra_credit3_f           = cfg_range_cos3_reg_f [31] ;

assign hqm_lsp_target_cfg_credit_sat_cos0_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_credit_sat_cos1_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_credit_sat_cos2_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_credit_sat_cos3_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_credit_sat_cos0_reg_nxt       = hqm_lsp_target_cfg_credit_sat_cos0_reg_f ;
assign hqm_lsp_target_cfg_credit_sat_cos1_reg_nxt       = hqm_lsp_target_cfg_credit_sat_cos1_reg_f ;
assign hqm_lsp_target_cfg_credit_sat_cos2_reg_nxt       = hqm_lsp_target_cfg_credit_sat_cos2_reg_f ;
assign hqm_lsp_target_cfg_credit_sat_cos3_reg_nxt       = hqm_lsp_target_cfg_credit_sat_cos3_reg_f ;
assign cfg_credit_sat_cos0_f    = hqm_lsp_target_cfg_credit_sat_cos0_reg_f [15:0] ;
assign cfg_credit_sat_cos1_f    = hqm_lsp_target_cfg_credit_sat_cos1_reg_f [15:0] ;
assign cfg_credit_sat_cos2_f    = hqm_lsp_target_cfg_credit_sat_cos2_reg_f [15:0] ;
assign cfg_credit_sat_cos3_f    = hqm_lsp_target_cfg_credit_sat_cos3_reg_f [15:0] ;

assign cfg_starv_avoid_enable_f         = hqm_lsp_target_cfg_cos_ctrl_reg_f [31] ;
assign cfg_starv_avoid_thresh_min_f     = hqm_lsp_target_cfg_cos_ctrl_reg_f [9:0] ;
assign cfg_starv_avoid_thresh_max_f     = hqm_lsp_target_cfg_cos_ctrl_reg_f [19:10] ;

assign hqm_lsp_target_cfg_credit_cnt_cos0_reg_nxt       = { 5'h0 , cfg_starv_avoid_cnt_cos0 , cfg_credit_cnt_cos0 } ;
assign hqm_lsp_target_cfg_credit_cnt_cos1_reg_nxt       = { 5'h0 , cfg_starv_avoid_cnt_cos1 , cfg_credit_cnt_cos1 } ;
assign hqm_lsp_target_cfg_credit_cnt_cos2_reg_nxt       = { 5'h0 , cfg_starv_avoid_cnt_cos2 , cfg_credit_cnt_cos2 } ;
assign hqm_lsp_target_cfg_credit_cnt_cos3_reg_nxt       = { 5'h0 , cfg_starv_avoid_cnt_cos3 , cfg_credit_cnt_cos3 } ;
assign hqm_lsp_target_cfg_credit_cnt_cos0_nc            = hqm_lsp_target_cfg_credit_cnt_cos0_reg_f ;
assign hqm_lsp_target_cfg_credit_cnt_cos1_nc            = hqm_lsp_target_cfg_credit_cnt_cos1_reg_f ;
assign hqm_lsp_target_cfg_credit_cnt_cos2_nc            = hqm_lsp_target_cfg_credit_cnt_cos2_reg_f ;
assign hqm_lsp_target_cfg_credit_cnt_cos3_nc            = hqm_lsp_target_cfg_credit_cnt_cos3_reg_f ;


// Self-clearing, RW/1S/V
assign hqm_lsp_target_cfg_shdw_ctrl_reg_nxt             = 32'h0 ;
assign cfg_shdw_ctrl_load                               = hqm_lsp_target_cfg_shdw_ctrl_reg_f [0] ;
assign cfg_shdw_ctrl_load_spare_nc                      = hqm_lsp_target_cfg_shdw_ctrl_reg_f [31:1] ;

// Only updated by config
assign hqm_lsp_target_cfg_shdw_range_cos0_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_shdw_range_cos1_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_shdw_range_cos2_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_shdw_range_cos3_reg_v         = 1'b0 ;
assign hqm_lsp_target_cfg_shdw_range_cos0_reg_nxt       = hqm_lsp_target_cfg_shdw_range_cos0_reg_f ;
assign hqm_lsp_target_cfg_shdw_range_cos1_reg_nxt       = hqm_lsp_target_cfg_shdw_range_cos1_reg_f ;
assign hqm_lsp_target_cfg_shdw_range_cos2_reg_nxt       = hqm_lsp_target_cfg_shdw_range_cos2_reg_f ;
assign hqm_lsp_target_cfg_shdw_range_cos3_reg_nxt       = hqm_lsp_target_cfg_shdw_range_cos3_reg_f ;

assign hqm_lsp_target_cfg_sch_rdy_inc                   = p0_lba_cq_arb_update ;
assign hqm_lsp_target_cfg_schd_cos0_inc                 = cfg_schd_cos [0] ;
assign hqm_lsp_target_cfg_schd_cos1_inc                 = cfg_schd_cos [1] ;
assign hqm_lsp_target_cfg_schd_cos2_inc                 = cfg_schd_cos [2] ;
assign hqm_lsp_target_cfg_schd_cos3_inc                 = cfg_schd_cos [3] ;
assign hqm_lsp_target_cfg_rdy_cos0_inc                  = cfg_rdy_cos [0] ;
assign hqm_lsp_target_cfg_rdy_cos1_inc                  = cfg_rdy_cos [1] ;
assign hqm_lsp_target_cfg_rdy_cos2_inc                  = cfg_rdy_cos [2] ;
assign hqm_lsp_target_cfg_rdy_cos3_inc                  = cfg_rdy_cos [3] ;
assign hqm_lsp_target_cfg_rnd_loss_cos0_inc             = cfg_rnd_loss_cos [0] ;
assign hqm_lsp_target_cfg_rnd_loss_cos1_inc             = cfg_rnd_loss_cos [1] ;
assign hqm_lsp_target_cfg_rnd_loss_cos2_inc             = cfg_rnd_loss_cos [2] ;
assign hqm_lsp_target_cfg_rnd_loss_cos3_inc             = cfg_rnd_loss_cos [3] ;
assign hqm_lsp_target_cfg_cnt_win_cos0_inc              = cfg_cnt_win_cos [0] ;
assign hqm_lsp_target_cfg_cnt_win_cos1_inc              = cfg_cnt_win_cos [1] ;
assign hqm_lsp_target_cfg_cnt_win_cos2_inc              = cfg_cnt_win_cos [2] ;
assign hqm_lsp_target_cfg_cnt_win_cos3_inc              = cfg_cnt_win_cos [3] ;

assign hqm_lsp_target_cfg_sch_rdy_en                    = 1'b1 ;
assign hqm_lsp_target_cfg_schd_cos0_en                  = 1'b1 ;
assign hqm_lsp_target_cfg_schd_cos1_en                  = 1'b1 ;
assign hqm_lsp_target_cfg_schd_cos2_en                  = 1'b1 ;
assign hqm_lsp_target_cfg_schd_cos3_en                  = 1'b1 ;
assign hqm_lsp_target_cfg_rdy_cos0_en                   = 1'b1 ;
assign hqm_lsp_target_cfg_rdy_cos1_en                   = 1'b1 ;
assign hqm_lsp_target_cfg_rdy_cos2_en                   = 1'b1 ;
assign hqm_lsp_target_cfg_rdy_cos3_en                   = 1'b1 ;
assign hqm_lsp_target_cfg_rnd_loss_cos0_en              = 1'b1 ;
assign hqm_lsp_target_cfg_rnd_loss_cos1_en              = 1'b1 ;
assign hqm_lsp_target_cfg_rnd_loss_cos2_en              = 1'b1 ;
assign hqm_lsp_target_cfg_rnd_loss_cos3_en              = 1'b1 ;
assign hqm_lsp_target_cfg_cnt_win_cos0_en               = 1'b1 ;
assign hqm_lsp_target_cfg_cnt_win_cos1_en               = 1'b1 ;
assign hqm_lsp_target_cfg_cnt_win_cos2_en               = 1'b1 ;
assign hqm_lsp_target_cfg_cnt_win_cos3_en               = 1'b1 ;

assign hqm_lsp_target_cfg_sch_rdy_clr                   = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos0_clr                 = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos1_clr                 = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos2_clr                 = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos3_clr                 = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos0_clr                  = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos1_clr                  = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos2_clr                  = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos3_clr                  = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos0_clr             = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos1_clr             = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos2_clr             = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos3_clr             = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos0_clr              = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos1_clr              = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos2_clr              = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos3_clr              = 1'b0 ;

assign hqm_lsp_target_cfg_sch_rdy_clrv                  = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos0_clrv                = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos1_clrv                = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos2_clrv                = 1'b0 ;
assign hqm_lsp_target_cfg_schd_cos3_clrv                = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos0_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos1_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos2_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_rdy_cos3_clrv                 = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos0_clrv            = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos1_clrv            = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos2_clrv            = 1'b0 ;
assign hqm_lsp_target_cfg_rnd_loss_cos3_clrv            = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos0_clrv             = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos1_clrv             = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos2_clrv             = 1'b0 ;
assign hqm_lsp_target_cfg_cnt_win_cos3_clrv             = 1'b0 ;

assign hqm_lsp_target_cfg_sch_rdy_count_nc              = hqm_lsp_target_cfg_sch_rdy_count ;
assign hqm_lsp_target_cfg_schd_cos0_count_nc            = hqm_lsp_target_cfg_schd_cos0_count ;
assign hqm_lsp_target_cfg_schd_cos1_count_nc            = hqm_lsp_target_cfg_schd_cos1_count ;
assign hqm_lsp_target_cfg_schd_cos2_count_nc            = hqm_lsp_target_cfg_schd_cos2_count ;
assign hqm_lsp_target_cfg_schd_cos3_count_nc            = hqm_lsp_target_cfg_schd_cos3_count ;
assign hqm_lsp_target_cfg_rdy_cos0_count_nc             = hqm_lsp_target_cfg_rdy_cos0_count ;
assign hqm_lsp_target_cfg_rdy_cos1_count_nc             = hqm_lsp_target_cfg_rdy_cos1_count ;
assign hqm_lsp_target_cfg_rdy_cos2_count_nc             = hqm_lsp_target_cfg_rdy_cos2_count ;
assign hqm_lsp_target_cfg_rdy_cos3_count_nc             = hqm_lsp_target_cfg_rdy_cos3_count ;
assign hqm_lsp_target_cfg_rnd_loss_cos0_count_nc        = hqm_lsp_target_cfg_rnd_loss_cos0_count ;
assign hqm_lsp_target_cfg_rnd_loss_cos1_count_nc        = hqm_lsp_target_cfg_rnd_loss_cos1_count ;
assign hqm_lsp_target_cfg_rnd_loss_cos2_count_nc        = hqm_lsp_target_cfg_rnd_loss_cos2_count ;
assign hqm_lsp_target_cfg_rnd_loss_cos3_count_nc        = hqm_lsp_target_cfg_rnd_loss_cos3_count ;
assign hqm_lsp_target_cfg_cnt_win_cos0_count_nc         = hqm_lsp_target_cfg_cnt_win_cos0_count ;
assign hqm_lsp_target_cfg_cnt_win_cos1_count_nc         = hqm_lsp_target_cfg_cnt_win_cos1_count ;
assign hqm_lsp_target_cfg_cnt_win_cos2_count_nc         = hqm_lsp_target_cfg_cnt_win_cos2_count ;
assign hqm_lsp_target_cfg_cnt_win_cos3_count_nc         = hqm_lsp_target_cfg_cnt_win_cos3_count ;

//-----------------------------------------------------------------------------------------------------
// New V25 registers

assign hqm_lsp_target_cfg_control_sched_slot_count_reg_v        = 1'b0 ;
assign hqm_lsp_target_cfg_control_sched_slot_count_reg_nxt      = hqm_lsp_target_cfg_control_sched_slot_count_reg_f ;

assign cfg_sched_slot_count_en                  = hqm_lsp_target_cfg_control_sched_slot_count_reg_f [0] ;
assign cfg_sched_slot_count_clr                 = hqm_lsp_target_cfg_control_sched_slot_count_reg_f [1] ;
assign cfg_sched_slot_count_cq                  = hqm_lsp_target_cfg_control_sched_slot_count_reg_f [15:8] ;

assign cfg_sched_slot_count_trigger             = p4_lba_ctrl_pipe_v_f & ~ p5_lba_ctrl_pipe.hold & p4_lba_ctrl_pipe_f.sch_v &
                                                  ( p4_lba_ctrl_pipe_f.sch_cq == cfg_sched_slot_count_cq [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ) ;

always_comb begin
  cfg_sched_slot_count_inc_nxt                                          = '0 ;
  cfg_sched_slot_count_prev_slot_v_nxt                                  = cfg_sched_slot_count_prev_slot_v_f ;
  cfg_sched_slot_count_prev_slot_nxt                                    = cfg_sched_slot_count_prev_slot_f ;
  if ( cfg_sched_slot_count_clr ) begin
    cfg_sched_slot_count_prev_slot_v_nxt                                = 1'b0 ;
    cfg_sched_slot_count_prev_slot_nxt                                  = '0 ;
  end
  else if ( cfg_sched_slot_count_trigger ) begin
    cfg_sched_slot_count_prev_slot_v_nxt                                = 1'b1 ;
    cfg_sched_slot_count_prev_slot_nxt                                  = p4_lba_sch_arb_winner_qidix ;
    if ( cfg_sched_slot_count_prev_slot_v_f & ( cfg_sched_slot_count_prev_slot_f == p4_lba_sch_arb_winner_qidix ) ) begin
      cfg_sched_slot_count_inc_nxt [ p4_lba_sch_arb_winner_qidix ]      = 1'b1 ;
    end
  end
end

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_sched_slot_count_inc_f          <= '0 ;
    cfg_sched_slot_count_prev_slot_v_f  <= 1'b0 ;
    cfg_sched_slot_count_prev_slot_f    <= '0 ;
  end
  else begin
    cfg_sched_slot_count_inc_f          <= cfg_sched_slot_count_inc_nxt ;
    cfg_sched_slot_count_prev_slot_v_f  <= cfg_sched_slot_count_prev_slot_v_nxt ;
    cfg_sched_slot_count_prev_slot_f    <= cfg_sched_slot_count_prev_slot_nxt ;
  end
end // always

assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_count ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count_nc    = hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_count ;

assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_inc         = cfg_sched_slot_count_inc_f [0] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_inc         = cfg_sched_slot_count_inc_f [1] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_inc         = cfg_sched_slot_count_inc_f [2] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_inc         = cfg_sched_slot_count_inc_f [3] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_inc         = cfg_sched_slot_count_inc_f [4] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_inc         = cfg_sched_slot_count_inc_f [5] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_inc         = cfg_sched_slot_count_inc_f [6] ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_inc         = cfg_sched_slot_count_inc_f [7] ;

assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_en          = cfg_sched_slot_count_en ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_en          = cfg_sched_slot_count_en ;

assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clr         = cfg_sched_slot_count_clr ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clr         = cfg_sched_slot_count_clr ;

assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_0_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_1_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_2_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_3_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_4_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_5_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_6_clrv        = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_sched_slot_count_7_clrv        = 1'b0 ;

//-----------------------------------------------------------------------------------------------------
// Detect conditions which should only be possible if logic bug, only for coverage/simulation, optimized out of hardware.
// Checked by eot_check task.
// Connect to debug config registers if necessary.

always_comb begin
  // Note, these errors should only occur if there is a logic bug
  hqm_lsp_target_cfg_debug_00_reg_nxt           = hqm_lsp_target_cfg_debug_00_reg_f ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [00]      = hqm_lsp_target_cfg_debug_00_reg_f [00] | p3_atq_enq_cnt_uflow_err_f ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [01]      = hqm_lsp_target_cfg_debug_00_reg_f [01] | p3_atq_enq_cnt_oflow_err_f ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [02]      = '0 ;                                   // spare
  hqm_lsp_target_cfg_debug_00_reg_nxt [03]      = hqm_lsp_target_cfg_debug_00_reg_f [03] | p4_atq_atm_active_oflow_err_f ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [04]      = hqm_lsp_target_cfg_debug_00_reg_f [04] | nalb_lsp_enq_rorply_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [05]      = hqm_lsp_target_cfg_debug_00_reg_f [05] | nalb_lsp_enq_rorply_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [06]      = hqm_lsp_target_cfg_debug_00_reg_f [06] | send_atm_to_cq_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [07]      = hqm_lsp_target_cfg_debug_00_reg_f [07] | send_atm_to_cq_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [08]      = hqm_lsp_target_cfg_debug_00_reg_f [08] | dp_lsp_enq_rorply_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [09]      = hqm_lsp_target_cfg_debug_00_reg_f [09] | dp_lsp_enq_rorply_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [10]      = hqm_lsp_target_cfg_debug_00_reg_f [10] | dp_lsp_enq_dir_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [11]      = hqm_lsp_target_cfg_debug_00_reg_f [11] | dp_lsp_enq_dir_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [12]      = hqm_lsp_target_cfg_debug_00_reg_f [12] | nalb_lsp_enq_lb_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [13]      = hqm_lsp_target_cfg_debug_00_reg_f [13] | nalb_lsp_enq_lb_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [14]      = hqm_lsp_target_cfg_debug_00_reg_f [14] | rop_lsp_reordercmp_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [15]      = hqm_lsp_target_cfg_debug_00_reg_f [15] | rop_lsp_reordercmp_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [16]      = hqm_lsp_target_cfg_debug_00_reg_f [16] | chp_lsp_cmp_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [17]      = hqm_lsp_target_cfg_debug_00_reg_f [17] | chp_lsp_cmp_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [18]      = hqm_lsp_target_cfg_debug_00_reg_f [18] | chp_lsp_token_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [19]      = hqm_lsp_target_cfg_debug_00_reg_f [19] | chp_lsp_token_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [20]      = hqm_lsp_target_cfg_debug_00_reg_f [20] | cfg_rx_sync_fifo_uf ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [21]      = hqm_lsp_target_cfg_debug_00_reg_f [21] | cfg_rx_sync_fifo_of ;
  hqm_lsp_target_cfg_debug_00_reg_nxt [31:22]   = '0 ;                                   // spare

// Note: Would be preferable to use parameter names here instead of literal values
// Note, these errors should only occur if there is a logic bug, possibly just with the detect_feature_0 settings
// Confirm that detect_feature_0 limits are correct, should never see a value greater than the max being detected
  hqm_lsp_target_cfg_debug_01_reg_nxt           = hqm_lsp_target_cfg_debug_01_reg_f ;
  hqm_lsp_target_cfg_debug_01_reg_nxt [00]      = '0 ;          // Bit 0 has dedicated hw error detect bit atq_fid_if_lim_err_f ( int_inf[6] bit 15 )
  hqm_lsp_target_cfg_debug_01_reg_nxt [01]      = '0 ;          // Bit 1 has dedicated hw error detect bit atq_tot_act_lim_err_f ( int_inf[6] bit 16 )
  hqm_lsp_target_cfg_debug_01_reg_nxt [02]      = hqm_lsp_target_cfg_debug_01_reg_f [02] | ( p2_direnq_enq_cnt_upd_v & ( p2_direnq_enq_cnt_upd.cnt > 15'h4000 ) ) ;             // Max V25 DIR credits = 16K
  hqm_lsp_target_cfg_debug_01_reg_nxt [03]      = hqm_lsp_target_cfg_debug_01_reg_f [03] | ( p2_direnq_tok_cnt_upd_v & ( p2_direnq_tok_cnt_upd.cnt > 11'h400 ) ) ;              // Max V25 DIR CQ depth = 1K
  hqm_lsp_target_cfg_debug_01_reg_nxt [04]      = hqm_lsp_target_cfg_debug_01_reg_f [04] | ( p2_atq_enq_cnt_upd_v & ( p2_atq_enq_cnt_upd.cnt > 15'h4000 ) ) ;                   // Max V25 LDB credits = 16K
  hqm_lsp_target_cfg_debug_01_reg_nxt [05]      = hqm_lsp_target_cfg_debug_01_reg_f [05] | ( p2_atq_aqed_act_cnt_upd_v & ( p2_atq_aqed_act_cnt_upd.cnt > 12'h800 ) ) ;          // Max AQED active = 2K
  hqm_lsp_target_cfg_debug_01_reg_nxt [06]      = hqm_lsp_target_cfg_debug_01_reg_f [06] | ( p3_atq_fid_inflight_cnt_upd_v & ( cfg_fid_inflight_count_f.cnt > 12'h800 ) ) ;     // Max FID inflight = 2K
  hqm_lsp_target_cfg_debug_01_reg_nxt [07]      = hqm_lsp_target_cfg_debug_01_reg_f [07] | ( p2_dirrpl_enq_cnt_upd_v & ( p2_dirrpl_enq_cnt_upd.cnt > 15'h4000 ) ) ;             // Max V25 DIR credits = 16K
  hqm_lsp_target_cfg_debug_01_reg_nxt [08]      = hqm_lsp_target_cfg_debug_01_reg_f [08] | ( p2_lbrpl_enq_cnt_upd_v & ( p2_lbrpl_enq_cnt_upd.cnt > 15'h4000 ) ) ;               // Max V25 LDB credits = 16K
  hqm_lsp_target_cfg_debug_01_reg_nxt [09]      = hqm_lsp_target_cfg_debug_01_reg_f [09] | ( p7_lba_qid_enq_cnt_upd_v & ( p7_lba_qid_enq_cnt_upd.cnt > 15'h4000 ) ) ;           // Max V25 LDB credits = 16K
  hqm_lsp_target_cfg_debug_01_reg_nxt [10]      = hqm_lsp_target_cfg_debug_01_reg_f [10] | ( p7_lba_cq_tok_cnt_upd_v & ( p7_lba_cq_tok_cnt_upd_cnt.cnt > 11'h400 ) ) ;          // Max LDB CQ depth = 1K
  hqm_lsp_target_cfg_debug_01_reg_nxt [11]      = hqm_lsp_target_cfg_debug_01_reg_f [11] | ( p7_lba_cq_if_cnt_upd_v & ( p7_lba_cq_if_cnt_upd_cnt.cnt > 12'h800 ) ) ;            // Hist list depth = 2K
  hqm_lsp_target_cfg_debug_01_reg_nxt [12]      = hqm_lsp_target_cfg_debug_01_reg_f [12] | ( p7_lba_qid_if_cnt_upd_v & ( p7_lba_qid_if_cnt_upd.cnt > 12'h800 ) ) ;              // Max SN = 2K
  hqm_lsp_target_cfg_debug_01_reg_nxt [31:13]   = '0 ;          //spare
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    hqm_lsp_target_cfg_debug_00_reg_f   <= 32'h0 ;
    hqm_lsp_target_cfg_debug_01_reg_f   <= 32'h0 ;
  end
  else begin
    hqm_lsp_target_cfg_debug_00_reg_f   <= hqm_lsp_target_cfg_debug_00_reg_nxt ;
    hqm_lsp_target_cfg_debug_01_reg_f   <= hqm_lsp_target_cfg_debug_01_reg_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
// Detect feature regs, only for coverage/simulation, optimized out of hardware

assign p3_atq_qid_v_any                 = | p3_atq_qid_v_f ;

always_comb begin
  cfg_detect_feature_0_set      = 32'h0 ;
  cfg_detect_feature_0_set [0]  = p3_atq_qid_v_any & p3_atq_fid_inflight_cnt_eq_lim ;
  cfg_detect_feature_0_set [1]  = p3_atq_qid_v_any & p3_atq_tot_act_cnt_eq_lim ;
  cfg_detect_feature_0_set [2]  = p2_direnq_enq_cnt_upd_v & p2_direnq_enq_cnt_upd.cnt[14] ;     // Max limit enforced by CHP = 15'h4000 = 16K
  cfg_detect_feature_0_set [3]  = p2_direnq_tok_cnt_upd_v & p2_direnq_tok_cnt_upd.cnt[10] ;     // Max LSP DIR CQ depth cfg limit = 11'h400 = 1K
  cfg_detect_feature_0_set [4]  = p2_atq_enq_cnt_upd_v & p2_atq_enq_cnt_upd.cnt[14] ;           // Max LB credits (QED depth) = 15'h4000 = 16K

  // Would be good to test that both per-qid and tot limits take effect (cfg_qid_aqed_active_limit and cfg_aqed_tot_enqueue_limit )
  cfg_detect_feature_0_set [5]  = p2_atq_aqed_act_cnt_upd_v & p2_atq_aqed_act_cnt_upd.cnt[11] ; // Max LSP cfg limit = 12'h800 = 2K
  cfg_detect_feature_0_set [6]  = p3_atq_fid_inflight_cnt_upd_v & cfg_fid_inflight_count_f.cnt[11] ;    // Max LSP cfg limit = 12'h800 = 2K
  cfg_detect_feature_0_set [7]  = p2_dirrpl_enq_cnt_upd_v & p2_dirrpl_enq_cnt_upd.cnt[13] ;     // Limited by 16K shared credits, can't quite get all in one QID and LSP starts sending out immediately, so max is 16K minus delta = bit 13 (count RAM has 15 count bits HQM_LSP_DIRRPL_ENQ_CNT_WIDTH)
  cfg_detect_feature_0_set [8]  = p2_lbrpl_enq_cnt_upd_v & p2_lbrpl_enq_cnt_upd.cnt[13] ;       // Limited by 16K shared credits, can't quite get all in one QID and LSP starts sending out immediately, so max is 16K minus delta = bit 13 (count RAM has 15 count bits HQM_LSP_LBRPL_ENQ_CNT_WIDTH)
  cfg_detect_feature_0_set [9]  = p7_lba_qid_enq_cnt_upd_v & p7_lba_qid_enq_cnt_upd.cnt[14] ;   // Max limit enforced by CHP = 15'h4000 = 16K
  cfg_detect_feature_0_set [10] = p7_lba_cq_tok_cnt_upd_v & p7_lba_cq_tok_cnt_upd_cnt.cnt[10] ; // Max LSP LB CQ depth cfg limit = 11'h400 = 1K
  cfg_detect_feature_0_set [11] = p7_lba_cq_if_cnt_upd_v & p7_lba_cq_if_cnt_upd_cnt.cnt[11] ;   // Max LSP cfg limit = 12'h800 = 2K (hist list)
  cfg_detect_feature_0_set [12] = p7_lba_qid_if_cnt_upd_v & p7_lba_qid_if_cnt_upd.cnt[11] ;     // Max LSP cfg limit = 12'h800 = 2K (max SN)
  // Coverpoint for LB total if count

  cfg_detect_feature_1_set      = 32'h0 ;
  cfg_detect_feature_1_set [0]  = p0_direnq_ctrl_pipe.en & p0_direnq_ctrl_pipe_nxt.blast_enq & ~ p0_direnq_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [1]  = p1_direnq_ctrl_pipe.en & p1_direnq_ctrl_pipe_nxt.blast_enq & ~ p1_direnq_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [2]  = p2_direnq_ctrl_pipe.en & p2_direnq_ctrl_pipe_nxt.blast_enq & ~ p2_direnq_ctrl_pipe_f.blast_enq ;
// Coverpoint for DIR blast_enq at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [3]  = p0_direnq_ctrl_pipe.en & p0_direnq_ctrl_pipe_nxt.blast_tok & ~ p0_direnq_ctrl_pipe_f.blast_tok ;
  cfg_detect_feature_1_set [4]  = p1_direnq_ctrl_pipe.en & p1_direnq_ctrl_pipe_nxt.blast_tok & ~ p1_direnq_ctrl_pipe_f.blast_tok ;
  cfg_detect_feature_1_set [5]  = p2_direnq_ctrl_pipe.en & p2_direnq_ctrl_pipe_nxt.blast_tok & ~ p2_direnq_ctrl_pipe_f.blast_tok ;
// Coverpoint for DIR blast_tok at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [6]  = p0_atq_ctrl_pipe.en & p0_atq_ctrl_pipe_nxt.blast_enq & ~ p0_atq_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [7]  = p1_atq_ctrl_pipe.en & p1_atq_ctrl_pipe_nxt.blast_enq & ~ p1_atq_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [8]  = p2_atq_ctrl_pipe.en & p2_atq_ctrl_pipe_nxt.blast_enq & ~ p2_atq_ctrl_pipe_f.blast_enq ;
// Coverpoint for ATQ blast_enq at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [9]  = p0_atq_ctrl_pipe.en & p0_atq_ctrl_pipe_nxt.blast_cmp & ~ p0_atq_ctrl_pipe_f.blast_cmp ;
  cfg_detect_feature_1_set [10] = p1_atq_ctrl_pipe.en & p1_atq_ctrl_pipe_nxt.blast_cmp & ~ p1_atq_ctrl_pipe_f.blast_cmp ;
  cfg_detect_feature_1_set [11] = p2_atq_ctrl_pipe.en & p2_atq_ctrl_pipe_nxt.blast_cmp & ~ p2_atq_ctrl_pipe_f.blast_cmp ;
// Coverpoint for ATQ blast_cmp at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [12] = p0_lbrpl_ctrl_pipe.en & p0_lbrpl_ctrl_pipe_nxt.blast_enq & ~ p0_lbrpl_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [13] = p1_lbrpl_ctrl_pipe.en & p1_lbrpl_ctrl_pipe_nxt.blast_enq & ~ p1_lbrpl_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [14] = p2_lbrpl_ctrl_pipe.en & p2_lbrpl_ctrl_pipe_nxt.blast_enq & ~ p2_lbrpl_ctrl_pipe_f.blast_enq ;
// Coverpoint for LBRPL blast_enq at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [15] = p0_dirrpl_ctrl_pipe.en & p0_dirrpl_ctrl_pipe_nxt.blast_enq & ~ p0_dirrpl_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [16] = p1_dirrpl_ctrl_pipe.en & p1_dirrpl_ctrl_pipe_nxt.blast_enq & ~ p1_dirrpl_ctrl_pipe_f.blast_enq ;
  cfg_detect_feature_1_set [17] = p2_dirrpl_ctrl_pipe.en & p2_dirrpl_ctrl_pipe_nxt.blast_enq & ~ p2_dirrpl_ctrl_pipe_f.blast_enq ;
// Coverpoint for DIRRPL blast_enq at p2 having an effect - too expensive for feature bit

  cfg_detect_feature_1_set [18] = p0_lba_ctrl_pipe_cmpblast_cond ;
  cfg_detect_feature_1_set [19] = p1_lba_ctrl_pipe_cmpblast_cond &   p1_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p1_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [20] = p1_lba_ctrl_pipe_cmpblast_cond & ~ p1_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p2_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [21] = p2_lba_ctrl_pipe_cmpblast_cond &   p2_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p2_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [22] = p2_lba_ctrl_pipe_cmpblast_cond & ~ p2_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p3_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [23] = p3_lba_ctrl_pipe_cmpblast_cond &   p3_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p3_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [24] = p3_lba_ctrl_pipe_cmpblast_cond & ~ p3_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p4_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [25] = p4_lba_ctrl_pipe_cmpblast_cond &   p4_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p4_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [26] = p4_lba_ctrl_pipe_cmpblast_cond & ~ p4_lba_ctrl_pipe.hold & ~ ( ap_lsp_qidixv == p5_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [27] = p5_lba_ctrl_pipe_cmpblast_cond &                           ~ ( ap_lsp_qidixv == p6_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [28] = p6_lba_ctrl_pipe_cmpblast_cond &                           ~ ( ap_lsp_qidixv == p7_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
  cfg_detect_feature_1_set [29] = p7_lba_ctrl_pipe_cmpblast_cond &                           ~ ( ap_lsp_qidixv == p8_lba_ctrl_pipe_f.sch_cmpblast_qidixv ) ;
end //always

always_comb begin
  cfg_detect_feature_0_nxt              = cfg_detect_feature_0_f | cfg_detect_feature_0_set ;
  cfg_detect_feature_1_nxt              = cfg_detect_feature_1_f | cfg_detect_feature_1_set ;
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    cfg_detect_feature_0_f              <= 32'h0 ;
    cfg_detect_feature_1_f              <= 32'h0 ;
  end
  else begin
    cfg_detect_feature_0_f              <= cfg_detect_feature_0_nxt ;
    cfg_detect_feature_1_f              <= cfg_detect_feature_1_nxt ;
  end
end // always

//-----------------------------------------------------------------------------------------------------
//----
assign cfg_cq_dir_disable_nxt                                   = cfg_cq_dir_disable_f ;
assign hqm_lsp_target_cfg_cq_dir_disable_reg_load               = 1'b0 ;

assign hqm_lsp_target_cfg_cq_dir_disable_reg_nxt                = cfg_cq_dir_disable_nxt ;
assign cfg_cq_dir_disable_f                                     = hqm_lsp_target_cfg_cq_dir_disable_reg_f ;

always_comb begin
  for ( int i = 0 ; i < HQM_NUM_LB_CQ ; i = i + 1 ) begin
    cfg_cq_ldb_disable_f [i]   = hqm_lsp_target_cfg_cq_ldb_disable_reg_f [ ( i * 2 ) +: 1 ] ;                         // TKM
    cfg_cq_ldb_enable_pcm_f [i]   = hqm_lsp_target_cfg_cq_ldb_disable_reg_f [ ( ( i * 2 ) + 1 ) +: 1 ] ;              // TKM
  end // for
end 

assign hqm_lsp_target_cfg_cq_ldb_disable_reg_load               = 1'b0 ;
assign hqm_lsp_target_cfg_cq_ldb_disable_reg_nxt                = hqm_lsp_target_cfg_cq_ldb_disable_reg_f ;
//----
assign p2_lba_inp_tok_cq_disable        = cfg_cq_ldb_disable_f [ p2_lba_ctrl_pipe_f.tok_cq [HQM_NUM_LB_CQB2-1:0] ] |
                                          core_chp_lsp_ldb_cq_off_f [ p2_lba_ctrl_pipe_f.tok_cq [HQM_NUM_LB_CQB2-1:0] ] ;
assign p3_lba_cq2qid_cq_disable         = cfg_cq_ldb_disable_f [ p3_lba_ctrl_pipe_f.sch_cq [HQM_NUM_LB_CQB2-1:0] ] |
                                          core_chp_lsp_ldb_cq_off_f [ p3_lba_ctrl_pipe_f.sch_cq [HQM_NUM_LB_CQB2-1:0] ] ;
assign p7_lba_if_cnt_cq_disable         = cfg_cq_ldb_disable_f [ p7_lba_cq_if_cnt_rmw_pipe_f.cq [HQM_NUM_LB_CQB2-1:0] ] |
                                          core_chp_lsp_ldb_cq_off_f [ p7_lba_cq_if_cnt_rmw_pipe_f.cq [HQM_NUM_LB_CQB2-1:0] ] ;
assign p7_lba_tok_cnt_cq_disable        = cfg_cq_ldb_disable_f [ p7_lba_cq_tok_cnt_rmw_pipe_f.cq [HQM_NUM_LB_CQB2-1:0] ] |
                                          core_chp_lsp_ldb_cq_off_f [ p7_lba_cq_tok_cnt_rmw_pipe_f.cq [HQM_NUM_LB_CQB2-1:0] ] ;

assign p0_direnq_inp_tok_cq_disable     = cfg_cq_dir_disable_f [ p0_direnq_tok_cnt_rmw_pipe_f_pnc.cq [HQM_NUM_DIR_CQB2-1:0] ] ;
assign p2_direnq_enq_cnt_cq_disable     = cfg_cq_dir_disable_f [ p2_direnq_enq_cnt_rmw_pipe_f.qid [HQM_NUM_DIR_CQB2-1:0] ] ;      // Direct mapping of qid to cq
assign p2_direnq_tok_cnt_cq_disable     = cfg_cq_dir_disable_f [ p2_direnq_tok_cnt_rmw_pipe_f.cq [HQM_NUM_DIR_CQB2-1:0] ] ;

//-----------------------------------------------------------------------------------------------------
// SMON

//----
assign hqm_lsp_target_cfg_smon0_disable_smon    = disable_smon ;
assign hqm_lsp_target_cfg_smon0_smon_v          = smon0_v ;
assign hqm_lsp_target_cfg_smon0_smon_comp       = smon0_comp ;
assign hqm_lsp_target_cfg_smon0_smon_val        = smon0_value ;
assign smon_enabled                             = hqm_lsp_target_cfg_smon0_smon_enabled ;
assign smon_interrupt_nc                        = hqm_lsp_target_cfg_smon0_smon_interrupt ;
//----

assign smon_enabled_any                         = smon_enabled ;

always_comb begin
  smon_lsp_dp_sch_dir_v_nxt                     = smon_lsp_dp_sch_dir_v_f ;
  smon_lsp_ap_atm_taken_nxt                     = smon_lsp_ap_atm_taken_f ;
  smon_lsp_ap_atm_stall_nxt                     = smon_lsp_ap_atm_stall_f ;
  smon_atq_sel_ap_stall_nxt                     = smon_atq_sel_ap_stall_f ;
  smon_rpl_dir_dp_stall_nxt                     = smon_rpl_dir_dp_stall_f ;
  smon_rpl_ldb_nalb_stall_nxt                   = smon_rpl_ldb_nalb_stall_f ;
  smon_chp_lsp_token_v_nxt                      = smon_chp_lsp_token_v_f ;
  smon_chp_lsp_cmp_v_nxt                        = smon_chp_lsp_cmp_v_f ;
  smon_rop_lsp_reordercmp_v_nxt                 = smon_rop_lsp_reordercmp_v_f ;
  smon_nalb_lsp_enq_lb_v_nxt                    = smon_nalb_lsp_enq_lb_v_f ;
  smon_dp_lsp_enq_dir_v_nxt                     = smon_dp_lsp_enq_dir_v_f ;
  smon_dp_lsp_enq_rorply_v_nxt                  = smon_dp_lsp_enq_rorply_v_f ;
  smon_send_atm_to_cq_v_nxt                     = smon_send_atm_to_cq_v_f ;
  smon_nalb_lsp_enq_rorply_v_nxt                = smon_nalb_lsp_enq_rorply_v_f ;
  smon_qed_lsp_deq_v_nxt                        = smon_qed_lsp_deq_v_f ;
  smon_aqed_lsp_deq_v_nxt                       = smon_aqed_lsp_deq_v_f ;
  smon_chp_lsp_token_ready_nxt                  = smon_chp_lsp_token_ready_f ;
  smon_chp_lsp_cmp_ready_nxt                    = smon_chp_lsp_cmp_ready_f ;
  smon_rop_lsp_reordercmp_ready_nxt             = smon_rop_lsp_reordercmp_ready_f ;
  smon_nalb_lsp_enq_lb_ready_nxt                = smon_nalb_lsp_enq_lb_ready_f ;
  smon_dp_lsp_enq_dir_ready_nxt                 = smon_dp_lsp_enq_dir_ready_f ;
  smon_dp_lsp_enq_rorply_ready_nxt              = smon_dp_lsp_enq_rorply_ready_f ;
  smon_send_atm_to_cq_ready_nxt                 = smon_send_atm_to_cq_ready_f ;
  smon_nalb_lsp_enq_rorply_ready_nxt            = smon_nalb_lsp_enq_rorply_ready_f ;

  smon_lsp_dp_sch_dir_rdy_nxt                   = smon_lsp_dp_sch_dir_rdy_f ;
  smon_lsp_dp_sch_dir_cm_nxt                    = smon_lsp_dp_sch_dir_cm_f ;
  smon_lsp_dp_sch_dir_wbo_nxt                   = smon_lsp_dp_sch_dir_wbo_f ;
  smon_lsp_dp_sch_dir_cq_nxt                    = smon_lsp_dp_sch_dir_cq_f ;
  smon_lsp_ap_atm_cmd_nxt                       = smon_lsp_ap_atm_cmd_f ;
  smon_lsp_ap_atm_cq_nxt                        = smon_lsp_ap_atm_cq_f ;
  smon_lsp_ap_atm_qid_nxt                       = smon_lsp_ap_atm_qid_f ;
  smon_lsp_ap_atm_fid_nxt                       = smon_lsp_ap_atm_fid_f ;
  smon_lsp_nalb_sch_unoord_cq_nxt               = smon_lsp_nalb_sch_unoord_cq_f ;
  smon_lsp_nalb_sch_unoord_qid_nxt              = smon_lsp_nalb_sch_unoord_qid_f ;
  smon_atq_sel_ap_qid_nxt                       = smon_atq_sel_ap_qid_f ;
  smon_rpl_dir_dp_qid_nxt                       = smon_rpl_dir_dp_qid_f ;
  smon_rpl_ldb_nalb_qid_nxt                     = smon_rpl_ldb_nalb_qid_f ;
  smon_dp_lsp_enq_dir_data_qid_nxt              = smon_dp_lsp_enq_dir_data_qid_f ;
  smon_chp_lsp_token_data_is_ldb_nxt            = smon_chp_lsp_token_data_is_ldb_f ;
  smon_chp_lsp_token_data_cq_nxt                = smon_chp_lsp_token_data_cq_f ;
  smon_chp_lsp_token_data_count_nxt             = smon_chp_lsp_token_data_count_f ;
  smon_nalb_lsp_enq_lb_data_qtype_nxt           = smon_nalb_lsp_enq_lb_data_qtype_f ;
  smon_nalb_lsp_enq_lb_data_qid_nxt             = smon_nalb_lsp_enq_lb_data_qid_f ;
  smon_chp_lsp_cmp_data_qid_nxt                 = smon_chp_lsp_cmp_data_qid_f ;
  smon_chp_lsp_cmp_data_cq_nxt                  = smon_chp_lsp_cmp_data_cq_f ;
  smon_chp_lsp_cmp_data_qtype_nxt               = smon_chp_lsp_cmp_data_qtype_f ;
  smon_chp_lsp_cmp_data_fid_nxt                 = smon_chp_lsp_cmp_data_fid_f ;
  smon_rop_lsp_reordercmp_data_qid_nxt          = smon_rop_lsp_reordercmp_data_qid_f ;
  smon_rop_lsp_reordercmp_data_cq_nxt           = smon_rop_lsp_reordercmp_data_cq_f ;
  smon_dp_lsp_enq_rorply_data_qid_nxt           = smon_dp_lsp_enq_rorply_data_qid_f ;
  smon_nalb_lsp_enq_rorply_data_qid_nxt         = smon_nalb_lsp_enq_rorply_data_qid_f ;
  smon_dp_lsp_enq_rorply_data_frag_cnt_nxt      = smon_dp_lsp_enq_rorply_data_frag_cnt_f ;
  smon_nalb_lsp_enq_rorply_data_frag_cnt_nxt    = smon_nalb_lsp_enq_rorply_data_frag_cnt_f ;
  smon_qed_lsp_deq_data_cq_nxt                  = smon_qed_lsp_deq_data_cq_f ;
  smon_aqed_lsp_deq_data_cq_nxt                 = smon_aqed_lsp_deq_data_cq_f ;

  if ( smon_enabled_any ) begin
    smon_lsp_dp_sch_dir_v_nxt                   = lsp_dp_sch_dir_v ;
    smon_lsp_ap_atm_taken_nxt                   = lsp_ap_atm_v & lsp_ap_atm_ready ;
    smon_lsp_ap_atm_stall_nxt                   = lsp_ap_atm_v & ~ lsp_ap_atm_ready ;
    smon_atq_sel_ap_stall_nxt                   = p3_atq_sch_stall_smon ;
    smon_rpl_dir_dp_stall_nxt                   = p3_dirrpl_sch_stall_smon ;
    smon_rpl_ldb_nalb_stall_nxt                 = p3_lbrpl_sch_stall_smon ;
    smon_chp_lsp_token_v_nxt                    = core_chp_lsp_token_v ;
    smon_chp_lsp_cmp_v_nxt                      = core_chp_lsp_cmp_v ;
    smon_rop_lsp_reordercmp_v_nxt               = core_rop_lsp_reordercmp_v ;
    smon_nalb_lsp_enq_lb_v_nxt                  = core_nalb_lsp_enq_lb_v ;
    smon_dp_lsp_enq_dir_v_nxt                   = core_dp_lsp_enq_dir_v ;
    smon_dp_lsp_enq_rorply_v_nxt                = core_dp_lsp_enq_rorply_v ;
    smon_send_atm_to_cq_v_nxt                   = send_atm_to_cq_v ;
    smon_nalb_lsp_enq_rorply_v_nxt              = core_nalb_lsp_enq_rorply_v ;
    smon_qed_lsp_deq_v_nxt                      = smon_qed_lsp_deq_v ;
    smon_aqed_lsp_deq_v_nxt                     = smon_aqed_lsp_deq_v ;
    smon_chp_lsp_token_ready_nxt                = core_chp_lsp_token_ready ;
    smon_chp_lsp_cmp_ready_nxt                  = core_chp_lsp_cmp_ready ;
    smon_rop_lsp_reordercmp_ready_nxt           = core_rop_lsp_reordercmp_ready ;
    smon_nalb_lsp_enq_lb_ready_nxt              = core_nalb_lsp_enq_lb_ready ;
    smon_dp_lsp_enq_dir_ready_nxt               = core_dp_lsp_enq_dir_ready ;
    smon_dp_lsp_enq_rorply_ready_nxt            = core_dp_lsp_enq_rorply_ready ;
    smon_send_atm_to_cq_ready_nxt               = send_atm_to_cq_ready ;
    smon_nalb_lsp_enq_rorply_ready_nxt          = core_nalb_lsp_enq_rorply_ready ;

    smon_lsp_dp_sch_dir_rdy_nxt                 = lsp_dp_sch_dir_ready ;
    smon_lsp_dp_sch_dir_cm_nxt                  = lsp_dp_sch_dir_data.hqm_core_flags.congestion_management ;
    smon_lsp_dp_sch_dir_wbo_nxt                 = lsp_dp_sch_dir_data.hqm_core_flags.write_buffer_optimization ;
    smon_lsp_dp_sch_dir_cq_nxt                  = lsp_dp_sch_dir_data.cq ;
    smon_lsp_ap_atm_cmd_nxt                     = lsp_ap_atm_data.cmd ;
    smon_lsp_ap_atm_cq_nxt                      = lsp_ap_atm_data.cq [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
    smon_lsp_ap_atm_qid_nxt                     = lsp_ap_atm_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    smon_lsp_ap_atm_fid_nxt                     = lsp_ap_atm_data.fid [HQM_LSP_ARCH_NUM_FIDB2-1:0] ;
    smon_lsp_nalb_sch_unoord_cq_nxt             = nalb_sel_nalb_fifo_pop_data.cq [HQM_LSP_ARCH_NUM_LB_CQB2-1:0] ;
    smon_lsp_nalb_sch_unoord_qid_nxt            = nalb_sel_nalb_fifo_pop_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    smon_atq_sel_ap_qid_nxt                     = atq_sel_ap_db_in_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    smon_rpl_dir_dp_qid_nxt                     = rpl_dir_dp_db_in_data.qid [HQM_LSP_ARCH_NUM_DIR_QIDB2-1:0] ;
    smon_rpl_ldb_nalb_qid_nxt                   = rpl_ldb_nalb_db_in_data.qid [HQM_LSP_ARCH_NUM_LB_QIDB2-1:0] ;
    smon_dp_lsp_enq_dir_data_qid_nxt            = core_dp_lsp_enq_dir_data.qid ;
    smon_chp_lsp_token_data_is_ldb_nxt          = core_chp_lsp_token_data.is_ldb ;
    smon_chp_lsp_token_data_cq_nxt              = core_chp_lsp_token_data.cq ;
    smon_chp_lsp_token_data_count_nxt           = core_chp_lsp_token_data.count ;
    smon_nalb_lsp_enq_lb_data_qtype_nxt         = core_nalb_lsp_enq_lb_data.qtype ;
    smon_nalb_lsp_enq_lb_data_qid_nxt           = core_nalb_lsp_enq_lb_data.qid ;
    smon_chp_lsp_cmp_data_qid_nxt               = core_chp_lsp_cmp_data.qid ;
    smon_chp_lsp_cmp_data_cq_nxt                = core_chp_lsp_cmp_data.pp ;
    smon_chp_lsp_cmp_data_qtype_nxt             = core_chp_lsp_cmp_data.hist_list_info.qtype ;
    smon_chp_lsp_cmp_data_fid_nxt               = core_chp_lsp_cmp_data.hist_list_info.sn_fid.fid ;
    smon_rop_lsp_reordercmp_data_qid_nxt        = core_rop_lsp_reordercmp_data.qid ;
    smon_rop_lsp_reordercmp_data_cq_nxt         = core_rop_lsp_reordercmp_data.cq ;
    smon_dp_lsp_enq_rorply_data_qid_nxt         = core_dp_lsp_enq_rorply_data.qid ;
    smon_nalb_lsp_enq_rorply_data_qid_nxt       = core_nalb_lsp_enq_rorply_data.qid ;
    smon_dp_lsp_enq_rorply_data_frag_cnt_nxt    = core_dp_lsp_enq_rorply_data.frag_cnt ;
    smon_nalb_lsp_enq_rorply_data_frag_cnt_nxt  = core_nalb_lsp_enq_rorply_data.frag_cnt ;
    smon_qed_lsp_deq_data_cq_nxt                = smon_qed_lsp_deq_data_cq ;
    smon_aqed_lsp_deq_data_cq_nxt               = smon_aqed_lsp_deq_data_cq ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    smon_lsp_dp_sch_dir_v_f                     <= 1'b0 ;
    smon_lsp_ap_atm_taken_f                     <= 1'b0 ;
    smon_lsp_ap_atm_stall_f                     <= 1'b0 ;
    smon_atq_sel_ap_stall_f                     <= 1'b0 ;
    smon_rpl_dir_dp_stall_f                     <= 1'b0 ;
    smon_rpl_ldb_nalb_stall_f                   <= 1'b0 ;
    smon_chp_lsp_token_v_f                      <= 1'b0 ;
    smon_chp_lsp_cmp_v_f                        <= 1'b0 ;
    smon_rop_lsp_reordercmp_v_f                 <= 1'b0 ;
    smon_nalb_lsp_enq_lb_v_f                    <= 1'b0 ;
    smon_dp_lsp_enq_dir_v_f                     <= 1'b0 ;
    smon_dp_lsp_enq_rorply_v_f                  <= 1'b0 ;
    smon_send_atm_to_cq_v_f                     <= 1'b0 ;
    smon_nalb_lsp_enq_rorply_v_f                <= 1'b0 ;
    smon_qed_lsp_deq_v_f                        <= 1'b0 ;
    smon_aqed_lsp_deq_v_f                       <= 1'b0 ;
    smon_chp_lsp_token_ready_f                  <= 1'b0 ;
    smon_chp_lsp_cmp_ready_f                    <= 1'b0 ;
    smon_rop_lsp_reordercmp_ready_f             <= 1'b0 ;
    smon_nalb_lsp_enq_lb_ready_f                <= 1'b0 ;
    smon_dp_lsp_enq_dir_ready_f                 <= 1'b0 ;
    smon_dp_lsp_enq_rorply_ready_f              <= 1'b0 ;
    smon_send_atm_to_cq_ready_f                 <= 1'b0 ;
    smon_nalb_lsp_enq_rorply_ready_f            <= 1'b0 ;
  end
  else begin
    smon_lsp_dp_sch_dir_v_f                     <= smon_lsp_dp_sch_dir_v_nxt ;
    smon_lsp_ap_atm_taken_f                     <= smon_lsp_ap_atm_taken_nxt ;
    smon_lsp_ap_atm_stall_f                     <= smon_lsp_ap_atm_stall_nxt ;
    smon_atq_sel_ap_stall_f                     <= smon_atq_sel_ap_stall_nxt ;
    smon_rpl_dir_dp_stall_f                     <= smon_rpl_dir_dp_stall_nxt ;
    smon_rpl_ldb_nalb_stall_f                   <= smon_rpl_ldb_nalb_stall_nxt ;
    smon_chp_lsp_token_v_f                      <= smon_chp_lsp_token_v_nxt ;
    smon_chp_lsp_cmp_v_f                        <= smon_chp_lsp_cmp_v_nxt ;
    smon_rop_lsp_reordercmp_v_f                 <= smon_rop_lsp_reordercmp_v_nxt ;
    smon_nalb_lsp_enq_lb_v_f                    <= smon_nalb_lsp_enq_lb_v_nxt ;
    smon_dp_lsp_enq_dir_v_f                     <= smon_dp_lsp_enq_dir_v_nxt ;
    smon_dp_lsp_enq_rorply_v_f                  <= smon_dp_lsp_enq_rorply_v_nxt ;
    smon_send_atm_to_cq_v_f                     <= smon_send_atm_to_cq_v_nxt ;
    smon_nalb_lsp_enq_rorply_v_f                <= smon_nalb_lsp_enq_rorply_v_nxt ;
    smon_qed_lsp_deq_v_f                        <= smon_qed_lsp_deq_v_nxt ;
    smon_aqed_lsp_deq_v_f                       <= smon_aqed_lsp_deq_v_nxt ;
    smon_chp_lsp_token_ready_f                  <= smon_chp_lsp_token_ready_nxt ;
    smon_chp_lsp_cmp_ready_f                    <= smon_chp_lsp_cmp_ready_nxt ;
    smon_rop_lsp_reordercmp_ready_f             <= smon_rop_lsp_reordercmp_ready_nxt ;
    smon_nalb_lsp_enq_lb_ready_f                <= smon_nalb_lsp_enq_lb_ready_nxt ;
    smon_dp_lsp_enq_dir_ready_f                 <= smon_dp_lsp_enq_dir_ready_nxt ;
    smon_dp_lsp_enq_rorply_ready_f              <= smon_dp_lsp_enq_rorply_ready_nxt ;
    smon_send_atm_to_cq_ready_f                 <= smon_send_atm_to_cq_ready_nxt ;
    smon_nalb_lsp_enq_rorply_ready_f            <= smon_nalb_lsp_enq_rorply_ready_nxt ;
  end
end // always

always_ff @ ( posedge hqm_gated_clk ) begin
  smon_lsp_dp_sch_dir_rdy_f                     <= smon_lsp_dp_sch_dir_rdy_nxt ;
  smon_lsp_dp_sch_dir_cm_f                      <= smon_lsp_dp_sch_dir_cm_nxt ;
  smon_lsp_dp_sch_dir_wbo_f                     <= smon_lsp_dp_sch_dir_wbo_nxt ;
  smon_lsp_dp_sch_dir_cq_f                      <= smon_lsp_dp_sch_dir_cq_nxt ;
  smon_lsp_ap_atm_cmd_f                         <= smon_lsp_ap_atm_cmd_nxt ;
  smon_lsp_ap_atm_cq_f                          <= smon_lsp_ap_atm_cq_nxt ;
  smon_lsp_ap_atm_qid_f                         <= smon_lsp_ap_atm_qid_nxt ;
  smon_lsp_ap_atm_fid_f                         <= smon_lsp_ap_atm_fid_nxt ;
  smon_lsp_nalb_sch_unoord_cq_f                 <= smon_lsp_nalb_sch_unoord_cq_nxt ;
  smon_lsp_nalb_sch_unoord_qid_f                <= smon_lsp_nalb_sch_unoord_qid_nxt ;
  smon_atq_sel_ap_qid_f                         <= smon_atq_sel_ap_qid_nxt ;
  smon_rpl_dir_dp_qid_f                         <= smon_rpl_dir_dp_qid_nxt ;
  smon_rpl_ldb_nalb_qid_f                       <= smon_rpl_ldb_nalb_qid_nxt ;
  smon_dp_lsp_enq_dir_data_qid_f                <= smon_dp_lsp_enq_dir_data_qid_nxt ;
  smon_chp_lsp_token_data_is_ldb_f              <= smon_chp_lsp_token_data_is_ldb_nxt ;
  smon_chp_lsp_token_data_cq_f                  <= smon_chp_lsp_token_data_cq_nxt ;
  smon_chp_lsp_token_data_count_f               <= smon_chp_lsp_token_data_count_nxt ;
  smon_nalb_lsp_enq_lb_data_qtype_f             <= smon_nalb_lsp_enq_lb_data_qtype_nxt ;
  smon_nalb_lsp_enq_lb_data_qid_f               <= smon_nalb_lsp_enq_lb_data_qid_nxt ;
  smon_chp_lsp_cmp_data_qid_f                   <= smon_chp_lsp_cmp_data_qid_nxt ;
  smon_chp_lsp_cmp_data_cq_f                    <= smon_chp_lsp_cmp_data_cq_nxt ;
  smon_chp_lsp_cmp_data_qtype_f                 <= smon_chp_lsp_cmp_data_qtype_nxt ;
  smon_chp_lsp_cmp_data_fid_f                   <= smon_chp_lsp_cmp_data_fid_nxt ;
  smon_rop_lsp_reordercmp_data_qid_f            <= smon_rop_lsp_reordercmp_data_qid_nxt ;
  smon_rop_lsp_reordercmp_data_cq_f             <= smon_rop_lsp_reordercmp_data_cq_nxt ;
  smon_dp_lsp_enq_rorply_data_qid_f             <= smon_dp_lsp_enq_rorply_data_qid_nxt ;
  smon_nalb_lsp_enq_rorply_data_qid_f           <= smon_nalb_lsp_enq_rorply_data_qid_nxt ;
  smon_dp_lsp_enq_rorply_data_frag_cnt_f        <= smon_dp_lsp_enq_rorply_data_frag_cnt_nxt ;
  smon_nalb_lsp_enq_rorply_data_frag_cnt_f      <= smon_nalb_lsp_enq_rorply_data_frag_cnt_nxt ;
  smon_qed_lsp_deq_data_cq_f                    <= smon_qed_lsp_deq_data_cq_nxt ;
  smon_aqed_lsp_deq_data_cq_f                   <= smon_aqed_lsp_deq_data_cq_nxt ;
end // always

assign smon_lsp_ap_atm_sch_rlist        = smon_lsp_ap_atm_taken_f & ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_SCH_RLST ) ;
assign smon_lsp_ap_atm_sch_slist        = smon_lsp_ap_atm_taken_f & ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_SCH_SLST ) ;
assign smon_lsp_ap_atm_sch_stall        = smon_lsp_ap_atm_stall_f & ( ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_SCH_RLST ) |
                                                                      ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_SCH_SLST ) ) ;

assign smon_lsp_dp_sch_dir_taken        = smon_lsp_dp_sch_dir_v_f & smon_lsp_dp_sch_dir_rdy_f ;
assign smon_lsp_dp_sch_dir_stalled      = smon_lsp_dp_sch_dir_v_f & ~ smon_lsp_dp_sch_dir_rdy_f ;

assign smon_chp_lsp_token_taken         = smon_chp_lsp_token_v_f & smon_chp_lsp_token_ready_f ;
assign smon_chp_lsp_cmp_taken           = smon_chp_lsp_cmp_v_f & smon_chp_lsp_cmp_ready_f ;
assign smon_rop_lsp_reordercmp_taken    = smon_rop_lsp_reordercmp_v_f & smon_rop_lsp_reordercmp_ready_f ;
assign smon_nalb_lsp_enq_lb_taken       = smon_nalb_lsp_enq_lb_v_f & smon_nalb_lsp_enq_lb_ready_f ;
assign smon_dp_lsp_enq_dir_taken        = smon_dp_lsp_enq_dir_v_f & smon_dp_lsp_enq_dir_ready_f ;
assign smon_dp_lsp_enq_rorply_taken     = smon_dp_lsp_enq_rorply_v_f & smon_dp_lsp_enq_rorply_ready_f ;
assign smon_send_atm_to_cq_taken        = smon_send_atm_to_cq_v_f & smon_send_atm_to_cq_ready_f ;
assign smon_nalb_lsp_enq_rorply_taken   = smon_nalb_lsp_enq_rorply_v_f & smon_nalb_lsp_enq_rorply_ready_f ;
assign smon_chp_lsp_token_stalled       = smon_chp_lsp_token_v_f & ~ smon_chp_lsp_token_ready_f ;
assign smon_chp_lsp_cmp_stalled         = smon_chp_lsp_cmp_v_f & ~ smon_chp_lsp_cmp_ready_f ;
assign smon_rop_lsp_reordercmp_stalled  = smon_rop_lsp_reordercmp_v_f & ~ smon_rop_lsp_reordercmp_ready_f ;
assign smon_nalb_lsp_enq_lb_stalled     = smon_nalb_lsp_enq_lb_v_f & ~ smon_nalb_lsp_enq_lb_ready_f ;
assign smon_dp_lsp_enq_dir_stalled      = smon_dp_lsp_enq_dir_v_f & ~ smon_dp_lsp_enq_dir_ready_f ;
assign smon_dp_lsp_enq_rorply_stalled   = smon_dp_lsp_enq_rorply_v_f & ~ smon_dp_lsp_enq_rorply_ready_f ;
assign smon_send_atm_to_cq_stalled      = smon_send_atm_to_cq_v_f & ~ smon_send_atm_to_cq_ready_f ;
assign smon_nalb_lsp_enq_rorply_stalled = smon_nalb_lsp_enq_rorply_v_f & ~ smon_nalb_lsp_enq_rorply_ready_f ;

// Note: DB status is registered, so anything conditioned by DB "data" output needs to look at a registered copy of the data
// in order to stay in sync with the DB status trigger condition.
always_comb begin
  smon0_v                               = '0 ;
  smon0_comp                            = '0 ;
  smon0_value                           = '0 ;

  //--------
  // DIR Enqueue
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 0 ]                        = smon_dp_lsp_enq_dir_taken ;
    1'b1 : smon0_v [ 0 ]                        = smon_dp_lsp_enq_dir_stalled ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 0 * 32 +: 32 ]                   = { 25'h0 , smon_dp_lsp_enq_dir_data_qid_f } ;
  smon0_value [ 0 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // Token return
  case ( cfg_smon0_v_sel [1:0] )
    2'h0 : smon0_v [ 1 ]                        = smon_chp_lsp_token_taken ;
    2'h1 : smon0_v [ 1 ]                        = smon_chp_lsp_token_stalled ;
    2'h2 : smon0_v [ 1 ]                        = smon_chp_lsp_token_taken & ( smon_chp_lsp_token_data_is_ldb_f == 1'b0 ) ;
    2'h3 : smon0_v [ 1 ]                        = smon_chp_lsp_token_taken & ( smon_chp_lsp_token_data_is_ldb_f == 1'b1 ) ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 1 * 32 +: 32 ]                   = { 24'h0 , smon_chp_lsp_token_data_cq_f } ;
  case ( cfg_smon0_value_sel )
    1'b0 : smon0_value [ 1 * 32 +: 32 ]         = { 19'h0 , smon_chp_lsp_token_data_count_f } ;
    1'b1 : smon0_value [ 1 * 32 +: 32 ]         = 32'h1 ;
  endcase // cfg_smon0_value_sel
  //--------
  // LB Enqueue
  case ( cfg_smon0_v_sel [1:0] )
    2'h0 : smon0_v [ 2 ]                        = smon_nalb_lsp_enq_lb_taken & ~ ( smon_nalb_lsp_enq_lb_data_qtype_f == DIRECT ) ;
    2'h1 : smon0_v [ 2 ]                        = smon_nalb_lsp_enq_lb_stalled ;
    2'h2 : smon0_v [ 2 ]                        = smon_nalb_lsp_enq_lb_taken & ( ( smon_nalb_lsp_enq_lb_data_qtype_f == ORDERED ) |
                                                                                 ( smon_nalb_lsp_enq_lb_data_qtype_f == UNORDERED ) ) ;
    2'h3 : smon0_v [ 2 ]                        = smon_nalb_lsp_enq_lb_taken & ( smon_nalb_lsp_enq_lb_data_qtype_f == ATOMIC ) ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 2 * 32 +: 32 ]                   = { 25'h0 , smon_nalb_lsp_enq_lb_data_qid_f } ;
  smon0_value [ 2 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // LB Completion
  case ( cfg_smon0_v_sel [1:0] )
    2'h0 : smon0_v [ 3 ]                        = smon_chp_lsp_cmp_taken ;
    2'h1 : smon0_v [ 3 ]                        = smon_chp_lsp_cmp_stalled ;
    2'h2 : smon0_v [ 3 ]                        = smon_chp_lsp_cmp_taken & ( ( smon_chp_lsp_cmp_data_qtype_f == ORDERED ) |
                                                                             ( smon_chp_lsp_cmp_data_qtype_f == UNORDERED ) ) ;
    2'h3 : smon0_v [ 3 ]                        = smon_chp_lsp_cmp_taken &   ( smon_chp_lsp_cmp_data_qtype_f == ATOMIC ) ;
  endcase // cfg_smon0_v_sel
  case ( cfg_smon0_comp_sel [1:0] )
    2'h0 : smon0_comp [ 3 * 32 +: 32 ]          = { 25'h0 , smon_chp_lsp_cmp_data_qid_f } ;
    2'h1 : smon0_comp [ 3 * 32 +: 32 ]          = { 24'h0 , smon_chp_lsp_cmp_data_cq_f } ;
    2'h2 : smon0_comp [ 3 * 32 +: 32 ]          = { 20'h0 , smon_chp_lsp_cmp_data_fid_f } ;
    2'h3 : smon0_comp [ 3 * 32 +: 32 ]          = 32'h0 ;
  endcase // cfg_smon0_comp_sel
  smon0_value [ 3 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // Send ATM to CQ (ATQ -> ATM)
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 4 ]                        = smon_send_atm_to_cq_taken ;
    1'b1 : smon0_v [ 4 ]                        = smon_send_atm_to_cq_stalled ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 4 * 32 +: 32 ]                   = { 25'h0 , send_atm_to_cq_data.qid } ;
  smon0_value [ 4 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // ORD QID Completion
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 5 ]                        = smon_rop_lsp_reordercmp_taken ;
    1'b1 : smon0_v [ 5 ]                        = smon_rop_lsp_reordercmp_stalled ;
  endcase // cfg_smon0_v_sel
  case ( cfg_smon0_comp_sel [0] )
    1'b0 : smon0_comp [ 5 * 32 +: 32 ]          = { 25'h0 , smon_rop_lsp_reordercmp_data_qid_f } ;
    1'b1 : smon0_comp [ 5 * 32 +: 32 ]          = { 24'h0 , smon_rop_lsp_reordercmp_data_cq_f } ;
  endcase // cfg_smon0_comp_sel
  smon0_value [ 5 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // DIR Replay Enqueue
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 6 ]                        = smon_dp_lsp_enq_rorply_taken ;
    1'b1 : smon0_v [ 6 ]                        = smon_dp_lsp_enq_rorply_stalled ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 6 * 32 +: 32 ]                   = { 25'h0 , smon_dp_lsp_enq_rorply_data_qid_f } ;
  case ( cfg_smon0_value_sel )
    1'b0 : smon0_value [ 6 * 32 +: 32 ]         = { 19'h0 , smon_dp_lsp_enq_rorply_data_frag_cnt_f } ;
    1'b1 : smon0_value [ 6 * 32 +: 32 ]         = 32'h1 ;
  endcase // cfg_smon0_value_sel
  //--------
  // LB Replay Enqueue
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 7 ]                        = smon_nalb_lsp_enq_rorply_taken ;
    1'b1 : smon0_v [ 7 ]                        = smon_nalb_lsp_enq_rorply_stalled ;
  endcase // cfg_smon0_v_sel
  smon0_comp [ 7 * 32 +: 32 ]                   = { 25'h0 , smon_nalb_lsp_enq_rorply_data_qid_f } ;
  case ( cfg_smon0_value_sel )
    1'b0 : smon0_value [ 7 * 32 +: 32 ]         = { 17'h0 , smon_nalb_lsp_enq_rorply_data_frag_cnt_f } ;
    1'b1 : smon0_value [ 7 * 32 +: 32 ]         = 32'h1 ;
  endcase // cfg_smon0_value_sel
  //--------
  // NALB Dequeue
  smon0_v [ 8 ]                                 = smon_qed_lsp_deq_v_f ;
  smon0_comp [ 8 * 32 +: 32 ]                   = { 26'h0 , smon_qed_lsp_deq_data_cq_f } ;
  smon0_value [ 8 * 32 +: 32 ]                  = 32'h1 ;
  //--------
  // DIR Schedule
  // Need to do on DB output since wbo function is performed there
  case ( cfg_smon0_v_sel [1:0] )
    2'h0 : smon0_v [ 9 ]                        = smon_lsp_dp_sch_dir_taken ;                                                           // output taken
    2'h1 : smon0_v [ 9 ]                        = smon_lsp_dp_sch_dir_stalled ;                                                         // output stall
    2'h2 : smon0_v [ 9 ]                        = smon_lsp_dp_sch_dir_taken & ( | smon_lsp_dp_sch_dir_wbo_f ) ;                         // any extra beats
    2'h3 : smon0_v [ 9 ]                        = smon_lsp_dp_sch_dir_taken & ( | smon_lsp_dp_sch_dir_cm_f ) ;                          // any type of congestion detected
  endcase // cfg_smon0_v_sel
  smon0_comp [ 9 * 32 +: 32 ]                   = { 24'h0 , smon_lsp_dp_sch_dir_cq_f } ;
  case ( cfg_smon0_value_sel )
    1'b0 : smon0_value [ 9 * 32 +: 32 ]         = 32'h1 ;
    1'b1 : smon0_value [ 9 * 32 +: 32 ]         = { 30'h0 , smon_lsp_dp_sch_dir_wbo_f } ;                                               // total extra beats
  endcase // cfg_smon0_value_sel
  //--------
  // LB Schedule (UNO, ORD, ATM)
  // Combining signals from two independent interfaces - increment amount could be 1 or 2.  No simple way to provide compare, so don't.
  case ( cfg_smon0_v_sel [0] )
    1'b0 : begin
      smon0_v [ 10 ]                            = lsp_nalb_sch_unoord_status_pnc [ 5 ] | smon_lsp_ap_atm_sch_rlist | smon_lsp_ap_atm_sch_slist ;
      smon0_value [ 10 * 32 +: 32 ]             = { 30'h0 , ( { 1'b0 , lsp_nalb_sch_unoord_status_pnc [ 5 ] } + { 1'b0 , ( smon_lsp_ap_atm_sch_rlist | smon_lsp_ap_atm_sch_slist ) } ) } ;
    end
    1'b1 : begin
      smon0_v [ 10 ]                            = lsp_nalb_sch_unoord_status_pnc [ 6 ] | smon_lsp_ap_atm_sch_stall ;
      smon0_value [ 10 * 32 +: 32 ]             = { 30'h0 , ( { 1'b0 , lsp_nalb_sch_unoord_status_pnc [ 6 ] } + { 1'b0 , smon_lsp_ap_atm_sch_stall } ) } ;
    end
  endcase // cfg_smon0_v_sel
  smon0_comp [ 10 * 32 +: 32 ]                  = 32'h0 ;
  //--------
  // ATQ "Schedule" (to AQED qid)
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 11 ]                       = atq_sel_ap_db_status_pnc [ 5 ] ;                                              // Core output taken
    1'b1 : smon0_v [ 11 ]                       = smon_atq_sel_ap_stall_f ;                                                     // Core output stall (v before masked with !rdy)
  endcase // cfg_smon0_v_sel
  smon0_comp [ 11 * 32 +: 32 ]                  = { 25'h0 , smon_atq_sel_ap_qid_f } ;
  smon0_value [ 11 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // ATM Schedule
  case ( cfg_smon0_v_sel [1:0] )
    2'h0 : smon0_v [ 12 ]                       = smon_lsp_ap_atm_sch_rlist | smon_lsp_ap_atm_sch_slist ;
    2'h1 : smon0_v [ 12 ]                       = smon_lsp_ap_atm_sch_stall ;
    2'h2 : smon0_v [ 12 ]                       = smon_lsp_ap_atm_sch_rlist ;
    2'h3 : smon0_v [ 12 ]                       = smon_lsp_ap_atm_sch_slist ;
  endcase // cfg_smon0_v_sel
  case ( cfg_smon0_comp_sel [1:0] )
    2'h0 : smon0_comp [ 12 * 32 +: 32 ]         = { 26'h0 , smon_lsp_ap_atm_cq_f } ;
    2'h1 : smon0_comp [ 12 * 32 +: 32 ]         = { 25'h0 , smon_lsp_ap_atm_qid_f } ;
    2'h2 : smon0_comp [ 12 * 32 +: 32 ]         = 32'h0 ;
    2'h3 : smon0_comp [ 12 * 32 +: 32 ]         = 32'h0 ;
  endcase // cfg_smon0_comp_sel
  smon0_value [ 12 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // ATM Completion
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 13 ]                       = smon_lsp_ap_atm_taken_f & ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_CMP ) ;
    1'b1 : smon0_v [ 13 ]                       = smon_lsp_ap_atm_stall_f & ( smon_lsp_ap_atm_cmd_f == LSP_AP_ATM_CMP ) ;
  endcase // cfg_smon0_v_sel
  case ( cfg_smon0_comp_sel [1:0] )
    2'h0 : smon0_comp [ 13 * 32 +: 32 ]         = { 26'h0 , smon_lsp_ap_atm_cq_f } ;
    2'h1 : smon0_comp [ 13 * 32 +: 32 ]         = { 25'h0 , smon_lsp_ap_atm_qid_f } ;
    2'h2 : smon0_comp [ 13 * 32 +: 32 ]         = { 20'h0 , smon_lsp_ap_atm_fid_f } ;
    2'h3 : smon0_comp [ 13 * 32 +: 32 ]         = 32'h0 ;
  endcase // cfg_smon0_comp_sel
  smon0_value [ 13 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // NALB Schedule (UNO, ORD)
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 14 ]                       = lsp_nalb_sch_unoord_status_pnc [ 5 ] ;                                        // Core output taken
    1'b1 : smon0_v [ 14 ]                       = lsp_nalb_sch_unoord_status_pnc [ 6 ] ;                                        // Core output stall
  endcase // cfg_smon0_v_sel
  case ( cfg_smon0_comp_sel [0] )
    1'b0 : smon0_comp [ 14 * 32 +: 32 ]         = { 26'h0 , smon_lsp_nalb_sch_unoord_cq_f } ;
    1'b1 : smon0_comp [ 14 * 32 +: 32 ]         = { 25'h0 , smon_lsp_nalb_sch_unoord_qid_f } ;
  endcase // cfg_smon0_comp_sel
  smon0_value [ 14 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // DIR Replay Schedule
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 15 ]                       = rpl_dir_dp_db_status_pnc [ 5 ] ;                                              // Core output taken
    1'b1 : smon0_v [ 15 ]                       = smon_rpl_dir_dp_stall_f ;                                                     // Core output stall (v before masked with !rdy)
  endcase // cfg_smon0_v_sel
  smon0_comp [ 15 * 32 +: 32 ]                  = { 25'h0 , smon_rpl_dir_dp_qid_f } ;
  smon0_value [ 15 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // LB Replay Schedule
  case ( cfg_smon0_v_sel [0] )
    1'b0 : smon0_v [ 16 ]                       = rpl_ldb_nalb_db_status_pnc [ 5 ] ;                                            // Core output taken
    1'b1 : smon0_v [ 16 ]                       = smon_rpl_ldb_nalb_stall_f ;                                                   // Core output stall (v before masked with !rdy)
  endcase // cfg_smon0_v_sel
  smon0_comp [ 16 * 32 +: 32 ]                  = { 25'h0 , smon_rpl_ldb_nalb_qid_f } ;
  smon0_value [ 16 * 32 +: 32 ]                 = 32'h1 ;
  //--------
  // ATM Dequeue
  smon0_v [ 17 ]                                = smon_aqed_lsp_deq_v_f ;
  smon0_comp [ 17 * 32 +: 32 ]                  = { 26'h0 , smon_aqed_lsp_deq_data_cq_f } ;
  smon0_value [ 17 * 32 +: 32 ]                 = 32'h1 ;

end // always

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: Agitate
//-----------------------------------------------------------------------------------------------------

assign cfg_agitate_control_nxt                  = cfg_agitate_control_f ;
assign cfg_agitate_select_nxt                   = cfg_agitate_select_f ;

//----
assign hqm_lsp_target_cfg_hw_agitate_control_reg_v              = 1'b0 ;
assign hqm_lsp_target_cfg_hw_agitate_control_reg_nxt            = cfg_agitate_control_nxt ;
assign cfg_agitate_control_f                                    = hqm_lsp_target_cfg_hw_agitate_control_reg_f ;

assign hqm_lsp_target_cfg_hw_agitate_select_reg_v               = 1'b0 ;
assign hqm_lsp_target_cfg_hw_agitate_select_reg_nxt             = cfg_agitate_select_nxt ;
assign cfg_agitate_select_f                                     = hqm_lsp_target_cfg_hw_agitate_select_reg_f ;
//----

// Removed agitator in potential critical path for p0_lba_cq_arb_winner_v and p0_lba_sch_state_ready_for_work.
// May want to reinstate if plenty of margin.  Previous bit 12 of agitate_select

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: To be deleted / renamed
//-----------------------------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: Config regs reserved for future use
//-----------------------------------------------------------------------------------------------------

//*****************************************************************************************************
//*****************************************************************************************************
// SECTION: Misc
//*****************************************************************************************************
//*****************************************************************************************************

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: lsp_atm_pipe
//-----------------------------------------------------------------------------------------------------

hqm_lsp_atm_pipe i_hqm_lsp_atm_pipe (

// lsp_atm_pipe top level interface
  .hqm_gated_clk ( hqm_gated_clk )
, .hqm_gated_rst_b ( hqm_gated_rst_b_atm )
, .hqm_inp_gated_clk ( hqm_inp_gated_clk )
, .hqm_inp_gated_rst_b ( hqm_inp_gated_rst_b_atm )
, .hqm_flr_prep ( hqm_rst_prep_atm )
, .hqm_proc_clk_en ( ap_hqm_proc_clk_en_nc )    // Would only be needed if lsp_atm_pipe had its own clock controller

, .hqm_gated_rst_b_start_atm ( hqm_gated_rst_b_start_atm )
, .hqm_gated_rst_b_active_atm ( hqm_gated_rst_b_active_atm )
, .hqm_gated_rst_b_done_atm ( hqm_gated_rst_b_done_atm )

, .atm_clk_idle ( atm_clk_idle )                // Includes AP input idle (unlike ap_unit_idle, which does not)
, .atm_clk_enable ( atm_clk_enable )

, .ap_unit_idle ( ap_unit_idle )
, .ap_unit_pipeidle ( ap_unit_pipeidle )
, .ap_reset_done ( ap_reset_done )

, .ap_cfg_req_up_read ( ap_cfg_req_up_read )
, .ap_cfg_req_up_write ( ap_cfg_req_up_write )
, .ap_cfg_req_up ( ap_cfg_req_up )
, .ap_cfg_rsp_up_ack ( ap_cfg_rsp_up_ack )
, .ap_cfg_rsp_up ( ap_cfg_rsp_up )
, .ap_cfg_req_down_read ( ap_cfg_req_down_read )
, .ap_cfg_req_down_write ( ap_cfg_req_down_write )
, .ap_cfg_req_down ( ap_cfg_req_down )
, .ap_cfg_rsp_down_ack ( ap_cfg_rsp_down_ack )
, .ap_cfg_rsp_down ( ap_cfg_rsp_down )

, .ap_alarm_up_v ( ap_alarm_up_v )
, .ap_alarm_up_ready ( ap_alarm_up_ready )
, .ap_alarm_up_data ( ap_alarm_up_data )

, .ap_alarm_down_v ( ap_alarm_down_v )
, .ap_alarm_down_ready ( ap_alarm_down_ready )
, .ap_alarm_down_data ( ap_alarm_down_data )

, .lsp_aqed_cmp_v ( lsp_aqed_cmp_v )
, .lsp_aqed_cmp_ready ( lsp_aqed_cmp_ready )
, .lsp_aqed_cmp_data ( lsp_aqed_cmp_data )

, .ap_aqed_v ( ap_aqed_v )
, .ap_aqed_ready ( ap_aqed_ready )
, .ap_aqed_data ( ap_aqed_data )

, .aqed_ap_enq_v ( aqed_ap_enq_v )
, .aqed_ap_enq_ready ( aqed_ap_enq_ready )
, .aqed_ap_enq_data ( aqed_ap_enq_data )

// lsp_atm_pipe to list_sel_pipe interface - no longer used, but extremely useful for debugging / accounting
, .ap_lsp_enq_v ( ap_lsp_enq_v_nc )
, .ap_lsp_enq_ready ( 1'b1 )
, .ap_lsp_enq_data ( ap_lsp_enq_data_nc )

, .lsp_ap_atm_v ( lsp_ap_atm_v )
, .lsp_ap_atm_ready ( lsp_ap_atm_ready )
, .lsp_ap_atm_data ( lsp_ap_atm_data )

, .ap_lsp_freeze ( ap_lsp_freeze )
, .lsp_ap_idle ( cfg_unit_idle_f.pipe_idle )

, .credit_fifo_ap_aqed_dec_sch ( credit_fifo_ap_aqed_dec_sch )
, .credit_fifo_ap_aqed_dec_cmp ( credit_fifo_ap_aqed_dec_cmp )

, .ap_lsp_haswork_slst_v ( ap_lsp_haswork_slst_v )
, .ap_lsp_haswork_slst_func ( ap_lsp_haswork_slst_func )

, .ap_lsp_haswork_rlst_v ( ap_lsp_haswork_rlst_v )
, .ap_lsp_haswork_rlst_func ( ap_lsp_haswork_rlst_func )

, .ap_lsp_cmpblast_v ( ap_lsp_cmpblast_v )
, .ap_lsp_dec_fid_cnt_v ( ap_lsp_dec_fid_cnt_v_nc )

, .ap_lsp_cmd_v ( ap_lsp_cmd_v )
, .ap_lsp_cmd ( ap_lsp_cmd )

, .ap_lsp_qidix_msb ( ap_lsp_qidix_msb )
, .ap_lsp_qidix ( ap_lsp_qidix )
, .ap_lsp_cq ( ap_lsp_cq )
, .ap_lsp_qid ( ap_lsp_qid_nc )
, .ap_lsp_qid2cqqidix ( ap_lsp_qid2cqqidix )

// lsp_atm_pipe top level RAM interface

// BEGIN HQM_MEMPORT_INST hqm_lsp_atm_pipe
    ,.rf_aqed_qid2cqidix_re                             (rf_aqed_qid2cqidix_re)
    ,.rf_aqed_qid2cqidix_rclk                           (rf_aqed_qid2cqidix_rclk)
    ,.rf_aqed_qid2cqidix_rclk_rst_n                     (rf_aqed_qid2cqidix_rclk_rst_n)
    ,.rf_aqed_qid2cqidix_raddr                          (rf_aqed_qid2cqidix_raddr)
    ,.rf_aqed_qid2cqidix_waddr                          (rf_aqed_qid2cqidix_waddr)
    ,.rf_aqed_qid2cqidix_we                             (rf_aqed_qid2cqidix_we)
    ,.rf_aqed_qid2cqidix_wclk                           (rf_aqed_qid2cqidix_wclk)
    ,.rf_aqed_qid2cqidix_wclk_rst_n                     (rf_aqed_qid2cqidix_wclk_rst_n)
    ,.rf_aqed_qid2cqidix_wdata                          (rf_aqed_qid2cqidix_wdata)
    ,.rf_aqed_qid2cqidix_rdata                          (rf_aqed_qid2cqidix_rdata)

    ,.rf_atm_fifo_ap_aqed_re                            (rf_atm_fifo_ap_aqed_re)
    ,.rf_atm_fifo_ap_aqed_rclk                          (rf_atm_fifo_ap_aqed_rclk)
    ,.rf_atm_fifo_ap_aqed_rclk_rst_n                    (rf_atm_fifo_ap_aqed_rclk_rst_n)
    ,.rf_atm_fifo_ap_aqed_raddr                         (rf_atm_fifo_ap_aqed_raddr)
    ,.rf_atm_fifo_ap_aqed_waddr                         (rf_atm_fifo_ap_aqed_waddr)
    ,.rf_atm_fifo_ap_aqed_we                            (rf_atm_fifo_ap_aqed_we)
    ,.rf_atm_fifo_ap_aqed_wclk                          (rf_atm_fifo_ap_aqed_wclk)
    ,.rf_atm_fifo_ap_aqed_wclk_rst_n                    (rf_atm_fifo_ap_aqed_wclk_rst_n)
    ,.rf_atm_fifo_ap_aqed_wdata                         (rf_atm_fifo_ap_aqed_wdata)
    ,.rf_atm_fifo_ap_aqed_rdata                         (rf_atm_fifo_ap_aqed_rdata)

    ,.rf_atm_fifo_aqed_ap_enq_re                        (rf_atm_fifo_aqed_ap_enq_re)
    ,.rf_atm_fifo_aqed_ap_enq_rclk                      (rf_atm_fifo_aqed_ap_enq_rclk)
    ,.rf_atm_fifo_aqed_ap_enq_rclk_rst_n                (rf_atm_fifo_aqed_ap_enq_rclk_rst_n)
    ,.rf_atm_fifo_aqed_ap_enq_raddr                     (rf_atm_fifo_aqed_ap_enq_raddr)
    ,.rf_atm_fifo_aqed_ap_enq_waddr                     (rf_atm_fifo_aqed_ap_enq_waddr)
    ,.rf_atm_fifo_aqed_ap_enq_we                        (rf_atm_fifo_aqed_ap_enq_we)
    ,.rf_atm_fifo_aqed_ap_enq_wclk                      (rf_atm_fifo_aqed_ap_enq_wclk)
    ,.rf_atm_fifo_aqed_ap_enq_wclk_rst_n                (rf_atm_fifo_aqed_ap_enq_wclk_rst_n)
    ,.rf_atm_fifo_aqed_ap_enq_wdata                     (rf_atm_fifo_aqed_ap_enq_wdata)
    ,.rf_atm_fifo_aqed_ap_enq_rdata                     (rf_atm_fifo_aqed_ap_enq_rdata)

    ,.rf_fid2cqqidix_re                                 (rf_fid2cqqidix_re)
    ,.rf_fid2cqqidix_rclk                               (rf_fid2cqqidix_rclk)
    ,.rf_fid2cqqidix_rclk_rst_n                         (rf_fid2cqqidix_rclk_rst_n)
    ,.rf_fid2cqqidix_raddr                              (rf_fid2cqqidix_raddr)
    ,.rf_fid2cqqidix_waddr                              (rf_fid2cqqidix_waddr)
    ,.rf_fid2cqqidix_we                                 (rf_fid2cqqidix_we)
    ,.rf_fid2cqqidix_wclk                               (rf_fid2cqqidix_wclk)
    ,.rf_fid2cqqidix_wclk_rst_n                         (rf_fid2cqqidix_wclk_rst_n)
    ,.rf_fid2cqqidix_wdata                              (rf_fid2cqqidix_wdata)
    ,.rf_fid2cqqidix_rdata                              (rf_fid2cqqidix_rdata)

    ,.rf_ll_enq_cnt_r_bin0_dup0_re                      (rf_ll_enq_cnt_r_bin0_dup0_re)
    ,.rf_ll_enq_cnt_r_bin0_dup0_rclk                    (rf_ll_enq_cnt_r_bin0_dup0_rclk)
    ,.rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup0_raddr                   (rf_ll_enq_cnt_r_bin0_dup0_raddr)
    ,.rf_ll_enq_cnt_r_bin0_dup0_waddr                   (rf_ll_enq_cnt_r_bin0_dup0_waddr)
    ,.rf_ll_enq_cnt_r_bin0_dup0_we                      (rf_ll_enq_cnt_r_bin0_dup0_we)
    ,.rf_ll_enq_cnt_r_bin0_dup0_wclk                    (rf_ll_enq_cnt_r_bin0_dup0_wclk)
    ,.rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup0_wdata                   (rf_ll_enq_cnt_r_bin0_dup0_wdata)
    ,.rf_ll_enq_cnt_r_bin0_dup0_rdata                   (rf_ll_enq_cnt_r_bin0_dup0_rdata)

    ,.rf_ll_enq_cnt_r_bin0_dup1_re                      (rf_ll_enq_cnt_r_bin0_dup1_re)
    ,.rf_ll_enq_cnt_r_bin0_dup1_rclk                    (rf_ll_enq_cnt_r_bin0_dup1_rclk)
    ,.rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup1_raddr                   (rf_ll_enq_cnt_r_bin0_dup1_raddr)
    ,.rf_ll_enq_cnt_r_bin0_dup1_waddr                   (rf_ll_enq_cnt_r_bin0_dup1_waddr)
    ,.rf_ll_enq_cnt_r_bin0_dup1_we                      (rf_ll_enq_cnt_r_bin0_dup1_we)
    ,.rf_ll_enq_cnt_r_bin0_dup1_wclk                    (rf_ll_enq_cnt_r_bin0_dup1_wclk)
    ,.rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup1_wdata                   (rf_ll_enq_cnt_r_bin0_dup1_wdata)
    ,.rf_ll_enq_cnt_r_bin0_dup1_rdata                   (rf_ll_enq_cnt_r_bin0_dup1_rdata)

    ,.rf_ll_enq_cnt_r_bin0_dup2_re                      (rf_ll_enq_cnt_r_bin0_dup2_re)
    ,.rf_ll_enq_cnt_r_bin0_dup2_rclk                    (rf_ll_enq_cnt_r_bin0_dup2_rclk)
    ,.rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup2_raddr                   (rf_ll_enq_cnt_r_bin0_dup2_raddr)
    ,.rf_ll_enq_cnt_r_bin0_dup2_waddr                   (rf_ll_enq_cnt_r_bin0_dup2_waddr)
    ,.rf_ll_enq_cnt_r_bin0_dup2_we                      (rf_ll_enq_cnt_r_bin0_dup2_we)
    ,.rf_ll_enq_cnt_r_bin0_dup2_wclk                    (rf_ll_enq_cnt_r_bin0_dup2_wclk)
    ,.rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup2_wdata                   (rf_ll_enq_cnt_r_bin0_dup2_wdata)
    ,.rf_ll_enq_cnt_r_bin0_dup2_rdata                   (rf_ll_enq_cnt_r_bin0_dup2_rdata)

    ,.rf_ll_enq_cnt_r_bin0_dup3_re                      (rf_ll_enq_cnt_r_bin0_dup3_re)
    ,.rf_ll_enq_cnt_r_bin0_dup3_rclk                    (rf_ll_enq_cnt_r_bin0_dup3_rclk)
    ,.rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup3_raddr                   (rf_ll_enq_cnt_r_bin0_dup3_raddr)
    ,.rf_ll_enq_cnt_r_bin0_dup3_waddr                   (rf_ll_enq_cnt_r_bin0_dup3_waddr)
    ,.rf_ll_enq_cnt_r_bin0_dup3_we                      (rf_ll_enq_cnt_r_bin0_dup3_we)
    ,.rf_ll_enq_cnt_r_bin0_dup3_wclk                    (rf_ll_enq_cnt_r_bin0_dup3_wclk)
    ,.rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n              (rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin0_dup3_wdata                   (rf_ll_enq_cnt_r_bin0_dup3_wdata)
    ,.rf_ll_enq_cnt_r_bin0_dup3_rdata                   (rf_ll_enq_cnt_r_bin0_dup3_rdata)

    ,.rf_ll_enq_cnt_r_bin1_dup0_re                      (rf_ll_enq_cnt_r_bin1_dup0_re)
    ,.rf_ll_enq_cnt_r_bin1_dup0_rclk                    (rf_ll_enq_cnt_r_bin1_dup0_rclk)
    ,.rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup0_raddr                   (rf_ll_enq_cnt_r_bin1_dup0_raddr)
    ,.rf_ll_enq_cnt_r_bin1_dup0_waddr                   (rf_ll_enq_cnt_r_bin1_dup0_waddr)
    ,.rf_ll_enq_cnt_r_bin1_dup0_we                      (rf_ll_enq_cnt_r_bin1_dup0_we)
    ,.rf_ll_enq_cnt_r_bin1_dup0_wclk                    (rf_ll_enq_cnt_r_bin1_dup0_wclk)
    ,.rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup0_wdata                   (rf_ll_enq_cnt_r_bin1_dup0_wdata)
    ,.rf_ll_enq_cnt_r_bin1_dup0_rdata                   (rf_ll_enq_cnt_r_bin1_dup0_rdata)

    ,.rf_ll_enq_cnt_r_bin1_dup1_re                      (rf_ll_enq_cnt_r_bin1_dup1_re)
    ,.rf_ll_enq_cnt_r_bin1_dup1_rclk                    (rf_ll_enq_cnt_r_bin1_dup1_rclk)
    ,.rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup1_raddr                   (rf_ll_enq_cnt_r_bin1_dup1_raddr)
    ,.rf_ll_enq_cnt_r_bin1_dup1_waddr                   (rf_ll_enq_cnt_r_bin1_dup1_waddr)
    ,.rf_ll_enq_cnt_r_bin1_dup1_we                      (rf_ll_enq_cnt_r_bin1_dup1_we)
    ,.rf_ll_enq_cnt_r_bin1_dup1_wclk                    (rf_ll_enq_cnt_r_bin1_dup1_wclk)
    ,.rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup1_wdata                   (rf_ll_enq_cnt_r_bin1_dup1_wdata)
    ,.rf_ll_enq_cnt_r_bin1_dup1_rdata                   (rf_ll_enq_cnt_r_bin1_dup1_rdata)

    ,.rf_ll_enq_cnt_r_bin1_dup2_re                      (rf_ll_enq_cnt_r_bin1_dup2_re)
    ,.rf_ll_enq_cnt_r_bin1_dup2_rclk                    (rf_ll_enq_cnt_r_bin1_dup2_rclk)
    ,.rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup2_raddr                   (rf_ll_enq_cnt_r_bin1_dup2_raddr)
    ,.rf_ll_enq_cnt_r_bin1_dup2_waddr                   (rf_ll_enq_cnt_r_bin1_dup2_waddr)
    ,.rf_ll_enq_cnt_r_bin1_dup2_we                      (rf_ll_enq_cnt_r_bin1_dup2_we)
    ,.rf_ll_enq_cnt_r_bin1_dup2_wclk                    (rf_ll_enq_cnt_r_bin1_dup2_wclk)
    ,.rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup2_wdata                   (rf_ll_enq_cnt_r_bin1_dup2_wdata)
    ,.rf_ll_enq_cnt_r_bin1_dup2_rdata                   (rf_ll_enq_cnt_r_bin1_dup2_rdata)

    ,.rf_ll_enq_cnt_r_bin1_dup3_re                      (rf_ll_enq_cnt_r_bin1_dup3_re)
    ,.rf_ll_enq_cnt_r_bin1_dup3_rclk                    (rf_ll_enq_cnt_r_bin1_dup3_rclk)
    ,.rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup3_raddr                   (rf_ll_enq_cnt_r_bin1_dup3_raddr)
    ,.rf_ll_enq_cnt_r_bin1_dup3_waddr                   (rf_ll_enq_cnt_r_bin1_dup3_waddr)
    ,.rf_ll_enq_cnt_r_bin1_dup3_we                      (rf_ll_enq_cnt_r_bin1_dup3_we)
    ,.rf_ll_enq_cnt_r_bin1_dup3_wclk                    (rf_ll_enq_cnt_r_bin1_dup3_wclk)
    ,.rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n              (rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin1_dup3_wdata                   (rf_ll_enq_cnt_r_bin1_dup3_wdata)
    ,.rf_ll_enq_cnt_r_bin1_dup3_rdata                   (rf_ll_enq_cnt_r_bin1_dup3_rdata)

    ,.rf_ll_enq_cnt_r_bin2_dup0_re                      (rf_ll_enq_cnt_r_bin2_dup0_re)
    ,.rf_ll_enq_cnt_r_bin2_dup0_rclk                    (rf_ll_enq_cnt_r_bin2_dup0_rclk)
    ,.rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup0_raddr                   (rf_ll_enq_cnt_r_bin2_dup0_raddr)
    ,.rf_ll_enq_cnt_r_bin2_dup0_waddr                   (rf_ll_enq_cnt_r_bin2_dup0_waddr)
    ,.rf_ll_enq_cnt_r_bin2_dup0_we                      (rf_ll_enq_cnt_r_bin2_dup0_we)
    ,.rf_ll_enq_cnt_r_bin2_dup0_wclk                    (rf_ll_enq_cnt_r_bin2_dup0_wclk)
    ,.rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup0_wdata                   (rf_ll_enq_cnt_r_bin2_dup0_wdata)
    ,.rf_ll_enq_cnt_r_bin2_dup0_rdata                   (rf_ll_enq_cnt_r_bin2_dup0_rdata)

    ,.rf_ll_enq_cnt_r_bin2_dup1_re                      (rf_ll_enq_cnt_r_bin2_dup1_re)
    ,.rf_ll_enq_cnt_r_bin2_dup1_rclk                    (rf_ll_enq_cnt_r_bin2_dup1_rclk)
    ,.rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup1_raddr                   (rf_ll_enq_cnt_r_bin2_dup1_raddr)
    ,.rf_ll_enq_cnt_r_bin2_dup1_waddr                   (rf_ll_enq_cnt_r_bin2_dup1_waddr)
    ,.rf_ll_enq_cnt_r_bin2_dup1_we                      (rf_ll_enq_cnt_r_bin2_dup1_we)
    ,.rf_ll_enq_cnt_r_bin2_dup1_wclk                    (rf_ll_enq_cnt_r_bin2_dup1_wclk)
    ,.rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup1_wdata                   (rf_ll_enq_cnt_r_bin2_dup1_wdata)
    ,.rf_ll_enq_cnt_r_bin2_dup1_rdata                   (rf_ll_enq_cnt_r_bin2_dup1_rdata)

    ,.rf_ll_enq_cnt_r_bin2_dup2_re                      (rf_ll_enq_cnt_r_bin2_dup2_re)
    ,.rf_ll_enq_cnt_r_bin2_dup2_rclk                    (rf_ll_enq_cnt_r_bin2_dup2_rclk)
    ,.rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup2_raddr                   (rf_ll_enq_cnt_r_bin2_dup2_raddr)
    ,.rf_ll_enq_cnt_r_bin2_dup2_waddr                   (rf_ll_enq_cnt_r_bin2_dup2_waddr)
    ,.rf_ll_enq_cnt_r_bin2_dup2_we                      (rf_ll_enq_cnt_r_bin2_dup2_we)
    ,.rf_ll_enq_cnt_r_bin2_dup2_wclk                    (rf_ll_enq_cnt_r_bin2_dup2_wclk)
    ,.rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup2_wdata                   (rf_ll_enq_cnt_r_bin2_dup2_wdata)
    ,.rf_ll_enq_cnt_r_bin2_dup2_rdata                   (rf_ll_enq_cnt_r_bin2_dup2_rdata)

    ,.rf_ll_enq_cnt_r_bin2_dup3_re                      (rf_ll_enq_cnt_r_bin2_dup3_re)
    ,.rf_ll_enq_cnt_r_bin2_dup3_rclk                    (rf_ll_enq_cnt_r_bin2_dup3_rclk)
    ,.rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup3_raddr                   (rf_ll_enq_cnt_r_bin2_dup3_raddr)
    ,.rf_ll_enq_cnt_r_bin2_dup3_waddr                   (rf_ll_enq_cnt_r_bin2_dup3_waddr)
    ,.rf_ll_enq_cnt_r_bin2_dup3_we                      (rf_ll_enq_cnt_r_bin2_dup3_we)
    ,.rf_ll_enq_cnt_r_bin2_dup3_wclk                    (rf_ll_enq_cnt_r_bin2_dup3_wclk)
    ,.rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n              (rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin2_dup3_wdata                   (rf_ll_enq_cnt_r_bin2_dup3_wdata)
    ,.rf_ll_enq_cnt_r_bin2_dup3_rdata                   (rf_ll_enq_cnt_r_bin2_dup3_rdata)

    ,.rf_ll_enq_cnt_r_bin3_dup0_re                      (rf_ll_enq_cnt_r_bin3_dup0_re)
    ,.rf_ll_enq_cnt_r_bin3_dup0_rclk                    (rf_ll_enq_cnt_r_bin3_dup0_rclk)
    ,.rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup0_raddr                   (rf_ll_enq_cnt_r_bin3_dup0_raddr)
    ,.rf_ll_enq_cnt_r_bin3_dup0_waddr                   (rf_ll_enq_cnt_r_bin3_dup0_waddr)
    ,.rf_ll_enq_cnt_r_bin3_dup0_we                      (rf_ll_enq_cnt_r_bin3_dup0_we)
    ,.rf_ll_enq_cnt_r_bin3_dup0_wclk                    (rf_ll_enq_cnt_r_bin3_dup0_wclk)
    ,.rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup0_wdata                   (rf_ll_enq_cnt_r_bin3_dup0_wdata)
    ,.rf_ll_enq_cnt_r_bin3_dup0_rdata                   (rf_ll_enq_cnt_r_bin3_dup0_rdata)

    ,.rf_ll_enq_cnt_r_bin3_dup1_re                      (rf_ll_enq_cnt_r_bin3_dup1_re)
    ,.rf_ll_enq_cnt_r_bin3_dup1_rclk                    (rf_ll_enq_cnt_r_bin3_dup1_rclk)
    ,.rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup1_raddr                   (rf_ll_enq_cnt_r_bin3_dup1_raddr)
    ,.rf_ll_enq_cnt_r_bin3_dup1_waddr                   (rf_ll_enq_cnt_r_bin3_dup1_waddr)
    ,.rf_ll_enq_cnt_r_bin3_dup1_we                      (rf_ll_enq_cnt_r_bin3_dup1_we)
    ,.rf_ll_enq_cnt_r_bin3_dup1_wclk                    (rf_ll_enq_cnt_r_bin3_dup1_wclk)
    ,.rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup1_wdata                   (rf_ll_enq_cnt_r_bin3_dup1_wdata)
    ,.rf_ll_enq_cnt_r_bin3_dup1_rdata                   (rf_ll_enq_cnt_r_bin3_dup1_rdata)

    ,.rf_ll_enq_cnt_r_bin3_dup2_re                      (rf_ll_enq_cnt_r_bin3_dup2_re)
    ,.rf_ll_enq_cnt_r_bin3_dup2_rclk                    (rf_ll_enq_cnt_r_bin3_dup2_rclk)
    ,.rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup2_raddr                   (rf_ll_enq_cnt_r_bin3_dup2_raddr)
    ,.rf_ll_enq_cnt_r_bin3_dup2_waddr                   (rf_ll_enq_cnt_r_bin3_dup2_waddr)
    ,.rf_ll_enq_cnt_r_bin3_dup2_we                      (rf_ll_enq_cnt_r_bin3_dup2_we)
    ,.rf_ll_enq_cnt_r_bin3_dup2_wclk                    (rf_ll_enq_cnt_r_bin3_dup2_wclk)
    ,.rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup2_wdata                   (rf_ll_enq_cnt_r_bin3_dup2_wdata)
    ,.rf_ll_enq_cnt_r_bin3_dup2_rdata                   (rf_ll_enq_cnt_r_bin3_dup2_rdata)

    ,.rf_ll_enq_cnt_r_bin3_dup3_re                      (rf_ll_enq_cnt_r_bin3_dup3_re)
    ,.rf_ll_enq_cnt_r_bin3_dup3_rclk                    (rf_ll_enq_cnt_r_bin3_dup3_rclk)
    ,.rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup3_raddr                   (rf_ll_enq_cnt_r_bin3_dup3_raddr)
    ,.rf_ll_enq_cnt_r_bin3_dup3_waddr                   (rf_ll_enq_cnt_r_bin3_dup3_waddr)
    ,.rf_ll_enq_cnt_r_bin3_dup3_we                      (rf_ll_enq_cnt_r_bin3_dup3_we)
    ,.rf_ll_enq_cnt_r_bin3_dup3_wclk                    (rf_ll_enq_cnt_r_bin3_dup3_wclk)
    ,.rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n              (rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n)
    ,.rf_ll_enq_cnt_r_bin3_dup3_wdata                   (rf_ll_enq_cnt_r_bin3_dup3_wdata)
    ,.rf_ll_enq_cnt_r_bin3_dup3_rdata                   (rf_ll_enq_cnt_r_bin3_dup3_rdata)

    ,.rf_ll_enq_cnt_s_bin0_re                           (rf_ll_enq_cnt_s_bin0_re)
    ,.rf_ll_enq_cnt_s_bin0_rclk                         (rf_ll_enq_cnt_s_bin0_rclk)
    ,.rf_ll_enq_cnt_s_bin0_rclk_rst_n                   (rf_ll_enq_cnt_s_bin0_rclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin0_raddr                        (rf_ll_enq_cnt_s_bin0_raddr)
    ,.rf_ll_enq_cnt_s_bin0_waddr                        (rf_ll_enq_cnt_s_bin0_waddr)
    ,.rf_ll_enq_cnt_s_bin0_we                           (rf_ll_enq_cnt_s_bin0_we)
    ,.rf_ll_enq_cnt_s_bin0_wclk                         (rf_ll_enq_cnt_s_bin0_wclk)
    ,.rf_ll_enq_cnt_s_bin0_wclk_rst_n                   (rf_ll_enq_cnt_s_bin0_wclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin0_wdata                        (rf_ll_enq_cnt_s_bin0_wdata)
    ,.rf_ll_enq_cnt_s_bin0_rdata                        (rf_ll_enq_cnt_s_bin0_rdata)

    ,.rf_ll_enq_cnt_s_bin1_re                           (rf_ll_enq_cnt_s_bin1_re)
    ,.rf_ll_enq_cnt_s_bin1_rclk                         (rf_ll_enq_cnt_s_bin1_rclk)
    ,.rf_ll_enq_cnt_s_bin1_rclk_rst_n                   (rf_ll_enq_cnt_s_bin1_rclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin1_raddr                        (rf_ll_enq_cnt_s_bin1_raddr)
    ,.rf_ll_enq_cnt_s_bin1_waddr                        (rf_ll_enq_cnt_s_bin1_waddr)
    ,.rf_ll_enq_cnt_s_bin1_we                           (rf_ll_enq_cnt_s_bin1_we)
    ,.rf_ll_enq_cnt_s_bin1_wclk                         (rf_ll_enq_cnt_s_bin1_wclk)
    ,.rf_ll_enq_cnt_s_bin1_wclk_rst_n                   (rf_ll_enq_cnt_s_bin1_wclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin1_wdata                        (rf_ll_enq_cnt_s_bin1_wdata)
    ,.rf_ll_enq_cnt_s_bin1_rdata                        (rf_ll_enq_cnt_s_bin1_rdata)

    ,.rf_ll_enq_cnt_s_bin2_re                           (rf_ll_enq_cnt_s_bin2_re)
    ,.rf_ll_enq_cnt_s_bin2_rclk                         (rf_ll_enq_cnt_s_bin2_rclk)
    ,.rf_ll_enq_cnt_s_bin2_rclk_rst_n                   (rf_ll_enq_cnt_s_bin2_rclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin2_raddr                        (rf_ll_enq_cnt_s_bin2_raddr)
    ,.rf_ll_enq_cnt_s_bin2_waddr                        (rf_ll_enq_cnt_s_bin2_waddr)
    ,.rf_ll_enq_cnt_s_bin2_we                           (rf_ll_enq_cnt_s_bin2_we)
    ,.rf_ll_enq_cnt_s_bin2_wclk                         (rf_ll_enq_cnt_s_bin2_wclk)
    ,.rf_ll_enq_cnt_s_bin2_wclk_rst_n                   (rf_ll_enq_cnt_s_bin2_wclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin2_wdata                        (rf_ll_enq_cnt_s_bin2_wdata)
    ,.rf_ll_enq_cnt_s_bin2_rdata                        (rf_ll_enq_cnt_s_bin2_rdata)

    ,.rf_ll_enq_cnt_s_bin3_re                           (rf_ll_enq_cnt_s_bin3_re)
    ,.rf_ll_enq_cnt_s_bin3_rclk                         (rf_ll_enq_cnt_s_bin3_rclk)
    ,.rf_ll_enq_cnt_s_bin3_rclk_rst_n                   (rf_ll_enq_cnt_s_bin3_rclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin3_raddr                        (rf_ll_enq_cnt_s_bin3_raddr)
    ,.rf_ll_enq_cnt_s_bin3_waddr                        (rf_ll_enq_cnt_s_bin3_waddr)
    ,.rf_ll_enq_cnt_s_bin3_we                           (rf_ll_enq_cnt_s_bin3_we)
    ,.rf_ll_enq_cnt_s_bin3_wclk                         (rf_ll_enq_cnt_s_bin3_wclk)
    ,.rf_ll_enq_cnt_s_bin3_wclk_rst_n                   (rf_ll_enq_cnt_s_bin3_wclk_rst_n)
    ,.rf_ll_enq_cnt_s_bin3_wdata                        (rf_ll_enq_cnt_s_bin3_wdata)
    ,.rf_ll_enq_cnt_s_bin3_rdata                        (rf_ll_enq_cnt_s_bin3_rdata)

    ,.rf_ll_rdylst_hp_bin0_re                           (rf_ll_rdylst_hp_bin0_re)
    ,.rf_ll_rdylst_hp_bin0_rclk                         (rf_ll_rdylst_hp_bin0_rclk)
    ,.rf_ll_rdylst_hp_bin0_rclk_rst_n                   (rf_ll_rdylst_hp_bin0_rclk_rst_n)
    ,.rf_ll_rdylst_hp_bin0_raddr                        (rf_ll_rdylst_hp_bin0_raddr)
    ,.rf_ll_rdylst_hp_bin0_waddr                        (rf_ll_rdylst_hp_bin0_waddr)
    ,.rf_ll_rdylst_hp_bin0_we                           (rf_ll_rdylst_hp_bin0_we)
    ,.rf_ll_rdylst_hp_bin0_wclk                         (rf_ll_rdylst_hp_bin0_wclk)
    ,.rf_ll_rdylst_hp_bin0_wclk_rst_n                   (rf_ll_rdylst_hp_bin0_wclk_rst_n)
    ,.rf_ll_rdylst_hp_bin0_wdata                        (rf_ll_rdylst_hp_bin0_wdata)
    ,.rf_ll_rdylst_hp_bin0_rdata                        (rf_ll_rdylst_hp_bin0_rdata)

    ,.rf_ll_rdylst_hp_bin1_re                           (rf_ll_rdylst_hp_bin1_re)
    ,.rf_ll_rdylst_hp_bin1_rclk                         (rf_ll_rdylst_hp_bin1_rclk)
    ,.rf_ll_rdylst_hp_bin1_rclk_rst_n                   (rf_ll_rdylst_hp_bin1_rclk_rst_n)
    ,.rf_ll_rdylst_hp_bin1_raddr                        (rf_ll_rdylst_hp_bin1_raddr)
    ,.rf_ll_rdylst_hp_bin1_waddr                        (rf_ll_rdylst_hp_bin1_waddr)
    ,.rf_ll_rdylst_hp_bin1_we                           (rf_ll_rdylst_hp_bin1_we)
    ,.rf_ll_rdylst_hp_bin1_wclk                         (rf_ll_rdylst_hp_bin1_wclk)
    ,.rf_ll_rdylst_hp_bin1_wclk_rst_n                   (rf_ll_rdylst_hp_bin1_wclk_rst_n)
    ,.rf_ll_rdylst_hp_bin1_wdata                        (rf_ll_rdylst_hp_bin1_wdata)
    ,.rf_ll_rdylst_hp_bin1_rdata                        (rf_ll_rdylst_hp_bin1_rdata)

    ,.rf_ll_rdylst_hp_bin2_re                           (rf_ll_rdylst_hp_bin2_re)
    ,.rf_ll_rdylst_hp_bin2_rclk                         (rf_ll_rdylst_hp_bin2_rclk)
    ,.rf_ll_rdylst_hp_bin2_rclk_rst_n                   (rf_ll_rdylst_hp_bin2_rclk_rst_n)
    ,.rf_ll_rdylst_hp_bin2_raddr                        (rf_ll_rdylst_hp_bin2_raddr)
    ,.rf_ll_rdylst_hp_bin2_waddr                        (rf_ll_rdylst_hp_bin2_waddr)
    ,.rf_ll_rdylst_hp_bin2_we                           (rf_ll_rdylst_hp_bin2_we)
    ,.rf_ll_rdylst_hp_bin2_wclk                         (rf_ll_rdylst_hp_bin2_wclk)
    ,.rf_ll_rdylst_hp_bin2_wclk_rst_n                   (rf_ll_rdylst_hp_bin2_wclk_rst_n)
    ,.rf_ll_rdylst_hp_bin2_wdata                        (rf_ll_rdylst_hp_bin2_wdata)
    ,.rf_ll_rdylst_hp_bin2_rdata                        (rf_ll_rdylst_hp_bin2_rdata)

    ,.rf_ll_rdylst_hp_bin3_re                           (rf_ll_rdylst_hp_bin3_re)
    ,.rf_ll_rdylst_hp_bin3_rclk                         (rf_ll_rdylst_hp_bin3_rclk)
    ,.rf_ll_rdylst_hp_bin3_rclk_rst_n                   (rf_ll_rdylst_hp_bin3_rclk_rst_n)
    ,.rf_ll_rdylst_hp_bin3_raddr                        (rf_ll_rdylst_hp_bin3_raddr)
    ,.rf_ll_rdylst_hp_bin3_waddr                        (rf_ll_rdylst_hp_bin3_waddr)
    ,.rf_ll_rdylst_hp_bin3_we                           (rf_ll_rdylst_hp_bin3_we)
    ,.rf_ll_rdylst_hp_bin3_wclk                         (rf_ll_rdylst_hp_bin3_wclk)
    ,.rf_ll_rdylst_hp_bin3_wclk_rst_n                   (rf_ll_rdylst_hp_bin3_wclk_rst_n)
    ,.rf_ll_rdylst_hp_bin3_wdata                        (rf_ll_rdylst_hp_bin3_wdata)
    ,.rf_ll_rdylst_hp_bin3_rdata                        (rf_ll_rdylst_hp_bin3_rdata)

    ,.rf_ll_rdylst_hpnxt_bin0_re                        (rf_ll_rdylst_hpnxt_bin0_re)
    ,.rf_ll_rdylst_hpnxt_bin0_rclk                      (rf_ll_rdylst_hpnxt_bin0_rclk)
    ,.rf_ll_rdylst_hpnxt_bin0_rclk_rst_n                (rf_ll_rdylst_hpnxt_bin0_rclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin0_raddr                     (rf_ll_rdylst_hpnxt_bin0_raddr)
    ,.rf_ll_rdylst_hpnxt_bin0_waddr                     (rf_ll_rdylst_hpnxt_bin0_waddr)
    ,.rf_ll_rdylst_hpnxt_bin0_we                        (rf_ll_rdylst_hpnxt_bin0_we)
    ,.rf_ll_rdylst_hpnxt_bin0_wclk                      (rf_ll_rdylst_hpnxt_bin0_wclk)
    ,.rf_ll_rdylst_hpnxt_bin0_wclk_rst_n                (rf_ll_rdylst_hpnxt_bin0_wclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin0_wdata                     (rf_ll_rdylst_hpnxt_bin0_wdata)
    ,.rf_ll_rdylst_hpnxt_bin0_rdata                     (rf_ll_rdylst_hpnxt_bin0_rdata)

    ,.rf_ll_rdylst_hpnxt_bin1_re                        (rf_ll_rdylst_hpnxt_bin1_re)
    ,.rf_ll_rdylst_hpnxt_bin1_rclk                      (rf_ll_rdylst_hpnxt_bin1_rclk)
    ,.rf_ll_rdylst_hpnxt_bin1_rclk_rst_n                (rf_ll_rdylst_hpnxt_bin1_rclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin1_raddr                     (rf_ll_rdylst_hpnxt_bin1_raddr)
    ,.rf_ll_rdylst_hpnxt_bin1_waddr                     (rf_ll_rdylst_hpnxt_bin1_waddr)
    ,.rf_ll_rdylst_hpnxt_bin1_we                        (rf_ll_rdylst_hpnxt_bin1_we)
    ,.rf_ll_rdylst_hpnxt_bin1_wclk                      (rf_ll_rdylst_hpnxt_bin1_wclk)
    ,.rf_ll_rdylst_hpnxt_bin1_wclk_rst_n                (rf_ll_rdylst_hpnxt_bin1_wclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin1_wdata                     (rf_ll_rdylst_hpnxt_bin1_wdata)
    ,.rf_ll_rdylst_hpnxt_bin1_rdata                     (rf_ll_rdylst_hpnxt_bin1_rdata)

    ,.rf_ll_rdylst_hpnxt_bin2_re                        (rf_ll_rdylst_hpnxt_bin2_re)
    ,.rf_ll_rdylst_hpnxt_bin2_rclk                      (rf_ll_rdylst_hpnxt_bin2_rclk)
    ,.rf_ll_rdylst_hpnxt_bin2_rclk_rst_n                (rf_ll_rdylst_hpnxt_bin2_rclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin2_raddr                     (rf_ll_rdylst_hpnxt_bin2_raddr)
    ,.rf_ll_rdylst_hpnxt_bin2_waddr                     (rf_ll_rdylst_hpnxt_bin2_waddr)
    ,.rf_ll_rdylst_hpnxt_bin2_we                        (rf_ll_rdylst_hpnxt_bin2_we)
    ,.rf_ll_rdylst_hpnxt_bin2_wclk                      (rf_ll_rdylst_hpnxt_bin2_wclk)
    ,.rf_ll_rdylst_hpnxt_bin2_wclk_rst_n                (rf_ll_rdylst_hpnxt_bin2_wclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin2_wdata                     (rf_ll_rdylst_hpnxt_bin2_wdata)
    ,.rf_ll_rdylst_hpnxt_bin2_rdata                     (rf_ll_rdylst_hpnxt_bin2_rdata)

    ,.rf_ll_rdylst_hpnxt_bin3_re                        (rf_ll_rdylst_hpnxt_bin3_re)
    ,.rf_ll_rdylst_hpnxt_bin3_rclk                      (rf_ll_rdylst_hpnxt_bin3_rclk)
    ,.rf_ll_rdylst_hpnxt_bin3_rclk_rst_n                (rf_ll_rdylst_hpnxt_bin3_rclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin3_raddr                     (rf_ll_rdylst_hpnxt_bin3_raddr)
    ,.rf_ll_rdylst_hpnxt_bin3_waddr                     (rf_ll_rdylst_hpnxt_bin3_waddr)
    ,.rf_ll_rdylst_hpnxt_bin3_we                        (rf_ll_rdylst_hpnxt_bin3_we)
    ,.rf_ll_rdylst_hpnxt_bin3_wclk                      (rf_ll_rdylst_hpnxt_bin3_wclk)
    ,.rf_ll_rdylst_hpnxt_bin3_wclk_rst_n                (rf_ll_rdylst_hpnxt_bin3_wclk_rst_n)
    ,.rf_ll_rdylst_hpnxt_bin3_wdata                     (rf_ll_rdylst_hpnxt_bin3_wdata)
    ,.rf_ll_rdylst_hpnxt_bin3_rdata                     (rf_ll_rdylst_hpnxt_bin3_rdata)

    ,.rf_ll_rdylst_tp_bin0_re                           (rf_ll_rdylst_tp_bin0_re)
    ,.rf_ll_rdylst_tp_bin0_rclk                         (rf_ll_rdylst_tp_bin0_rclk)
    ,.rf_ll_rdylst_tp_bin0_rclk_rst_n                   (rf_ll_rdylst_tp_bin0_rclk_rst_n)
    ,.rf_ll_rdylst_tp_bin0_raddr                        (rf_ll_rdylst_tp_bin0_raddr)
    ,.rf_ll_rdylst_tp_bin0_waddr                        (rf_ll_rdylst_tp_bin0_waddr)
    ,.rf_ll_rdylst_tp_bin0_we                           (rf_ll_rdylst_tp_bin0_we)
    ,.rf_ll_rdylst_tp_bin0_wclk                         (rf_ll_rdylst_tp_bin0_wclk)
    ,.rf_ll_rdylst_tp_bin0_wclk_rst_n                   (rf_ll_rdylst_tp_bin0_wclk_rst_n)
    ,.rf_ll_rdylst_tp_bin0_wdata                        (rf_ll_rdylst_tp_bin0_wdata)
    ,.rf_ll_rdylst_tp_bin0_rdata                        (rf_ll_rdylst_tp_bin0_rdata)

    ,.rf_ll_rdylst_tp_bin1_re                           (rf_ll_rdylst_tp_bin1_re)
    ,.rf_ll_rdylst_tp_bin1_rclk                         (rf_ll_rdylst_tp_bin1_rclk)
    ,.rf_ll_rdylst_tp_bin1_rclk_rst_n                   (rf_ll_rdylst_tp_bin1_rclk_rst_n)
    ,.rf_ll_rdylst_tp_bin1_raddr                        (rf_ll_rdylst_tp_bin1_raddr)
    ,.rf_ll_rdylst_tp_bin1_waddr                        (rf_ll_rdylst_tp_bin1_waddr)
    ,.rf_ll_rdylst_tp_bin1_we                           (rf_ll_rdylst_tp_bin1_we)
    ,.rf_ll_rdylst_tp_bin1_wclk                         (rf_ll_rdylst_tp_bin1_wclk)
    ,.rf_ll_rdylst_tp_bin1_wclk_rst_n                   (rf_ll_rdylst_tp_bin1_wclk_rst_n)
    ,.rf_ll_rdylst_tp_bin1_wdata                        (rf_ll_rdylst_tp_bin1_wdata)
    ,.rf_ll_rdylst_tp_bin1_rdata                        (rf_ll_rdylst_tp_bin1_rdata)

    ,.rf_ll_rdylst_tp_bin2_re                           (rf_ll_rdylst_tp_bin2_re)
    ,.rf_ll_rdylst_tp_bin2_rclk                         (rf_ll_rdylst_tp_bin2_rclk)
    ,.rf_ll_rdylst_tp_bin2_rclk_rst_n                   (rf_ll_rdylst_tp_bin2_rclk_rst_n)
    ,.rf_ll_rdylst_tp_bin2_raddr                        (rf_ll_rdylst_tp_bin2_raddr)
    ,.rf_ll_rdylst_tp_bin2_waddr                        (rf_ll_rdylst_tp_bin2_waddr)
    ,.rf_ll_rdylst_tp_bin2_we                           (rf_ll_rdylst_tp_bin2_we)
    ,.rf_ll_rdylst_tp_bin2_wclk                         (rf_ll_rdylst_tp_bin2_wclk)
    ,.rf_ll_rdylst_tp_bin2_wclk_rst_n                   (rf_ll_rdylst_tp_bin2_wclk_rst_n)
    ,.rf_ll_rdylst_tp_bin2_wdata                        (rf_ll_rdylst_tp_bin2_wdata)
    ,.rf_ll_rdylst_tp_bin2_rdata                        (rf_ll_rdylst_tp_bin2_rdata)

    ,.rf_ll_rdylst_tp_bin3_re                           (rf_ll_rdylst_tp_bin3_re)
    ,.rf_ll_rdylst_tp_bin3_rclk                         (rf_ll_rdylst_tp_bin3_rclk)
    ,.rf_ll_rdylst_tp_bin3_rclk_rst_n                   (rf_ll_rdylst_tp_bin3_rclk_rst_n)
    ,.rf_ll_rdylst_tp_bin3_raddr                        (rf_ll_rdylst_tp_bin3_raddr)
    ,.rf_ll_rdylst_tp_bin3_waddr                        (rf_ll_rdylst_tp_bin3_waddr)
    ,.rf_ll_rdylst_tp_bin3_we                           (rf_ll_rdylst_tp_bin3_we)
    ,.rf_ll_rdylst_tp_bin3_wclk                         (rf_ll_rdylst_tp_bin3_wclk)
    ,.rf_ll_rdylst_tp_bin3_wclk_rst_n                   (rf_ll_rdylst_tp_bin3_wclk_rst_n)
    ,.rf_ll_rdylst_tp_bin3_wdata                        (rf_ll_rdylst_tp_bin3_wdata)
    ,.rf_ll_rdylst_tp_bin3_rdata                        (rf_ll_rdylst_tp_bin3_rdata)

    ,.rf_ll_rlst_cnt_re                                 (rf_ll_rlst_cnt_re)
    ,.rf_ll_rlst_cnt_rclk                               (rf_ll_rlst_cnt_rclk)
    ,.rf_ll_rlst_cnt_rclk_rst_n                         (rf_ll_rlst_cnt_rclk_rst_n)
    ,.rf_ll_rlst_cnt_raddr                              (rf_ll_rlst_cnt_raddr)
    ,.rf_ll_rlst_cnt_waddr                              (rf_ll_rlst_cnt_waddr)
    ,.rf_ll_rlst_cnt_we                                 (rf_ll_rlst_cnt_we)
    ,.rf_ll_rlst_cnt_wclk                               (rf_ll_rlst_cnt_wclk)
    ,.rf_ll_rlst_cnt_wclk_rst_n                         (rf_ll_rlst_cnt_wclk_rst_n)
    ,.rf_ll_rlst_cnt_wdata                              (rf_ll_rlst_cnt_wdata)
    ,.rf_ll_rlst_cnt_rdata                              (rf_ll_rlst_cnt_rdata)

    ,.rf_ll_sch_cnt_dup0_re                             (rf_ll_sch_cnt_dup0_re)
    ,.rf_ll_sch_cnt_dup0_rclk                           (rf_ll_sch_cnt_dup0_rclk)
    ,.rf_ll_sch_cnt_dup0_rclk_rst_n                     (rf_ll_sch_cnt_dup0_rclk_rst_n)
    ,.rf_ll_sch_cnt_dup0_raddr                          (rf_ll_sch_cnt_dup0_raddr)
    ,.rf_ll_sch_cnt_dup0_waddr                          (rf_ll_sch_cnt_dup0_waddr)
    ,.rf_ll_sch_cnt_dup0_we                             (rf_ll_sch_cnt_dup0_we)
    ,.rf_ll_sch_cnt_dup0_wclk                           (rf_ll_sch_cnt_dup0_wclk)
    ,.rf_ll_sch_cnt_dup0_wclk_rst_n                     (rf_ll_sch_cnt_dup0_wclk_rst_n)
    ,.rf_ll_sch_cnt_dup0_wdata                          (rf_ll_sch_cnt_dup0_wdata)
    ,.rf_ll_sch_cnt_dup0_rdata                          (rf_ll_sch_cnt_dup0_rdata)

    ,.rf_ll_sch_cnt_dup1_re                             (rf_ll_sch_cnt_dup1_re)
    ,.rf_ll_sch_cnt_dup1_rclk                           (rf_ll_sch_cnt_dup1_rclk)
    ,.rf_ll_sch_cnt_dup1_rclk_rst_n                     (rf_ll_sch_cnt_dup1_rclk_rst_n)
    ,.rf_ll_sch_cnt_dup1_raddr                          (rf_ll_sch_cnt_dup1_raddr)
    ,.rf_ll_sch_cnt_dup1_waddr                          (rf_ll_sch_cnt_dup1_waddr)
    ,.rf_ll_sch_cnt_dup1_we                             (rf_ll_sch_cnt_dup1_we)
    ,.rf_ll_sch_cnt_dup1_wclk                           (rf_ll_sch_cnt_dup1_wclk)
    ,.rf_ll_sch_cnt_dup1_wclk_rst_n                     (rf_ll_sch_cnt_dup1_wclk_rst_n)
    ,.rf_ll_sch_cnt_dup1_wdata                          (rf_ll_sch_cnt_dup1_wdata)
    ,.rf_ll_sch_cnt_dup1_rdata                          (rf_ll_sch_cnt_dup1_rdata)

    ,.rf_ll_sch_cnt_dup2_re                             (rf_ll_sch_cnt_dup2_re)
    ,.rf_ll_sch_cnt_dup2_rclk                           (rf_ll_sch_cnt_dup2_rclk)
    ,.rf_ll_sch_cnt_dup2_rclk_rst_n                     (rf_ll_sch_cnt_dup2_rclk_rst_n)
    ,.rf_ll_sch_cnt_dup2_raddr                          (rf_ll_sch_cnt_dup2_raddr)
    ,.rf_ll_sch_cnt_dup2_waddr                          (rf_ll_sch_cnt_dup2_waddr)
    ,.rf_ll_sch_cnt_dup2_we                             (rf_ll_sch_cnt_dup2_we)
    ,.rf_ll_sch_cnt_dup2_wclk                           (rf_ll_sch_cnt_dup2_wclk)
    ,.rf_ll_sch_cnt_dup2_wclk_rst_n                     (rf_ll_sch_cnt_dup2_wclk_rst_n)
    ,.rf_ll_sch_cnt_dup2_wdata                          (rf_ll_sch_cnt_dup2_wdata)
    ,.rf_ll_sch_cnt_dup2_rdata                          (rf_ll_sch_cnt_dup2_rdata)

    ,.rf_ll_sch_cnt_dup3_re                             (rf_ll_sch_cnt_dup3_re)
    ,.rf_ll_sch_cnt_dup3_rclk                           (rf_ll_sch_cnt_dup3_rclk)
    ,.rf_ll_sch_cnt_dup3_rclk_rst_n                     (rf_ll_sch_cnt_dup3_rclk_rst_n)
    ,.rf_ll_sch_cnt_dup3_raddr                          (rf_ll_sch_cnt_dup3_raddr)
    ,.rf_ll_sch_cnt_dup3_waddr                          (rf_ll_sch_cnt_dup3_waddr)
    ,.rf_ll_sch_cnt_dup3_we                             (rf_ll_sch_cnt_dup3_we)
    ,.rf_ll_sch_cnt_dup3_wclk                           (rf_ll_sch_cnt_dup3_wclk)
    ,.rf_ll_sch_cnt_dup3_wclk_rst_n                     (rf_ll_sch_cnt_dup3_wclk_rst_n)
    ,.rf_ll_sch_cnt_dup3_wdata                          (rf_ll_sch_cnt_dup3_wdata)
    ,.rf_ll_sch_cnt_dup3_rdata                          (rf_ll_sch_cnt_dup3_rdata)

    ,.rf_ll_schlst_hp_bin0_re                           (rf_ll_schlst_hp_bin0_re)
    ,.rf_ll_schlst_hp_bin0_rclk                         (rf_ll_schlst_hp_bin0_rclk)
    ,.rf_ll_schlst_hp_bin0_rclk_rst_n                   (rf_ll_schlst_hp_bin0_rclk_rst_n)
    ,.rf_ll_schlst_hp_bin0_raddr                        (rf_ll_schlst_hp_bin0_raddr)
    ,.rf_ll_schlst_hp_bin0_waddr                        (rf_ll_schlst_hp_bin0_waddr)
    ,.rf_ll_schlst_hp_bin0_we                           (rf_ll_schlst_hp_bin0_we)
    ,.rf_ll_schlst_hp_bin0_wclk                         (rf_ll_schlst_hp_bin0_wclk)
    ,.rf_ll_schlst_hp_bin0_wclk_rst_n                   (rf_ll_schlst_hp_bin0_wclk_rst_n)
    ,.rf_ll_schlst_hp_bin0_wdata                        (rf_ll_schlst_hp_bin0_wdata)
    ,.rf_ll_schlst_hp_bin0_rdata                        (rf_ll_schlst_hp_bin0_rdata)

    ,.rf_ll_schlst_hp_bin1_re                           (rf_ll_schlst_hp_bin1_re)
    ,.rf_ll_schlst_hp_bin1_rclk                         (rf_ll_schlst_hp_bin1_rclk)
    ,.rf_ll_schlst_hp_bin1_rclk_rst_n                   (rf_ll_schlst_hp_bin1_rclk_rst_n)
    ,.rf_ll_schlst_hp_bin1_raddr                        (rf_ll_schlst_hp_bin1_raddr)
    ,.rf_ll_schlst_hp_bin1_waddr                        (rf_ll_schlst_hp_bin1_waddr)
    ,.rf_ll_schlst_hp_bin1_we                           (rf_ll_schlst_hp_bin1_we)
    ,.rf_ll_schlst_hp_bin1_wclk                         (rf_ll_schlst_hp_bin1_wclk)
    ,.rf_ll_schlst_hp_bin1_wclk_rst_n                   (rf_ll_schlst_hp_bin1_wclk_rst_n)
    ,.rf_ll_schlst_hp_bin1_wdata                        (rf_ll_schlst_hp_bin1_wdata)
    ,.rf_ll_schlst_hp_bin1_rdata                        (rf_ll_schlst_hp_bin1_rdata)

    ,.rf_ll_schlst_hp_bin2_re                           (rf_ll_schlst_hp_bin2_re)
    ,.rf_ll_schlst_hp_bin2_rclk                         (rf_ll_schlst_hp_bin2_rclk)
    ,.rf_ll_schlst_hp_bin2_rclk_rst_n                   (rf_ll_schlst_hp_bin2_rclk_rst_n)
    ,.rf_ll_schlst_hp_bin2_raddr                        (rf_ll_schlst_hp_bin2_raddr)
    ,.rf_ll_schlst_hp_bin2_waddr                        (rf_ll_schlst_hp_bin2_waddr)
    ,.rf_ll_schlst_hp_bin2_we                           (rf_ll_schlst_hp_bin2_we)
    ,.rf_ll_schlst_hp_bin2_wclk                         (rf_ll_schlst_hp_bin2_wclk)
    ,.rf_ll_schlst_hp_bin2_wclk_rst_n                   (rf_ll_schlst_hp_bin2_wclk_rst_n)
    ,.rf_ll_schlst_hp_bin2_wdata                        (rf_ll_schlst_hp_bin2_wdata)
    ,.rf_ll_schlst_hp_bin2_rdata                        (rf_ll_schlst_hp_bin2_rdata)

    ,.rf_ll_schlst_hp_bin3_re                           (rf_ll_schlst_hp_bin3_re)
    ,.rf_ll_schlst_hp_bin3_rclk                         (rf_ll_schlst_hp_bin3_rclk)
    ,.rf_ll_schlst_hp_bin3_rclk_rst_n                   (rf_ll_schlst_hp_bin3_rclk_rst_n)
    ,.rf_ll_schlst_hp_bin3_raddr                        (rf_ll_schlst_hp_bin3_raddr)
    ,.rf_ll_schlst_hp_bin3_waddr                        (rf_ll_schlst_hp_bin3_waddr)
    ,.rf_ll_schlst_hp_bin3_we                           (rf_ll_schlst_hp_bin3_we)
    ,.rf_ll_schlst_hp_bin3_wclk                         (rf_ll_schlst_hp_bin3_wclk)
    ,.rf_ll_schlst_hp_bin3_wclk_rst_n                   (rf_ll_schlst_hp_bin3_wclk_rst_n)
    ,.rf_ll_schlst_hp_bin3_wdata                        (rf_ll_schlst_hp_bin3_wdata)
    ,.rf_ll_schlst_hp_bin3_rdata                        (rf_ll_schlst_hp_bin3_rdata)

    ,.rf_ll_schlst_hpnxt_bin0_re                        (rf_ll_schlst_hpnxt_bin0_re)
    ,.rf_ll_schlst_hpnxt_bin0_rclk                      (rf_ll_schlst_hpnxt_bin0_rclk)
    ,.rf_ll_schlst_hpnxt_bin0_rclk_rst_n                (rf_ll_schlst_hpnxt_bin0_rclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin0_raddr                     (rf_ll_schlst_hpnxt_bin0_raddr)
    ,.rf_ll_schlst_hpnxt_bin0_waddr                     (rf_ll_schlst_hpnxt_bin0_waddr)
    ,.rf_ll_schlst_hpnxt_bin0_we                        (rf_ll_schlst_hpnxt_bin0_we)
    ,.rf_ll_schlst_hpnxt_bin0_wclk                      (rf_ll_schlst_hpnxt_bin0_wclk)
    ,.rf_ll_schlst_hpnxt_bin0_wclk_rst_n                (rf_ll_schlst_hpnxt_bin0_wclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin0_wdata                     (rf_ll_schlst_hpnxt_bin0_wdata)
    ,.rf_ll_schlst_hpnxt_bin0_rdata                     (rf_ll_schlst_hpnxt_bin0_rdata)

    ,.rf_ll_schlst_hpnxt_bin1_re                        (rf_ll_schlst_hpnxt_bin1_re)
    ,.rf_ll_schlst_hpnxt_bin1_rclk                      (rf_ll_schlst_hpnxt_bin1_rclk)
    ,.rf_ll_schlst_hpnxt_bin1_rclk_rst_n                (rf_ll_schlst_hpnxt_bin1_rclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin1_raddr                     (rf_ll_schlst_hpnxt_bin1_raddr)
    ,.rf_ll_schlst_hpnxt_bin1_waddr                     (rf_ll_schlst_hpnxt_bin1_waddr)
    ,.rf_ll_schlst_hpnxt_bin1_we                        (rf_ll_schlst_hpnxt_bin1_we)
    ,.rf_ll_schlst_hpnxt_bin1_wclk                      (rf_ll_schlst_hpnxt_bin1_wclk)
    ,.rf_ll_schlst_hpnxt_bin1_wclk_rst_n                (rf_ll_schlst_hpnxt_bin1_wclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin1_wdata                     (rf_ll_schlst_hpnxt_bin1_wdata)
    ,.rf_ll_schlst_hpnxt_bin1_rdata                     (rf_ll_schlst_hpnxt_bin1_rdata)

    ,.rf_ll_schlst_hpnxt_bin2_re                        (rf_ll_schlst_hpnxt_bin2_re)
    ,.rf_ll_schlst_hpnxt_bin2_rclk                      (rf_ll_schlst_hpnxt_bin2_rclk)
    ,.rf_ll_schlst_hpnxt_bin2_rclk_rst_n                (rf_ll_schlst_hpnxt_bin2_rclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin2_raddr                     (rf_ll_schlst_hpnxt_bin2_raddr)
    ,.rf_ll_schlst_hpnxt_bin2_waddr                     (rf_ll_schlst_hpnxt_bin2_waddr)
    ,.rf_ll_schlst_hpnxt_bin2_we                        (rf_ll_schlst_hpnxt_bin2_we)
    ,.rf_ll_schlst_hpnxt_bin2_wclk                      (rf_ll_schlst_hpnxt_bin2_wclk)
    ,.rf_ll_schlst_hpnxt_bin2_wclk_rst_n                (rf_ll_schlst_hpnxt_bin2_wclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin2_wdata                     (rf_ll_schlst_hpnxt_bin2_wdata)
    ,.rf_ll_schlst_hpnxt_bin2_rdata                     (rf_ll_schlst_hpnxt_bin2_rdata)

    ,.rf_ll_schlst_hpnxt_bin3_re                        (rf_ll_schlst_hpnxt_bin3_re)
    ,.rf_ll_schlst_hpnxt_bin3_rclk                      (rf_ll_schlst_hpnxt_bin3_rclk)
    ,.rf_ll_schlst_hpnxt_bin3_rclk_rst_n                (rf_ll_schlst_hpnxt_bin3_rclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin3_raddr                     (rf_ll_schlst_hpnxt_bin3_raddr)
    ,.rf_ll_schlst_hpnxt_bin3_waddr                     (rf_ll_schlst_hpnxt_bin3_waddr)
    ,.rf_ll_schlst_hpnxt_bin3_we                        (rf_ll_schlst_hpnxt_bin3_we)
    ,.rf_ll_schlst_hpnxt_bin3_wclk                      (rf_ll_schlst_hpnxt_bin3_wclk)
    ,.rf_ll_schlst_hpnxt_bin3_wclk_rst_n                (rf_ll_schlst_hpnxt_bin3_wclk_rst_n)
    ,.rf_ll_schlst_hpnxt_bin3_wdata                     (rf_ll_schlst_hpnxt_bin3_wdata)
    ,.rf_ll_schlst_hpnxt_bin3_rdata                     (rf_ll_schlst_hpnxt_bin3_rdata)

    ,.rf_ll_schlst_tp_bin0_re                           (rf_ll_schlst_tp_bin0_re)
    ,.rf_ll_schlst_tp_bin0_rclk                         (rf_ll_schlst_tp_bin0_rclk)
    ,.rf_ll_schlst_tp_bin0_rclk_rst_n                   (rf_ll_schlst_tp_bin0_rclk_rst_n)
    ,.rf_ll_schlst_tp_bin0_raddr                        (rf_ll_schlst_tp_bin0_raddr)
    ,.rf_ll_schlst_tp_bin0_waddr                        (rf_ll_schlst_tp_bin0_waddr)
    ,.rf_ll_schlst_tp_bin0_we                           (rf_ll_schlst_tp_bin0_we)
    ,.rf_ll_schlst_tp_bin0_wclk                         (rf_ll_schlst_tp_bin0_wclk)
    ,.rf_ll_schlst_tp_bin0_wclk_rst_n                   (rf_ll_schlst_tp_bin0_wclk_rst_n)
    ,.rf_ll_schlst_tp_bin0_wdata                        (rf_ll_schlst_tp_bin0_wdata)
    ,.rf_ll_schlst_tp_bin0_rdata                        (rf_ll_schlst_tp_bin0_rdata)

    ,.rf_ll_schlst_tp_bin1_re                           (rf_ll_schlst_tp_bin1_re)
    ,.rf_ll_schlst_tp_bin1_rclk                         (rf_ll_schlst_tp_bin1_rclk)
    ,.rf_ll_schlst_tp_bin1_rclk_rst_n                   (rf_ll_schlst_tp_bin1_rclk_rst_n)
    ,.rf_ll_schlst_tp_bin1_raddr                        (rf_ll_schlst_tp_bin1_raddr)
    ,.rf_ll_schlst_tp_bin1_waddr                        (rf_ll_schlst_tp_bin1_waddr)
    ,.rf_ll_schlst_tp_bin1_we                           (rf_ll_schlst_tp_bin1_we)
    ,.rf_ll_schlst_tp_bin1_wclk                         (rf_ll_schlst_tp_bin1_wclk)
    ,.rf_ll_schlst_tp_bin1_wclk_rst_n                   (rf_ll_schlst_tp_bin1_wclk_rst_n)
    ,.rf_ll_schlst_tp_bin1_wdata                        (rf_ll_schlst_tp_bin1_wdata)
    ,.rf_ll_schlst_tp_bin1_rdata                        (rf_ll_schlst_tp_bin1_rdata)

    ,.rf_ll_schlst_tp_bin2_re                           (rf_ll_schlst_tp_bin2_re)
    ,.rf_ll_schlst_tp_bin2_rclk                         (rf_ll_schlst_tp_bin2_rclk)
    ,.rf_ll_schlst_tp_bin2_rclk_rst_n                   (rf_ll_schlst_tp_bin2_rclk_rst_n)
    ,.rf_ll_schlst_tp_bin2_raddr                        (rf_ll_schlst_tp_bin2_raddr)
    ,.rf_ll_schlst_tp_bin2_waddr                        (rf_ll_schlst_tp_bin2_waddr)
    ,.rf_ll_schlst_tp_bin2_we                           (rf_ll_schlst_tp_bin2_we)
    ,.rf_ll_schlst_tp_bin2_wclk                         (rf_ll_schlst_tp_bin2_wclk)
    ,.rf_ll_schlst_tp_bin2_wclk_rst_n                   (rf_ll_schlst_tp_bin2_wclk_rst_n)
    ,.rf_ll_schlst_tp_bin2_wdata                        (rf_ll_schlst_tp_bin2_wdata)
    ,.rf_ll_schlst_tp_bin2_rdata                        (rf_ll_schlst_tp_bin2_rdata)

    ,.rf_ll_schlst_tp_bin3_re                           (rf_ll_schlst_tp_bin3_re)
    ,.rf_ll_schlst_tp_bin3_rclk                         (rf_ll_schlst_tp_bin3_rclk)
    ,.rf_ll_schlst_tp_bin3_rclk_rst_n                   (rf_ll_schlst_tp_bin3_rclk_rst_n)
    ,.rf_ll_schlst_tp_bin3_raddr                        (rf_ll_schlst_tp_bin3_raddr)
    ,.rf_ll_schlst_tp_bin3_waddr                        (rf_ll_schlst_tp_bin3_waddr)
    ,.rf_ll_schlst_tp_bin3_we                           (rf_ll_schlst_tp_bin3_we)
    ,.rf_ll_schlst_tp_bin3_wclk                         (rf_ll_schlst_tp_bin3_wclk)
    ,.rf_ll_schlst_tp_bin3_wclk_rst_n                   (rf_ll_schlst_tp_bin3_wclk_rst_n)
    ,.rf_ll_schlst_tp_bin3_wdata                        (rf_ll_schlst_tp_bin3_wdata)
    ,.rf_ll_schlst_tp_bin3_rdata                        (rf_ll_schlst_tp_bin3_rdata)

    ,.rf_ll_schlst_tpprv_bin0_re                        (rf_ll_schlst_tpprv_bin0_re)
    ,.rf_ll_schlst_tpprv_bin0_rclk                      (rf_ll_schlst_tpprv_bin0_rclk)
    ,.rf_ll_schlst_tpprv_bin0_rclk_rst_n                (rf_ll_schlst_tpprv_bin0_rclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin0_raddr                     (rf_ll_schlst_tpprv_bin0_raddr)
    ,.rf_ll_schlst_tpprv_bin0_waddr                     (rf_ll_schlst_tpprv_bin0_waddr)
    ,.rf_ll_schlst_tpprv_bin0_we                        (rf_ll_schlst_tpprv_bin0_we)
    ,.rf_ll_schlst_tpprv_bin0_wclk                      (rf_ll_schlst_tpprv_bin0_wclk)
    ,.rf_ll_schlst_tpprv_bin0_wclk_rst_n                (rf_ll_schlst_tpprv_bin0_wclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin0_wdata                     (rf_ll_schlst_tpprv_bin0_wdata)
    ,.rf_ll_schlst_tpprv_bin0_rdata                     (rf_ll_schlst_tpprv_bin0_rdata)

    ,.rf_ll_schlst_tpprv_bin1_re                        (rf_ll_schlst_tpprv_bin1_re)
    ,.rf_ll_schlst_tpprv_bin1_rclk                      (rf_ll_schlst_tpprv_bin1_rclk)
    ,.rf_ll_schlst_tpprv_bin1_rclk_rst_n                (rf_ll_schlst_tpprv_bin1_rclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin1_raddr                     (rf_ll_schlst_tpprv_bin1_raddr)
    ,.rf_ll_schlst_tpprv_bin1_waddr                     (rf_ll_schlst_tpprv_bin1_waddr)
    ,.rf_ll_schlst_tpprv_bin1_we                        (rf_ll_schlst_tpprv_bin1_we)
    ,.rf_ll_schlst_tpprv_bin1_wclk                      (rf_ll_schlst_tpprv_bin1_wclk)
    ,.rf_ll_schlst_tpprv_bin1_wclk_rst_n                (rf_ll_schlst_tpprv_bin1_wclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin1_wdata                     (rf_ll_schlst_tpprv_bin1_wdata)
    ,.rf_ll_schlst_tpprv_bin1_rdata                     (rf_ll_schlst_tpprv_bin1_rdata)

    ,.rf_ll_schlst_tpprv_bin2_re                        (rf_ll_schlst_tpprv_bin2_re)
    ,.rf_ll_schlst_tpprv_bin2_rclk                      (rf_ll_schlst_tpprv_bin2_rclk)
    ,.rf_ll_schlst_tpprv_bin2_rclk_rst_n                (rf_ll_schlst_tpprv_bin2_rclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin2_raddr                     (rf_ll_schlst_tpprv_bin2_raddr)
    ,.rf_ll_schlst_tpprv_bin2_waddr                     (rf_ll_schlst_tpprv_bin2_waddr)
    ,.rf_ll_schlst_tpprv_bin2_we                        (rf_ll_schlst_tpprv_bin2_we)
    ,.rf_ll_schlst_tpprv_bin2_wclk                      (rf_ll_schlst_tpprv_bin2_wclk)
    ,.rf_ll_schlst_tpprv_bin2_wclk_rst_n                (rf_ll_schlst_tpprv_bin2_wclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin2_wdata                     (rf_ll_schlst_tpprv_bin2_wdata)
    ,.rf_ll_schlst_tpprv_bin2_rdata                     (rf_ll_schlst_tpprv_bin2_rdata)

    ,.rf_ll_schlst_tpprv_bin3_re                        (rf_ll_schlst_tpprv_bin3_re)
    ,.rf_ll_schlst_tpprv_bin3_rclk                      (rf_ll_schlst_tpprv_bin3_rclk)
    ,.rf_ll_schlst_tpprv_bin3_rclk_rst_n                (rf_ll_schlst_tpprv_bin3_rclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin3_raddr                     (rf_ll_schlst_tpprv_bin3_raddr)
    ,.rf_ll_schlst_tpprv_bin3_waddr                     (rf_ll_schlst_tpprv_bin3_waddr)
    ,.rf_ll_schlst_tpprv_bin3_we                        (rf_ll_schlst_tpprv_bin3_we)
    ,.rf_ll_schlst_tpprv_bin3_wclk                      (rf_ll_schlst_tpprv_bin3_wclk)
    ,.rf_ll_schlst_tpprv_bin3_wclk_rst_n                (rf_ll_schlst_tpprv_bin3_wclk_rst_n)
    ,.rf_ll_schlst_tpprv_bin3_wdata                     (rf_ll_schlst_tpprv_bin3_wdata)
    ,.rf_ll_schlst_tpprv_bin3_rdata                     (rf_ll_schlst_tpprv_bin3_rdata)

    ,.rf_ll_slst_cnt_re                                 (rf_ll_slst_cnt_re)
    ,.rf_ll_slst_cnt_rclk                               (rf_ll_slst_cnt_rclk)
    ,.rf_ll_slst_cnt_rclk_rst_n                         (rf_ll_slst_cnt_rclk_rst_n)
    ,.rf_ll_slst_cnt_raddr                              (rf_ll_slst_cnt_raddr)
    ,.rf_ll_slst_cnt_waddr                              (rf_ll_slst_cnt_waddr)
    ,.rf_ll_slst_cnt_we                                 (rf_ll_slst_cnt_we)
    ,.rf_ll_slst_cnt_wclk                               (rf_ll_slst_cnt_wclk)
    ,.rf_ll_slst_cnt_wclk_rst_n                         (rf_ll_slst_cnt_wclk_rst_n)
    ,.rf_ll_slst_cnt_wdata                              (rf_ll_slst_cnt_wdata)
    ,.rf_ll_slst_cnt_rdata                              (rf_ll_slst_cnt_rdata)

    ,.rf_qid_rdylst_clamp_re                            (rf_qid_rdylst_clamp_re)
    ,.rf_qid_rdylst_clamp_rclk                          (rf_qid_rdylst_clamp_rclk)
    ,.rf_qid_rdylst_clamp_rclk_rst_n                    (rf_qid_rdylst_clamp_rclk_rst_n)
    ,.rf_qid_rdylst_clamp_raddr                         (rf_qid_rdylst_clamp_raddr)
    ,.rf_qid_rdylst_clamp_waddr                         (rf_qid_rdylst_clamp_waddr)
    ,.rf_qid_rdylst_clamp_we                            (rf_qid_rdylst_clamp_we)
    ,.rf_qid_rdylst_clamp_wclk                          (rf_qid_rdylst_clamp_wclk)
    ,.rf_qid_rdylst_clamp_wclk_rst_n                    (rf_qid_rdylst_clamp_wclk_rst_n)
    ,.rf_qid_rdylst_clamp_wdata                         (rf_qid_rdylst_clamp_wdata)
    ,.rf_qid_rdylst_clamp_rdata                         (rf_qid_rdylst_clamp_rdata)

// END HQM_MEMPORT_INST hqm_lsp_atm_pipe
) ; 

always_ff @ ( posedge hqm_gated_clk or negedge hqm_gated_rst_n ) begin
  if ( ~ hqm_gated_rst_n ) begin
    core_chp_lsp_ldb_cq_off_f <= { HQM_NUM_LB_CQ { 1'b0 } } ;
  end
  else begin
    core_chp_lsp_ldb_cq_off_f <= chp_lsp_ldb_cq_off ;
  end
end

//-----------------------------------------------------------------------------------------------------
// Spares

hqm_AW_spare_ports i_spare_ports_qed (

     .clk                       (hqm_inp_gated_clk)
    ,.rst_n                     (hqm_inp_gated_rst_b_lsp)
    ,.spare_in                  (spare_qed_lsp)
    ,.spare_out                 (spare_lsp_qed)
);

hqm_AW_spare_ports i_spare_ports_sys (

     .clk                       (hqm_inp_gated_clk)
    ,.rst_n                     (hqm_inp_gated_rst_b_lsp)
    ,.spare_in                  (spare_sys_lsp)
    ,.spare_out                 (spare_lsp_sys)
);

//-----------------------------------------------------------------------------------------------------
// SUBSECTION: Debug
//-----------------------------------------------------------------------------------------------------




//-----------------------------------------------------------------------------------------------------
// SUBSECTION: To be deleted
//-----------------------------------------------------------------------------------------------------
endmodule // hqm_list_sel_pipe_core
