module ctech_lib_latch_async_rst (clk, d, rb, o);
   input clk, d, rb;
   output o;
   logic o;
   d04lyn03ld0b0 ctech_lib_dcszo (.clk(clk),.d(d),.rb(rb),.o(o));
endmodule
