//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr1 : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr1
(
  // Synchronous Clock/Reset
  iosf_idf_side_clk,
  iosf_idf_side_rst_b,

  // Asynchronous Clock/Reset(s)
  iosf_fust_side_clk,
  iosf_swf_side_clk,

  // Power Well Isolation Input Signals
  crp_sbr1_xu_en,
  crp_sbr1_scu1_en,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  p3_fab_init_idle_exit,
  p3_fab_init_idle_exit_ack,
  p4_fab_init_idle_exit,
  p4_fab_init_idle_exit_ack,
  p5_fab_init_idle_exit,
  p5_fab_init_idle_exit_ack,
  p6_fab_init_idle_exit,
  p6_fab_init_idle_exit_ack,
  p7_fab_init_idle_exit,
  p7_fab_init_idle_exit_ack,
  p8_fab_init_idle_exit,
  p8_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_iosf_idf_side_clk,
  visa_vp_iosf_idf_side_clk,
  visa_p0_tier1_iosf_idf_side_clk,
  visa_p0_tier2_iosf_idf_side_clk,
  visa_p1_tier1_iosf_fust_side_clk,
  visa_p1_tier2_iosf_fust_side_clk,
  visa_p1_ififo_tier1_iosf_idf_side_clk,
  visa_p1_ififo_tier2_iosf_idf_side_clk,
  visa_p1_efifo_tier1_iosf_idf_side_clk,
  visa_p1_efifo_tier2_iosf_idf_side_clk,
  visa_p2_tier1_iosf_swf_side_clk,
  visa_p2_tier2_iosf_swf_side_clk,
  visa_p2_ififo_tier1_iosf_idf_side_clk,
  visa_p2_ififo_tier2_iosf_idf_side_clk,
  visa_p2_efifo_tier1_iosf_idf_side_clk,
  visa_p2_efifo_tier2_iosf_idf_side_clk,
  visa_p3_tier1_iosf_idf_side_clk,
  visa_p3_tier2_iosf_idf_side_clk,
  visa_p4_tier1_iosf_idf_side_clk,
  visa_p4_tier2_iosf_idf_side_clk,
  visa_p5_tier1_iosf_idf_side_clk,
  visa_p5_tier2_iosf_idf_side_clk,
  visa_p6_tier1_iosf_idf_side_clk,
  visa_p6_tier2_iosf_idf_side_clk,
  visa_p7_tier1_iosf_idf_side_clk,
  visa_p7_tier2_iosf_idf_side_clk,
  visa_p8_tier1_iosf_idf_side_clk,
  visa_p8_tier2_iosf_idf_side_clk,


  // Register wires
  dfxa_sbr1_cgovrd,
  dfxa_sbr1_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  ccsb_sbr1_side_ism_agent,
  sbr1_ccsb_side_ism_fabric,
  ccsb_sbr1_pccup,
  ccsb_sbr1_npcup,
  sbr1_ccsb_pcput,
  sbr1_ccsb_npput,
  sbr1_ccsb_eom,
  sbr1_ccsb_payload,
  sbr1_ccsb_pccup,
  sbr1_ccsb_npcup,
  ccsb_sbr1_pcput,
  ccsb_sbr1_npput,
  ccsb_sbr1_eom,
  ccsb_sbr1_payload,

  // Port 1 declarations
  fust_sbr1_side_ism_agent,
  sbr1_fust_side_ism_fabric,
  fust_sbr1_pccup,
  fust_sbr1_npcup,
  sbr1_fust_pcput,
  sbr1_fust_npput,
  sbr1_fust_eom,
  sbr1_fust_payload,
  sbr1_fust_pccup,
  sbr1_fust_npcup,
  fust_sbr1_pcput,
  fust_sbr1_npput,
  fust_sbr1_eom,
  fust_sbr1_payload,

  // Port 2 declarations
  sbr2_sbr1_side_ism_fabric,
  sbr1_sbr2_side_ism_agent,
  sbr2_sbr1_pccup,
  sbr2_sbr1_npcup,
  sbr1_sbr2_pcput,
  sbr1_sbr2_npput,
  sbr1_sbr2_eom,
  sbr1_sbr2_payload,
  sbr1_sbr2_pccup,
  sbr1_sbr2_npcup,
  sbr2_sbr1_pcput,
  sbr2_sbr1_npput,
  sbr2_sbr1_eom,
  sbr2_sbr1_payload,

  // Port 3 declarations
  isa_sbr1_side_ism_agent,
  sbr1_isa_side_ism_fabric,
  isa_sbr1_pccup,
  isa_sbr1_npcup,
  sbr1_isa_pcput,
  sbr1_isa_npput,
  sbr1_isa_eom,
  sbr1_isa_payload,
  sbr1_isa_pccup,
  sbr1_isa_npcup,
  isa_sbr1_pcput,
  isa_sbr1_npput,
  isa_sbr1_eom,
  isa_sbr1_payload,

  // Port 4 declarations
  dfxa_sbr1_side_ism_agent,
  sbr1_dfxa_side_ism_fabric,
  dfxa_sbr1_pccup,
  dfxa_sbr1_npcup,
  sbr1_dfxa_pcput,
  sbr1_dfxa_npput,
  sbr1_dfxa_eom,
  sbr1_dfxa_payload,
  sbr1_dfxa_pccup,
  sbr1_dfxa_npcup,
  dfxa_sbr1_pcput,
  dfxa_sbr1_npput,
  dfxa_sbr1_eom,
  dfxa_sbr1_payload,

  // Port 5 declarations
  scu0_sbr1_side_ism_agent,
  sbr1_scu0_side_ism_fabric,
  scu0_sbr1_pccup,
  scu0_sbr1_npcup,
  sbr1_scu0_pcput,
  sbr1_scu0_npput,
  sbr1_scu0_eom,
  sbr1_scu0_payload,
  sbr1_scu0_pccup,
  sbr1_scu0_npcup,
  scu0_sbr1_pcput,
  scu0_sbr1_npput,
  scu0_sbr1_eom,
  scu0_sbr1_payload,

  // Port 6 declarations
  scu1_sbr1_side_ism_agent,
  sbr1_scu1_side_ism_fabric,
  scu1_sbr1_pccup,
  scu1_sbr1_npcup,
  sbr1_scu1_pcput,
  sbr1_scu1_npput,
  sbr1_scu1_eom,
  sbr1_scu1_payload,
  sbr1_scu1_pccup,
  sbr1_scu1_npcup,
  scu1_sbr1_pcput,
  scu1_sbr1_npput,
  scu1_sbr1_eom,
  scu1_sbr1_payload,

  // Port 7 declarations
  idf_sbr1_side_ism_agent,
  sbr1_idf_side_ism_fabric,
  idf_sbr1_pccup,
  idf_sbr1_npcup,
  sbr1_idf_pcput,
  sbr1_idf_npput,
  sbr1_idf_eom,
  sbr1_idf_payload,
  sbr1_idf_pccup,
  sbr1_idf_npcup,
  idf_sbr1_pcput,
  idf_sbr1_npput,
  idf_sbr1_eom,
  idf_sbr1_payload,

  // Port 8 declarations
  rsp_sbr1_side_ism_agent,
  sbr1_rsp_side_ism_fabric,
  rsp_sbr1_pccup,
  rsp_sbr1_npcup,
  sbr1_rsp_pcput,
  sbr1_rsp_npput,
  sbr1_rsp_eom,
  sbr1_rsp_payload,
  sbr1_rsp_pccup,
  sbr1_rsp_npcup,
  rsp_sbr1_pcput,
  rsp_sbr1_npput,
  rsp_sbr1_eom,
  rsp_sbr1_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic iosf_idf_side_clk;
  input logic iosf_idf_side_rst_b;

  // Asynchronous Clock/Reset(s)
  input logic iosf_fust_side_clk;
  input logic iosf_swf_side_clk;

  // Power Well Isolation Input Signals
  input logic crp_sbr1_xu_en;
  input logic crp_sbr1_scu1_en;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic p3_fab_init_idle_exit;
  input logic p3_fab_init_idle_exit_ack;
  output logic p4_fab_init_idle_exit;
  input logic p4_fab_init_idle_exit_ack;
  output logic p5_fab_init_idle_exit;
  input logic p5_fab_init_idle_exit_ack;
  output logic p6_fab_init_idle_exit;
  input logic p6_fab_init_idle_exit_ack;
  output logic p7_fab_init_idle_exit;
  input logic p7_fab_init_idle_exit_ack;
  output logic p8_fab_init_idle_exit;
  input logic p8_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_iosf_idf_side_clk;
  output visa_vp  visa_vp_iosf_idf_side_clk;
  output visa_port_tier1 visa_p0_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p0_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p1_tier1_iosf_fust_side_clk;
  output visa_port_tier2 visa_p1_tier2_iosf_fust_side_clk;
  output visa_ififo_tier1 visa_p1_ififo_tier1_iosf_idf_side_clk;
  output visa_ififo_tier2 visa_p1_ififo_tier2_iosf_idf_side_clk;
  output visa_efifo_tier1 visa_p1_efifo_tier1_iosf_idf_side_clk;
  output visa_efifo_tier2 visa_p1_efifo_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p2_tier1_iosf_swf_side_clk;
  output visa_port_tier2 visa_p2_tier2_iosf_swf_side_clk;
  output visa_ififo_tier1 visa_p2_ififo_tier1_iosf_idf_side_clk;
  output visa_ififo_tier2 visa_p2_ififo_tier2_iosf_idf_side_clk;
  output visa_efifo_tier1 visa_p2_efifo_tier1_iosf_idf_side_clk;
  output visa_efifo_tier2 visa_p2_efifo_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p3_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p3_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p4_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p4_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p5_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p5_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p6_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p6_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p7_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p7_tier2_iosf_idf_side_clk;
  output visa_port_tier1 visa_p8_tier1_iosf_idf_side_clk;
  output visa_port_tier2 visa_p8_tier2_iosf_idf_side_clk;

  // Register wires
  input logic [4:0]  dfxa_sbr1_cgovrd;
  input logic [15:0] dfxa_sbr1_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic [1:0] fscan_rstbypen;
  input logic [1:0] fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] ccsb_sbr1_side_ism_agent;
  output logic [2:0] sbr1_ccsb_side_ism_fabric;
  input logic ccsb_sbr1_pccup;
  input logic ccsb_sbr1_npcup;
  output logic sbr1_ccsb_pcput;
  output logic sbr1_ccsb_npput;
  output logic sbr1_ccsb_eom;
  output logic [7:0] sbr1_ccsb_payload;
  output logic sbr1_ccsb_pccup;
  output logic sbr1_ccsb_npcup;
  input logic ccsb_sbr1_pcput;
  input logic ccsb_sbr1_npput;
  input logic ccsb_sbr1_eom;
  input logic [7:0] ccsb_sbr1_payload;

  // Port 1 declarations
  input logic [2:0] fust_sbr1_side_ism_agent;
  output logic [2:0] sbr1_fust_side_ism_fabric;
  input logic fust_sbr1_pccup;
  input logic fust_sbr1_npcup;
  output logic sbr1_fust_pcput;
  output logic sbr1_fust_npput;
  output logic sbr1_fust_eom;
  output logic [7:0] sbr1_fust_payload;
  output logic sbr1_fust_pccup;
  output logic sbr1_fust_npcup;
  input logic fust_sbr1_pcput;
  input logic fust_sbr1_npput;
  input logic fust_sbr1_eom;
  input logic [7:0] fust_sbr1_payload;

  // Port 2 declarations
  input logic [2:0] sbr2_sbr1_side_ism_fabric;
  output logic [2:0] sbr1_sbr2_side_ism_agent;
  input logic sbr2_sbr1_pccup;
  input logic sbr2_sbr1_npcup;
  output logic sbr1_sbr2_pcput;
  output logic sbr1_sbr2_npput;
  output logic sbr1_sbr2_eom;
  output logic [7:0] sbr1_sbr2_payload;
  output logic sbr1_sbr2_pccup;
  output logic sbr1_sbr2_npcup;
  input logic sbr2_sbr1_pcput;
  input logic sbr2_sbr1_npput;
  input logic sbr2_sbr1_eom;
  input logic [7:0] sbr2_sbr1_payload;

  // Port 3 declarations
  input logic [2:0] isa_sbr1_side_ism_agent;
  output logic [2:0] sbr1_isa_side_ism_fabric;
  input logic isa_sbr1_pccup;
  input logic isa_sbr1_npcup;
  output logic sbr1_isa_pcput;
  output logic sbr1_isa_npput;
  output logic sbr1_isa_eom;
  output logic [7:0] sbr1_isa_payload;
  output logic sbr1_isa_pccup;
  output logic sbr1_isa_npcup;
  input logic isa_sbr1_pcput;
  input logic isa_sbr1_npput;
  input logic isa_sbr1_eom;
  input logic [7:0] isa_sbr1_payload;

  // Port 4 declarations
  input logic [2:0] dfxa_sbr1_side_ism_agent;
  output logic [2:0] sbr1_dfxa_side_ism_fabric;
  input logic dfxa_sbr1_pccup;
  input logic dfxa_sbr1_npcup;
  output logic sbr1_dfxa_pcput;
  output logic sbr1_dfxa_npput;
  output logic sbr1_dfxa_eom;
  output logic [7:0] sbr1_dfxa_payload;
  output logic sbr1_dfxa_pccup;
  output logic sbr1_dfxa_npcup;
  input logic dfxa_sbr1_pcput;
  input logic dfxa_sbr1_npput;
  input logic dfxa_sbr1_eom;
  input logic [7:0] dfxa_sbr1_payload;

  // Port 5 declarations
  input logic [2:0] scu0_sbr1_side_ism_agent;
  output logic [2:0] sbr1_scu0_side_ism_fabric;
  input logic scu0_sbr1_pccup;
  input logic scu0_sbr1_npcup;
  output logic sbr1_scu0_pcput;
  output logic sbr1_scu0_npput;
  output logic sbr1_scu0_eom;
  output logic [7:0] sbr1_scu0_payload;
  output logic sbr1_scu0_pccup;
  output logic sbr1_scu0_npcup;
  input logic scu0_sbr1_pcput;
  input logic scu0_sbr1_npput;
  input logic scu0_sbr1_eom;
  input logic [7:0] scu0_sbr1_payload;

  // Port 6 declarations
  input logic [2:0] scu1_sbr1_side_ism_agent;
  output logic [2:0] sbr1_scu1_side_ism_fabric;
  input logic scu1_sbr1_pccup;
  input logic scu1_sbr1_npcup;
  output logic sbr1_scu1_pcput;
  output logic sbr1_scu1_npput;
  output logic sbr1_scu1_eom;
  output logic [7:0] sbr1_scu1_payload;
  output logic sbr1_scu1_pccup;
  output logic sbr1_scu1_npcup;
  input logic scu1_sbr1_pcput;
  input logic scu1_sbr1_npput;
  input logic scu1_sbr1_eom;
  input logic [7:0] scu1_sbr1_payload;

  // Port 7 declarations
  input logic [2:0] idf_sbr1_side_ism_agent;
  output logic [2:0] sbr1_idf_side_ism_fabric;
  input logic idf_sbr1_pccup;
  input logic idf_sbr1_npcup;
  output logic sbr1_idf_pcput;
  output logic sbr1_idf_npput;
  output logic sbr1_idf_eom;
  output logic [7:0] sbr1_idf_payload;
  output logic sbr1_idf_pccup;
  output logic sbr1_idf_npcup;
  input logic idf_sbr1_pcput;
  input logic idf_sbr1_npput;
  input logic idf_sbr1_eom;
  input logic [7:0] idf_sbr1_payload;

  // Port 8 declarations
  input logic [2:0] rsp_sbr1_side_ism_agent;
  output logic [2:0] sbr1_rsp_side_ism_fabric;
  input logic rsp_sbr1_pccup;
  input logic rsp_sbr1_npcup;
  output logic sbr1_rsp_pcput;
  output logic sbr1_rsp_npput;
  output logic sbr1_rsp_eom;
  output logic [7:0] sbr1_rsp_payload;
  output logic sbr1_rsp_pccup;
  output logic sbr1_rsp_npcup;
  input logic rsp_sbr1_pcput;
  input logic rsp_sbr1_npput;
  input logic rsp_sbr1_eom;
  input logic [7:0] rsp_sbr1_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr1_sbcportmap;
always_comb sbr1_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr1 (sbr1)                                   SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {   15 { 17'b0_0000_0000_0000_0000 }},   //   254:240      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //   239:238      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   237          SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //   236:234      SBCPORTMAPTABLE
      {  224 { 17'b0_0000_0000_0000_0000 }},   //   233: 10      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0100 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //     7          SBCPORTMAPTABLE
               17'b0_0000_0001_0000_0000,      //     6          SBCPORTMAPTABLE
               17'b0_0000_0000_1000_0000,      //     5          SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //     4          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //     3          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //     2          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //     1          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010       //     0          SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  8;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;
logic                              p6_pcdstvld;
logic                              p7_pcdstvld;
logic                              p8_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic                              p6_npfence;
logic                              p7_npfence;
logic                              p8_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;
logic                              p6_npdstvld;
logic                              p7_npdstvld;
logic                              p8_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              p3_ism_idle;
logic                              p3_cg_inprogress;
logic                              p3_credit_reinit;
logic                              p4_ism_idle;
logic                              p4_cg_inprogress;
logic                              p4_credit_reinit;
logic                              p5_ism_idle;
logic                              p5_cg_inprogress;
logic                              p5_credit_reinit;
logic                              p6_ism_idle;
logic                              p6_cg_inprogress;
logic                              p6_credit_reinit;
logic                              p7_ism_idle;
logic                              p7_cg_inprogress;
logic                              p7_credit_reinit;
logic                              p8_ism_idle;
logic                              p8_cg_inprogress;
logic                              p8_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              crp_sbr1_xu_en_ff2;
logic                              crp_sbr1_scu1_en_ff2;
logic                              iosf_swf_side_clk_crp_sbr1_xu_en_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = dfxa_sbr1_cgctrl[15];
always_comb cfg_clkgatedef    = dfxa_sbr1_cgctrl[14];
always_comb cfg_idlecnt       = dfxa_sbr1_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = dfxa_sbr1_cgovrd[3];
always_comb jta_force_idle    = dfxa_sbr1_cgovrd[1];
always_comb jta_force_notidle = dfxa_sbr1_cgovrd[0];
always_comb jta_force_creditreq = dfxa_sbr1_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

// Asynchronous port signals
logic                              p1_clkgaten;
logic                              p1_clkgatedef;
logic                              p1_clkgate_ovrd;
logic                              p1_force_idle;
logic                              p1_force_notidle;
logic                              p1_force_creditreq;
logic                              p1_clken;
logic                              p1_gated_clk;
logic                              p1_agent_idle;
logic                              p1_eagent_idle;
logic                              p1_port_idle;
logic                              p1_ififo_idle;
logic                              p1_efifo_idle;
logic                              p1_pctrdy;
logic                              p1_pcirdy;
logic             [INTMAXPLDBIT:0] p1_pcdata;
logic                              p1_pceom;
logic                              p1_nptrdy;
logic                              p1_npirdy;
logic                              p1_npfence;
logic             [INTMAXPLDBIT:0] p1_npdata;
logic                              p1_npeom;
logic                              p1_enpstall;
logic                              p1_epctrdy;
logic                              p1_enptrdy;
logic                              p1_epcirdy;
logic                              p1_enpirdy;
logic                              p1_eom;
logic             [INTMAXPLDBIT:0] p1_data;

logic                              p2_clkgaten;
logic                              p2_clkgatedef;
logic                              p2_clkgate_ovrd;
logic                              p2_force_idle;
logic                              p2_force_notidle;
logic                              p2_force_creditreq;
logic                              p2_clken;
logic                              p2_gated_clk;
logic                              p2_agent_idle;
logic                              p2_eagent_idle;
logic                              p2_port_idle;
logic                              p2_ififo_idle;
logic                              p2_efifo_idle;
logic                              p2_pctrdy;
logic                              p2_pcirdy;
logic             [INTMAXPLDBIT:0] p2_pcdata;
logic                              p2_pceom;
logic                              p2_nptrdy;
logic                              p2_npirdy;
logic                              p2_npfence;
logic             [INTMAXPLDBIT:0] p2_npdata;
logic                              p2_npeom;
logic                              p2_enpstall;
logic                              p2_epctrdy;
logic                              p2_enptrdy;
logic                              p2_epcirdy;
logic                              p2_enpirdy;
logic                              p2_eom;
logic             [INTMAXPLDBIT:0] p2_data;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr1_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr1_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// Async clock reset synchronization
//
//------------------------------------------------------------------------------
logic iosf_fust_side_clk_rst_b, iosf_fust_side_clk_rst_b_pre;
sbc_doublesync sync_rst_iosf_fust_side_clk (
  .d     ( 1'b1 ),
  .clr_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_fust_side_clk ),
  .q     ( iosf_fust_side_clk_rst_b_pre ));

always_comb iosf_fust_side_clk_rst_b = fscan_rstbypen[0] ? fscan_byprst_b[0] : iosf_fust_side_clk_rst_b_pre;

logic iosf_swf_side_clk_rst_b, iosf_swf_side_clk_rst_b_pre;
sbc_doublesync sync_rst_iosf_swf_side_clk (
  .d     ( 1'b1 ),
  .clr_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_swf_side_clk ),
  .q     ( iosf_swf_side_clk_rst_b_pre ));

always_comb iosf_swf_side_clk_rst_b = fscan_rstbypen[1] ? fscan_byprst_b[1] : iosf_swf_side_clk_rst_b_pre;


//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( iosf_idf_side_rst_b           ),
  .clk                 ( iosf_idf_side_clk             ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( iosf_idf_side_rst_b           ),
  .clk                 ( iosf_idf_side_clk             ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( iosf_idf_side_rst_b           ),
  .clk                 ( iosf_idf_side_clk             ),
  .q                   ( force_creditreq               )
);

sbc_doublesync sync_p2_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_force_idle                 )
);

sbc_doublesync sync_p2_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_force_notidle              )
);

sbc_doublesync sync_p2_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_force_creditreq            )
);

sbc_doublesync sync_p1_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_force_idle                 )
);

sbc_doublesync sync_p1_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_force_notidle              )
);

sbc_doublesync sync_p1_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_force_creditreq            )
);

//------------------------------------------------------------------------------
//
// Asynchronous port local clock gating
//
//------------------------------------------------------------------------------
// Port 2
sbc_doublesync sync_p2_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_clkgaten                   )
);

sbc_doublesync sync_p2_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_clkgatedef                 )
);

sbc_doublesync sync_p2_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( p2_clkgate_ovrd               )
);

always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_clk_rst_b)
  if (~iosf_swf_side_clk_rst_b)
    p2_clken <= '1;
  else
    p2_clken <= ~p2_clkgate_ovrd &
    iosf_swf_side_clk_crp_sbr1_xu_en_ff2 &
      (p2_clkgatedef | ~p2_clkgaten | ~p2_cg_inprogress |
       ((sbr1_sbr2_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr2_sbr1_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (sbr1_sbr2_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((sbr1_sbr2_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr2_sbr1_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p2_clkgate  (
  .en                  ( p2_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( iosf_swf_side_clk             ),
  .enclk               ( p2_gated_clk                  )
);

// Port 1
sbc_doublesync sync_p1_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_clkgaten                   )
);

sbc_doublesync sync_p1_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_clkgatedef                 )
);

sbc_doublesync sync_p1_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk                 ( iosf_fust_side_clk            ),
  .q                   ( p1_clkgate_ovrd               )
);

always_ff @(posedge iosf_fust_side_clk or negedge iosf_fust_side_clk_rst_b)
  if (~iosf_fust_side_clk_rst_b)
    p1_clken <= '1;
  else
    p1_clken <= ~p1_clkgate_ovrd &
      (p1_clkgatedef | ~p1_clkgaten | ~p1_cg_inprogress |
       ((fust_sbr1_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr1_fust_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (fust_sbr1_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((fust_sbr1_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr1_fust_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p1_clkgate  (
  .en                  ( p1_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( iosf_fust_side_clk            ),
  .enclk               ( p1_gated_clk                  )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_crp_sbr1_xu_en (
  .d                   ( crp_sbr1_xu_en                ),
  .clr_b               ( iosf_idf_side_rst_b           ),
  .clk                 ( iosf_idf_side_clk             ),
  .q                   ( crp_sbr1_xu_en_ff2            )
);

sbc_doublesync sync_crp_sbr1_scu1_en (
  .d                   ( crp_sbr1_scu1_en              ),
  .clr_b               ( iosf_idf_side_rst_b           ),
  .clk                 ( iosf_idf_side_clk             ),
  .q                   ( crp_sbr1_scu1_en_ff2          )
);

sbc_doublesync sync_crp_sbr1_xu_en_iosf_swf_side_clk (
  .d                   ( crp_sbr1_xu_en                ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( iosf_swf_side_clk_crp_sbr1_xu_en_ff2 )
);


always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          crp_sbr1_scu1_en_ff2,
                          1'b1,
                          1'b1,
                          1'b1,
                          crp_sbr1_xu_en_ff2,
                          1'b1,
                          1'b1
                        };

logic p6_gated_clk;
sbc_clock_gate p6_pwr_clkgate  (
  .en ( endpoint_pwrgd[6] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p6_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p8_ism_idle | ~endpoint_pwrgd[8])
                  &  (p7_ism_idle | ~endpoint_pwrgd[7])
                  &  (p6_ism_idle | ~endpoint_pwrgd[6])
                  &  (p5_ism_idle | ~endpoint_pwrgd[5])
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  &  p2_efifo_idle
                  &  p1_efifo_idle
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
logic p1_ism_idle_ff2, p1_ism_idle_pre;
always_ff @(posedge iosf_fust_side_clk or negedge iosf_fust_side_clk_rst_b)
  if ( ~iosf_fust_side_clk_rst_b)
    p1_ism_idle_pre <= '1;
  else
    p1_ism_idle_pre <= p1_ism_idle;

sbc_doublesync sync_idle_p1 (
  .d ( p1_ism_idle_pre ),
  .clr_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_idf_side_clk ),
  .q     ( p1_ism_idle_ff2 ));

logic p2_ism_idle_ff2, p2_ism_idle_pre;
always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_clk_rst_b)
  if ( ~iosf_swf_side_clk_rst_b)
    p2_ism_idle_pre <= '1;
  else
    p2_ism_idle_pre <= p2_ism_idle;

sbc_doublesync sync_idle_p2 (
  .d ( p2_ism_idle_pre ),
  .clr_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_idf_side_clk ),
  .q     ( p2_ism_idle_ff2 ));

// SBR_IDLE signal for PMU
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle_ff2 &
                  p2_ism_idle_ff2 &
                  p3_ism_idle &
                  p4_ism_idle &
                  p5_ism_idle &
                  p6_ism_idle &
                  p7_ism_idle &
                  p8_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p8_npfence,
                 p7_npfence,
                 p6_npfence,
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 1'b0,
                 1'b0,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p8_pcdstvld,
                 p7_pcdstvld,
                 p6_pcdstvld,
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 pcirdy[2],
                 pcirdy[1],
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p8_npdstvld,
                 p7_npdstvld,
                 p6_npdstvld,
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 npirdy[2],
                 npirdy[1],
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_iosf_idf_side_clk = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( iosf_idf_side_clk             ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_iosf_idf_side_clk = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle & agent_idle[0] & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle & p0_side_clk_valid )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_iosf_idf_side_clk = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_iosf_idf_side_clk = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( ccsb_sbr1_side_ism_agent      ),
  .side_ism_out        ( sbr1_ccsb_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr1_ccsb_pccup               ),
  .tnpcup              ( sbr1_ccsb_npcup               ),
  .tpcput              ( ccsb_sbr1_pcput               ),
  .tnpput              ( ccsb_sbr1_npput               ),
  .teom                ( ccsb_sbr1_eom                 ),
  .tpayload            ( ccsb_sbr1_payload             ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( ccsb_sbr1_pccup               ),
  .mnpcup              ( ccsb_sbr1_npcup               ),
  .mpcput              ( sbr1_ccsb_pcput               ),
  .mnpput              ( sbr1_ccsb_npput               ),
  .meom                ( sbr1_ccsb_eom                 ),
  .mpayload            ( sbr1_ccsb_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1 (Asynchronous port)
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  logic p1_credit_reinit_ff2;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit_ff2 & p1_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & (~agent_idle[1] || ~p1_efifo_idle) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & agent_idle[1] & p1_efifo_idle & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle_ff2 & p1_side_clk_valid & ~p1_fab_init_idle_exit )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle_ff2 )
          p1_side_clk_valid <= '1;
      end

logic p1_side_clk_valid_ff2;
sbc_doublesync sync_p1_clk_valid (
  .d     ( p1_side_clk_valid ),
  .clr_b ( iosf_fust_side_clk_rst_b ),
  .clk   ( iosf_fust_side_clk ),
  .q     ( p1_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p1_credit_reinit (
  .d     ( p1_credit_reinit ),
  .set_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_idf_side_clk ),
  .q     ( p1_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

logic [15:0] p1_dbgbus_ing;
logic [15:0] p1_dbgbus_egr;
  always_comb
    begin
      visa_p1_tier1_iosf_fust_side_clk = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_iosf_fust_side_clk = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
      visa_p1_ififo_tier1_iosf_idf_side_clk = { p1_dbgbus_ing[15:14],
                             p1_dbgbus_ing[5:0]};
      visa_p1_ififo_tier2_iosf_idf_side_clk = { p1_dbgbus_ing[13:6] };
      visa_p1_efifo_tier1_iosf_idf_side_clk = { p1_dbgbus_egr[7:0] };
      visa_p1_efifo_tier2_iosf_idf_side_clk = { p1_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( iosf_fust_side_clk            ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b ( iosf_fust_side_clk_rst_b ),
  .side_clk_valid      ( p1_side_clk_valid_ff2         ),
  .side_ism_in         ( fust_sbr1_side_ism_agent      ),
  .side_ism_out        ( sbr1_fust_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( p1_agent_idle                 ),
  .port_idle           ( p1_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr1_fust_pccup               ),
  .tnpcup              ( sbr1_fust_npcup               ),
  .tpcput              ( fust_sbr1_pcput               ),
  .tnpput              ( fust_sbr1_npput               ),
  .teom                ( fust_sbr1_eom                 ),
  .tpayload            ( fust_sbr1_payload             ),
  .pctrdy              ( p1_pctrdy                     ),
  .pcirdy              ( p1_pcirdy                     ),
  .pcdata              ( p1_pcdata                     ),
  .pceom               ( p1_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p1_nptrdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( p1_npdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( fust_sbr1_pccup               ),
  .mnpcup              ( fust_sbr1_npcup               ),
  .mpcput              ( sbr1_fust_pcput               ),
  .mnpput              ( sbr1_fust_npput               ),
  .meom                ( sbr1_fust_eom                 ),
  .mpayload            ( sbr1_fust_payload             ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .data                ( p1_data                       ),
  .eom                 ( p1_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p1_clkgaten                   ),
  .force_idle          ( p1_force_idle                 ),
  .force_notidle       ( p1_force_notidle              ),
  .force_creditreq     ( p1_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress1 (
  .ing_side_clk        ( p1_gated_clk                  ),
  .ing_side_rst_b ( iosf_fust_side_clk_rst_b ),
  .port_idle           ( p1_port_idle                  ),
  .pcirdy              ( p1_pcirdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .pceom               ( p1_pceom                      ),
  .pcdata              ( p1_pcdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdata              ( p1_npdata                     ),
  .pctrdy              ( p1_pctrdy                     ),
  .nptrdy              ( p1_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p1_ififo_idle                 ),
  .egr_side_clk        ( iosf_idf_side_clk             ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( iosf_idf_side_rst_b           ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[1]                     ),
  .enptrdy             ( nptrdy[1]                     ),
  .epcirdy             ( pcirdy[1]                     ),
  .enpirdy             ( npirdy[1]                     ),
  .eom                 ( npeom[1]                      ),
  .data                ( npdata[1]                     ),
  .opceom              ( pceom[1]                      ),
  .opcdata             ( pcdata[1]                     ),
  .agent_idle          ( port_idle[1]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p1_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress1 (
  .ing_side_clk        ( iosf_idf_side_clk             ),
  .ing_side_rst_b      ( iosf_idf_side_rst_b           ),
  .port_idle           ( agent_idle[1]                 ),
  .pcirdy              ( epcirdy[1]                    ),
  .npirdy              ( enpirdy[1]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[1]                    ),
  .nptrdy              ( enptrdy[1]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p1_efifo_idle                 ),
  .egr_side_clk        ( iosf_fust_side_clk            ),
  .gated_egr_side_clk  ( p1_gated_clk                  ),
  .egr_side_rst_b ( iosf_fust_side_clk_rst_b ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .eom                 ( p1_eom                        ),
  .data                ( p1_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p1_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p1_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p1_agent_idle  = p1_eagent_idle & p1_ififo_idle;

// Port 2 (Asynchronous port)
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  logic p2_credit_reinit_ff2;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit_ff2 & p2_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle_ff2 & (~agent_idle[2] || ~p2_efifo_idle) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle_ff2 & agent_idle[2] & p2_efifo_idle & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle_ff2 & p2_side_clk_valid & ~p2_fab_init_idle_exit )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle_ff2 )
          p2_side_clk_valid <= '1;
      end

logic p2_side_clk_valid_ff2;
sbc_doublesync sync_p2_clk_valid (
  .d     ( p2_side_clk_valid ),
  .clr_b ( iosf_swf_side_clk_rst_b ),
  .clk   ( iosf_swf_side_clk ),
  .q     ( p2_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p2_credit_reinit (
  .d     ( p2_credit_reinit ),
  .set_b ( iosf_idf_side_rst_b ),
  .clk   ( iosf_idf_side_clk ),
  .q     ( p2_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

logic [15:0] p2_dbgbus_ing;
logic [15:0] p2_dbgbus_egr;
  always_comb
    begin
      visa_p2_tier1_iosf_swf_side_clk = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_iosf_swf_side_clk = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
      visa_p2_ififo_tier1_iosf_idf_side_clk = { p2_dbgbus_ing[15:14],
                             p2_dbgbus_ing[5:0]};
      visa_p2_ififo_tier2_iosf_idf_side_clk = { p2_dbgbus_ing[13:6] };
      visa_p2_efifo_tier1_iosf_idf_side_clk = { p2_dbgbus_egr[7:0] };
      visa_p2_efifo_tier2_iosf_idf_side_clk = { p2_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  1                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( iosf_swf_side_clk             ),
  .gated_side_clk      ( p2_gated_clk                  ),
  .side_rst_b ( iosf_swf_side_clk_rst_b ),
  .side_clk_valid      ( p2_side_clk_valid_ff2         ),
  .side_ism_in         ( sbr2_sbr1_side_ism_fabric     ),
  .side_ism_out        ( sbr1_sbr2_side_ism_agent      ),
  .int_pok             (  iosf_swf_side_clk_crp_sbr1_xu_en_ff2 ), 
  .agent_idle          ( p2_agent_idle                 ),
  .port_idle           ( p2_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr1_sbr2_pccup               ),
  .tnpcup              ( sbr1_sbr2_npcup               ),
  .tpcput              ( sbr2_sbr1_pcput               ),
  .tnpput              ( sbr2_sbr1_npput               ),
  .teom                ( sbr2_sbr1_eom                 ),
  .tpayload            ( sbr2_sbr1_payload             ),
  .pctrdy              ( p2_pctrdy                     ),
  .pcirdy              ( p2_pcirdy                     ),
  .pcdata              ( p2_pcdata                     ),
  .pceom               ( p2_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p2_nptrdy                     ),
  .npirdy              ( p2_npirdy                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( p2_npdata                     ),
  .npeom               ( p2_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( sbr2_sbr1_pccup               ),
  .mnpcup              ( sbr2_sbr1_npcup               ),
  .mpcput              ( sbr1_sbr2_pcput               ),
  .mnpput              ( sbr1_sbr2_npput               ),
  .meom                ( sbr1_sbr2_eom                 ),
  .mpayload            ( sbr1_sbr2_payload             ),
  .enpstall            ( p2_enpstall                   ),
  .epctrdy             ( p2_epctrdy                    ),
  .enptrdy             ( p2_enptrdy                    ),
  .epcirdy             ( p2_epcirdy                    ),
  .enpirdy             ( p2_enpirdy                    ),
  .data                ( p2_data                       ),
  .eom                 ( p2_eom                        ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .cfg_clkgaten        ( p2_clkgaten                   ),
  .force_idle          ( p2_force_idle                 ),
  .force_notidle       ( p2_force_notidle              ),
  .force_creditreq     ( p2_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress2 (
  .ing_side_clk        ( p2_gated_clk                  ),
  .ing_side_rst_b ( iosf_swf_side_clk_rst_b ),
  .port_idle           ( p2_port_idle                  ),
  .pcirdy              ( p2_pcirdy                     ),
  .npirdy              ( p2_npirdy                     ),
  .npfence             ( p2_npfence                    ),
  .pceom               ( p2_pceom                      ),
  .pcdata              ( p2_pcdata                     ),
  .npeom               ( p2_npeom                      ),
  .npdata              ( p2_npdata                     ),
  .pctrdy              ( p2_pctrdy                     ),
  .nptrdy              ( p2_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p2_ififo_idle                 ),
  .egr_side_clk        ( iosf_idf_side_clk             ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( iosf_idf_side_rst_b           ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[2]                     ),
  .enptrdy             ( nptrdy[2]                     ),
  .epcirdy             ( pcirdy[2]                     ),
  .enpirdy             ( npirdy[2]                     ),
  .eom                 ( npeom[2]                      ),
  .data                ( npdata[2]                     ),
  .opceom              ( pceom[2]                      ),
  .opcdata             ( pcdata[2]                     ),
  .agent_idle          ( port_idle[2]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p2_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress2 (
  .ing_side_clk        ( iosf_idf_side_clk             ),
  .ing_side_rst_b      ( iosf_idf_side_rst_b           ),
  .port_idle           ( agent_idle[2]                 ),
  .pcirdy              ( epcirdy[2]                    ),
  .npirdy              ( enpirdy[2]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[2]                    ),
  .nptrdy              ( enptrdy[2]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p2_efifo_idle                 ),
  .egr_side_clk        ( iosf_swf_side_clk             ),
  .gated_egr_side_clk  ( p2_gated_clk                  ),
  .egr_side_rst_b ( iosf_swf_side_clk_rst_b ),
  .enpstall            ( p2_enpstall                   ),
  .epctrdy             ( p2_epctrdy                    ),
  .enptrdy             ( p2_enptrdy                    ),
  .epcirdy             ( p2_epcirdy                    ),
  .enpirdy             ( p2_enpirdy                    ),
  .eom                 ( p2_eom                        ),
  .data                ( p2_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p2_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p2_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p2_agent_idle  = p2_eagent_idle & p2_ififo_idle;

// Port 3
logic p3_side_clk_valid, p3_idle_egress, p3_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p3_rst_suppress <= 1'b1;
    else
      p3_rst_suppress <= p3_credit_reinit & p3_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p3_fab_init_idle_exit <= '1;
    else
      if ( ~p3_rst_suppress & (p3_ism_idle & (~agent_idle[3] || ~p3_idle_egress) & ~p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '1;
      else if ( ~p3_rst_suppress & (p3_ism_idle & agent_idle[3] & p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( p3_ism_idle & p3_side_clk_valid )
          p3_side_clk_valid <= '0;
        else if ( (p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack) || ~p3_ism_idle )
          p3_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

  always_comb
    begin
      visa_p3_tier1_iosf_idf_side_clk = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_iosf_idf_side_clk = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( isa_sbr1_side_ism_agent       ),
  .side_ism_out        ( sbr1_isa_side_ism_fabric      ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .idle_egress         ( p3_idle_egress                ),
  .ism_idle            ( p3_ism_idle                   ),
  .credit_reinit       ( p3_credit_reinit              ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr1_isa_pccup                ),
  .tnpcup              ( sbr1_isa_npcup                ),
  .tpcput              ( isa_sbr1_pcput                ),
  .tnpput              ( isa_sbr1_npput                ),
  .teom                ( isa_sbr1_eom                  ),
  .tpayload            ( isa_sbr1_payload              ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( isa_sbr1_pccup                ),
  .mnpcup              ( isa_sbr1_npcup                ),
  .mpcput              ( sbr1_isa_pcput                ),
  .mnpput              ( sbr1_isa_npput                ),
  .meom                ( sbr1_isa_eom                  ),
  .mpayload            ( sbr1_isa_payload              ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
logic p4_side_clk_valid, p4_idle_egress, p4_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p4_rst_suppress <= 1'b1;
    else
      p4_rst_suppress <= p4_credit_reinit & p4_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p4_fab_init_idle_exit <= '1;
    else
      if ( ~p4_rst_suppress & (p4_ism_idle & (~agent_idle[4] || ~p4_idle_egress) & ~p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '1;
      else if ( ~p4_rst_suppress & (p4_ism_idle & agent_idle[4] & p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( p4_ism_idle & p4_side_clk_valid )
          p4_side_clk_valid <= '0;
        else if ( (p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack) || ~p4_ism_idle )
          p4_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

  always_comb
    begin
      visa_p4_tier1_iosf_idf_side_clk = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_iosf_idf_side_clk = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( dfxa_sbr1_side_ism_agent      ),
  .side_ism_out        ( sbr1_dfxa_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .idle_egress         ( p4_idle_egress                ),
  .ism_idle            ( p4_ism_idle                   ),
  .credit_reinit       ( p4_credit_reinit              ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr1_dfxa_pccup               ),
  .tnpcup              ( sbr1_dfxa_npcup               ),
  .tpcput              ( dfxa_sbr1_pcput               ),
  .tnpput              ( dfxa_sbr1_npput               ),
  .teom                ( dfxa_sbr1_eom                 ),
  .tpayload            ( dfxa_sbr1_payload             ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( dfxa_sbr1_pccup               ),
  .mnpcup              ( dfxa_sbr1_npcup               ),
  .mpcput              ( sbr1_dfxa_pcput               ),
  .mnpput              ( sbr1_dfxa_npput               ),
  .meom                ( sbr1_dfxa_eom                 ),
  .mpayload            ( sbr1_dfxa_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

// Port 5
logic p5_side_clk_valid, p5_idle_egress, p5_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p5_rst_suppress <= 1'b1;
    else
      p5_rst_suppress <= p5_credit_reinit & p5_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p5_fab_init_idle_exit <= '1;
    else
      if ( ~p5_rst_suppress & (p5_ism_idle & (~agent_idle[5] || ~p5_idle_egress) & ~p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '1;
      else if ( ~p5_rst_suppress & (p5_ism_idle & agent_idle[5] & p5_fab_init_idle_exit_ack ))
        p5_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p5_side_clk_valid <= 1'b0;
    else
      begin
        if ( p5_ism_idle & p5_side_clk_valid )
          p5_side_clk_valid <= '0;
        else if ( (p5_fab_init_idle_exit & p5_fab_init_idle_exit_ack) || ~p5_ism_idle )
          p5_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p5_dbgbus;

  always_comb
    begin
      visa_p5_tier1_iosf_idf_side_clk = { p5_dbgbus[31],
                            p5_dbgbus[27:24],
                            p5_dbgbus[21:19],
                            p5_dbgbus[15:12],
                            p5_dbgbus[7:4] };
      visa_p5_tier2_iosf_idf_side_clk = { p5_dbgbus[30:28],
                            p5_dbgbus[23:22],
                            p5_dbgbus[18:16],
                            p5_dbgbus[11:8],
                            p5_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport5 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( scu0_sbr1_side_ism_agent      ),
  .side_ism_out        ( sbr1_scu0_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[5] ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .idle_egress         ( p5_idle_egress                ),
  .ism_idle            ( p5_ism_idle                   ),
  .credit_reinit       ( p5_credit_reinit              ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr1_scu0_pccup               ),
  .tnpcup              ( sbr1_scu0_npcup               ),
  .tpcput              ( scu0_sbr1_pcput               ),
  .tnpput              ( scu0_sbr1_npput               ),
  .teom                ( scu0_sbr1_eom                 ),
  .tpayload            ( scu0_sbr1_payload             ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( scu0_sbr1_pccup               ),
  .mnpcup              ( scu0_sbr1_npcup               ),
  .mpcput              ( sbr1_scu0_pcput               ),
  .mnpput              ( sbr1_scu0_npput               ),
  .meom                ( sbr1_scu0_eom                 ),
  .mpayload            ( sbr1_scu0_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p5_dbgbus                     )
);

// Port 6
logic p6_side_clk_valid, p6_idle_egress, p6_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p6_rst_suppress <= 1'b1;
    else
      p6_rst_suppress <= p6_credit_reinit & p6_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p6_fab_init_idle_exit <= '1;
    else
      if ( ~p6_rst_suppress & (p6_ism_idle & (~agent_idle[6] || ~p6_idle_egress) & ~p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '1;
      else if ( ~p6_rst_suppress & (p6_ism_idle & agent_idle[6] & p6_fab_init_idle_exit_ack ))
        p6_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p6_side_clk_valid <= 1'b0;
    else
      begin
        if ( p6_ism_idle & p6_side_clk_valid )
          p6_side_clk_valid <= '0;
        else if ( (p6_fab_init_idle_exit & p6_fab_init_idle_exit_ack) || ~p6_ism_idle )
          p6_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p6_dbgbus;

  always_comb
    begin
      visa_p6_tier1_iosf_idf_side_clk = { p6_dbgbus[31],
                            p6_dbgbus[27:24],
                            p6_dbgbus[21:19],
                            p6_dbgbus[15:12],
                            p6_dbgbus[7:4] };
      visa_p6_tier2_iosf_idf_side_clk = { p6_dbgbus[30:28],
                            p6_dbgbus[23:22],
                            p6_dbgbus[18:16],
                            p6_dbgbus[11:8],
                            p6_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport6 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( p6_gated_clk                  ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p6_side_clk_valid             ),
  .side_ism_in         ( scu1_sbr1_side_ism_agent      ),
  .side_ism_out        ( sbr1_scu1_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[6] ),
  .agent_idle          ( agent_idle[6]                 ),
  .port_idle           ( port_idle[6]                  ),
  .idle_egress         ( p6_idle_egress                ),
  .ism_idle            ( p6_ism_idle                   ),
  .credit_reinit       ( p6_credit_reinit              ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr1_scu1_pccup               ),
  .tnpcup              ( sbr1_scu1_npcup               ),
  .tpcput              ( scu1_sbr1_pcput               ),
  .tnpput              ( scu1_sbr1_npput               ),
  .teom                ( scu1_sbr1_eom                 ),
  .tpayload            ( scu1_sbr1_payload             ),
  .pctrdy              ( pctrdy[6]                     ),
  .pcirdy              ( pcirdy[6]                     ),
  .pcdata              ( pcdata[6]                     ),
  .pceom               ( pceom[6]                      ),
  .pcdstvld            ( p6_pcdstvld                   ),
  .nptrdy              ( nptrdy[6]                     ),
  .npirdy              ( npirdy[6]                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( npdata[6]                     ),
  .npeom               ( npeom[6]                      ),
  .npdstvld            ( p6_npdstvld                   ),
  .mpccup              ( scu1_sbr1_pccup               ),
  .mnpcup              ( scu1_sbr1_npcup               ),
  .mpcput              ( sbr1_scu1_pcput               ),
  .mnpput              ( sbr1_scu1_npput               ),
  .meom                ( sbr1_scu1_eom                 ),
  .mpayload            ( sbr1_scu1_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[6]                    ),
  .enptrdy             ( enptrdy[6]                    ),
  .epcirdy             ( epcirdy[6]                    ),
  .enpirdy             ( enpirdy[6]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p6_dbgbus                     )
);

// Port 7
logic p7_side_clk_valid, p7_idle_egress, p7_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p7_rst_suppress <= 1'b1;
    else
      p7_rst_suppress <= p7_credit_reinit & p7_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p7_fab_init_idle_exit <= '1;
    else
      if ( ~p7_rst_suppress & (p7_ism_idle & (~agent_idle[7] || ~p7_idle_egress) & ~p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '1;
      else if ( ~p7_rst_suppress & (p7_ism_idle & agent_idle[7] & p7_fab_init_idle_exit_ack ))
        p7_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p7_side_clk_valid <= 1'b0;
    else
      begin
        if ( p7_ism_idle & p7_side_clk_valid )
          p7_side_clk_valid <= '0;
        else if ( (p7_fab_init_idle_exit & p7_fab_init_idle_exit_ack) || ~p7_ism_idle )
          p7_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p7_dbgbus;

  always_comb
    begin
      visa_p7_tier1_iosf_idf_side_clk = { p7_dbgbus[31],
                            p7_dbgbus[27:24],
                            p7_dbgbus[21:19],
                            p7_dbgbus[15:12],
                            p7_dbgbus[7:4] };
      visa_p7_tier2_iosf_idf_side_clk = { p7_dbgbus[30:28],
                            p7_dbgbus[23:22],
                            p7_dbgbus[18:16],
                            p7_dbgbus[11:8],
                            p7_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport7 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( idf_sbr1_side_ism_agent       ),
  .side_ism_out        ( sbr1_idf_side_ism_fabric      ),
  .int_pok             ( endpoint_pwrgd[7] ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .idle_egress         ( p7_idle_egress                ),
  .ism_idle            ( p7_ism_idle                   ),
  .credit_reinit       ( p7_credit_reinit              ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr1_idf_pccup                ),
  .tnpcup              ( sbr1_idf_npcup                ),
  .tpcput              ( idf_sbr1_pcput                ),
  .tnpput              ( idf_sbr1_npput                ),
  .teom                ( idf_sbr1_eom                  ),
  .tpayload            ( idf_sbr1_payload              ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( idf_sbr1_pccup                ),
  .mnpcup              ( idf_sbr1_npcup                ),
  .mpcput              ( sbr1_idf_pcput                ),
  .mnpput              ( sbr1_idf_npput                ),
  .meom                ( sbr1_idf_eom                  ),
  .mpayload            ( sbr1_idf_payload              ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p7_dbgbus                     )
);

// Port 8
logic p8_side_clk_valid, p8_idle_egress, p8_rst_suppress;
  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p8_rst_suppress <= 1'b1;
    else
      p8_rst_suppress <= p8_credit_reinit & p8_rst_suppress;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if (~iosf_idf_side_rst_b)
      p8_fab_init_idle_exit <= '1;
    else
      if ( ~p8_rst_suppress & (p8_ism_idle & (~agent_idle[8] || ~p8_idle_egress) & ~p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '1;
      else if ( ~p8_rst_suppress & (p8_ism_idle & agent_idle[8] & p8_fab_init_idle_exit_ack ))
        p8_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)
    if ( ~iosf_idf_side_rst_b )
      p8_side_clk_valid <= 1'b0;
    else
      begin
        if ( p8_ism_idle & p8_side_clk_valid )
          p8_side_clk_valid <= '0;
        else if ( (p8_fab_init_idle_exit & p8_fab_init_idle_exit_ack) || ~p8_ism_idle )
          p8_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p8_dbgbus;

  always_comb
    begin
      visa_p8_tier1_iosf_idf_side_clk = { p8_dbgbus[31],
                            p8_dbgbus[27:24],
                            p8_dbgbus[21:19],
                            p8_dbgbus[15:12],
                            p8_dbgbus[7:4] };
      visa_p8_tier2_iosf_idf_side_clk = { p8_dbgbus[30:28],
                            p8_dbgbus[23:22],
                            p8_dbgbus[18:16],
                            p8_dbgbus[11:8],
                            p8_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport8 (
  .side_clk            ( iosf_idf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_idf_side_rst_b           ),
  .side_clk_valid      ( p8_side_clk_valid             ),
  .side_ism_in         ( rsp_sbr1_side_ism_agent       ),
  .side_ism_out        ( sbr1_rsp_side_ism_fabric      ),
  .int_pok             ( endpoint_pwrgd[8] ),
  .agent_idle          ( agent_idle[8]                 ),
  .port_idle           ( port_idle[8]                  ),
  .idle_egress         ( p8_idle_egress                ),
  .ism_idle            ( p8_ism_idle                   ),
  .credit_reinit       ( p8_credit_reinit              ),
  .cg_inprogress       ( p8_cg_inprogress              ),
  .tpccup              ( sbr1_rsp_pccup                ),
  .tnpcup              ( sbr1_rsp_npcup                ),
  .tpcput              ( rsp_sbr1_pcput                ),
  .tnpput              ( rsp_sbr1_npput                ),
  .teom                ( rsp_sbr1_eom                  ),
  .tpayload            ( rsp_sbr1_payload              ),
  .pctrdy              ( pctrdy[8]                     ),
  .pcirdy              ( pcirdy[8]                     ),
  .pcdata              ( pcdata[8]                     ),
  .pceom               ( pceom[8]                      ),
  .pcdstvld            ( p8_pcdstvld                   ),
  .nptrdy              ( nptrdy[8]                     ),
  .npirdy              ( npirdy[8]                     ),
  .npfence             ( p8_npfence                    ),
  .npdata              ( npdata[8]                     ),
  .npeom               ( npeom[8]                      ),
  .npdstvld            ( p8_npdstvld                   ),
  .mpccup              ( rsp_sbr1_pccup                ),
  .mnpcup              ( rsp_sbr1_npcup                ),
  .mpcput              ( sbr1_rsp_pcput                ),
  .mnpput              ( sbr1_rsp_npput                ),
  .meom                ( sbr1_rsp_eom                  ),
  .mpayload            ( sbr1_rsp_payload              ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[8]                    ),
  .enptrdy             ( enptrdy[8]                    ),
  .epcirdy             ( epcirdy[8]                    ),
  .enpirdy             ( enpirdy[8]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p8_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr1_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr1_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge iosf_idf_side_clk or negedge iosf_idf_side_rst_b)

      if (~iosf_idf_side_rst_b) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge iosf_idf_side_clk) disable iff (iosf_idf_side_rst_b !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge iosf_idf_side_clk) disable iff (iosf_idf_side_rst_b !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 0, bb_cclk, bb_rst_b, 0, , 4ns
ClockReset, 3, iosf_fust_side_clk, iosf_fust_side_rst_b, 0, , 2ns
ClockReset, 4, iosf_idf_side_clk, iosf_idf_side_rst_b, 0, cgc0, 2ns
ClockReset, 5, iosf_swf_side_clk, iosf_swf_side_rst_b, 0, cgc1, 2ns
ClockReset, 1, sosc_125_clk_core, sbi_rst_125_core_b, 0, , 4ns
ClockReset, 2, sosc_25_clk_core, sbi_rst_25_core_b, 0, , 40ns
SyncRouter, ccsb, ccsb,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 2, sbra, sbr1, , , , , , , , , , , , , , , 
RouterAgentPort, ccsb, 0
RouterAgentPort, ccsb, 1
Endpoint, dfxa,1, 1, 4, 0, 3, 3, 1, 2, 3, 3, 
Endpoint, fust,1, 1, 3, 0, 3, 3, 1, 0, 3, 3, 
Endpoint, idf,1, 1, 4, 0, 3, 3, 1, 5, 3, 3, 
Endpoint, io_dmi,0, 1, 2, 0, 1, 1, 1, 235, 3, 3, 
Endpoint, io_pxp,0, 1, 2, 0, 1, 1, 1, 236, 3, 3, 
Endpoint, io_st,0, 1, 2, 0, 1, 1, 1, 234, 3, 3, 
Endpoint, isa,1, 1, 4, 0, 3, 3, 1, 1, 3, 3, 
Endpoint, npsb,0, 1, 0, 0, 1, 1, 1, 239, 3, 3, 
Endpoint, rsp,1, 1, 4, 0, 3, 3, 1, 6, 3, 3, 
SyncRouter, sbr1, sbr1,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 9, ccsb, fust, sbr2, isa, dfxa, scu0, scu1, idf, rsp, , , , , , , , 
RouterAgentPort, sbr1, 2
SyncRouter, sbr2, sbr2,2, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 5, 3, sbr1, xut, swf, , , , , , , , , , , , , , 
SyncRouter, sbra, sbra,0, 0, 0, 1, 4, 1, 0, 1, noa, dfxa, 2, 6, npsb, xpsb, ccsb, io_pxp, io_dmi, io_st, , , , , , , , , , , 
Endpoint, scu0,1, 1, 4, 0, 3, 3, 1, 3, 3, 3, 
Endpoint, scu1,3, 1, 4, 0, 3, 3, 1, 4, 3, 3, 
Endpoint, swf,2, 1, 5, 0, 3, 3, 1, 9, 3, 3, 
Endpoint, xpsb,0, 1, 1, 0, 1, 1, 1, 238, 3, 3, 
Endpoint, xut,2, 1, 5, 0, 3, 3, 1, 8, 3, 3, 
AsyncPort, ccsb, 0, 4, 4, 0, 
AsyncPort, sbr1, 1, 4, 4, 0, 
AsyncPort, sbr1, 2, 4, 4, 0, 
AsyncPort, sbra, 0, 2, 2, 0, 
AsyncPort, sbra, 1, 2, 2, 0, 
PowerWell, 0, 
PowerWell, 1, eva_present
PowerWell, 2, crp_sbr1_xu_en
PowerWell, 3, crp_sbr1_scu1_en
*/
//------------------------------------------------------------------------------
