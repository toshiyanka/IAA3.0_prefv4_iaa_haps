VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf156b040e2r2w0cbbehbaa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf156b040e2r2w0cbbehbaa4acw 0 0 ;
  SIZE 37.8 BY 46.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 23.64 13.628 24.84 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.444 23.64 17.488 24.84 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 20.76 13.628 21.96 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.612 20.76 17.656 21.96 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 23.64 15.428 24.84 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.644 23.64 15.688 24.84 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 23.64 15.856 24.84 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 23.64 16.116 24.84 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 23.64 16.416 24.84 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 23.64 17.228 24.84 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 23.64 14.316 24.84 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.64 14.616 24.84 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 23.64 19.028 24.84 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 23.64 19.288 24.84 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 23.64 19.716 24.84 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 23.64 20.016 24.84 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 23.64 20.828 24.84 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 23.64 21.088 24.84 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.612 23.64 17.656 24.84 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 23.64 18.216 24.84 ;
    END
  END rdaddrp1_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 0.36 13.628 1.56 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 30.6 15.128 31.8 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 30.6 15.216 31.8 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 30.6 21.516 31.8 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 30.6 21.728 31.8 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 31.56 13.888 32.76 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 31.56 13.972 32.76 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 31.56 20.528 32.76 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 31.56 20.616 32.76 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 32.52 15.128 33.72 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 32.52 15.216 33.72 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 2.28 21.428 3.48 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 32.52 21.516 33.72 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 32.52 21.728 33.72 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 33.48 13.888 34.68 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 33.48 13.972 34.68 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 33.48 20.528 34.68 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 33.48 20.616 34.68 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 34.44 15.128 35.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 34.44 15.216 35.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 34.44 21.516 35.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 34.44 21.728 35.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 2.28 21.516 3.48 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 35.4 13.888 36.6 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 35.4 13.972 36.6 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 35.4 20.528 36.6 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 35.4 20.616 36.6 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 36.36 15.128 37.56 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 36.36 15.216 37.56 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 36.36 21.516 37.56 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 36.36 21.728 37.56 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 37.32 13.888 38.52 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 37.32 13.972 38.52 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.24 13.716 4.44 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 37.32 20.528 38.52 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 37.32 20.616 38.52 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 38.28 15.128 39.48 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 38.28 15.216 39.48 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 38.28 21.516 39.48 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 38.28 21.728 39.48 ;
    END
  END rddatap0[135]
  PIN rddatap0[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 39.24 13.888 40.44 ;
    END
  END rddatap0[136]
  PIN rddatap0[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 39.24 13.972 40.44 ;
    END
  END rddatap0[137]
  PIN rddatap0[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 39.24 20.528 40.44 ;
    END
  END rddatap0[138]
  PIN rddatap0[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 39.24 20.616 40.44 ;
    END
  END rddatap0[139]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 3.24 13.888 4.44 ;
    END
  END rddatap0[13]
  PIN rddatap0[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 40.2 15.128 41.4 ;
    END
  END rddatap0[140]
  PIN rddatap0[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 40.2 15.216 41.4 ;
    END
  END rddatap0[141]
  PIN rddatap0[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 40.2 21.516 41.4 ;
    END
  END rddatap0[142]
  PIN rddatap0[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 40.2 21.728 41.4 ;
    END
  END rddatap0[143]
  PIN rddatap0[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 41.16 13.888 42.36 ;
    END
  END rddatap0[144]
  PIN rddatap0[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 41.16 13.972 42.36 ;
    END
  END rddatap0[145]
  PIN rddatap0[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 41.16 20.528 42.36 ;
    END
  END rddatap0[146]
  PIN rddatap0[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 41.16 20.616 42.36 ;
    END
  END rddatap0[147]
  PIN rddatap0[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 42.12 15.128 43.32 ;
    END
  END rddatap0[148]
  PIN rddatap0[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 42.12 15.216 43.32 ;
    END
  END rddatap0[149]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 3.24 20.272 4.44 ;
    END
  END rddatap0[14]
  PIN rddatap0[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 42.12 21.516 43.32 ;
    END
  END rddatap0[150]
  PIN rddatap0[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 42.12 21.728 43.32 ;
    END
  END rddatap0[151]
  PIN rddatap0[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 43.08 13.888 44.28 ;
    END
  END rddatap0[152]
  PIN rddatap0[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 43.08 13.972 44.28 ;
    END
  END rddatap0[153]
  PIN rddatap0[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 43.08 20.528 44.28 ;
    END
  END rddatap0[154]
  PIN rddatap0[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 43.08 20.616 44.28 ;
    END
  END rddatap0[155]
  PIN rddatap0[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 44.04 15.128 45.24 ;
    END
  END rddatap0[156]
  PIN rddatap0[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 44.04 15.216 45.24 ;
    END
  END rddatap0[157]
  PIN rddatap0[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 44.04 21.516 45.24 ;
    END
  END rddatap0[158]
  PIN rddatap0[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 44.04 21.728 45.24 ;
    END
  END rddatap0[159]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 3.24 20.356 4.44 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 4.2 14.956 5.4 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 4.2 15.128 5.4 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 4.2 21.428 5.4 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 4.2 21.516 5.4 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.36 13.716 1.56 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 5.16 13.716 6.36 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 5.16 13.888 6.36 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 5.16 20.272 6.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 5.16 20.356 6.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 6.12 14.956 7.32 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 6.12 15.128 7.32 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 6.12 21.428 7.32 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 6.12 21.516 7.32 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 7.08 13.716 8.28 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 7.08 13.888 8.28 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 0.36 21.428 1.56 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 7.08 20.272 8.28 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 7.08 20.356 8.28 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 8.04 14.956 9.24 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 8.04 15.128 9.24 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 8.04 21.428 9.24 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 8.04 21.516 9.24 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 9 13.716 10.2 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 9 13.888 10.2 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 9 20.272 10.2 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 9 20.356 10.2 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 0.36 21.516 1.56 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 9.96 14.956 11.16 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 9.96 15.128 11.16 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 9.96 21.428 11.16 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 9.96 21.516 11.16 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 10.92 13.716 12.12 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 10.92 13.888 12.12 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 10.92 20.272 12.12 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 10.92 20.356 12.12 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 11.88 14.956 13.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 11.88 15.128 13.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 1.32 14.228 2.52 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 11.88 21.428 13.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 11.88 21.516 13.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 12.84 13.716 14.04 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 12.84 13.888 14.04 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 12.84 20.272 14.04 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 12.84 20.356 14.04 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 13.8 14.956 15 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 13.8 15.128 15 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 13.8 21.428 15 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 13.8 21.516 15 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 1.32 14.316 2.52 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 14.76 13.716 15.96 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 14.76 13.888 15.96 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 14.76 20.272 15.96 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 14.76 20.356 15.96 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 15.72 14.956 16.92 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 15.72 15.128 16.92 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 15.72 21.428 16.92 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 15.72 21.516 16.92 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 16.68 13.716 17.88 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 16.68 13.888 17.88 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 1.32 20.272 2.52 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 16.68 20.272 17.88 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 16.68 20.356 17.88 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 17.64 14.956 18.84 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 17.64 15.128 18.84 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.384 17.64 21.428 18.84 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 17.64 21.516 18.84 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 18.6 13.716 19.8 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 18.6 13.888 19.8 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.228 18.6 20.272 19.8 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 18.6 20.356 19.8 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.312 1.32 20.356 2.52 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 25.8 13.888 27 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 25.8 13.972 27 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 25.8 20.528 27 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 25.8 20.616 27 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 26.76 15.128 27.96 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 26.76 15.216 27.96 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 26.76 21.516 27.96 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 26.76 21.728 27.96 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 27.72 13.888 28.92 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 27.72 13.972 28.92 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.912 2.28 14.956 3.48 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 27.72 20.528 28.92 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 27.72 20.616 28.92 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 28.68 15.128 29.88 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 28.68 15.216 29.88 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 28.68 21.516 29.88 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 28.68 21.728 29.88 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 29.64 13.888 30.84 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 29.64 13.972 30.84 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 29.64 20.528 30.84 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 29.64 20.616 30.84 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 2.28 15.128 3.48 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 0.36 13.888 1.56 ;
    END
  END rddatap1[0]
  PIN rddatap1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 30.6 15.428 31.8 ;
    END
  END rddatap1[100]
  PIN rddatap1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 30.6 15.516 31.8 ;
    END
  END rddatap1[101]
  PIN rddatap1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 30.6 21.816 31.8 ;
    END
  END rddatap1[102]
  PIN rddatap1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 30.6 20.016 31.8 ;
    END
  END rddatap1[103]
  PIN rddatap1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 31.56 14.056 32.76 ;
    END
  END rddatap1[104]
  PIN rddatap1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 31.56 14.228 32.76 ;
    END
  END rddatap1[105]
  PIN rddatap1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 31.56 20.828 32.76 ;
    END
  END rddatap1[106]
  PIN rddatap1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 31.56 20.916 32.76 ;
    END
  END rddatap1[107]
  PIN rddatap1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 32.52 15.428 33.72 ;
    END
  END rddatap1[108]
  PIN rddatap1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 32.52 15.516 33.72 ;
    END
  END rddatap1[109]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 2.28 21.728 3.48 ;
    END
  END rddatap1[10]
  PIN rddatap1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 32.52 21.816 33.72 ;
    END
  END rddatap1[110]
  PIN rddatap1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 32.52 20.016 33.72 ;
    END
  END rddatap1[111]
  PIN rddatap1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 33.48 14.056 34.68 ;
    END
  END rddatap1[112]
  PIN rddatap1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 33.48 14.228 34.68 ;
    END
  END rddatap1[113]
  PIN rddatap1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 33.48 20.828 34.68 ;
    END
  END rddatap1[114]
  PIN rddatap1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 33.48 20.916 34.68 ;
    END
  END rddatap1[115]
  PIN rddatap1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 34.44 15.428 35.64 ;
    END
  END rddatap1[116]
  PIN rddatap1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 34.44 15.516 35.64 ;
    END
  END rddatap1[117]
  PIN rddatap1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 34.44 21.816 35.64 ;
    END
  END rddatap1[118]
  PIN rddatap1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 34.44 20.016 35.64 ;
    END
  END rddatap1[119]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 2.28 21.816 3.48 ;
    END
  END rddatap1[11]
  PIN rddatap1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 35.4 14.056 36.6 ;
    END
  END rddatap1[120]
  PIN rddatap1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 35.4 14.228 36.6 ;
    END
  END rddatap1[121]
  PIN rddatap1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 35.4 20.828 36.6 ;
    END
  END rddatap1[122]
  PIN rddatap1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 35.4 20.916 36.6 ;
    END
  END rddatap1[123]
  PIN rddatap1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 36.36 15.428 37.56 ;
    END
  END rddatap1[124]
  PIN rddatap1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 36.36 15.516 37.56 ;
    END
  END rddatap1[125]
  PIN rddatap1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 36.36 21.816 37.56 ;
    END
  END rddatap1[126]
  PIN rddatap1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 36.36 20.016 37.56 ;
    END
  END rddatap1[127]
  PIN rddatap1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 37.32 14.056 38.52 ;
    END
  END rddatap1[128]
  PIN rddatap1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 37.32 14.228 38.52 ;
    END
  END rddatap1[129]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.24 13.972 4.44 ;
    END
  END rddatap1[12]
  PIN rddatap1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 37.32 20.828 38.52 ;
    END
  END rddatap1[130]
  PIN rddatap1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 37.32 20.916 38.52 ;
    END
  END rddatap1[131]
  PIN rddatap1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 38.28 15.428 39.48 ;
    END
  END rddatap1[132]
  PIN rddatap1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 38.28 15.516 39.48 ;
    END
  END rddatap1[133]
  PIN rddatap1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 38.28 21.816 39.48 ;
    END
  END rddatap1[134]
  PIN rddatap1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 38.28 20.016 39.48 ;
    END
  END rddatap1[135]
  PIN rddatap1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 39.24 14.056 40.44 ;
    END
  END rddatap1[136]
  PIN rddatap1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 39.24 14.228 40.44 ;
    END
  END rddatap1[137]
  PIN rddatap1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 39.24 20.828 40.44 ;
    END
  END rddatap1[138]
  PIN rddatap1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 39.24 20.916 40.44 ;
    END
  END rddatap1[139]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 3.24 14.056 4.44 ;
    END
  END rddatap1[13]
  PIN rddatap1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 40.2 15.428 41.4 ;
    END
  END rddatap1[140]
  PIN rddatap1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 40.2 15.516 41.4 ;
    END
  END rddatap1[141]
  PIN rddatap1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 40.2 21.816 41.4 ;
    END
  END rddatap1[142]
  PIN rddatap1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 40.2 20.016 41.4 ;
    END
  END rddatap1[143]
  PIN rddatap1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 41.16 14.056 42.36 ;
    END
  END rddatap1[144]
  PIN rddatap1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 41.16 14.228 42.36 ;
    END
  END rddatap1[145]
  PIN rddatap1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 41.16 20.828 42.36 ;
    END
  END rddatap1[146]
  PIN rddatap1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 41.16 20.916 42.36 ;
    END
  END rddatap1[147]
  PIN rddatap1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 42.12 15.428 43.32 ;
    END
  END rddatap1[148]
  PIN rddatap1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 42.12 15.516 43.32 ;
    END
  END rddatap1[149]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 3.24 20.528 4.44 ;
    END
  END rddatap1[14]
  PIN rddatap1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 42.12 21.816 43.32 ;
    END
  END rddatap1[150]
  PIN rddatap1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 42.12 20.016 43.32 ;
    END
  END rddatap1[151]
  PIN rddatap1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 43.08 14.056 44.28 ;
    END
  END rddatap1[152]
  PIN rddatap1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 43.08 14.228 44.28 ;
    END
  END rddatap1[153]
  PIN rddatap1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 43.08 20.828 44.28 ;
    END
  END rddatap1[154]
  PIN rddatap1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 43.08 20.916 44.28 ;
    END
  END rddatap1[155]
  PIN rddatap1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 44.04 15.428 45.24 ;
    END
  END rddatap1[156]
  PIN rddatap1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 44.04 15.516 45.24 ;
    END
  END rddatap1[157]
  PIN rddatap1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 44.04 21.816 45.24 ;
    END
  END rddatap1[158]
  PIN rddatap1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 44.04 20.016 45.24 ;
    END
  END rddatap1[159]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 3.24 20.616 4.44 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 4.2 15.216 5.4 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.2 15.428 5.4 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 4.2 21.728 5.4 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 4.2 21.816 5.4 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.36 13.972 1.56 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 5.16 13.972 6.36 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 5.16 14.056 6.36 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 5.16 20.528 6.36 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 5.16 20.616 6.36 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 6.12 15.216 7.32 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6.12 15.428 7.32 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 6.12 21.728 7.32 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 6.12 21.816 7.32 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 7.08 13.972 8.28 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 7.08 14.056 8.28 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 0.36 21.728 1.56 ;
    END
  END rddatap1[2]
  PIN rddatap1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 7.08 20.528 8.28 ;
    END
  END rddatap1[30]
  PIN rddatap1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 7.08 20.616 8.28 ;
    END
  END rddatap1[31]
  PIN rddatap1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 8.04 15.216 9.24 ;
    END
  END rddatap1[32]
  PIN rddatap1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.04 15.428 9.24 ;
    END
  END rddatap1[33]
  PIN rddatap1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 8.04 21.728 9.24 ;
    END
  END rddatap1[34]
  PIN rddatap1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 8.04 21.816 9.24 ;
    END
  END rddatap1[35]
  PIN rddatap1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 9 13.972 10.2 ;
    END
  END rddatap1[36]
  PIN rddatap1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 9 14.056 10.2 ;
    END
  END rddatap1[37]
  PIN rddatap1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 9 20.528 10.2 ;
    END
  END rddatap1[38]
  PIN rddatap1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 9 20.616 10.2 ;
    END
  END rddatap1[39]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 0.36 21.816 1.56 ;
    END
  END rddatap1[3]
  PIN rddatap1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 9.96 15.216 11.16 ;
    END
  END rddatap1[40]
  PIN rddatap1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 9.96 15.428 11.16 ;
    END
  END rddatap1[41]
  PIN rddatap1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 9.96 21.728 11.16 ;
    END
  END rddatap1[42]
  PIN rddatap1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 9.96 21.816 11.16 ;
    END
  END rddatap1[43]
  PIN rddatap1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 10.92 13.972 12.12 ;
    END
  END rddatap1[44]
  PIN rddatap1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 10.92 14.056 12.12 ;
    END
  END rddatap1[45]
  PIN rddatap1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 10.92 20.528 12.12 ;
    END
  END rddatap1[46]
  PIN rddatap1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 10.92 20.616 12.12 ;
    END
  END rddatap1[47]
  PIN rddatap1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 11.88 15.216 13.08 ;
    END
  END rddatap1[48]
  PIN rddatap1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 11.88 15.428 13.08 ;
    END
  END rddatap1[49]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 1.32 14.528 2.52 ;
    END
  END rddatap1[4]
  PIN rddatap1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 11.88 21.728 13.08 ;
    END
  END rddatap1[50]
  PIN rddatap1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 11.88 21.816 13.08 ;
    END
  END rddatap1[51]
  PIN rddatap1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 12.84 13.972 14.04 ;
    END
  END rddatap1[52]
  PIN rddatap1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 12.84 14.056 14.04 ;
    END
  END rddatap1[53]
  PIN rddatap1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 12.84 20.528 14.04 ;
    END
  END rddatap1[54]
  PIN rddatap1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 12.84 20.616 14.04 ;
    END
  END rddatap1[55]
  PIN rddatap1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 13.8 15.216 15 ;
    END
  END rddatap1[56]
  PIN rddatap1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 13.8 15.428 15 ;
    END
  END rddatap1[57]
  PIN rddatap1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 13.8 21.728 15 ;
    END
  END rddatap1[58]
  PIN rddatap1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 13.8 21.816 15 ;
    END
  END rddatap1[59]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 1.32 14.616 2.52 ;
    END
  END rddatap1[5]
  PIN rddatap1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 14.76 13.972 15.96 ;
    END
  END rddatap1[60]
  PIN rddatap1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 14.76 14.056 15.96 ;
    END
  END rddatap1[61]
  PIN rddatap1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 14.76 20.528 15.96 ;
    END
  END rddatap1[62]
  PIN rddatap1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 14.76 20.616 15.96 ;
    END
  END rddatap1[63]
  PIN rddatap1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 15.72 15.216 16.92 ;
    END
  END rddatap1[64]
  PIN rddatap1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 15.72 15.428 16.92 ;
    END
  END rddatap1[65]
  PIN rddatap1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 15.72 21.728 16.92 ;
    END
  END rddatap1[66]
  PIN rddatap1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 15.72 21.816 16.92 ;
    END
  END rddatap1[67]
  PIN rddatap1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 16.68 13.972 17.88 ;
    END
  END rddatap1[68]
  PIN rddatap1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 16.68 14.056 17.88 ;
    END
  END rddatap1[69]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 1.32 20.528 2.52 ;
    END
  END rddatap1[6]
  PIN rddatap1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 16.68 20.528 17.88 ;
    END
  END rddatap1[70]
  PIN rddatap1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 16.68 20.616 17.88 ;
    END
  END rddatap1[71]
  PIN rddatap1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 17.64 15.216 18.84 ;
    END
  END rddatap1[72]
  PIN rddatap1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 17.64 15.428 18.84 ;
    END
  END rddatap1[73]
  PIN rddatap1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.684 17.64 21.728 18.84 ;
    END
  END rddatap1[74]
  PIN rddatap1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 17.64 21.816 18.84 ;
    END
  END rddatap1[75]
  PIN rddatap1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 18.6 13.972 19.8 ;
    END
  END rddatap1[76]
  PIN rddatap1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 18.6 14.056 19.8 ;
    END
  END rddatap1[77]
  PIN rddatap1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.484 18.6 20.528 19.8 ;
    END
  END rddatap1[78]
  PIN rddatap1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 18.6 20.616 19.8 ;
    END
  END rddatap1[79]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.572 1.32 20.616 2.52 ;
    END
  END rddatap1[7]
  PIN rddatap1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 25.8 14.056 27 ;
    END
  END rddatap1[80]
  PIN rddatap1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 25.8 14.228 27 ;
    END
  END rddatap1[81]
  PIN rddatap1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 25.8 20.916 27 ;
    END
  END rddatap1[82]
  PIN rddatap1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.128 25.8 21.172 27 ;
    END
  END rddatap1[83]
  PIN rddatap1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 26.76 15.428 27.96 ;
    END
  END rddatap1[84]
  PIN rddatap1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 26.76 15.516 27.96 ;
    END
  END rddatap1[85]
  PIN rddatap1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 26.76 21.816 27.96 ;
    END
  END rddatap1[86]
  PIN rddatap1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 26.76 20.016 27.96 ;
    END
  END rddatap1[87]
  PIN rddatap1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 27.72 14.056 28.92 ;
    END
  END rddatap1[88]
  PIN rddatap1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 27.72 14.228 28.92 ;
    END
  END rddatap1[89]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 2.28 15.216 3.48 ;
    END
  END rddatap1[8]
  PIN rddatap1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 27.72 20.828 28.92 ;
    END
  END rddatap1[90]
  PIN rddatap1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 27.72 20.916 28.92 ;
    END
  END rddatap1[91]
  PIN rddatap1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 28.68 15.428 29.88 ;
    END
  END rddatap1[92]
  PIN rddatap1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 28.68 15.516 29.88 ;
    END
  END rddatap1[93]
  PIN rddatap1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.772 28.68 21.816 29.88 ;
    END
  END rddatap1[94]
  PIN rddatap1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 28.68 20.016 29.88 ;
    END
  END rddatap1[95]
  PIN rddatap1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 29.64 14.056 30.84 ;
    END
  END rddatap1[96]
  PIN rddatap1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 29.64 14.228 30.84 ;
    END
  END rddatap1[97]
  PIN rddatap1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 29.64 20.828 30.84 ;
    END
  END rddatap1[98]
  PIN rddatap1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.872 29.64 20.916 30.84 ;
    END
  END rddatap1[99]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 2.28 15.428 3.48 ;
    END
  END rddatap1[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 23.64 14.872 24.84 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 23.64 18.472 24.84 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 23.64 15.128 24.84 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 23.64 18.728 24.84 ;
    END
  END sdl_initp1
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 36.862 0.06 36.938 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.062 0.06 35.138 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 33.262 0.06 33.338 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.462 0.06 31.538 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.662 0.06 29.738 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 27.862 0.06 27.938 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.062 0.06 26.138 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.262 0.06 24.338 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 22.462 0.06 22.538 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.662 0.06 20.738 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.862 0.06 18.938 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.062 0.06 17.138 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.262 0.06 15.338 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 46.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 35.962 0.06 36.038 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 34.162 0.06 34.238 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 32.362 0.06 32.438 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.562 0.06 30.638 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 28.762 0.06 28.838 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.962 0.06 27.038 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.162 0.06 25.238 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.362 0.06 23.438 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 21.562 0.06 21.638 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 19.762 0.06 19.838 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.962 0.06 18.038 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 16.162 0.06 16.238 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.362 0.06 14.438 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 46.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 46.02 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.644 20.76 15.688 21.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 20.76 15.856 21.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 20.76 16.116 21.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 20.76 16.416 21.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 20.76 17.228 21.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.444 20.76 17.488 21.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 20.76 14.316 21.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 20.76 14.616 21.96 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.672 20.76 19.716 21.96 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.972 20.76 20.016 21.96 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 20.784 20.76 20.828 21.96 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.044 20.76 21.088 21.96 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.212 20.76 21.256 21.96 ;
    END
  END wraddrp1[4]
  PIN wraddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 21.472 20.76 21.516 21.96 ;
    END
  END wraddrp1[5]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 20.76 18.216 21.96 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 20.76 18.472 21.96 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 0.36 16.116 1.56 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 30.6 15.772 31.8 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 30.6 15.856 31.8 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 30.6 18.816 31.8 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 30.6 19.028 31.8 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 31.56 16.928 32.76 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 31.56 17.016 32.76 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 31.56 19.628 32.76 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 31.56 17.916 32.76 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 32.52 15.772 33.72 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 32.52 15.856 33.72 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 2.28 18.556 3.48 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 32.52 18.816 33.72 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 32.52 19.028 33.72 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 33.48 16.928 34.68 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 33.48 17.016 34.68 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 33.48 19.628 34.68 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 33.48 17.916 34.68 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 34.44 15.772 35.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 34.44 15.856 35.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 34.44 18.816 35.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 34.44 19.028 35.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 2.28 18.728 3.48 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 35.4 16.928 36.6 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 35.4 17.016 36.6 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 35.4 19.628 36.6 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 35.4 17.916 36.6 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 36.36 15.772 37.56 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 36.36 15.856 37.56 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 36.36 18.816 37.56 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 36.36 19.028 37.56 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 37.32 16.928 38.52 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 37.32 17.016 38.52 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 3.24 16.672 4.44 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 37.32 19.628 38.52 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 37.32 17.916 38.52 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 38.28 15.772 39.48 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 38.28 15.856 39.48 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 38.28 18.816 39.48 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 38.28 19.028 39.48 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 39.24 16.928 40.44 ;
    END
  END wrdatap0[136]
  PIN wrdatap0[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 39.24 17.016 40.44 ;
    END
  END wrdatap0[137]
  PIN wrdatap0[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 39.24 19.628 40.44 ;
    END
  END wrdatap0[138]
  PIN wrdatap0[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 39.24 17.916 40.44 ;
    END
  END wrdatap0[139]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 3.24 16.756 4.44 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 40.2 15.772 41.4 ;
    END
  END wrdatap0[140]
  PIN wrdatap0[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 40.2 15.856 41.4 ;
    END
  END wrdatap0[141]
  PIN wrdatap0[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 40.2 18.816 41.4 ;
    END
  END wrdatap0[142]
  PIN wrdatap0[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 40.2 19.028 41.4 ;
    END
  END wrdatap0[143]
  PIN wrdatap0[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 41.16 16.928 42.36 ;
    END
  END wrdatap0[144]
  PIN wrdatap0[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 41.16 17.016 42.36 ;
    END
  END wrdatap0[145]
  PIN wrdatap0[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 41.16 19.628 42.36 ;
    END
  END wrdatap0[146]
  PIN wrdatap0[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 41.16 17.916 42.36 ;
    END
  END wrdatap0[147]
  PIN wrdatap0[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 42.12 15.772 43.32 ;
    END
  END wrdatap0[148]
  PIN wrdatap0[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 42.12 15.856 43.32 ;
    END
  END wrdatap0[149]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 3.24 19.456 4.44 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 42.12 18.816 43.32 ;
    END
  END wrdatap0[150]
  PIN wrdatap0[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 42.12 19.028 43.32 ;
    END
  END wrdatap0[151]
  PIN wrdatap0[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 43.08 16.928 44.28 ;
    END
  END wrdatap0[152]
  PIN wrdatap0[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 43.08 17.016 44.28 ;
    END
  END wrdatap0[153]
  PIN wrdatap0[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 43.08 19.628 44.28 ;
    END
  END wrdatap0[154]
  PIN wrdatap0[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 43.08 17.916 44.28 ;
    END
  END wrdatap0[155]
  PIN wrdatap0[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 44.04 15.772 45.24 ;
    END
  END wrdatap0[156]
  PIN wrdatap0[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 44.04 15.856 45.24 ;
    END
  END wrdatap0[157]
  PIN wrdatap0[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 44.04 18.816 45.24 ;
    END
  END wrdatap0[158]
  PIN wrdatap0[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 44.04 19.028 45.24 ;
    END
  END wrdatap0[159]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 3.24 19.628 4.44 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 4.2 17.572 5.4 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 4.2 15.772 5.4 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 4.2 18.556 5.4 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 4.2 18.728 5.4 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 0.36 16.328 1.56 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 5.16 16.672 6.36 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 5.16 16.756 6.36 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 5.16 19.456 6.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 5.16 19.628 6.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 6.12 17.572 7.32 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 6.12 15.772 7.32 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 6.12 18.556 7.32 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 6.12 18.728 7.32 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 7.08 16.672 8.28 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 7.08 16.756 8.28 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.36 18.816 1.56 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 7.08 19.456 8.28 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 7.08 19.628 8.28 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 8.04 17.572 9.24 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 8.04 15.772 9.24 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 8.04 18.556 9.24 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 8.04 18.728 9.24 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 9 16.672 10.2 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 9 16.756 10.2 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 9 19.456 10.2 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 9 19.628 10.2 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.36 19.028 1.56 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 9.96 17.572 11.16 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 9.96 15.772 11.16 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 9.96 18.556 11.16 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 9.96 18.728 11.16 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 10.92 16.672 12.12 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 10.92 16.756 12.12 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 10.92 19.456 12.12 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 10.92 19.628 12.12 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 11.88 17.572 13.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 11.88 15.772 13.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 1.32 16.756 2.52 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 11.88 18.556 13.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 11.88 18.728 13.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 12.84 16.672 14.04 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 12.84 16.756 14.04 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 12.84 19.456 14.04 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 12.84 19.628 14.04 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 13.8 17.572 15 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 13.8 15.772 15 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 13.8 18.556 15 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 13.8 18.728 15 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 1.32 16.928 2.52 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 14.76 16.672 15.96 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 14.76 16.756 15.96 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 14.76 19.456 15.96 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 14.76 19.628 15.96 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 15.72 17.572 16.92 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 15.72 15.772 16.92 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 15.72 18.556 16.92 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 15.72 18.728 16.92 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 16.68 16.672 17.88 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 16.68 16.756 17.88 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 1.32 19.456 2.52 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 16.68 19.456 17.88 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 16.68 19.628 17.88 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 17.64 17.572 18.84 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 17.64 15.772 18.84 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.512 17.64 18.556 18.84 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 17.64 18.728 18.84 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 18.6 16.672 19.8 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 18.6 16.756 19.8 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.412 18.6 19.456 19.8 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 18.6 19.628 19.8 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 1.32 19.628 2.52 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.712 25.8 16.756 27 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 25.8 16.928 27 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 25.8 19.628 27 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 25.8 17.916 27 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 26.76 15.772 27.96 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 26.76 15.856 27.96 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.76 18.816 27.96 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.76 19.028 27.96 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 27.72 16.928 28.92 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 27.72 17.016 28.92 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 2.28 17.572 3.48 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 27.72 19.628 28.92 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 27.72 17.916 28.92 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 28.68 15.772 29.88 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 28.68 15.856 29.88 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 28.68 18.816 29.88 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 28.68 19.028 29.88 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 29.64 16.928 30.84 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 29.64 17.016 30.84 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.584 29.64 19.628 30.84 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 29.64 17.916 30.84 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 2.28 15.772 3.48 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 20.76 15.128 21.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 20.76 15.428 21.96 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 0.36 16.416 1.56 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 30.6 16.028 31.8 ;
    END
  END wrdatap1[100]
  PIN wrdatap1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 30.6 16.116 31.8 ;
    END
  END wrdatap1[101]
  PIN wrdatap1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 30.6 19.116 31.8 ;
    END
  END wrdatap1[102]
  PIN wrdatap1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 30.6 19.288 31.8 ;
    END
  END wrdatap1[103]
  PIN wrdatap1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 31.56 17.228 32.76 ;
    END
  END wrdatap1[104]
  PIN wrdatap1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 31.56 17.316 32.76 ;
    END
  END wrdatap1[105]
  PIN wrdatap1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 31.56 18.128 32.76 ;
    END
  END wrdatap1[106]
  PIN wrdatap1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 31.56 18.216 32.76 ;
    END
  END wrdatap1[107]
  PIN wrdatap1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 32.52 16.028 33.72 ;
    END
  END wrdatap1[108]
  PIN wrdatap1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 32.52 16.116 33.72 ;
    END
  END wrdatap1[109]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 2.28 18.816 3.48 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 32.52 19.116 33.72 ;
    END
  END wrdatap1[110]
  PIN wrdatap1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 32.52 19.288 33.72 ;
    END
  END wrdatap1[111]
  PIN wrdatap1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 33.48 17.228 34.68 ;
    END
  END wrdatap1[112]
  PIN wrdatap1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 33.48 17.316 34.68 ;
    END
  END wrdatap1[113]
  PIN wrdatap1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 33.48 18.128 34.68 ;
    END
  END wrdatap1[114]
  PIN wrdatap1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 33.48 18.216 34.68 ;
    END
  END wrdatap1[115]
  PIN wrdatap1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 34.44 16.028 35.64 ;
    END
  END wrdatap1[116]
  PIN wrdatap1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 34.44 16.116 35.64 ;
    END
  END wrdatap1[117]
  PIN wrdatap1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 34.44 19.116 35.64 ;
    END
  END wrdatap1[118]
  PIN wrdatap1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 34.44 19.288 35.64 ;
    END
  END wrdatap1[119]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 2.28 19.028 3.48 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 35.4 17.228 36.6 ;
    END
  END wrdatap1[120]
  PIN wrdatap1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 35.4 17.316 36.6 ;
    END
  END wrdatap1[121]
  PIN wrdatap1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 35.4 18.128 36.6 ;
    END
  END wrdatap1[122]
  PIN wrdatap1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 35.4 18.216 36.6 ;
    END
  END wrdatap1[123]
  PIN wrdatap1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 36.36 16.028 37.56 ;
    END
  END wrdatap1[124]
  PIN wrdatap1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 36.36 16.116 37.56 ;
    END
  END wrdatap1[125]
  PIN wrdatap1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 36.36 19.116 37.56 ;
    END
  END wrdatap1[126]
  PIN wrdatap1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 36.36 19.288 37.56 ;
    END
  END wrdatap1[127]
  PIN wrdatap1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 37.32 17.228 38.52 ;
    END
  END wrdatap1[128]
  PIN wrdatap1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 37.32 17.316 38.52 ;
    END
  END wrdatap1[129]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 3.24 16.928 4.44 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 37.32 18.128 38.52 ;
    END
  END wrdatap1[130]
  PIN wrdatap1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 37.32 18.216 38.52 ;
    END
  END wrdatap1[131]
  PIN wrdatap1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 38.28 16.028 39.48 ;
    END
  END wrdatap1[132]
  PIN wrdatap1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 38.28 16.116 39.48 ;
    END
  END wrdatap1[133]
  PIN wrdatap1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 38.28 19.116 39.48 ;
    END
  END wrdatap1[134]
  PIN wrdatap1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 38.28 19.288 39.48 ;
    END
  END wrdatap1[135]
  PIN wrdatap1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 39.24 17.228 40.44 ;
    END
  END wrdatap1[136]
  PIN wrdatap1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 39.24 17.316 40.44 ;
    END
  END wrdatap1[137]
  PIN wrdatap1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 39.24 18.128 40.44 ;
    END
  END wrdatap1[138]
  PIN wrdatap1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 39.24 18.216 40.44 ;
    END
  END wrdatap1[139]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 3.24 17.016 4.44 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 40.2 16.028 41.4 ;
    END
  END wrdatap1[140]
  PIN wrdatap1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 40.2 16.116 41.4 ;
    END
  END wrdatap1[141]
  PIN wrdatap1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 40.2 19.116 41.4 ;
    END
  END wrdatap1[142]
  PIN wrdatap1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 40.2 19.288 41.4 ;
    END
  END wrdatap1[143]
  PIN wrdatap1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 41.16 17.228 42.36 ;
    END
  END wrdatap1[144]
  PIN wrdatap1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 41.16 17.316 42.36 ;
    END
  END wrdatap1[145]
  PIN wrdatap1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 41.16 18.128 42.36 ;
    END
  END wrdatap1[146]
  PIN wrdatap1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 41.16 18.216 42.36 ;
    END
  END wrdatap1[147]
  PIN wrdatap1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 42.12 16.028 43.32 ;
    END
  END wrdatap1[148]
  PIN wrdatap1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 42.12 16.116 43.32 ;
    END
  END wrdatap1[149]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 3.24 17.916 4.44 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 42.12 19.116 43.32 ;
    END
  END wrdatap1[150]
  PIN wrdatap1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 42.12 19.288 43.32 ;
    END
  END wrdatap1[151]
  PIN wrdatap1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 43.08 17.228 44.28 ;
    END
  END wrdatap1[152]
  PIN wrdatap1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 43.08 17.316 44.28 ;
    END
  END wrdatap1[153]
  PIN wrdatap1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 43.08 18.128 44.28 ;
    END
  END wrdatap1[154]
  PIN wrdatap1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 43.08 18.216 44.28 ;
    END
  END wrdatap1[155]
  PIN wrdatap1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 44.04 16.028 45.24 ;
    END
  END wrdatap1[156]
  PIN wrdatap1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 44.04 16.116 45.24 ;
    END
  END wrdatap1[157]
  PIN wrdatap1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 44.04 19.116 45.24 ;
    END
  END wrdatap1[158]
  PIN wrdatap1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 44.04 19.288 45.24 ;
    END
  END wrdatap1[159]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 3.24 18.128 4.44 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 4.2 15.856 5.4 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 4.2 16.028 5.4 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 4.2 18.816 5.4 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 4.2 19.028 5.4 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.544 0.36 16.588 1.56 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 5.16 16.928 6.36 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 5.16 17.016 6.36 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 5.16 17.916 6.36 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 5.16 18.128 6.36 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 6.12 15.856 7.32 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 6.12 16.028 7.32 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 6.12 18.816 7.32 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 6.12 19.028 7.32 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 7.08 16.928 8.28 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 7.08 17.016 8.28 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 0.36 19.116 1.56 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 7.08 17.916 8.28 ;
    END
  END wrdatap1[30]
  PIN wrdatap1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 7.08 18.128 8.28 ;
    END
  END wrdatap1[31]
  PIN wrdatap1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 8.04 15.856 9.24 ;
    END
  END wrdatap1[32]
  PIN wrdatap1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 8.04 16.028 9.24 ;
    END
  END wrdatap1[33]
  PIN wrdatap1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.04 18.816 9.24 ;
    END
  END wrdatap1[34]
  PIN wrdatap1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.04 19.028 9.24 ;
    END
  END wrdatap1[35]
  PIN wrdatap1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 9 16.928 10.2 ;
    END
  END wrdatap1[36]
  PIN wrdatap1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 9 17.016 10.2 ;
    END
  END wrdatap1[37]
  PIN wrdatap1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 9 17.916 10.2 ;
    END
  END wrdatap1[38]
  PIN wrdatap1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 9 18.128 10.2 ;
    END
  END wrdatap1[39]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 0.36 19.288 1.56 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 9.96 15.856 11.16 ;
    END
  END wrdatap1[40]
  PIN wrdatap1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 9.96 16.028 11.16 ;
    END
  END wrdatap1[41]
  PIN wrdatap1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 9.96 18.816 11.16 ;
    END
  END wrdatap1[42]
  PIN wrdatap1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 9.96 19.028 11.16 ;
    END
  END wrdatap1[43]
  PIN wrdatap1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 10.92 16.928 12.12 ;
    END
  END wrdatap1[44]
  PIN wrdatap1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 10.92 17.016 12.12 ;
    END
  END wrdatap1[45]
  PIN wrdatap1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 10.92 17.916 12.12 ;
    END
  END wrdatap1[46]
  PIN wrdatap1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 10.92 18.128 12.12 ;
    END
  END wrdatap1[47]
  PIN wrdatap1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 11.88 15.856 13.08 ;
    END
  END wrdatap1[48]
  PIN wrdatap1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 11.88 16.028 13.08 ;
    END
  END wrdatap1[49]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 1.32 17.016 2.52 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 11.88 18.816 13.08 ;
    END
  END wrdatap1[50]
  PIN wrdatap1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 11.88 19.028 13.08 ;
    END
  END wrdatap1[51]
  PIN wrdatap1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 12.84 16.928 14.04 ;
    END
  END wrdatap1[52]
  PIN wrdatap1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 12.84 17.016 14.04 ;
    END
  END wrdatap1[53]
  PIN wrdatap1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 12.84 17.916 14.04 ;
    END
  END wrdatap1[54]
  PIN wrdatap1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 12.84 18.128 14.04 ;
    END
  END wrdatap1[55]
  PIN wrdatap1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 13.8 15.856 15 ;
    END
  END wrdatap1[56]
  PIN wrdatap1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 13.8 16.028 15 ;
    END
  END wrdatap1[57]
  PIN wrdatap1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 13.8 18.816 15 ;
    END
  END wrdatap1[58]
  PIN wrdatap1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 13.8 19.028 15 ;
    END
  END wrdatap1[59]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 1.32 17.228 2.52 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 14.76 16.928 15.96 ;
    END
  END wrdatap1[60]
  PIN wrdatap1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 14.76 17.016 15.96 ;
    END
  END wrdatap1[61]
  PIN wrdatap1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 14.76 17.916 15.96 ;
    END
  END wrdatap1[62]
  PIN wrdatap1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 14.76 18.128 15.96 ;
    END
  END wrdatap1[63]
  PIN wrdatap1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 15.72 15.856 16.92 ;
    END
  END wrdatap1[64]
  PIN wrdatap1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 15.72 16.028 16.92 ;
    END
  END wrdatap1[65]
  PIN wrdatap1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 15.72 18.816 16.92 ;
    END
  END wrdatap1[66]
  PIN wrdatap1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 15.72 19.028 16.92 ;
    END
  END wrdatap1[67]
  PIN wrdatap1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 16.68 16.928 17.88 ;
    END
  END wrdatap1[68]
  PIN wrdatap1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 16.68 17.016 17.88 ;
    END
  END wrdatap1[69]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 1.32 17.916 2.52 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 16.68 17.916 17.88 ;
    END
  END wrdatap1[70]
  PIN wrdatap1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 16.68 18.128 17.88 ;
    END
  END wrdatap1[71]
  PIN wrdatap1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 17.64 15.856 18.84 ;
    END
  END wrdatap1[72]
  PIN wrdatap1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 17.64 16.028 18.84 ;
    END
  END wrdatap1[73]
  PIN wrdatap1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 17.64 18.816 18.84 ;
    END
  END wrdatap1[74]
  PIN wrdatap1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 17.64 19.028 18.84 ;
    END
  END wrdatap1[75]
  PIN wrdatap1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 18.6 16.928 19.8 ;
    END
  END wrdatap1[76]
  PIN wrdatap1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 18.6 17.016 19.8 ;
    END
  END wrdatap1[77]
  PIN wrdatap1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 18.6 17.916 19.8 ;
    END
  END wrdatap1[78]
  PIN wrdatap1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 18.6 18.128 19.8 ;
    END
  END wrdatap1[79]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 1.32 18.128 2.52 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 25.8 17.016 27 ;
    END
  END wrdatap1[80]
  PIN wrdatap1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 25.8 17.316 27 ;
    END
  END wrdatap1[81]
  PIN wrdatap1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 25.8 18.128 27 ;
    END
  END wrdatap1[82]
  PIN wrdatap1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.344 25.8 18.388 27 ;
    END
  END wrdatap1[83]
  PIN wrdatap1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 26.76 16.028 27.96 ;
    END
  END wrdatap1[84]
  PIN wrdatap1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 26.76 16.116 27.96 ;
    END
  END wrdatap1[85]
  PIN wrdatap1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 26.76 19.116 27.96 ;
    END
  END wrdatap1[86]
  PIN wrdatap1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 26.76 19.288 27.96 ;
    END
  END wrdatap1[87]
  PIN wrdatap1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 27.72 17.228 28.92 ;
    END
  END wrdatap1[88]
  PIN wrdatap1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 27.72 17.316 28.92 ;
    END
  END wrdatap1[89]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.812 2.28 15.856 3.48 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 27.72 18.128 28.92 ;
    END
  END wrdatap1[90]
  PIN wrdatap1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 27.72 18.216 28.92 ;
    END
  END wrdatap1[91]
  PIN wrdatap1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 28.68 16.028 29.88 ;
    END
  END wrdatap1[92]
  PIN wrdatap1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 28.68 16.116 29.88 ;
    END
  END wrdatap1[93]
  PIN wrdatap1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 28.68 19.116 29.88 ;
    END
  END wrdatap1[94]
  PIN wrdatap1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 28.68 19.288 29.88 ;
    END
  END wrdatap1[95]
  PIN wrdatap1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 29.64 17.228 30.84 ;
    END
  END wrdatap1[96]
  PIN wrdatap1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 29.64 17.316 30.84 ;
    END
  END wrdatap1[97]
  PIN wrdatap1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 29.64 18.128 30.84 ;
    END
  END wrdatap1[98]
  PIN wrdatap1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 29.64 18.216 30.84 ;
    END
  END wrdatap1[99]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 2.28 16.028 3.48 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 20.76 19.028 21.96 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.244 20.76 19.288 21.96 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 20.76 14.872 21.96 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 20.76 18.728 21.96 ;
    END
  END wrenp1
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 37.8 46.08 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 37.8 46.08 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 37.8705 46.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 37.835 46.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 37.87 46.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 37.859 46.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 37.89 46.142 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 37.892 46.14 ;
  END
END arf156b040e2r2w0cbbehbaa4acw
END LIBRARY
