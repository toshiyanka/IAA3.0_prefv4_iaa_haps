VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf132b192e1r1w0cbbehcaa4acw
  CLASS BLOCK ;
  FOREIGN arf132b192e1r1w0cbbehcaa4acw ;
  ORIGIN 0 0 ;
  SIZE 70.2 BY 29.76 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.372 16.68 34.416 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.728 14.76 33.772 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.272 16.68 35.316 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.728 16.68 33.772 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.984 16.68 34.028 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.072 16.68 34.116 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.284 16.68 34.328 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.372 18.6 34.416 19.8 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.628 18.6 34.672 19.8 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.884 18.6 34.928 19.8 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.628 16.68 34.672 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.884 16.68 34.928 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.972 16.68 35.016 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.184 16.68 35.228 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.884 14.76 34.928 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.972 14.76 35.016 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.184 14.76 35.228 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 35.272 14.76 35.316 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.728 12.84 33.772 14.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.984 12.84 34.028 14.04 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.072 12.84 34.116 14.04 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.284 12.84 34.328 14.04 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 33.984 14.76 34.028 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.072 14.76 34.116 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 22.56 12.728 23.76 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 22.56 12.816 23.76 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 22.56 47.916 23.76 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 22.56 48.172 23.76 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 23.28 14.228 24.48 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 23.28 14.316 24.48 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 23.28 44.572 24.48 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 23.28 44.828 24.48 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 24 10.716 25.2 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 24 10.928 25.2 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 1.68 48.816 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 24 46.716 25.2 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 24 46.928 25.2 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 24.72 12.816 25.92 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 24.72 13.072 25.92 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 24.72 48.172 25.92 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 24.72 48.428 25.92 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 25.44 14.316 26.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 25.44 14.528 26.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 25.44 44.828 26.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 25.44 44.916 26.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 1.68 49.072 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 26.16 11.016 27.36 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 26.16 11.272 27.36 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 26.16 46.928 27.36 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 26.16 47.016 27.36 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 26.88 13.072 28.08 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 26.88 13.328 28.08 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 26.88 48.428 28.08 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 26.88 48.516 28.08 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 27.6 14.528 28.8 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 27.6 14.616 28.8 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 2.4 10.372 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 27.6 44.916 28.8 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 27.6 45.128 28.8 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 28.32 11.528 29.52 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 28.32 11.616 29.52 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 28.32 47.016 29.52 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 28.32 47.272 29.52 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 2.4 10.628 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 2.4 46.028 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.072 2.4 46.116 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 3.12 12.516 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 3.12 12.728 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 3.12 47.828 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 3.12 47.916 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 3.84 13.972 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 3.84 14.228 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 3.84 44.572 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 3.84 44.828 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 4.56 10.716 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 4.56 10.928 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 4.56 46.716 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 4.56 46.928 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 5.28 12.816 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 5.28 13.072 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 0.24 45.216 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 5.28 48.172 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 5.28 48.428 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 6 14.316 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 6 14.528 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 6 44.828 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 6 44.916 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 6.72 11.016 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 6.72 11.272 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 6.72 46.928 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 6.72 47.016 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.428 0.24 45.472 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 7.44 13.072 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 7.44 13.328 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 7.44 48.428 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 7.44 48.516 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 8.16 14.528 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.16 14.616 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 8.16 44.916 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 8.16 45.128 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 8.88 11.528 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 8.88 11.616 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 0.96 12.172 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 8.88 47.016 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 8.88 47.272 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 9.6 13.328 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 9.6 13.416 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 9.6 48.516 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 9.6 48.728 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 10.32 14.616 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 10.32 10.028 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 10.32 45.128 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 10.32 45.216 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 0.96 12.428 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 11.04 11.828 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 11.04 11.916 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 11.04 47.272 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 11.04 47.528 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 11.76 13.416 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.76 13.628 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 11.76 48.728 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 11.76 48.816 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 12.48 10.116 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 12.48 10.372 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 0.96 47.528 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 12.48 45.728 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 12.48 45.816 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 13.2 12.428 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 13.2 12.516 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 13.2 47.616 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 13.2 47.828 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 18.24 11.272 19.44 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 18.24 11.528 19.44 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 18.24 46.628 19.44 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 18.24 46.716 19.44 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 0.96 47.616 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 18.96 13.416 20.16 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 18.96 13.628 20.16 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 18.96 48.728 20.16 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 18.96 48.816 20.16 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 19.68 10.116 20.88 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 19.68 10.372 20.88 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 19.68 45.728 20.88 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 19.68 45.816 20.88 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 20.4 12.428 21.6 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 20.4 12.516 21.6 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 1.68 13.628 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 20.4 47.616 21.6 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 20.4 47.828 21.6 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 21.12 13.716 22.32 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 21.12 13.972 22.32 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 21.12 49.072 22.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 21.12 44.572 22.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 21.84 10.628 23.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 21.84 10.716 23.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.328 21.84 46.372 23.04 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 21.84 46.628 23.04 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 1.68 13.716 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.372 14.76 34.416 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.628 14.76 34.672 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 34.284 14.76 34.328 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.24 10.372 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 22.56 13.072 23.76 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 22.56 13.328 23.76 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 22.56 48.428 23.76 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 22.56 48.516 23.76 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 23.28 14.528 24.48 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.28 14.616 24.48 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 23.28 44.916 24.48 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 23.28 45.128 24.48 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 24 11.016 25.2 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 24 11.272 25.2 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 1.68 44.572 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 24 47.016 25.2 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 24 47.272 25.2 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 24.72 13.328 25.92 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 24.72 13.416 25.92 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 24.72 48.516 25.92 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 24.72 48.728 25.92 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 25.44 14.616 26.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 25.44 10.028 26.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 25.44 45.128 26.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 25.44 45.216 26.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 1.68 44.828 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 26.16 11.528 27.36 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 26.16 11.616 27.36 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 26.16 47.272 27.36 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 26.16 47.528 27.36 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 26.88 13.416 28.08 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 26.88 13.628 28.08 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 26.88 48.728 28.08 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 26.88 48.816 28.08 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 27.6 10.028 28.8 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 27.6 10.116 28.8 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 2.4 10.716 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 27.6 45.216 28.8 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.428 27.6 45.472 28.8 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 28.32 11.828 29.52 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 28.32 11.916 29.52 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 28.32 47.528 29.52 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 28.32 47.616 29.52 ;
    END
  END rddatap0[135]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 2.4 10.928 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.328 2.4 46.372 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.584 2.4 46.628 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 3.12 12.816 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 3.12 13.072 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 3.12 48.172 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.384 3.12 48.428 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 0.24 10.628 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 3.84 14.316 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 3.84 14.528 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 3.84 44.916 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 3.84 45.128 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 4.56 11.016 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 4.56 11.272 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 4.56 47.016 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 4.56 47.272 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 5.28 13.328 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 5.28 13.416 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 0.24 45.728 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.472 5.28 48.516 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 5.28 48.728 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6 14.616 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 6 10.028 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.084 6 45.128 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 6 45.216 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 6.72 11.528 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 6.72 11.616 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.228 6.72 47.272 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 6.72 47.528 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.772 0.24 45.816 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 7.44 13.416 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 7.44 13.628 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.684 7.44 48.728 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 7.44 48.816 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 8.16 10.028 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.16 10.116 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.172 8.16 45.216 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.428 8.16 45.472 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 8.88 11.828 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 8.88 11.916 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 0.96 12.516 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.484 8.88 47.528 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 8.88 47.616 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 9.6 13.628 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 9.6 13.716 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.772 9.6 48.816 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 9.6 49.072 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 10.32 10.116 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 10.32 10.372 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.428 10.32 45.472 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.684 10.32 45.728 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 0.96 12.728 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 11.04 12.172 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 11.04 12.428 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.572 11.04 47.616 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 11.04 47.828 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 11.76 13.716 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 11.76 13.972 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 11.76 49.072 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 11.76 44.572 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 12.48 10.628 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 12.48 10.716 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.784 0.96 47.828 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 12.48 46.028 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.072 12.48 46.116 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 13.2 12.728 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 13.2 12.816 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 13.2 47.916 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 13.2 48.172 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 18.24 11.616 19.44 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 18.24 11.828 19.44 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 18.24 46.928 19.44 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.972 18.24 47.016 19.44 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 0.96 47.916 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 18.96 13.716 20.16 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 18.96 13.972 20.16 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 49.028 18.96 49.072 20.16 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.528 18.96 44.572 20.16 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 19.68 10.628 20.88 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 19.68 10.716 20.88 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 45.984 19.68 46.028 20.88 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.072 19.68 46.116 20.88 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 20.4 12.728 21.6 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 20.4 12.816 21.6 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 1.68 13.972 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 47.872 20.4 47.916 21.6 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 48.128 20.4 48.172 21.6 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 21.12 14.228 22.32 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 21.12 14.316 22.32 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.784 21.12 44.828 22.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 44.872 21.12 44.916 22.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 21.84 10.928 23.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 21.84 11.016 23.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.672 21.84 46.716 23.04 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 46.884 21.84 46.928 23.04 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 1.68 14.228 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 29.7 ;
        RECT 2.662 0.06 2.738 29.7 ;
        RECT 4.462 0.06 4.538 29.7 ;
        RECT 6.262 0.06 6.338 29.7 ;
        RECT 8.062 0.06 8.138 29.7 ;
        RECT 9.862 0.06 9.938 29.7 ;
        RECT 11.662 0.06 11.738 29.7 ;
        RECT 13.462 0.06 13.538 29.7 ;
        RECT 15.262 0.06 15.338 29.7 ;
        RECT 17.062 0.06 17.138 29.7 ;
        RECT 18.862 0.06 18.938 29.7 ;
        RECT 20.662 0.06 20.738 29.7 ;
        RECT 22.462 0.06 22.538 29.7 ;
        RECT 24.262 0.06 24.338 29.7 ;
        RECT 26.062 0.06 26.138 29.7 ;
        RECT 27.862 0.06 27.938 29.7 ;
        RECT 29.662 0.06 29.738 29.7 ;
        RECT 31.462 0.06 31.538 29.7 ;
        RECT 33.262 0.06 33.338 29.7 ;
        RECT 35.062 0.06 35.138 29.7 ;
        RECT 36.862 0.06 36.938 29.7 ;
        RECT 38.662 0.06 38.738 29.7 ;
        RECT 40.462 0.06 40.538 29.7 ;
        RECT 42.262 0.06 42.338 29.7 ;
        RECT 44.062 0.06 44.138 29.7 ;
        RECT 45.862 0.06 45.938 29.7 ;
        RECT 47.662 0.06 47.738 29.7 ;
        RECT 49.462 0.06 49.538 29.7 ;
        RECT 51.262 0.06 51.338 29.7 ;
        RECT 53.062 0.06 53.138 29.7 ;
        RECT 54.862 0.06 54.938 29.7 ;
        RECT 56.662 0.06 56.738 29.7 ;
        RECT 58.462 0.06 58.538 29.7 ;
        RECT 60.262 0.06 60.338 29.7 ;
        RECT 62.062 0.06 62.138 29.7 ;
        RECT 63.862 0.06 63.938 29.7 ;
        RECT 65.662 0.06 65.738 29.7 ;
        RECT 67.462 0.06 67.538 29.7 ;
        RECT 69.262 0.06 69.338 29.7 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 29.7 ;
        RECT 3.562 0.06 3.638 29.7 ;
        RECT 5.362 0.06 5.438 29.7 ;
        RECT 7.162 0.06 7.238 29.7 ;
        RECT 8.962 0.06 9.038 29.7 ;
        RECT 10.762 0.06 10.838 29.7 ;
        RECT 12.562 0.06 12.638 29.7 ;
        RECT 14.362 0.06 14.438 29.7 ;
        RECT 16.162 0.06 16.238 29.7 ;
        RECT 17.962 0.06 18.038 29.7 ;
        RECT 19.762 0.06 19.838 29.7 ;
        RECT 21.562 0.06 21.638 29.7 ;
        RECT 23.362 0.06 23.438 29.7 ;
        RECT 25.162 0.06 25.238 29.7 ;
        RECT 26.962 0.06 27.038 29.7 ;
        RECT 28.762 0.06 28.838 29.7 ;
        RECT 30.562 0.06 30.638 29.7 ;
        RECT 32.362 0.06 32.438 29.7 ;
        RECT 34.162 0.06 34.238 29.7 ;
        RECT 35.962 0.06 36.038 29.7 ;
        RECT 37.762 0.06 37.838 29.7 ;
        RECT 39.562 0.06 39.638 29.7 ;
        RECT 41.362 0.06 41.438 29.7 ;
        RECT 43.162 0.06 43.238 29.7 ;
        RECT 44.962 0.06 45.038 29.7 ;
        RECT 46.762 0.06 46.838 29.7 ;
        RECT 48.562 0.06 48.638 29.7 ;
        RECT 50.362 0.06 50.438 29.7 ;
        RECT 52.162 0.06 52.238 29.7 ;
        RECT 53.962 0.06 54.038 29.7 ;
        RECT 55.762 0.06 55.838 29.7 ;
        RECT 57.562 0.06 57.638 29.7 ;
        RECT 59.362 0.06 59.438 29.7 ;
        RECT 61.162 0.06 61.238 29.7 ;
        RECT 62.962 0.06 63.038 29.7 ;
        RECT 64.762 0.06 64.838 29.7 ;
        RECT 66.562 0.06 66.638 29.7 ;
        RECT 68.362 0.06 68.438 29.7 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 70.216 29.774 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 70.22 29.78 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 70.2705 29.798 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 70.235 29.83 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 70.27 29.798 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 70.259 29.85 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 70.29 29.822 ;
    LAYER m7 SPACING 0 ;
      RECT 69.338 29.82 70.24 29.88 ;
      RECT 69.338 -0.06 70.292 29.82 ;
      RECT 69.338 -0.12 70.24 -0.06 ;
      RECT 68.438 -0.12 69.262 29.88 ;
      RECT 67.538 -0.12 68.362 29.88 ;
      RECT 66.638 -0.12 67.462 29.88 ;
      RECT 65.738 -0.12 66.562 29.88 ;
      RECT 64.838 -0.12 65.662 29.88 ;
      RECT 63.938 -0.12 64.762 29.88 ;
      RECT 63.038 -0.12 63.862 29.88 ;
      RECT 62.138 -0.12 62.962 29.88 ;
      RECT 61.238 -0.12 62.062 29.88 ;
      RECT 60.338 -0.12 61.162 29.88 ;
      RECT 59.438 -0.12 60.262 29.88 ;
      RECT 58.538 -0.12 59.362 29.88 ;
      RECT 57.638 -0.12 58.462 29.88 ;
      RECT 56.738 -0.12 57.562 29.88 ;
      RECT 55.838 -0.12 56.662 29.88 ;
      RECT 54.938 -0.12 55.762 29.88 ;
      RECT 54.038 -0.12 54.862 29.88 ;
      RECT 53.138 -0.12 53.962 29.88 ;
      RECT 52.238 -0.12 53.062 29.88 ;
      RECT 51.338 -0.12 52.162 29.88 ;
      RECT 50.438 -0.12 51.262 29.88 ;
      RECT 49.538 -0.12 50.362 29.88 ;
      RECT 48.638 28.08 49.462 29.88 ;
      RECT 48.638 26.88 48.684 28.08 ;
      RECT 48.728 26.88 48.772 28.08 ;
      RECT 48.816 26.88 49.462 28.08 ;
      RECT 48.638 25.92 49.462 26.88 ;
      RECT 48.638 24.72 48.684 25.92 ;
      RECT 48.728 24.72 49.462 25.92 ;
      RECT 48.638 22.32 49.462 24.72 ;
      RECT 48.638 21.12 49.028 22.32 ;
      RECT 49.072 21.12 49.462 22.32 ;
      RECT 48.638 20.16 49.462 21.12 ;
      RECT 48.638 18.96 48.684 20.16 ;
      RECT 48.728 18.96 48.772 20.16 ;
      RECT 48.816 18.96 49.028 20.16 ;
      RECT 49.072 18.96 49.462 20.16 ;
      RECT 48.638 12.96 49.462 18.96 ;
      RECT 48.638 11.76 48.684 12.96 ;
      RECT 48.728 11.76 48.772 12.96 ;
      RECT 48.816 11.76 49.028 12.96 ;
      RECT 49.072 11.76 49.462 12.96 ;
      RECT 48.638 10.8 49.462 11.76 ;
      RECT 48.638 9.6 48.684 10.8 ;
      RECT 48.728 9.6 48.772 10.8 ;
      RECT 48.816 9.6 49.028 10.8 ;
      RECT 49.072 9.6 49.462 10.8 ;
      RECT 48.638 8.64 49.462 9.6 ;
      RECT 48.638 7.44 48.684 8.64 ;
      RECT 48.728 7.44 48.772 8.64 ;
      RECT 48.816 7.44 49.462 8.64 ;
      RECT 48.638 6.48 49.462 7.44 ;
      RECT 48.638 5.28 48.684 6.48 ;
      RECT 48.728 5.28 49.462 6.48 ;
      RECT 48.638 2.88 49.462 5.28 ;
      RECT 48.638 1.68 48.772 2.88 ;
      RECT 48.816 1.68 49.028 2.88 ;
      RECT 49.072 1.68 49.462 2.88 ;
      RECT 48.638 -0.12 49.462 1.68 ;
      RECT 47.738 28.08 48.562 29.88 ;
      RECT 47.738 26.88 48.384 28.08 ;
      RECT 48.428 26.88 48.472 28.08 ;
      RECT 48.516 26.88 48.562 28.08 ;
      RECT 47.738 25.92 48.562 26.88 ;
      RECT 47.738 24.72 48.128 25.92 ;
      RECT 48.172 24.72 48.384 25.92 ;
      RECT 48.428 24.72 48.472 25.92 ;
      RECT 48.516 24.72 48.562 25.92 ;
      RECT 47.738 23.76 48.562 24.72 ;
      RECT 47.738 22.56 47.872 23.76 ;
      RECT 47.916 22.56 48.128 23.76 ;
      RECT 48.172 22.56 48.384 23.76 ;
      RECT 48.428 22.56 48.472 23.76 ;
      RECT 48.516 22.56 48.562 23.76 ;
      RECT 47.738 21.6 48.562 22.56 ;
      RECT 47.738 20.4 47.784 21.6 ;
      RECT 47.828 20.4 47.872 21.6 ;
      RECT 47.916 20.4 48.128 21.6 ;
      RECT 48.172 20.4 48.562 21.6 ;
      RECT 47.738 14.4 48.562 20.4 ;
      RECT 47.738 13.2 47.784 14.4 ;
      RECT 47.828 13.2 47.872 14.4 ;
      RECT 47.916 13.2 48.128 14.4 ;
      RECT 48.172 13.2 48.562 14.4 ;
      RECT 47.738 12.24 48.562 13.2 ;
      RECT 47.738 11.04 47.784 12.24 ;
      RECT 47.828 11.04 48.562 12.24 ;
      RECT 47.738 10.8 48.562 11.04 ;
      RECT 47.738 9.6 48.472 10.8 ;
      RECT 48.516 9.6 48.562 10.8 ;
      RECT 47.738 8.64 48.562 9.6 ;
      RECT 47.738 7.44 48.384 8.64 ;
      RECT 48.428 7.44 48.472 8.64 ;
      RECT 48.516 7.44 48.562 8.64 ;
      RECT 47.738 6.48 48.562 7.44 ;
      RECT 47.738 5.28 48.128 6.48 ;
      RECT 48.172 5.28 48.384 6.48 ;
      RECT 48.428 5.28 48.472 6.48 ;
      RECT 48.516 5.28 48.562 6.48 ;
      RECT 47.738 4.32 48.562 5.28 ;
      RECT 47.738 3.12 47.784 4.32 ;
      RECT 47.828 3.12 47.872 4.32 ;
      RECT 47.916 3.12 48.128 4.32 ;
      RECT 48.172 3.12 48.384 4.32 ;
      RECT 48.428 3.12 48.562 4.32 ;
      RECT 47.738 2.16 48.562 3.12 ;
      RECT 47.738 0.96 47.784 2.16 ;
      RECT 47.828 0.96 47.872 2.16 ;
      RECT 47.916 0.96 48.562 2.16 ;
      RECT 47.738 -0.12 48.562 0.96 ;
      RECT 46.838 29.52 47.662 29.88 ;
      RECT 46.838 28.32 46.972 29.52 ;
      RECT 47.016 28.32 47.228 29.52 ;
      RECT 47.272 28.32 47.484 29.52 ;
      RECT 47.528 28.32 47.572 29.52 ;
      RECT 47.616 28.32 47.662 29.52 ;
      RECT 46.838 27.36 47.662 28.32 ;
      RECT 46.838 26.16 46.884 27.36 ;
      RECT 46.928 26.16 46.972 27.36 ;
      RECT 47.016 26.16 47.228 27.36 ;
      RECT 47.272 26.16 47.484 27.36 ;
      RECT 47.528 26.16 47.662 27.36 ;
      RECT 46.838 25.2 47.662 26.16 ;
      RECT 46.838 24 46.884 25.2 ;
      RECT 46.928 24 46.972 25.2 ;
      RECT 47.016 24 47.228 25.2 ;
      RECT 47.272 24 47.662 25.2 ;
      RECT 46.838 23.04 47.662 24 ;
      RECT 46.838 21.84 46.884 23.04 ;
      RECT 46.928 21.84 47.662 23.04 ;
      RECT 46.838 21.6 47.662 21.84 ;
      RECT 46.838 20.4 47.572 21.6 ;
      RECT 47.616 20.4 47.662 21.6 ;
      RECT 46.838 19.44 47.662 20.4 ;
      RECT 46.838 18.24 46.884 19.44 ;
      RECT 46.928 18.24 46.972 19.44 ;
      RECT 47.016 18.24 47.662 19.44 ;
      RECT 46.838 14.4 47.662 18.24 ;
      RECT 46.838 13.2 47.572 14.4 ;
      RECT 47.616 13.2 47.662 14.4 ;
      RECT 46.838 12.24 47.662 13.2 ;
      RECT 46.838 11.04 47.228 12.24 ;
      RECT 47.272 11.04 47.484 12.24 ;
      RECT 47.528 11.04 47.572 12.24 ;
      RECT 47.616 11.04 47.662 12.24 ;
      RECT 46.838 10.08 47.662 11.04 ;
      RECT 46.838 8.88 46.972 10.08 ;
      RECT 47.016 8.88 47.228 10.08 ;
      RECT 47.272 8.88 47.484 10.08 ;
      RECT 47.528 8.88 47.572 10.08 ;
      RECT 47.616 8.88 47.662 10.08 ;
      RECT 46.838 7.92 47.662 8.88 ;
      RECT 46.838 6.72 46.884 7.92 ;
      RECT 46.928 6.72 46.972 7.92 ;
      RECT 47.016 6.72 47.228 7.92 ;
      RECT 47.272 6.72 47.484 7.92 ;
      RECT 47.528 6.72 47.662 7.92 ;
      RECT 46.838 5.76 47.662 6.72 ;
      RECT 46.838 4.56 46.884 5.76 ;
      RECT 46.928 4.56 46.972 5.76 ;
      RECT 47.016 4.56 47.228 5.76 ;
      RECT 47.272 4.56 47.662 5.76 ;
      RECT 46.838 2.16 47.662 4.56 ;
      RECT 46.838 0.96 47.484 2.16 ;
      RECT 47.528 0.96 47.572 2.16 ;
      RECT 47.616 0.96 47.662 2.16 ;
      RECT 46.838 -0.12 47.662 0.96 ;
      RECT 45.938 25.2 46.762 29.88 ;
      RECT 45.938 24 46.672 25.2 ;
      RECT 46.716 24 46.762 25.2 ;
      RECT 45.938 23.04 46.762 24 ;
      RECT 45.938 21.84 46.328 23.04 ;
      RECT 46.372 21.84 46.584 23.04 ;
      RECT 46.628 21.84 46.672 23.04 ;
      RECT 46.716 21.84 46.762 23.04 ;
      RECT 45.938 20.88 46.762 21.84 ;
      RECT 45.938 19.68 45.984 20.88 ;
      RECT 46.028 19.68 46.072 20.88 ;
      RECT 46.116 19.68 46.762 20.88 ;
      RECT 45.938 19.44 46.762 19.68 ;
      RECT 45.938 18.24 46.584 19.44 ;
      RECT 46.628 18.24 46.672 19.44 ;
      RECT 46.716 18.24 46.762 19.44 ;
      RECT 45.938 13.68 46.762 18.24 ;
      RECT 45.938 12.48 45.984 13.68 ;
      RECT 46.028 12.48 46.072 13.68 ;
      RECT 46.116 12.48 46.762 13.68 ;
      RECT 45.938 5.76 46.762 12.48 ;
      RECT 45.938 4.56 46.672 5.76 ;
      RECT 46.716 4.56 46.762 5.76 ;
      RECT 45.938 3.6 46.762 4.56 ;
      RECT 45.938 2.4 45.984 3.6 ;
      RECT 46.028 2.4 46.072 3.6 ;
      RECT 46.116 2.4 46.328 3.6 ;
      RECT 46.372 2.4 46.584 3.6 ;
      RECT 46.628 2.4 46.762 3.6 ;
      RECT 45.938 -0.12 46.762 2.4 ;
      RECT 45.038 28.8 45.862 29.88 ;
      RECT 45.038 27.6 45.084 28.8 ;
      RECT 45.128 27.6 45.172 28.8 ;
      RECT 45.216 27.6 45.428 28.8 ;
      RECT 45.472 27.6 45.862 28.8 ;
      RECT 45.038 26.64 45.862 27.6 ;
      RECT 45.038 25.44 45.084 26.64 ;
      RECT 45.128 25.44 45.172 26.64 ;
      RECT 45.216 25.44 45.862 26.64 ;
      RECT 45.038 24.48 45.862 25.44 ;
      RECT 45.038 23.28 45.084 24.48 ;
      RECT 45.128 23.28 45.862 24.48 ;
      RECT 45.038 20.88 45.862 23.28 ;
      RECT 45.038 19.68 45.684 20.88 ;
      RECT 45.728 19.68 45.772 20.88 ;
      RECT 45.816 19.68 45.862 20.88 ;
      RECT 45.038 13.68 45.862 19.68 ;
      RECT 45.038 12.48 45.684 13.68 ;
      RECT 45.728 12.48 45.772 13.68 ;
      RECT 45.816 12.48 45.862 13.68 ;
      RECT 45.038 11.52 45.862 12.48 ;
      RECT 45.038 10.32 45.084 11.52 ;
      RECT 45.128 10.32 45.172 11.52 ;
      RECT 45.216 10.32 45.428 11.52 ;
      RECT 45.472 10.32 45.684 11.52 ;
      RECT 45.728 10.32 45.862 11.52 ;
      RECT 45.038 9.36 45.862 10.32 ;
      RECT 45.038 8.16 45.084 9.36 ;
      RECT 45.128 8.16 45.172 9.36 ;
      RECT 45.216 8.16 45.428 9.36 ;
      RECT 45.472 8.16 45.862 9.36 ;
      RECT 45.038 7.2 45.862 8.16 ;
      RECT 45.038 6 45.084 7.2 ;
      RECT 45.128 6 45.172 7.2 ;
      RECT 45.216 6 45.862 7.2 ;
      RECT 45.038 5.04 45.862 6 ;
      RECT 45.038 3.84 45.084 5.04 ;
      RECT 45.128 3.84 45.862 5.04 ;
      RECT 45.038 1.44 45.862 3.84 ;
      RECT 45.038 0.24 45.172 1.44 ;
      RECT 45.216 0.24 45.428 1.44 ;
      RECT 45.472 0.24 45.684 1.44 ;
      RECT 45.728 0.24 45.772 1.44 ;
      RECT 45.816 0.24 45.862 1.44 ;
      RECT 45.038 -0.12 45.862 0.24 ;
      RECT 44.138 28.8 44.962 29.88 ;
      RECT 44.138 27.6 44.872 28.8 ;
      RECT 44.916 27.6 44.962 28.8 ;
      RECT 44.138 26.64 44.962 27.6 ;
      RECT 44.138 25.44 44.784 26.64 ;
      RECT 44.828 25.44 44.872 26.64 ;
      RECT 44.916 25.44 44.962 26.64 ;
      RECT 44.138 24.48 44.962 25.44 ;
      RECT 44.138 23.28 44.528 24.48 ;
      RECT 44.572 23.28 44.784 24.48 ;
      RECT 44.828 23.28 44.872 24.48 ;
      RECT 44.916 23.28 44.962 24.48 ;
      RECT 44.138 22.32 44.962 23.28 ;
      RECT 44.138 21.12 44.528 22.32 ;
      RECT 44.572 21.12 44.784 22.32 ;
      RECT 44.828 21.12 44.872 22.32 ;
      RECT 44.916 21.12 44.962 22.32 ;
      RECT 44.138 20.16 44.962 21.12 ;
      RECT 44.138 18.96 44.528 20.16 ;
      RECT 44.572 18.96 44.962 20.16 ;
      RECT 44.138 12.96 44.962 18.96 ;
      RECT 44.138 11.76 44.528 12.96 ;
      RECT 44.572 11.76 44.962 12.96 ;
      RECT 44.138 9.36 44.962 11.76 ;
      RECT 44.138 8.16 44.872 9.36 ;
      RECT 44.916 8.16 44.962 9.36 ;
      RECT 44.138 7.2 44.962 8.16 ;
      RECT 44.138 6 44.784 7.2 ;
      RECT 44.828 6 44.872 7.2 ;
      RECT 44.916 6 44.962 7.2 ;
      RECT 44.138 5.04 44.962 6 ;
      RECT 44.138 3.84 44.528 5.04 ;
      RECT 44.572 3.84 44.784 5.04 ;
      RECT 44.828 3.84 44.872 5.04 ;
      RECT 44.916 3.84 44.962 5.04 ;
      RECT 44.138 2.88 44.962 3.84 ;
      RECT 44.138 1.68 44.528 2.88 ;
      RECT 44.572 1.68 44.784 2.88 ;
      RECT 44.828 1.68 44.962 2.88 ;
      RECT 44.138 -0.12 44.962 1.68 ;
      RECT 43.238 -0.12 44.062 29.88 ;
      RECT 42.338 -0.12 43.162 29.88 ;
      RECT 41.438 -0.12 42.262 29.88 ;
      RECT 40.538 -0.12 41.362 29.88 ;
      RECT 39.638 -0.12 40.462 29.88 ;
      RECT 38.738 -0.12 39.562 29.88 ;
      RECT 37.838 -0.12 38.662 29.88 ;
      RECT 36.938 -0.12 37.762 29.88 ;
      RECT 36.038 -0.12 36.862 29.88 ;
      RECT 35.138 17.88 35.962 29.88 ;
      RECT 35.138 16.68 35.184 17.88 ;
      RECT 35.228 16.68 35.272 17.88 ;
      RECT 35.316 16.68 35.962 17.88 ;
      RECT 35.138 15.96 35.962 16.68 ;
      RECT 35.138 14.76 35.184 15.96 ;
      RECT 35.228 14.76 35.272 15.96 ;
      RECT 35.316 14.76 35.962 15.96 ;
      RECT 35.138 -0.12 35.962 14.76 ;
      RECT 34.238 19.8 35.062 29.88 ;
      RECT 34.238 18.6 34.372 19.8 ;
      RECT 34.416 18.6 34.628 19.8 ;
      RECT 34.672 18.6 34.884 19.8 ;
      RECT 34.928 18.6 35.062 19.8 ;
      RECT 34.238 17.88 35.062 18.6 ;
      RECT 34.238 16.68 34.284 17.88 ;
      RECT 34.328 16.68 34.372 17.88 ;
      RECT 34.416 16.68 34.628 17.88 ;
      RECT 34.672 16.68 34.884 17.88 ;
      RECT 34.928 16.68 34.972 17.88 ;
      RECT 35.016 16.68 35.062 17.88 ;
      RECT 34.238 15.96 35.062 16.68 ;
      RECT 34.238 14.76 34.284 15.96 ;
      RECT 34.328 14.76 34.372 15.96 ;
      RECT 34.416 14.76 34.628 15.96 ;
      RECT 34.672 14.76 34.884 15.96 ;
      RECT 34.928 14.76 34.972 15.96 ;
      RECT 35.016 14.76 35.062 15.96 ;
      RECT 34.238 14.04 35.062 14.76 ;
      RECT 34.238 12.84 34.284 14.04 ;
      RECT 34.328 12.84 35.062 14.04 ;
      RECT 34.238 -0.12 35.062 12.84 ;
      RECT 33.338 17.88 34.162 29.88 ;
      RECT 33.338 16.68 33.728 17.88 ;
      RECT 33.772 16.68 33.984 17.88 ;
      RECT 34.028 16.68 34.072 17.88 ;
      RECT 34.116 16.68 34.162 17.88 ;
      RECT 33.338 15.96 34.162 16.68 ;
      RECT 33.338 14.76 33.728 15.96 ;
      RECT 33.772 14.76 33.984 15.96 ;
      RECT 34.028 14.76 34.072 15.96 ;
      RECT 34.116 14.76 34.162 15.96 ;
      RECT 33.338 14.04 34.162 14.76 ;
      RECT 33.338 12.84 33.728 14.04 ;
      RECT 33.772 12.84 33.984 14.04 ;
      RECT 34.028 12.84 34.072 14.04 ;
      RECT 34.116 12.84 34.162 14.04 ;
      RECT 33.338 -0.12 34.162 12.84 ;
      RECT 32.438 -0.12 33.262 29.88 ;
      RECT 31.538 -0.12 32.362 29.88 ;
      RECT 30.638 -0.12 31.462 29.88 ;
      RECT 29.738 -0.12 30.562 29.88 ;
      RECT 28.838 -0.12 29.662 29.88 ;
      RECT 27.938 -0.12 28.762 29.88 ;
      RECT 27.038 -0.12 27.862 29.88 ;
      RECT 26.138 -0.12 26.962 29.88 ;
      RECT 25.238 -0.12 26.062 29.88 ;
      RECT 24.338 -0.12 25.162 29.88 ;
      RECT 23.438 -0.12 24.262 29.88 ;
      RECT 22.538 -0.12 23.362 29.88 ;
      RECT 21.638 -0.12 22.462 29.88 ;
      RECT 20.738 -0.12 21.562 29.88 ;
      RECT 19.838 -0.12 20.662 29.88 ;
      RECT 18.938 -0.12 19.762 29.88 ;
      RECT 18.038 -0.12 18.862 29.88 ;
      RECT 17.138 -0.12 17.962 29.88 ;
      RECT 16.238 -0.12 17.062 29.88 ;
      RECT 15.338 -0.12 16.162 29.88 ;
      RECT 14.438 28.8 15.262 29.88 ;
      RECT 14.438 27.6 14.484 28.8 ;
      RECT 14.528 27.6 14.572 28.8 ;
      RECT 14.616 27.6 15.262 28.8 ;
      RECT 14.438 26.64 15.262 27.6 ;
      RECT 14.438 25.44 14.484 26.64 ;
      RECT 14.528 25.44 14.572 26.64 ;
      RECT 14.616 25.44 15.262 26.64 ;
      RECT 14.438 24.48 15.262 25.44 ;
      RECT 14.438 23.28 14.484 24.48 ;
      RECT 14.528 23.28 14.572 24.48 ;
      RECT 14.616 23.28 15.262 24.48 ;
      RECT 14.438 11.52 15.262 23.28 ;
      RECT 14.438 10.32 14.572 11.52 ;
      RECT 14.616 10.32 15.262 11.52 ;
      RECT 14.438 9.36 15.262 10.32 ;
      RECT 14.438 8.16 14.484 9.36 ;
      RECT 14.528 8.16 14.572 9.36 ;
      RECT 14.616 8.16 15.262 9.36 ;
      RECT 14.438 7.2 15.262 8.16 ;
      RECT 14.438 6 14.484 7.2 ;
      RECT 14.528 6 14.572 7.2 ;
      RECT 14.616 6 15.262 7.2 ;
      RECT 14.438 5.04 15.262 6 ;
      RECT 14.438 3.84 14.484 5.04 ;
      RECT 14.528 3.84 15.262 5.04 ;
      RECT 14.438 -0.12 15.262 3.84 ;
      RECT 13.538 28.08 14.362 29.88 ;
      RECT 13.538 26.88 13.584 28.08 ;
      RECT 13.628 26.88 14.362 28.08 ;
      RECT 13.538 26.64 14.362 26.88 ;
      RECT 13.538 25.44 14.272 26.64 ;
      RECT 14.316 25.44 14.362 26.64 ;
      RECT 13.538 24.48 14.362 25.44 ;
      RECT 13.538 23.28 14.184 24.48 ;
      RECT 14.228 23.28 14.272 24.48 ;
      RECT 14.316 23.28 14.362 24.48 ;
      RECT 13.538 22.32 14.362 23.28 ;
      RECT 13.538 21.12 13.672 22.32 ;
      RECT 13.716 21.12 13.928 22.32 ;
      RECT 13.972 21.12 14.184 22.32 ;
      RECT 14.228 21.12 14.272 22.32 ;
      RECT 14.316 21.12 14.362 22.32 ;
      RECT 13.538 20.16 14.362 21.12 ;
      RECT 13.538 18.96 13.584 20.16 ;
      RECT 13.628 18.96 13.672 20.16 ;
      RECT 13.716 18.96 13.928 20.16 ;
      RECT 13.972 18.96 14.362 20.16 ;
      RECT 13.538 12.96 14.362 18.96 ;
      RECT 13.538 11.76 13.584 12.96 ;
      RECT 13.628 11.76 13.672 12.96 ;
      RECT 13.716 11.76 13.928 12.96 ;
      RECT 13.972 11.76 14.362 12.96 ;
      RECT 13.538 10.8 14.362 11.76 ;
      RECT 13.538 9.6 13.584 10.8 ;
      RECT 13.628 9.6 13.672 10.8 ;
      RECT 13.716 9.6 14.362 10.8 ;
      RECT 13.538 8.64 14.362 9.6 ;
      RECT 13.538 7.44 13.584 8.64 ;
      RECT 13.628 7.44 14.362 8.64 ;
      RECT 13.538 7.2 14.362 7.44 ;
      RECT 13.538 6 14.272 7.2 ;
      RECT 14.316 6 14.362 7.2 ;
      RECT 13.538 5.04 14.362 6 ;
      RECT 13.538 3.84 13.928 5.04 ;
      RECT 13.972 3.84 14.184 5.04 ;
      RECT 14.228 3.84 14.272 5.04 ;
      RECT 14.316 3.84 14.362 5.04 ;
      RECT 13.538 2.88 14.362 3.84 ;
      RECT 13.538 1.68 13.584 2.88 ;
      RECT 13.628 1.68 13.672 2.88 ;
      RECT 13.716 1.68 13.928 2.88 ;
      RECT 13.972 1.68 14.184 2.88 ;
      RECT 14.228 1.68 14.362 2.88 ;
      RECT 13.538 -0.12 14.362 1.68 ;
      RECT 12.638 28.08 13.462 29.88 ;
      RECT 12.638 26.88 13.028 28.08 ;
      RECT 13.072 26.88 13.284 28.08 ;
      RECT 13.328 26.88 13.372 28.08 ;
      RECT 13.416 26.88 13.462 28.08 ;
      RECT 12.638 25.92 13.462 26.88 ;
      RECT 12.638 24.72 12.772 25.92 ;
      RECT 12.816 24.72 13.028 25.92 ;
      RECT 13.072 24.72 13.284 25.92 ;
      RECT 13.328 24.72 13.372 25.92 ;
      RECT 13.416 24.72 13.462 25.92 ;
      RECT 12.638 23.76 13.462 24.72 ;
      RECT 12.638 22.56 12.684 23.76 ;
      RECT 12.728 22.56 12.772 23.76 ;
      RECT 12.816 22.56 13.028 23.76 ;
      RECT 13.072 22.56 13.284 23.76 ;
      RECT 13.328 22.56 13.462 23.76 ;
      RECT 12.638 21.6 13.462 22.56 ;
      RECT 12.638 20.4 12.684 21.6 ;
      RECT 12.728 20.4 12.772 21.6 ;
      RECT 12.816 20.4 13.462 21.6 ;
      RECT 12.638 20.16 13.462 20.4 ;
      RECT 12.638 18.96 13.372 20.16 ;
      RECT 13.416 18.96 13.462 20.16 ;
      RECT 12.638 14.4 13.462 18.96 ;
      RECT 12.638 13.2 12.684 14.4 ;
      RECT 12.728 13.2 12.772 14.4 ;
      RECT 12.816 13.2 13.462 14.4 ;
      RECT 12.638 12.96 13.462 13.2 ;
      RECT 12.638 11.76 13.372 12.96 ;
      RECT 13.416 11.76 13.462 12.96 ;
      RECT 12.638 10.8 13.462 11.76 ;
      RECT 12.638 9.6 13.284 10.8 ;
      RECT 13.328 9.6 13.372 10.8 ;
      RECT 13.416 9.6 13.462 10.8 ;
      RECT 12.638 8.64 13.462 9.6 ;
      RECT 12.638 7.44 13.028 8.64 ;
      RECT 13.072 7.44 13.284 8.64 ;
      RECT 13.328 7.44 13.372 8.64 ;
      RECT 13.416 7.44 13.462 8.64 ;
      RECT 12.638 6.48 13.462 7.44 ;
      RECT 12.638 5.28 12.772 6.48 ;
      RECT 12.816 5.28 13.028 6.48 ;
      RECT 13.072 5.28 13.284 6.48 ;
      RECT 13.328 5.28 13.372 6.48 ;
      RECT 13.416 5.28 13.462 6.48 ;
      RECT 12.638 4.32 13.462 5.28 ;
      RECT 12.638 3.12 12.684 4.32 ;
      RECT 12.728 3.12 12.772 4.32 ;
      RECT 12.816 3.12 13.028 4.32 ;
      RECT 13.072 3.12 13.462 4.32 ;
      RECT 12.638 2.16 13.462 3.12 ;
      RECT 12.638 0.96 12.684 2.16 ;
      RECT 12.728 0.96 13.462 2.16 ;
      RECT 12.638 -0.12 13.462 0.96 ;
      RECT 11.738 29.52 12.562 29.88 ;
      RECT 11.738 28.32 11.784 29.52 ;
      RECT 11.828 28.32 11.872 29.52 ;
      RECT 11.916 28.32 12.562 29.52 ;
      RECT 11.738 21.6 12.562 28.32 ;
      RECT 11.738 20.4 12.384 21.6 ;
      RECT 12.428 20.4 12.472 21.6 ;
      RECT 12.516 20.4 12.562 21.6 ;
      RECT 11.738 19.44 12.562 20.4 ;
      RECT 11.738 18.24 11.784 19.44 ;
      RECT 11.828 18.24 12.562 19.44 ;
      RECT 11.738 14.4 12.562 18.24 ;
      RECT 11.738 13.2 12.384 14.4 ;
      RECT 12.428 13.2 12.472 14.4 ;
      RECT 12.516 13.2 12.562 14.4 ;
      RECT 11.738 12.24 12.562 13.2 ;
      RECT 11.738 11.04 11.784 12.24 ;
      RECT 11.828 11.04 11.872 12.24 ;
      RECT 11.916 11.04 12.128 12.24 ;
      RECT 12.172 11.04 12.384 12.24 ;
      RECT 12.428 11.04 12.562 12.24 ;
      RECT 11.738 10.08 12.562 11.04 ;
      RECT 11.738 8.88 11.784 10.08 ;
      RECT 11.828 8.88 11.872 10.08 ;
      RECT 11.916 8.88 12.562 10.08 ;
      RECT 11.738 4.32 12.562 8.88 ;
      RECT 11.738 3.12 12.472 4.32 ;
      RECT 12.516 3.12 12.562 4.32 ;
      RECT 11.738 2.16 12.562 3.12 ;
      RECT 11.738 0.96 12.128 2.16 ;
      RECT 12.172 0.96 12.384 2.16 ;
      RECT 12.428 0.96 12.472 2.16 ;
      RECT 12.516 0.96 12.562 2.16 ;
      RECT 11.738 -0.12 12.562 0.96 ;
      RECT 10.838 29.52 11.662 29.88 ;
      RECT 10.838 28.32 11.484 29.52 ;
      RECT 11.528 28.32 11.572 29.52 ;
      RECT 11.616 28.32 11.662 29.52 ;
      RECT 10.838 27.36 11.662 28.32 ;
      RECT 10.838 26.16 10.972 27.36 ;
      RECT 11.016 26.16 11.228 27.36 ;
      RECT 11.272 26.16 11.484 27.36 ;
      RECT 11.528 26.16 11.572 27.36 ;
      RECT 11.616 26.16 11.662 27.36 ;
      RECT 10.838 25.2 11.662 26.16 ;
      RECT 10.838 24 10.884 25.2 ;
      RECT 10.928 24 10.972 25.2 ;
      RECT 11.016 24 11.228 25.2 ;
      RECT 11.272 24 11.662 25.2 ;
      RECT 10.838 23.04 11.662 24 ;
      RECT 10.838 21.84 10.884 23.04 ;
      RECT 10.928 21.84 10.972 23.04 ;
      RECT 11.016 21.84 11.662 23.04 ;
      RECT 10.838 19.44 11.662 21.84 ;
      RECT 10.838 18.24 11.228 19.44 ;
      RECT 11.272 18.24 11.484 19.44 ;
      RECT 11.528 18.24 11.572 19.44 ;
      RECT 11.616 18.24 11.662 19.44 ;
      RECT 10.838 10.08 11.662 18.24 ;
      RECT 10.838 8.88 11.484 10.08 ;
      RECT 11.528 8.88 11.572 10.08 ;
      RECT 11.616 8.88 11.662 10.08 ;
      RECT 10.838 7.92 11.662 8.88 ;
      RECT 10.838 6.72 10.972 7.92 ;
      RECT 11.016 6.72 11.228 7.92 ;
      RECT 11.272 6.72 11.484 7.92 ;
      RECT 11.528 6.72 11.572 7.92 ;
      RECT 11.616 6.72 11.662 7.92 ;
      RECT 10.838 5.76 11.662 6.72 ;
      RECT 10.838 4.56 10.884 5.76 ;
      RECT 10.928 4.56 10.972 5.76 ;
      RECT 11.016 4.56 11.228 5.76 ;
      RECT 11.272 4.56 11.662 5.76 ;
      RECT 10.838 3.6 11.662 4.56 ;
      RECT 10.838 2.4 10.884 3.6 ;
      RECT 10.928 2.4 11.662 3.6 ;
      RECT 10.838 -0.12 11.662 2.4 ;
      RECT 9.938 28.8 10.762 29.88 ;
      RECT 9.938 27.6 9.984 28.8 ;
      RECT 10.028 27.6 10.072 28.8 ;
      RECT 10.116 27.6 10.762 28.8 ;
      RECT 9.938 26.64 10.762 27.6 ;
      RECT 9.938 25.44 9.984 26.64 ;
      RECT 10.028 25.44 10.762 26.64 ;
      RECT 9.938 25.2 10.762 25.44 ;
      RECT 9.938 24 10.672 25.2 ;
      RECT 10.716 24 10.762 25.2 ;
      RECT 9.938 23.04 10.762 24 ;
      RECT 9.938 21.84 10.584 23.04 ;
      RECT 10.628 21.84 10.672 23.04 ;
      RECT 10.716 21.84 10.762 23.04 ;
      RECT 9.938 20.88 10.762 21.84 ;
      RECT 9.938 19.68 10.072 20.88 ;
      RECT 10.116 19.68 10.328 20.88 ;
      RECT 10.372 19.68 10.584 20.88 ;
      RECT 10.628 19.68 10.672 20.88 ;
      RECT 10.716 19.68 10.762 20.88 ;
      RECT 9.938 13.68 10.762 19.68 ;
      RECT 9.938 12.48 10.072 13.68 ;
      RECT 10.116 12.48 10.328 13.68 ;
      RECT 10.372 12.48 10.584 13.68 ;
      RECT 10.628 12.48 10.672 13.68 ;
      RECT 10.716 12.48 10.762 13.68 ;
      RECT 9.938 11.52 10.762 12.48 ;
      RECT 9.938 10.32 9.984 11.52 ;
      RECT 10.028 10.32 10.072 11.52 ;
      RECT 10.116 10.32 10.328 11.52 ;
      RECT 10.372 10.32 10.762 11.52 ;
      RECT 9.938 9.36 10.762 10.32 ;
      RECT 9.938 8.16 9.984 9.36 ;
      RECT 10.028 8.16 10.072 9.36 ;
      RECT 10.116 8.16 10.762 9.36 ;
      RECT 9.938 7.2 10.762 8.16 ;
      RECT 9.938 6 9.984 7.2 ;
      RECT 10.028 6 10.762 7.2 ;
      RECT 9.938 5.76 10.762 6 ;
      RECT 9.938 4.56 10.672 5.76 ;
      RECT 10.716 4.56 10.762 5.76 ;
      RECT 9.938 3.6 10.762 4.56 ;
      RECT 9.938 2.4 10.328 3.6 ;
      RECT 10.372 2.4 10.584 3.6 ;
      RECT 10.628 2.4 10.672 3.6 ;
      RECT 10.716 2.4 10.762 3.6 ;
      RECT 9.938 1.44 10.762 2.4 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.328 1.44 ;
      RECT 10.372 0.24 10.584 1.44 ;
      RECT 10.628 0.24 10.762 1.44 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 29.88 ;
      RECT 8.138 -0.12 8.962 29.88 ;
      RECT 7.238 -0.12 8.062 29.88 ;
      RECT 6.338 -0.12 7.162 29.88 ;
      RECT 5.438 -0.12 6.262 29.88 ;
      RECT 4.538 -0.12 5.362 29.88 ;
      RECT 3.638 -0.12 4.462 29.88 ;
      RECT 2.738 -0.12 3.562 29.88 ;
      RECT 1.838 -0.12 2.662 29.88 ;
      RECT 0.938 -0.12 1.762 29.88 ;
      RECT -0.04 29.82 0.862 29.88 ;
      RECT -0.092 -0.06 0.862 29.82 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 69.458 0 70.12 29.76 ;
      RECT 68.558 0 69.142 29.76 ;
      RECT 67.658 0 68.242 29.76 ;
      RECT 66.758 0 67.342 29.76 ;
      RECT 65.858 0 66.442 29.76 ;
      RECT 64.958 0 65.542 29.76 ;
      RECT 64.058 0 64.642 29.76 ;
      RECT 63.158 0 63.742 29.76 ;
      RECT 62.258 0 62.842 29.76 ;
      RECT 61.358 0 61.942 29.76 ;
      RECT 60.458 0 61.042 29.76 ;
      RECT 59.558 0 60.142 29.76 ;
      RECT 58.658 0 59.242 29.76 ;
      RECT 57.758 0 58.342 29.76 ;
      RECT 56.858 0 57.442 29.76 ;
      RECT 55.958 0 56.542 29.76 ;
      RECT 55.058 0 55.642 29.76 ;
      RECT 54.158 0 54.742 29.76 ;
      RECT 53.258 0 53.842 29.76 ;
      RECT 52.358 0 52.942 29.76 ;
      RECT 51.458 0 52.042 29.76 ;
      RECT 50.558 0 51.142 29.76 ;
      RECT 49.658 0 50.242 29.76 ;
      RECT 48.758 28.2 49.342 29.76 ;
      RECT 48.936 26.76 49.342 28.2 ;
      RECT 48.758 26.04 49.342 26.76 ;
      RECT 48.848 24.6 49.342 26.04 ;
      RECT 48.758 22.44 49.342 24.6 ;
      RECT 48.758 21 48.908 22.44 ;
      RECT 49.192 21 49.342 22.44 ;
      RECT 48.758 20.28 49.342 21 ;
      RECT 49.192 18.84 49.342 20.28 ;
      RECT 48.758 13.08 49.342 18.84 ;
      RECT 49.192 11.64 49.342 13.08 ;
      RECT 48.758 10.92 49.342 11.64 ;
      RECT 49.192 9.48 49.342 10.92 ;
      RECT 48.758 8.76 49.342 9.48 ;
      RECT 48.936 7.32 49.342 8.76 ;
      RECT 48.758 6.6 49.342 7.32 ;
      RECT 48.848 5.16 49.342 6.6 ;
      RECT 48.758 3 49.342 5.16 ;
      RECT 49.192 1.56 49.342 3 ;
      RECT 48.758 0 49.342 1.56 ;
      RECT 47.858 28.2 48.442 29.76 ;
      RECT 47.858 26.76 48.264 28.2 ;
      RECT 47.858 26.04 48.442 26.76 ;
      RECT 47.858 24.6 48.008 26.04 ;
      RECT 47.858 23.88 48.442 24.6 ;
      RECT 46.958 29.64 47.542 29.76 ;
      RECT 46.058 25.32 46.642 29.76 ;
      RECT 46.058 23.88 46.552 25.32 ;
      RECT 46.058 23.16 46.642 23.88 ;
      RECT 46.058 21.72 46.208 23.16 ;
      RECT 46.058 21 46.642 21.72 ;
      RECT 46.236 19.56 46.642 21 ;
      RECT 46.058 18.12 46.464 19.56 ;
      RECT 46.058 13.8 46.642 18.12 ;
      RECT 46.236 12.36 46.642 13.8 ;
      RECT 46.058 5.88 46.642 12.36 ;
      RECT 46.058 4.44 46.552 5.88 ;
      RECT 46.058 3.72 46.642 4.44 ;
      RECT 45.158 28.92 45.742 29.76 ;
      RECT 45.592 27.48 45.742 28.92 ;
      RECT 45.158 26.76 45.742 27.48 ;
      RECT 45.336 25.32 45.742 26.76 ;
      RECT 45.158 24.6 45.742 25.32 ;
      RECT 45.248 23.16 45.742 24.6 ;
      RECT 45.158 21 45.742 23.16 ;
      RECT 45.158 19.56 45.564 21 ;
      RECT 45.158 13.8 45.742 19.56 ;
      RECT 45.158 12.36 45.564 13.8 ;
      RECT 45.158 11.64 45.742 12.36 ;
      RECT 44.258 28.92 44.842 29.76 ;
      RECT 44.258 27.48 44.752 28.92 ;
      RECT 44.258 26.76 44.842 27.48 ;
      RECT 44.258 25.32 44.664 26.76 ;
      RECT 44.258 24.6 44.842 25.32 ;
      RECT 44.258 23.16 44.408 24.6 ;
      RECT 44.258 22.44 44.842 23.16 ;
      RECT 44.258 21 44.408 22.44 ;
      RECT 44.258 20.28 44.842 21 ;
      RECT 44.258 18.84 44.408 20.28 ;
      RECT 44.692 18.84 44.842 20.28 ;
      RECT 44.258 13.08 44.842 18.84 ;
      RECT 44.258 11.64 44.408 13.08 ;
      RECT 44.692 11.64 44.842 13.08 ;
      RECT 44.258 9.48 44.842 11.64 ;
      RECT 44.258 8.04 44.752 9.48 ;
      RECT 44.258 7.32 44.842 8.04 ;
      RECT 44.258 5.88 44.664 7.32 ;
      RECT 44.258 5.16 44.842 5.88 ;
      RECT 44.258 3.72 44.408 5.16 ;
      RECT 44.258 3 44.842 3.72 ;
      RECT 44.258 1.56 44.408 3 ;
      RECT 44.258 0 44.842 1.56 ;
      RECT 43.358 0 43.942 29.76 ;
      RECT 42.458 0 43.042 29.76 ;
      RECT 41.558 0 42.142 29.76 ;
      RECT 40.658 0 41.242 29.76 ;
      RECT 39.758 0 40.342 29.76 ;
      RECT 38.858 0 39.442 29.76 ;
      RECT 37.958 0 38.542 29.76 ;
      RECT 37.058 0 37.642 29.76 ;
      RECT 36.158 0 36.742 29.76 ;
      RECT 35.258 18 35.842 29.76 ;
      RECT 35.436 16.56 35.842 18 ;
      RECT 35.258 16.08 35.842 16.56 ;
      RECT 35.436 14.64 35.842 16.08 ;
      RECT 35.258 0 35.842 14.64 ;
      RECT 34.358 19.92 34.942 29.76 ;
      RECT 33.458 18 34.042 29.76 ;
      RECT 33.458 16.56 33.608 18 ;
      RECT 33.458 16.08 34.042 16.56 ;
      RECT 33.458 14.64 33.608 16.08 ;
      RECT 33.458 14.16 34.042 14.64 ;
      RECT 33.458 12.72 33.608 14.16 ;
      RECT 33.458 0 34.042 12.72 ;
      RECT 32.558 0 33.142 29.76 ;
      RECT 31.658 0 32.242 29.76 ;
      RECT 30.758 0 31.342 29.76 ;
      RECT 29.858 0 30.442 29.76 ;
      RECT 28.958 0 29.542 29.76 ;
      RECT 28.058 0 28.642 29.76 ;
      RECT 27.158 0 27.742 29.76 ;
      RECT 26.258 0 26.842 29.76 ;
      RECT 25.358 0 25.942 29.76 ;
      RECT 24.458 0 25.042 29.76 ;
      RECT 23.558 0 24.142 29.76 ;
      RECT 22.658 0 23.242 29.76 ;
      RECT 21.758 0 22.342 29.76 ;
      RECT 20.858 0 21.442 29.76 ;
      RECT 19.958 0 20.542 29.76 ;
      RECT 19.058 0 19.642 29.76 ;
      RECT 18.158 0 18.742 29.76 ;
      RECT 17.258 0 17.842 29.76 ;
      RECT 16.358 0 16.942 29.76 ;
      RECT 15.458 0 16.042 29.76 ;
      RECT 14.558 28.92 15.142 29.76 ;
      RECT 14.736 27.48 15.142 28.92 ;
      RECT 14.558 26.76 15.142 27.48 ;
      RECT 14.736 25.32 15.142 26.76 ;
      RECT 14.558 24.6 15.142 25.32 ;
      RECT 14.736 23.16 15.142 24.6 ;
      RECT 14.558 11.64 15.142 23.16 ;
      RECT 14.736 10.2 15.142 11.64 ;
      RECT 14.558 9.48 15.142 10.2 ;
      RECT 14.736 8.04 15.142 9.48 ;
      RECT 14.558 7.32 15.142 8.04 ;
      RECT 14.736 5.88 15.142 7.32 ;
      RECT 14.558 5.16 15.142 5.88 ;
      RECT 14.648 3.72 15.142 5.16 ;
      RECT 14.558 0 15.142 3.72 ;
      RECT 13.658 28.2 14.242 29.76 ;
      RECT 13.748 26.76 14.242 28.2 ;
      RECT 13.658 25.32 14.152 26.76 ;
      RECT 13.658 24.6 14.242 25.32 ;
      RECT 13.658 23.16 14.064 24.6 ;
      RECT 13.658 22.44 14.242 23.16 ;
      RECT 12.758 28.2 13.342 29.76 ;
      RECT 12.758 26.76 12.908 28.2 ;
      RECT 12.758 26.04 13.342 26.76 ;
      RECT 11.858 29.64 12.442 29.76 ;
      RECT 12.036 28.2 12.442 29.64 ;
      RECT 11.858 21.72 12.442 28.2 ;
      RECT 11.858 20.28 12.264 21.72 ;
      RECT 11.858 19.56 12.442 20.28 ;
      RECT 11.948 18.12 12.442 19.56 ;
      RECT 11.858 14.52 12.442 18.12 ;
      RECT 11.858 13.08 12.264 14.52 ;
      RECT 11.858 12.36 12.442 13.08 ;
      RECT 10.958 29.64 11.542 29.76 ;
      RECT 10.958 28.2 11.364 29.64 ;
      RECT 10.958 27.48 11.542 28.2 ;
      RECT 10.058 28.92 10.642 29.76 ;
      RECT 10.236 27.48 10.642 28.92 ;
      RECT 10.058 26.76 10.642 27.48 ;
      RECT 10.148 25.32 10.642 26.76 ;
      RECT 10.058 23.88 10.552 25.32 ;
      RECT 10.058 23.16 10.642 23.88 ;
      RECT 10.058 21.72 10.464 23.16 ;
      RECT 10.058 21 10.642 21.72 ;
      RECT 9.158 0 9.742 29.76 ;
      RECT 8.258 0 8.842 29.76 ;
      RECT 7.358 0 7.942 29.76 ;
      RECT 6.458 0 7.042 29.76 ;
      RECT 5.558 0 6.142 29.76 ;
      RECT 4.658 0 5.242 29.76 ;
      RECT 3.758 0 4.342 29.76 ;
      RECT 2.858 0 3.442 29.76 ;
      RECT 1.958 0 2.542 29.76 ;
      RECT 1.058 0 1.642 29.76 ;
      RECT 0.08 0 0.742 29.76 ;
      RECT 46.958 27.48 47.542 28.2 ;
      RECT 46.958 25.32 47.542 26.04 ;
      RECT 47.392 23.88 47.542 25.32 ;
      RECT 46.958 23.16 47.542 23.88 ;
      RECT 47.048 21.72 47.542 23.16 ;
      RECT 46.958 20.28 47.452 21.72 ;
      RECT 46.958 19.56 47.542 20.28 ;
      RECT 47.136 18.12 47.542 19.56 ;
      RECT 46.958 14.52 47.542 18.12 ;
      RECT 46.958 13.08 47.452 14.52 ;
      RECT 46.958 12.36 47.542 13.08 ;
      RECT 46.958 10.92 47.108 12.36 ;
      RECT 46.958 10.2 47.542 10.92 ;
      RECT 10.958 25.32 11.542 26.04 ;
      RECT 11.392 23.88 11.542 25.32 ;
      RECT 10.958 23.16 11.542 23.88 ;
      RECT 11.136 21.72 11.542 23.16 ;
      RECT 10.958 19.56 11.542 21.72 ;
      RECT 10.958 18.12 11.108 19.56 ;
      RECT 10.958 10.2 11.542 18.12 ;
      RECT 10.958 8.76 11.364 10.2 ;
      RECT 10.958 8.04 11.542 8.76 ;
      RECT 12.758 23.88 13.342 24.6 ;
      RECT 47.858 21.72 48.442 22.44 ;
      RECT 48.292 20.28 48.442 21.72 ;
      RECT 47.858 14.52 48.442 20.28 ;
      RECT 48.292 13.08 48.442 14.52 ;
      RECT 47.858 12.36 48.442 13.08 ;
      RECT 47.948 10.92 48.442 12.36 ;
      RECT 47.858 9.48 48.352 10.92 ;
      RECT 47.858 8.76 48.442 9.48 ;
      RECT 47.858 7.32 48.264 8.76 ;
      RECT 47.858 6.6 48.442 7.32 ;
      RECT 47.858 5.16 48.008 6.6 ;
      RECT 47.858 4.44 48.442 5.16 ;
      RECT 12.758 21.72 13.342 22.44 ;
      RECT 12.936 20.28 13.342 21.72 ;
      RECT 12.758 18.84 13.252 20.28 ;
      RECT 12.758 14.52 13.342 18.84 ;
      RECT 12.936 13.08 13.342 14.52 ;
      RECT 12.758 11.64 13.252 13.08 ;
      RECT 12.758 10.92 13.342 11.64 ;
      RECT 12.758 9.48 13.164 10.92 ;
      RECT 12.758 8.76 13.342 9.48 ;
      RECT 12.758 7.32 12.908 8.76 ;
      RECT 12.758 6.6 13.342 7.32 ;
      RECT 13.658 20.28 14.242 21 ;
      RECT 14.092 18.84 14.242 20.28 ;
      RECT 13.658 13.08 14.242 18.84 ;
      RECT 14.092 11.64 14.242 13.08 ;
      RECT 13.658 10.92 14.242 11.64 ;
      RECT 13.836 9.48 14.242 10.92 ;
      RECT 13.658 8.76 14.242 9.48 ;
      RECT 13.748 7.32 14.242 8.76 ;
      RECT 13.658 5.88 14.152 7.32 ;
      RECT 13.658 5.16 14.242 5.88 ;
      RECT 13.658 3.72 13.808 5.16 ;
      RECT 13.658 3 14.242 3.72 ;
      RECT 10.058 13.8 10.642 19.56 ;
      RECT 34.358 18 34.942 18.48 ;
      RECT 34.358 16.08 34.942 16.56 ;
      RECT 34.358 14.16 34.942 14.64 ;
      RECT 34.448 12.72 34.942 14.16 ;
      RECT 34.358 0 34.942 12.72 ;
      RECT 10.058 11.64 10.642 12.36 ;
      RECT 10.492 10.2 10.642 11.64 ;
      RECT 10.058 9.48 10.642 10.2 ;
      RECT 10.236 8.04 10.642 9.48 ;
      RECT 10.058 7.32 10.642 8.04 ;
      RECT 10.148 5.88 10.642 7.32 ;
      RECT 10.058 4.44 10.552 5.88 ;
      RECT 10.058 3.72 10.642 4.44 ;
      RECT 10.058 2.28 10.208 3.72 ;
      RECT 10.058 1.56 10.642 2.28 ;
      RECT 11.858 10.2 12.442 10.92 ;
      RECT 12.036 8.76 12.442 10.2 ;
      RECT 11.858 4.44 12.442 8.76 ;
      RECT 11.858 3 12.352 4.44 ;
      RECT 11.858 2.28 12.442 3 ;
      RECT 11.858 0.84 12.008 2.28 ;
      RECT 11.858 0 12.442 0.84 ;
      RECT 45.158 9.48 45.742 10.2 ;
      RECT 45.592 8.04 45.742 9.48 ;
      RECT 45.158 7.32 45.742 8.04 ;
      RECT 45.336 5.88 45.742 7.32 ;
      RECT 45.158 5.16 45.742 5.88 ;
      RECT 45.248 3.72 45.742 5.16 ;
      RECT 45.158 1.56 45.742 3.72 ;
      RECT 46.958 8.04 47.542 8.76 ;
      RECT 46.958 5.88 47.542 6.6 ;
      RECT 47.392 4.44 47.542 5.88 ;
      RECT 46.958 2.28 47.542 4.44 ;
      RECT 46.958 0.84 47.364 2.28 ;
      RECT 46.958 0 47.542 0.84 ;
      RECT 10.958 5.88 11.542 6.6 ;
      RECT 11.392 4.44 11.542 5.88 ;
      RECT 10.958 3.72 11.542 4.44 ;
      RECT 11.048 2.28 11.542 3.72 ;
      RECT 10.958 0 11.542 2.28 ;
      RECT 12.758 4.44 13.342 5.16 ;
      RECT 13.192 3 13.342 4.44 ;
      RECT 12.758 2.28 13.342 3 ;
      RECT 12.848 0.84 13.342 2.28 ;
      RECT 12.758 0 13.342 0.84 ;
      RECT 47.858 2.28 48.442 3 ;
      RECT 48.036 0.84 48.442 2.28 ;
      RECT 47.858 0 48.442 0.84 ;
      RECT 46.058 0 46.642 2.28 ;
      RECT 13.658 0 14.242 1.56 ;
      RECT 45.158 0 45.742 0.12 ;
      RECT 10.058 0 10.642 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 70.2 29.758 ;
    LAYER m1 ;
      RECT 0 0 70.2 29.76 ;
    LAYER m2 ;
      RECT 0 0.015 70.2 29.745 ;
    LAYER m3 ;
      RECT 0.015 0 70.185 29.76 ;
    LAYER m4 ;
      RECT 0 0.02 70.2 29.74 ;
    LAYER m5 ;
      RECT 0.012 0 70.188 29.76 ;
    LAYER m6 ;
      RECT 0 0.012 70.2 29.748 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf132b192e1r1w0cbbehcaa4acw

END LIBRARY
