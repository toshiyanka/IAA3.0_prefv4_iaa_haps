//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// These are the global parameters for the IOSF SideBand EndPoint that are ported to the top.
//-----------------------------------------------------------------------------------------------------

         parameter SBE_DATAWIDTH                = 8
        ,parameter SBE_NPQUEUEDEPTH             = 4
        ,parameter SBE_PCQUEUEDEPTH             = 4
        ,parameter SBE_ASYNCIQDEPTH             = 2
        ,parameter SBE_ASYNCEQDEPTH             = 2
        ,parameter SBE_PIPEISMS                 = 0
        ,parameter SBE_PIPEINPS                 = 0
        ,parameter SBE_CLKREQ_HYST_CNT          = 15
        ,parameter SBE_PARITY_REQUIRED          = 1
        ,parameter SBE_DO_SERR_MASTER           = 1

