`topo_picker_class_begin(rcfwl_picker, RCFWL )

`run_knobs_begin
 `run_knobs_end

  
 
`picker_class_end
