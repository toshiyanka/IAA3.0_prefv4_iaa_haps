//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/fpv_sbr/fpv_sbr.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr
(
  // Synchronous Clock/Reset
  clk,
  rstb,

  // Power Well Isolation Input Signals
  pd1_pwrgd,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_clk,
  visa_vp_clk,
  visa_p0_tier1_clk,
  visa_p0_tier2_clk,
  visa_p1_tier1_clk,
  visa_p1_tier2_clk,


  // DFx signals
  fscan_latchopen,
  fscan_latchclosed_b,
  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  ep0_sbr_side_ism_agent,
  sbr_ep0_side_ism_fabric,
  ep0_sbr_pccup,
  ep0_sbr_npcup,
  sbr_ep0_pcput,
  sbr_ep0_npput,
  sbr_ep0_eom,
  sbr_ep0_payload,
  sbr_ep0_pccup,
  sbr_ep0_npcup,
  ep0_sbr_pcput,
  ep0_sbr_npput,
  ep0_sbr_eom,
  ep0_sbr_payload,

  // Port 1 declarations
  ep1_sbr_side_ism_agent,
  sbr_ep1_side_ism_fabric,
  ep1_sbr_pccup,
  ep1_sbr_npcup,
  sbr_ep1_pcput,
  sbr_ep1_npput,
  sbr_ep1_eom,
  sbr_ep1_payload,
  sbr_ep1_pccup,
  sbr_ep1_npcup,
  ep1_sbr_pcput,
  ep1_sbr_npput,
  ep1_sbr_eom,
  ep1_sbr_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic clk;
  input logic rstb;

  // Power Well Isolation Input Signals
  input logic pd1_pwrgd;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_clk;
  output visa_vp  visa_vp_clk;
  output visa_port_tier1 visa_p0_tier1_clk;
  output visa_port_tier2 visa_p0_tier2_clk;
  output visa_port_tier1 visa_p1_tier1_clk;
  output visa_port_tier2 visa_p1_tier2_clk;

  // DFx signals
  input logic fscan_latchopen;
  input logic fscan_latchclosed_b;
  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic fscan_rstbypen;
  input logic fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] ep0_sbr_side_ism_agent;
  output logic [2:0] sbr_ep0_side_ism_fabric;
  input logic ep0_sbr_pccup;
  input logic ep0_sbr_npcup;
  output logic sbr_ep0_pcput;
  output logic sbr_ep0_npput;
  output logic sbr_ep0_eom;
  output logic [7:0] sbr_ep0_payload;
  output logic sbr_ep0_pccup;
  output logic sbr_ep0_npcup;
  input logic ep0_sbr_pcput;
  input logic ep0_sbr_npput;
  input logic ep0_sbr_eom;
  input logic [7:0] ep0_sbr_payload;

  // Port 1 declarations
  input logic [2:0] ep1_sbr_side_ism_agent;
  output logic [2:0] sbr_ep1_side_ism_fabric;
  input logic ep1_sbr_pccup;
  input logic ep1_sbr_npcup;
  output logic sbr_ep1_pcput;
  output logic sbr_ep1_npput;
  output logic sbr_ep1_eom;
  output logic [7:0] sbr_ep1_payload;
  output logic sbr_ep1_pccup;
  output logic sbr_ep1_npcup;
  input logic ep1_sbr_pcput;
  input logic ep1_sbr_npput;
  input logic ep1_sbr_eom;
  input logic [7:0] ep1_sbr_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_sbcportmap;
always_comb sbr_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr (sbr)                                     SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  250 { 17'b0_0000_0000_0000_0000 }},   //   254:  5      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //     4          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     3:  2      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //     1          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000       //     0          SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  1;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              pd1_pwrgd_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = '1;
always_comb cfg_clkgatedef    = '0;
always_comb cfg_idlecnt       = 8'h10;
always_comb jta_clkgate_ovrd  = '0;
always_comb jta_force_idle    = '0;
always_comb jta_force_notidle = '0;
always_comb jta_force_creditreq = '0;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_creditreq               )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_pd1_pwrgd (
  .d                   ( pd1_pwrgd                     ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( pd1_pwrgd_ff2                 )
);


always_comb endpoint_pwrgd = { pd1_pwrgd_ff2,
                          1'b1
                        };

logic p1_gated_clk;
sbc_clock_gate p1_pwr_clkgate  (
  .en ( endpoint_pwrgd[1] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p1_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
// SBR_IDLE signal for PMU
  logic [1:0] idle_suppress; // delay idle assertion till after power state is synchronized out of reset.

  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
       idle_suppress <= '0;
    else
       idle_suppress <= {idle_suppress[0], 1'b1};

  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      sbr_idle <= '0;
    else
      sbr_idle <= (&idle_suppress) & arbiter_idle & all_idle &
                  p0_ism_idle & ~p0_fab_init_idle_exit &
                  p1_ism_idle & ~p1_fab_init_idle_exit;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_clk = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk                           ),
  .side_rst_b          ( rstb                          ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_clk = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p0_fab_init_idle_exit <= '0;
    else
      if (~endpoint_pwrgd[0])
         p0_fab_init_idle_exit <= '0;
      else
         begin
          if ( p0_rst_suppress | (~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack )))
            p0_fab_init_idle_exit <= '1;
          else if ( p0_fab_init_idle_exit_ack & (~p0_rst_suppress & p0_ism_idle & agent_idle[0] ))
            p0_fab_init_idle_exit <= '0;
         end

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( (p0_ism_idle & p0_side_clk_valid) | ~endpoint_pwrgd[0] )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_clk = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_clk = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport0 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( ep0_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep0_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_ep0_pccup                 ),
  .tnpcup              ( sbr_ep0_npcup                 ),
  .tpcput              ( ep0_sbr_pcput                 ),
  .tnpput              ( ep0_sbr_npput                 ),
  .teom                ( ep0_sbr_eom                   ),
  .tpayload            ( ep0_sbr_payload               ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( ep0_sbr_pccup                 ),
  .mnpcup              ( ep0_sbr_npcup                 ),
  .mpcput              ( sbr_ep0_pcput                 ),
  .mnpput              ( sbr_ep0_npput                 ),
  .meom                ( sbr_ep0_eom                   ),
  .mpayload            ( sbr_ep0_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit & p1_rst_suppress;

  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p1_fab_init_idle_exit <= '0;
    else
      if (~endpoint_pwrgd[1])
         p1_fab_init_idle_exit <= '0;
      else
         begin
          if ( p1_rst_suppress | (~p1_rst_suppress & (p1_ism_idle & (~agent_idle[1] || ~p1_idle_egress) & ~p1_fab_init_idle_exit_ack )))
            p1_fab_init_idle_exit <= '1;
          else if ( p1_fab_init_idle_exit_ack & (~p1_rst_suppress & p1_ism_idle & agent_idle[1] ))
            p1_fab_init_idle_exit <= '0;
         end

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( (p1_ism_idle & p1_side_clk_valid) | ~endpoint_pwrgd[1] )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle )
          p1_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

  always_comb
    begin
      visa_p1_tier1_clk = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_clk = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport1 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( ep1_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep1_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .idle_egress         ( p1_idle_egress                ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_ep1_pccup                 ),
  .tnpcup              ( sbr_ep1_npcup                 ),
  .tpcput              ( ep1_sbr_pcput                 ),
  .tnpput              ( ep1_sbr_npput                 ),
  .teom                ( ep1_sbr_eom                   ),
  .tpayload            ( ep1_sbr_payload               ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( ep1_sbr_pccup                 ),
  .mnpcup              ( ep1_sbr_npcup                 ),
  .mpcput              ( sbr_ep1_pcput                 ),
  .mnpput              ( sbr_ep1_npput                 ),
  .meom                ( sbr_ep1_eom                   ),
  .mpayload            ( sbr_ep1_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk or negedge rstb)

      if (~rstb) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (rstb !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (rstb !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/fpv_sbr/fpv_sbr.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 0, clk, rstb, 0, , 1ns
Endpoint, ep0,0, 1, 0, 1, 3, 3, 1, 1, 1, 1, 
Endpoint, ep1,1, 1, 0, 1, 3, 3, 1, 4, 2, 2, 
SyncRouter, sbr, sbr,0, 1, 0, 3, 4, 4, 0, 1, , , 0, 2, ep0, ep1, , , , , , , , , , , , , , , 
PowerWell, 0, 
PowerWell, 1, pd1_pwrgd
*/
//------------------------------------------------------------------------------
