`ifndef HQM_TESTS__PKG
`define HQM_TESTS__PKG

package hqm_tests_pkg;

  `include "vip_layering_macros.svh"

  `import_base(ovm_pkg::*)
  `include_base("ovm_macros.svh")

  `import_base(sla_pkg::*)
  `include_base("sla_macros.svh")


  import hqm_saola_pkg::*;
  `import_mid(pcie_seqlib_pkg::*)
  `import_mid(hqm_tb_test_sequences_pkg::*)

  //-- test base
  `include_typ("hqm_base_test.sv")  //--`include_mid
  `include_typ("hqm_pwr_base_test.sv")
  `include_typ("hqm_iosf_base_test.sv")
  `include_typ("hqm_pcie_tests_list.sv")
  `include_typ("hqm_sciov_tests_list.sv")
  `include_typ("hqm_pcie_error_test.sv")
  `include_typ("hqm_pcie_interrupt_test.sv")
  `include_typ("hqm_iosf_sideband_file_test.sv")
  `include_typ("hqm_iosf_sideband_file_test.svh")
  `include_typ("hqm_iosf_prim_pf_dump_test.sv")
  `include_typ("hqm_iosf_prim_file_test.svh")
  `include_typ("hqm_base_iosf_test.sv")
  `include_typ("hqm_check_test.sv")
  //`include_typ("back2back_cfgrd_check_seq.sv")
  `include_typ("cfg_generic_test.svh")
  `include_typ("reset_test.sv")
  `include_typ("reset_test.svh")
  `include_typ("cfg_generic_test.sv")
  `include_typ("mem_generic_test.svh")
  `include_typ("mem_generic_test.sv")
  `include_typ("cfg_error_test.svh")
  `include_typ("cfg_error_test.sv")
  `include_typ("mem_error_test.svh")
  `include_typ("mem_error_test.sv")
  `include_typ("SAI_test.svh")
  `include_typ("SAI_test.sv")
  `include_typ("BE_test.svh")
  `include_typ("BE_test.sv")
  `include_typ("cpl_test.svh")
  `include_typ("cpl_test.sv")
  `include_typ("hqm_iosf_tb_file_test.sv")
  `include_typ("hqm_iosf_tb_file_test.svh")
  `include_typ("unsupport_cmd_test.svh")
  `include_typ("unsupport_cmd_test.sv")
  `include_typ("unsupport_cmd_sai_test.svh")
  `include_typ("unsupport_cmd_sai_test.sv")
  `include_typ("hqm_iosf_sideband_test.svh")
  `include_typ("hqm_iosf_sideband_test.sv")
  `include_typ("hqm_iosf_sideband_UC_test.svh")
  `include_typ("hqm_iosf_sideband_UC_test.sv")
  `include_typ("hqm_error_test.svh")
  `include_typ("hqm_error_test.sv")
  `include_typ("iosf_cg_test.svh")
  `include_typ("iosf_cg_test.sv")
  `include_typ("sideband_crdinit_test.svh")
  `include_typ("sideband_crdinit_test.sv")
  `include_typ("hqm_newTR_test.svh")
  `include_typ("hqm_newTR_test.sv")
  `include_typ("sb_error_test.svh")
  `include_typ("sb_error_test.sv")
  `include_typ("hqm_top_test.svh")
  `include_typ("hqm_top_test.sv")
  `include_typ("mix_test.svh")
  `include_typ("mix_test.sv")

   // new IOSF test implementation
  `include_typ("hqm_iosf_test.svh") 

  `include_typ("hqm_sb_test.sv") 
  `include_typ("hqm_prim_n_sb_error_test.sv") 
  `include_typ("hqm_ldb_qos_test.svh")
  `include_typ("hqm_arb_pri_test.svh")
  `include_typ("hqm_trf_test.svh")
  `include_typ("hqm_iosf_sb_file_test.svh")
  `include_typ("hqm_cfg_test.svh")
  `include_typ("hqm_raw_test.svh")
  `include_typ("hqm_idle_test.svh")
  `include_typ("hqm_pok_test.svh")
  `include_typ("hqm_system_burst_test.svh")
  `include_typ("hqm_system_error_burst_test/hqm_system_error_burst_test.svh")
  `include_typ("hqm_unimp_addr_test.svh")
  `include_typ("hqm_pfvf_space_acc_test.svh")
  `include_typ("hcw_pipeline_stress_test.svh")
  `include_typ("hqm_strap_chk_test.svh")
  `include_typ("hqm_mra_connect_chk_test.svh")
  `include_typ("hqm_pcie_msg_test.svh")
  `include_typ("hqm_survivability_test.svh")
  `include_typ("hcw_perf_test1.svh")
  `include_typ("hcw_perf_dir_test1.svh")
  `include_typ("hcw_dir_test.svh")
  `include_typ("hqm_ral_cfg_test.sv")
  `include_typ("hcw_ldb_test.sv")
  `include_typ("hcw_dir_traffic_test.sv")
  `include_typ("hcw_ldb_traffic_test.sv")
  `include_typ("hcw_perf_ldb_test1.svh")
  `include_typ("hcw_perf_atm_test.svh")
  `include_typ("hcw_perf_dir_ldb_test1.svh")
  `include_typ("hcw_perf_dir_ldb_test1_agi.svh")
  `include_typ("hcw_perf_dir_ldb_pkgc_vret_test.svh")
  `include_typ("hcw_sciov_test.svh")
  `include_typ("hcw_sciov_test2.svh")
  `include_typ("hcw_pf_test.svh") //--`include_mid
  `include_typ("hqmv30_pf_test.svh") 
  `include_typ("hqmv30_sciov_test.svh") 
  `include_typ("hcw_pf_vf_test.svh")
  `include_typ("hqm_hdr_log_cov_test.svh")
  `include_typ("hcw_processing_with_intermediate_flr_test.svh")
  `include_typ("hqm_cfg_with_intermediate_flr_test.svh")
  `include_typ("hqm_cfg_with_intermediate_primrst_test.svh")
  `include_typ("hcw_ingress_check_test.svh")
  `include_typ("hcw_ingress_token_error_test.svh")
  `include_typ("hcw_test0.svh")
  `include_typ("hcw_test1.svh")
  `include_typ("hcw_ldb_test1.svh")
  `include_typ("hqm_cfg_iosf_test.svh")
  `include_typ("hqm_reg_test.svh")
  `include_typ("hqm_reg_aliasing_test.svh")
  `include_typ("hqm_async_prim_rst_test.svh")
  `include_typ("hqm_visa_test.svh")
  `include_typ("hqm_pwr_test.svh")
  `include_typ("hqm_pcie_header_sweep_test.svh")
  `include_typ("cq_dead_wd_timer.svh")
  `include_typ("hqm_fuse_load_test.sv")
  `include_typ("hqm_trigger_test.sv")
  `include_typ("hqm_hvm_test.svh")
  `include_typ("hcw_enqtrf_hqmproc_test.svh")
  `include_typ("hcw_hqmproc_test.svh")
  `include_typ("hqm_config_master_test.svh")

  `include_typ("hqm_reset_cycle_test.sv")
  `include_typ("hcw_d0_d3_d0_test.svh")
  `include_typ("hqm_tap_rtdr_test.svh")

endpackage
`endif
