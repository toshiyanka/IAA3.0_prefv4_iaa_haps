module ctech_lib_tieoff_1 (out);
    output logic out;
   d04rid11nnz00 ctech_lib_dcszo (.o(out));
endmodule
