`ifdef EP_CFG0
`include "cfg0"
`endif
`ifdef EP_CFG1
`include "cfg1"
`endif
`ifdef EP_CFG2
`include "cfg2"
`endif
`ifdef EP_CFG3
`include "cfg3"
`endif
`ifdef EP_CFG4
`include "cfg4"
`endif
`ifdef EP_CFG5
`include "cfg5"
`endif
`ifdef EP_CFG6
`include "cfg6"
`endif
`ifdef EP_CFG7
`include "cfg7"
`endif
`ifdef EP_CFG8
`include "cfg8"
`endif
`ifdef EP_CFG9
`include "cfg9"
`endif
`ifdef EP_CFG10
`include "cfg10"
`endif
`ifdef EP_CFG11
`include "cfg11"
`endif
`ifdef EP_CFG12
`include "cfg12"
`endif
`ifdef EP_CFG13
`include "cfg13"
`endif
`ifdef EP_CFG14
`include "cfg14"
`endif
`ifdef EP_CFG15
`include "cfg15"
`endif
`ifdef EP_CFG16
`include "cfg16"
`endif
`ifdef EP_CFG17
`include "cfg17"
`endif
`ifdef EP_CFG18
`include "cfg18"
`endif
`ifdef EP_CFG19
`include "cfg19"
`endif
`ifdef EP_CFG20
`include "cfg20"
`endif
`ifdef EP_CFG21
`include "cfg21"
`endif
`ifdef EP_CFG22
`include "cfg22"
`endif
`ifdef EP_CFG23
`include "cfg23"
`endif
`ifdef EP_CFG24
`include "cfg24"
`endif
`ifdef EP_CFG25
`include "cfg25"
`endif
`ifdef EP_CFG26
`include "cfg26"
`endif
`ifdef EP_CFG27
`include "cfg27"
`endif
`ifdef EP_CFG28
`include "cfg28"
`endif
`ifdef EP_CFG29
`include "cfg29"
`endif
`ifdef EP_CFG30
`include "cfg30"
`endif
`ifdef EP_CFG31
`include "cfg31"
`endif
`ifdef EP_CFG32
`include "cfg32"
`endif
`ifdef EP_CFG33
`include "cfg33"
`endif
`ifdef EP_CFG34
`include "cfg34"
`endif
`ifdef EP_CFG35
`include "cfg35"
`endif
`ifdef EP_CFG36
`include "cfg36"
`endif
`ifdef EP_CFG37
`include "cfg37"
`endif
`ifdef EP_CFG38
`include "cfg38"
`endif
`ifdef EP_CFG39
`include "cfg39"
`endif
`ifdef EP_CFG40
`include "cfg40"
`endif
`ifdef EP_CFG41
`include "cfg41"
`endif
`ifdef EP_CFG42
`include "cfg42"
`endif
`ifdef EP_CFG43
`include "cfg43"
`endif
`ifdef EP_CFG44
`include "cfg44"
`endif
`ifdef EP_CFG45
`include "cfg45"
`endif
`ifdef EP_CFG46
`include "cfg46"
`endif
