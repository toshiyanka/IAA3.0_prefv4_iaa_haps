parameter NUMBER_OF_HIER  = 10;
parameter NUMBER_OF_STAPS  = 14;
parameter NUMBER_OF_TERTIARY_PORTS = 0;
