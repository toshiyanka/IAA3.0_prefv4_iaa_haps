package hqm_tap_rtdr_common_val_tb_pkg;

`include "ovm_macros.svh"
`include "sla_macros.svh"

import ovm_pkg::*;
import sla_pkg::*;

// DFT TB class includes here
/////////////////////////////////////////////////
`include "hqm_tap_rtdr_common_val_sim_component.svh"

endpackage : hqm_tap_rtdr_common_val_tb_pkg
