module ctech_lib_latch (clk, d, o);
  input logic clk, d;
  output logic o;
   d04ltn00ld0b0 ctech_lib_dcszo (.clk(clk),.d(d),.o(o));
endmodule
