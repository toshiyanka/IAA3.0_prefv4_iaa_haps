module ctech_lib_dq (
   input logic a,
   input logic b,
   output logic o
);
   d04ann02ln0b0 ctech_lib_dcszo (.a(a), .b(b), .o(o));
endmodule
