VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf066b128e2r1w0cbbehsaa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf066b128e2r1w0cbbehsaa4acw 0 0 ;
  SIZE 45 BY 22.08 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 11.16 0.388 12.36 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 11.16 4.156 12.36 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 9 0.388 10.2 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 11.16 1.928 12.36 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 11.16 2.188 12.36 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 11.16 2.356 12.36 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 11.16 2.616 12.36 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 11.16 2.916 12.36 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 11.16 3.172 12.36 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 11.16 3.988 12.36 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 11.16 0.556 12.36 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 11.16 0.816 12.36 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 11.16 5.528 12.36 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 11.16 5.788 12.36 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 11.16 5.956 12.36 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 11.16 6.216 12.36 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 11.16 6.516 12.36 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 11.16 0.472 12.36 ;
    END
  END rdaddrp1[5]
  PIN rdaddrp1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 11.16 0.728 12.36 ;
    END
  END rdaddrp1[6]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 11.16 4.416 12.36 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 11.16 4.716 12.36 ;
    END
  END rdaddrp1_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 0.12 3.256 1.32 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 2.52 4.716 3.72 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 2.52 4.888 3.72 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 3 3.988 4.2 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 3 4.072 4.2 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 3.48 5.228 4.68 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 3.48 5.316 4.68 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 3.96 3.428 5.16 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.96 3.516 5.16 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 4.44 4.716 5.64 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 4.44 4.888 5.64 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.12 3.428 1.32 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 4.92 3.988 6.12 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 4.92 4.072 6.12 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 5.4 5.228 6.6 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 5.4 5.316 6.6 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 5.88 3.428 7.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.88 3.516 7.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 6.36 4.716 7.56 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 6.36 4.888 7.56 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 6.84 3.988 8.04 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.84 4.072 8.04 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 0.6 4.628 1.8 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 7.32 5.228 8.52 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 7.32 5.316 8.52 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 7.8 3.428 9 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.8 3.516 9 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 13.08 4.072 14.28 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 13.08 4.328 14.28 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 13.56 3.516 14.76 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 13.56 3.728 14.76 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 14.04 5.228 15.24 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 14.04 5.316 15.24 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 0.6 4.716 1.8 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 14.52 3.428 15.72 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 14.52 3.988 15.72 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 15 4.716 16.2 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 15 4.888 16.2 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 15.48 3.516 16.68 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 15.48 3.728 16.68 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 15.96 5.228 17.16 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 15.96 5.316 17.16 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.44 3.428 17.64 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 16.44 3.988 17.64 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 1.08 3.988 2.28 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 16.92 4.716 18.12 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 16.92 4.888 18.12 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 17.4 3.516 18.6 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 17.4 3.728 18.6 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 17.88 5.228 19.08 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 17.88 5.316 19.08 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 18.36 3.428 19.56 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 18.36 3.988 19.56 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 18.84 4.716 20.04 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 18.84 4.888 20.04 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 1.08 4.072 2.28 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.32 3.516 20.52 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 19.32 3.728 20.52 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 19.8 5.228 21 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 19.8 5.316 21 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.28 3.428 21.48 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 20.28 3.988 21.48 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 20.76 4.716 21.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 20.76 4.888 21.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 1.56 5.228 2.76 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 1.56 5.316 2.76 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.04 3.428 3.24 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 2.04 3.516 3.24 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 0.12 3.516 1.32 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 2.52 4.972 3.72 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 2.52 5.056 3.72 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 3 4.156 4.2 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 3 4.328 4.2 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 3.48 5.528 4.68 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 3.48 5.616 4.68 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.96 3.728 5.16 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 3.96 3.816 5.16 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 4.44 4.972 5.64 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 4.44 5.056 5.64 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.12 3.728 1.32 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 4.92 4.156 6.12 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 4.92 4.328 6.12 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 5.4 5.528 6.6 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 5.4 5.616 6.6 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 5.88 3.728 7.08 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 5.88 3.816 7.08 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 6.36 4.972 7.56 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 6.36 5.056 7.56 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 6.84 4.156 8.04 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6.84 4.328 8.04 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 0.6 4.888 1.8 ;
    END
  END rddatap1[2]
  PIN rddatap1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 7.32 5.528 8.52 ;
    END
  END rddatap1[30]
  PIN rddatap1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 7.32 5.616 8.52 ;
    END
  END rddatap1[31]
  PIN rddatap1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 7.8 3.728 9 ;
    END
  END rddatap1[32]
  PIN rddatap1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 7.8 3.816 9 ;
    END
  END rddatap1[33]
  PIN rddatap1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 13.08 4.628 14.28 ;
    END
  END rddatap1[34]
  PIN rddatap1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 13.08 4.888 14.28 ;
    END
  END rddatap1[35]
  PIN rddatap1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 13.56 3.816 14.76 ;
    END
  END rddatap1[36]
  PIN rddatap1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 13.56 5.056 14.76 ;
    END
  END rddatap1[37]
  PIN rddatap1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 14.04 5.528 15.24 ;
    END
  END rddatap1[38]
  PIN rddatap1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 14.04 5.616 15.24 ;
    END
  END rddatap1[39]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 0.6 4.972 1.8 ;
    END
  END rddatap1[3]
  PIN rddatap1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 14.52 4.072 15.72 ;
    END
  END rddatap1[40]
  PIN rddatap1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 14.52 4.156 15.72 ;
    END
  END rddatap1[41]
  PIN rddatap1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 15 4.972 16.2 ;
    END
  END rddatap1[42]
  PIN rddatap1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 15 5.056 16.2 ;
    END
  END rddatap1[43]
  PIN rddatap1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 15.48 3.816 16.68 ;
    END
  END rddatap1[44]
  PIN rddatap1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 15.48 4.328 16.68 ;
    END
  END rddatap1[45]
  PIN rddatap1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 15.96 5.528 17.16 ;
    END
  END rddatap1[46]
  PIN rddatap1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 15.96 5.616 17.16 ;
    END
  END rddatap1[47]
  PIN rddatap1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.44 4.072 17.64 ;
    END
  END rddatap1[48]
  PIN rddatap1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 16.44 4.156 17.64 ;
    END
  END rddatap1[49]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 1.08 4.156 2.28 ;
    END
  END rddatap1[4]
  PIN rddatap1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 16.92 4.972 18.12 ;
    END
  END rddatap1[50]
  PIN rddatap1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 16.92 5.056 18.12 ;
    END
  END rddatap1[51]
  PIN rddatap1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 17.4 3.816 18.6 ;
    END
  END rddatap1[52]
  PIN rddatap1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 17.4 4.328 18.6 ;
    END
  END rddatap1[53]
  PIN rddatap1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 17.88 5.528 19.08 ;
    END
  END rddatap1[54]
  PIN rddatap1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 17.88 5.616 19.08 ;
    END
  END rddatap1[55]
  PIN rddatap1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 18.36 4.072 19.56 ;
    END
  END rddatap1[56]
  PIN rddatap1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 18.36 4.156 19.56 ;
    END
  END rddatap1[57]
  PIN rddatap1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 18.84 4.972 20.04 ;
    END
  END rddatap1[58]
  PIN rddatap1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 18.84 5.056 20.04 ;
    END
  END rddatap1[59]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 1.08 4.328 2.28 ;
    END
  END rddatap1[5]
  PIN rddatap1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 19.32 3.816 20.52 ;
    END
  END rddatap1[60]
  PIN rddatap1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 19.32 4.328 20.52 ;
    END
  END rddatap1[61]
  PIN rddatap1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 19.8 5.528 21 ;
    END
  END rddatap1[62]
  PIN rddatap1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 19.8 5.616 21 ;
    END
  END rddatap1[63]
  PIN rddatap1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 20.28 4.072 21.48 ;
    END
  END rddatap1[64]
  PIN rddatap1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 20.28 4.156 21.48 ;
    END
  END rddatap1[65]
  PIN rddatap1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 20.76 4.972 21.96 ;
    END
  END rddatap1[66]
  PIN rddatap1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.012 20.76 5.056 21.96 ;
    END
  END rddatap1[67]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 1.56 5.528 2.76 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 1.56 5.616 2.76 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 2.04 3.728 3.24 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 2.04 3.816 3.24 ;
    END
  END rddatap1[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 11.16 1.116 12.36 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 11.16 4.972 12.36 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 11.16 1.628 12.36 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 11.16 5.228 12.36 ;
    END
  END sdl_initp1
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 44.062 0.06 44.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 42.262 0.06 42.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 40.462 0.06 40.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 38.662 0.06 38.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 36.862 0.06 36.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.062 0.06 35.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 33.262 0.06 33.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.462 0.06 31.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.662 0.06 29.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 27.862 0.06 27.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.062 0.06 26.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.262 0.06 24.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 22.462 0.06 22.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.662 0.06 20.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.862 0.06 18.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.062 0.06 17.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.262 0.06 15.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 22.02 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 43.162 0.06 43.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 41.362 0.06 41.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 39.562 0.06 39.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 37.762 0.06 37.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.962 0.06 36.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 34.162 0.06 34.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 32.362 0.06 32.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.562 0.06 30.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 28.762 0.06 28.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.962 0.06 27.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.162 0.06 25.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.362 0.06 23.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 21.562 0.06 21.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 19.762 0.06 19.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.962 0.06 18.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 16.162 0.06 16.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.362 0.06 14.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 22.02 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 22.02 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 9 2.188 10.2 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 9 2.356 10.2 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 9 2.916 10.2 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 9 3.172 10.2 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 9 3.988 10.2 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 9 4.156 10.2 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 9 4.416 10.2 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 9 0.556 10.2 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 9 0.816 10.2 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.244 0.12 1.288 1.32 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 2.52 2.356 3.72 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.52 2.528 3.72 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 3 1.628 4.2 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 3 1.716 4.2 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.48 2.616 4.68 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 3.48 2.828 4.68 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 3.96 1.372 5.16 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 3.96 1.456 5.16 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 4.44 2.356 5.64 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 4.44 2.528 5.64 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 0.12 1.372 1.32 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 4.92 1.628 6.12 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 4.92 1.716 6.12 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.4 2.616 6.6 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.4 2.828 6.6 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 5.88 1.372 7.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 5.88 1.456 7.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 6.36 2.356 7.56 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6.36 2.528 7.56 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 6.84 1.628 8.04 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 6.84 1.716 8.04 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.6 2.272 1.8 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 7.32 2.616 8.52 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 7.32 2.828 8.52 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 7.8 1.372 9 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 7.8 1.456 9 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 13.08 2.828 14.28 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 13.08 1.716 14.28 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 13.56 1.372 14.76 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 13.56 1.456 14.76 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 14.04 2.528 15.24 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.04 2.616 15.24 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 0.6 2.356 1.8 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 14.52 1.628 15.72 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 14.52 1.716 15.72 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 15 2.356 16.2 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 15 2.828 16.2 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 15.48 1.372 16.68 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 15.48 1.456 16.68 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 15.96 2.528 17.16 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 15.96 2.616 17.16 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 16.44 1.628 17.64 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 16.44 1.716 17.64 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 1.08 1.628 2.28 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 16.92 2.356 18.12 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 16.92 2.828 18.12 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 17.4 1.372 18.6 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 17.4 1.456 18.6 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 17.88 2.528 19.08 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 17.88 2.616 19.08 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 18.36 1.628 19.56 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 18.36 1.716 19.56 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 18.84 2.356 20.04 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 18.84 2.828 20.04 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 1.08 1.716 2.28 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 19.32 1.372 20.52 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 19.32 1.456 20.52 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 19.8 2.528 21 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.8 2.616 21 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 20.28 1.628 21.48 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 20.28 1.716 21.48 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 20.76 2.356 21.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 20.76 2.828 21.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 1.56 2.616 2.76 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 1.56 2.828 2.76 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 2.04 1.372 3.24 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.412 2.04 1.456 3.24 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 9 1.628 10.2 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 9 1.928 10.2 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 9 1.116 10.2 ;
    END
  END wrenp0
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 45 22.08 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 45 22.08 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 45.0705 22.118 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 45.035 22.15 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 45.07 22.118 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 45.059 22.17 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 45.09 22.142 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 45.092 22.14 ;
  END
END arf066b128e2r1w0cbbehsaa4acw
END LIBRARY
