parameter NPQUEUEDEPTH=4; 
parameter PCQUEUEDEPTH=4;
parameter VALONLYMODEL=0; 
parameter MAXNPMSTR=0; 
parameter MAXPCMSTR=0; 
parameter MAXPCTRGT=0; 
parameter MAXNPTRGT=0;
parameter TARGETREG=1;
parameter MASTERREG=1;
parameter ASYNCEQDEPTH=32;
parameter ASYNCIQDEPTH=32;
parameter ASYNCENDPT=1;
parameter MAXTRGTADDR=31;
parameter MAXMSTRADDR=31;
parameter MAXMSTRDATA=63;
parameter MAXTRGTDATA=63;
parameter MAXPLDBIT=7;
parameter CUP2PUT1CYC=0;
parameter DUMMY_CLKBUF=0;
parameter TX_EXT_HEADER_SUPPORT=1;
parameter RX_EXT_HEADER_SUPPORT=1;
parameter NUM_RX_EXT_HEADERS=1;
parameter NUM_TX_EXT_HEADERS=1;
parameter RX_EXT_HEADER_IDS=7'h01;
parameter DISABLE_COMPLETION_FENCING=0;
parameter LATCHQUEUES=0;
parameter SKIP_ACTIVEREQ=1;
parameter AGT_CLK_PERIOD=0.7ns;
parameter FAB_CLK_PERIOD=1ns;
parameter PIPEISMS=0;
parameter PIPEINPS=0;
parameter USYNC_ENABLE = 1;
parameter IOSFSB_EP_SPEC_REV=1;
parameter IOSFSB_FBRC_SPEC_REV=1;
parameter AGT_EXT_HEADER_SUPPORT=1;
parameter FBRC_EXT_HEADER_SUPPORT=1;
