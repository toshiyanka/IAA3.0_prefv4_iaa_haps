  `include "hqm_pasid_disabled_test.sv"
  `include "hqm_pasid_enabled_test.sv"
  `include "hqm_addr_within_bar_chk_test.sv"
