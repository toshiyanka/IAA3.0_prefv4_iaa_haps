module dfxsecure_plugin_ctrl;

endmodule

