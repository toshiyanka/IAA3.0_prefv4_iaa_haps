// CCTypes begin

	typedef class PGCBAgent;
	typedef class PGCBAgentSequencer;
	typedef class PGCBAgentDriver;
	typedef class PGCBAgentSeqItem;
	typedef class PGCBAgentFabricResponder;
	typedef class PGCBAgentSIPResponder;

	typedef class PGCBAgentResponseSeqItem;
	typedef class PGCBAgentSIPFSM;
	typedef class PGCBAgentFabricFSM;
//	typedef class PGCBAgentAONFSM;

