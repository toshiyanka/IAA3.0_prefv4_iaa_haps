


	class ErrorPMCWakeTest extends PowerGatingBaseTest;
		SIPPMCWakeSequence sipPMCWake;
		SIPSWPGReqSequence sipSWPGReqSeq;

		SIPHWUGReqSequence sipHWUGReqSeq;
		SIPHWSaveReqSequence sipHWSaveReqSeq;
		DESIPPMCWakeSequence desipPMCWake;

		`ovm_component_utils(PowerGatingSaolaPkg::ErrorPMCWakeTest)
	
		function new(string name = "ErrorPMCWakeTest", ovm_component parent = null);
			super.new(name, parent);
		endfunction

		function void build();
			set_config_int("sla_env", "data_phase_mode", SLA_RANDOM_NONE );
			set_config_int("*", "count", 0);
			set_config_int("*","recording_detail", OVM_FULL);
	  		ovm_top.set_report_verbosity_level(OVM_FULL);   
			
			super.build();
		endfunction

		function void connect();
			super.connect();   
		endfunction  
  		task run();
			//exitIdleSeq = new();
			//enterIdleSeq = new();
			sipHWUGReqSeq = new();
			sipHWSaveReqSeq = new();
			sipSWPGReqSeq = new();
			sipPMCWake = new();
			desipPMCWake = new();

  			`ovm_info(get_type_name(),"RUNNING",OVM_LOW)
			#100us;
			//start test
			/*
1.	Wake up the SIP using PMC wake
2.	Make sure req and ack deassert
3.	Assert SW PG request
4.	Make sure req and ack assert
7.	Assert HW UG req
8.	Make sure req and ack assert
9.	Assert HW PG req
10.	Make sure req and ack deassert			
			*/
		   //PMC wake
		    sipPMCWake.start(sla_env.ccAgent.sequencer);
			wait(sla_env._vif.pmc_ip_pg_ack_b[0] == 1'b1);
			//desipPMCWake.start(sla_env.ccAgent.sequencer);		
			

			#100ns;
			//HW PG req
			//Aseert HW req and make sure an error is flagged
			sipHWSaveReqSeq.start(sla_env.pgcbAgent.sequencer);
			wait(sla_env._vif.pmc_ip_pg_ack_b[0] == 1'b0);
			

			#100us;
			global_stop_request();

  		endtask

		function void report();
			ovm_report_info("ErrorPMCWakeTest", "Test Passed!");
		endfunction

	endclass
	


		
