.DFX_NUM_OF_FEATURES_TO_SECURE         (STAP_DFX_NUM_OF_FEATURES_TO_SECURE),
.DFX_SECURE_WIDTH                      (STAP_DFX_SECURE_WIDTH),
.DFX_USE_SB_OVR                        (STAP_DFX_USE_SB_OVR),
.DFX_VISA_BLACK                        (STAP_DFX_VISA_BLACK),
.DFX_VISA_GREEN                        (STAP_DFX_VISA_GREEN),
.DFX_VISA_ORANGE                       (STAP_DFX_VISA_ORANGE),
.DFX_VISA_RED                          (STAP_DFX_VISA_RED),
.DFX_EARLYBOOT_FEATURE_ENABLE          (STAP_DFX_EARLYBOOT_FEATURE_ENABLE),
.DFX_SECURE_POLICY_MATRIX              (STAP_DFX_SECURE_POLICY_MATRIX)
