// File output was printed on: Saturday, January 19, 2013 2:59:29 PM
// Chassis TAP Tool version: 0.6.0.0
// ---------------------------------------------------- 
case (Node)
   'd0 : begin
            Tap_Info_Int.Next_Tap[0] = NOTAP;
        end
endcase


