interface sbr_mbp_intf();

logic fsta_dfxact;

endinterface
