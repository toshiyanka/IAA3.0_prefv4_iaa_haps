`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

(* inserted_by="VISA IT" *) logic     [24:0] visaPrbsFrom_hqm_visa_mux3;
(* inserted_by="VISA IT" *) logic      [0:0] visaSrcClk_i_hqm_visa_repeater_vcfn;
(* inserted_by="VISA IT" *) logic [4:0][7:0] visaLaneIn_i_hqm_visa_mux_top_vcfn;
(* inserted_by="VISA IT" *) logic      [0:0] visaSrcClk_i_hqm_visa_mux_top_vcfn;
(* inserted_by="VISA IT" *) logic      [2:0] visaRt_serial_cfg_in_local;
(* inserted_by="VISA IT" *) logic      [0:0] visaRt_bypass_cr_out_from_i_hqm_visa_mux_top_vcfn;
(* inserted_by="VISA IT" *) logic [0:0][7:0] visaRt_lane_out_from_i_hqm_visa_mux_top_vcfn;
(* inserted_by="VISA IT" *) logic      [2:0] visaRt_serial_cfg_in_from_i_hqm_visa_repeater_vcfn;



`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
