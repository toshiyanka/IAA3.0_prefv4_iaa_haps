//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2020 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//
//  Collateral Description:
//  IOSF - Sideband Channel IP
//
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//
//  Revision:
//  2020WW22_PICr33
//
//  Module <mTAP> :  < put your functional description here in plain text >
//
//------------------------------------------------------------------------------

//----------------------------------------------------------------------
// Intel Proprietary -- Copyright 2009 Intel -- All rights reserved
//----------------------------------------------------------------------
// NOTE: Log history is at end of file.
//----------------------------------------------------------------------
//
//    FILENAME    : mtap_irdecoder.sv
//    DESIGNER    : Sunjiv Sachan
//    PROJECT     : mTAP
//    
//    
//    PURPOSE     : MTAP IR Decoder Logic
//    DESCRIPTION :
//       This module generated decoder enable signals. This is generated by
//       comparing instruction address with address defined by parameter.
//----------------------------------------------------------------------
//    LOCAL PARAMETERS:
//
//    HIGH
//       This is 1 bit one value
//
//    LOW
//       This is 1 bit zero value
//
//    ONE
//       This is number 1 to and is declared just to avoid lint warnings
//
//    TWO
//       This is number 2 to and is declared just to avoid lint warnings
//
//    FOUR
//       This is number 4 to and is declared just to avoid lint warnings
//
//    SIX
//       This is number 6 to and is declared just to avoid lint warnings
//
//    SEVEN
//       This is number 7 to and is declared just to avoid lint warnings
//
//    EIGHT
//       This is number 8 to and is declared just to avoid lint warnings
//
//    IRDECODER_MTAP_ADDRESS_OF_USERCODE
//       This is address of optional USERCODE register.
//----------------------------------------------------------------------
module mtap_irdecoder #(
// *********************************************************************
// Parameters
// *********************************************************************
                        parameter IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION       = 8,
                        parameter IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS      = 0,
                        parameter IRDECODER_MTAP_INSTRUCTION_FOR_DATA_REGISTERS = 0,
                        parameter IRDECODER_MTAP_ADDRESS_OF_CLAMP               = 0,
                        parameter IRDECODER_MTAP_MINIMUM_SIZEOF_INSTRUCTION     = 0
                       )
                      (
                       input  logic                                                    powergoodrst_trst_b, // kbbhagwa cdc fix
                       input  logic                                                    atappris_tck, // kbbhagwa cdc fix
                       input  logic [(IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  mtap_irreg_ireg_nxt, // kbbhagwa cdc fix

                       input  logic [(IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  mtap_irreg_ireg,
                       output logic [(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] mtap_irdecoder_drselect,
                       output logic                                                    mtap_and_all_bits_irreg,
                       output logic                                                    mtap_or_all_bits_irreg
                      );

   // *********************************************************************
   // Local parameters
   // *********************************************************************
   localparam HIGH                               = 1'b1;
   localparam LOW                                = 1'b0;
   localparam ONE                                = 1;
   localparam TWO                                = 2;
   localparam FOUR                               = 4;
   localparam SIX                                = 6;
   localparam SEVEN                              = 7;
   localparam EIGHT                              = 8;
   localparam IRDECODER_MTAP_ADDRESS_OF_USERCODE = (IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION == 8) ? 8'h05 :
      {{(IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION - IRDECODER_MTAP_MINIMUM_SIZEOF_INSTRUCTION + 4){LOW}}, 4'h5};
   localparam DRREG_MTAP_POSITION_OF_BYPASS = 2; //kbbhagwa cdc fix

   // *********************************************************************
   // Internal signals
   // *********************************************************************

  //logic [(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - 1):0]  drselect_reset_value;
   logic [(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] decoder_drselect;
   logic                                                    decode_clamp;
   logic                                                    decode_usercode;

   logic [(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] irdecoder_drselect_nxt; //kbbhagwa cdc fix
   logic                                                    and_all_bits_irreg_nxt; //kbbhagwa cdc fix
   logic                                                    or_all_bits_irreg_nxt; //kbbhagwa cdc fix

   // *********************************************************************
   // Generate construct is used to generate number of decoded output lines
   // which is equal to IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS
   // *********************************************************************
   generate
      for (genvar i = 0; i < IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS; i = i + 1)
      begin
         mtap_decoder #(
                        .DECODER_INSTRUCTION_TO_DECODE
                           (IRDECODER_MTAP_INSTRUCTION_FOR_DATA_REGISTERS[
                              (((i * IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION) +
                                IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION) - 1):
                              (i * IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION)]),
                        .DECODER_MTAP_SIZE_OF_EACH_INSTRUCTION
                           (IRDECODER_MTAP_SIZE_OF_EACH_INSTRUCTION)
                       )
         i_mtap_decoder (
//                         .mtap_irreg_ireg  (mtap_irreg_ireg),
                         .mtap_irreg_ireg  (mtap_irreg_ireg_nxt), //kbbhagwa cdc fix
                         .decoder_drselect (decoder_drselect[i])
                        );
      end
   endgenerate

always_ff @(negedge atappris_tck or negedge powergoodrst_trst_b)
begin
  if ( ~ powergoodrst_trst_b )
  begin 
      for ( integer i = 0; i <= (IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS -1); i++ )
      begin
       if ( i == DRREG_MTAP_POSITION_OF_BYPASS )
        mtap_irdecoder_drselect[DRREG_MTAP_POSITION_OF_BYPASS] <= 1'b1;
       else
        mtap_irdecoder_drselect[i] <= 1'b0;
      end
  end
  else 
      mtap_irdecoder_drselect <= irdecoder_drselect_nxt;
end
//kbbhagwa cdc fix


   // *********************************************************************
   // Decoding of some of the Instructions
   // *********************************************************************
   assign mtap_and_all_bits_irreg = &(mtap_irreg_ireg);
   assign and_all_bits_irreg_nxt = &(mtap_irreg_ireg_nxt); //kbbhagwa cdc fix

   assign mtap_or_all_bits_irreg  = |(mtap_irreg_ireg);
   assign or_all_bits_irreg_nxt  = |(mtap_irreg_ireg_nxt); //kbbhagwa cdc fix

//kbbhagwa cdc fix   assign decode_clamp            = (mtap_irreg_ireg == IRDECODER_MTAP_ADDRESS_OF_CLAMP)    ? HIGH : LOW;
   assign decode_clamp            = (mtap_irreg_ireg_nxt == IRDECODER_MTAP_ADDRESS_OF_CLAMP)    ? HIGH : LOW;
//kbbhagwa cdc fix   assign decode_usercode         = (mtap_irreg_ireg == IRDECODER_MTAP_ADDRESS_OF_USERCODE) ? HIGH : LOW;
   assign decode_usercode         = (mtap_irreg_ireg_nxt == IRDECODER_MTAP_ADDRESS_OF_USERCODE) ? HIGH : LOW;

   // *********************************************************************
   // Default value of decoder select points to BYPASS register
   // *********************************************************************
//   assign mtap_irdecoder_drselect =
   assign irdecoder_drselect_nxt =
// kbbhagwa cdc fix      (mtap_and_all_bits_irreg     == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
      (and_all_bits_irreg_nxt     == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
// kbbhagwa cdc fix         (mtap_or_all_bits_irreg   == LOW ) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - TWO){LOW}}, HIGH, LOW} :
         (or_all_bits_irreg_nxt   == LOW ) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - TWO){LOW}}, HIGH, LOW} :
         (decode_clamp             == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         (decode_usercode          == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         (decoder_drselect         ==   {IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS{LOW}}) ?
                                      {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}              :
         (decoder_drselect [FOUR]  == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         //(decoder_drselect [SIX]   == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         //(decoder_drselect [SEVEN] == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         //(decoder_drselect [EIGHT] == HIGH) ? {{(IRDECODER_MTAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
          decoder_drselect;

endmodule
