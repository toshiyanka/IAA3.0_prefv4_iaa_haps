iosf_sb_compliance
            #(.MAX_AGENT_NP_CREDITS (1024),
              .MAX_AGENT_PC_CREDITS (1024),
              .MAX_FABRIC_NP_CREDITS (1024),
              .MAX_FABRIC_PC_CREDITS (1024),
              .PAYLOAD_BANDWIDTH (8),
              .AGENT_IS_DUT(1),
              .FABRIC_IS_DUT(0),
              .CHECKER_IS_DUT(0)
              )
