package hqm_picker_pkg;

import ovm_pkg::*;
import ConfigDB::*;
import systeminit::*;
import base_picker_pkg::*;

//`include "hqm_arch_picker.sv"
`include "hqm_agent_picker.sv"
//`include "hqm_chassis_picker.sv"
`include "hqm_ip_picker.sv"
`include "default_hqm_constraints.sv"
endpackage: hqm_picker_pkg
