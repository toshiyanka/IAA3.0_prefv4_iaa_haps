//Place any new sequences in the SeqLib directory & `include them here. This file `included in your main include file.
`include "SeqLib/CCAgentBaseSequence.svh"
`include "SeqLib/CCAgentDefaultSequence.svh"
//`include "SeqLib/CCAgentBaseResponseVSeq.svh"
