//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2020 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
// AW_unused_bits
//
// This module is used to identify bits of a vector as unused for lint. It takes an input vector
// and assigns it to an internal wire, which is then marked as unused bits for lint purposes.
//
// The following parameters are supported:
//
//	WIDTH	Width of the input.
//
//-----------------------------------------------------------------------------------------------------

module hqm_AW_unused_bits
#(

	 parameter WIDTH	= 1
) (
	 input	logic	[WIDTH-1:0]	a
);

generate
 if (WIDTH > 0) begin: g_unused
   logic [WIDTH-1:0] a_unused_nc;

   assign a_unused_nc = a;
 end
endgenerate

endmodule // AW_unused_bits

