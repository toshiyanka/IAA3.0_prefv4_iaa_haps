`constraint_begin(default_rcfwl_constraints, rcfwl_picker, rcfwl)
  
`constraint_end

