// File output was printed on: Saturday, January 19, 2013 2:59:29 PM
// Chassis TAP Tool version: 0.6.0.0
//----------------------------------------------------------------------
//             TAP                SlvIDcode       IDcode      IR_Width  Node  Sec_connections  Hybrid_en  Dfx_Security  Hierarchy_Level  PositionOfTap  IsIdcode_eq0C
Create_TAP_LUT (IPLEVEL_STAP,  32'h1234_5679,  32'h0000_0001,   'h8,     'd0,       'd0,         'd0,       GREEN,           1,               0,             1);
