//-----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright (2013) (2013) Intel Corporation All Rights Reserved. 
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors. The
// Material is protected by worldwide copyright and trade secret laws and 
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or disclosed
// in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual 
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be 
// express and approved by Intel in writing.
//------------------------------------------------------------------------------
// File   : intr_transaction.sv
//
// Description :
//
// This class is derived form uvm_sequence_item and it represents the transaction 
// object being generated by sequence/sequencer and sent to the DUT through driver
//------------------------------------------------------------------------------
`ifndef INTR_TRANSACTION__SV
`define INTR_TRANSACTION__SV

class intr_transaction extends uvm_sequence_item;



 //------------------------- 
 //-- intr_fields
 //------------------------- 	 
 

 bit            cq_is_ldb;
 logic [7:0]    cq_occ_cq;
 int            cq_occ_cnt;


 bit                    is_done; //- 
 rand bit               is_vf;                  // identifies if the hcw is associated with a VF or PF
 rand bit [3:0]         vf_num;                 // VF number if HCW associated with a VF


 //-------------------------  
 //Constraints
 //-------------------------  
 
constraint c_vf {
                  soft is_vf == 1'b0;
                }


 //-------------------------  
 //static constraint if any
 //-------------------------  
 //static constraint disable_type {xxx == 0;};
  
 

 //------------------------- 
 //-------------------------    
  `uvm_object_utils_begin(intr_transaction)
     `uvm_field_int(cq_is_ldb,   UVM_ALL_ON)
     `uvm_field_int(cq_occ_cq,   UVM_ALL_ON)
     `uvm_field_int(cq_occ_cnt,  UVM_ALL_ON)
     `uvm_field_int(is_vf,           UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(vf_num,          UVM_ALL_ON | UVM_NOCOMPARE)
  `uvm_object_utils_end
  
  
 
 //------------------------- 
 // Function: new 
 // Class constructor
 //------------------------- 
  function new (string name = "intr_xaction_inst");
    super.new(name);

    is_vf = 1'b0;
  endfunction : new


 //------------------------- 
 // Function: post_randomize
 // SV function overload for randomizing this class
 //------------------------- 
 function void post_randomize();
   super.post_randomize();
 endfunction
   
 


  //---------------------------------------------------------------------------- 
  //---------------------------------------------------------------------------- 
  //-- other supporting functions 
  //----------------------------------------------------------------------------   
  extern   virtual         function   void         do_copy(uvm_object rhs);
  extern   virtual         function   bit          do_compare(uvm_object rhs, uvm_comparer comparer);
                                
endclass : intr_transaction


//----------------------------------------------------------------------------
//-- do_copy
//----------------------------------------------------------------------------
function void intr_transaction::do_copy(uvm_object rhs);
    intr_transaction rhs_;
    
    if (!$cast(rhs_, rhs)) begin
       uvm_report_error(get_full_name(), $psprintf("input is not a intr_transaction"));
    end 

    super.do_copy(this);

    cq_is_ldb  = rhs_.cq_is_ldb;
    cq_occ_cq  = rhs_.cq_occ_cq;
    
    cq_occ_cnt = rhs_.cq_occ_cnt;
    is_done    = rhs_.is_done;
 
endfunction

  
 
 
//----------------------------------------------------------------------------
//-- do_compare
//----------------------------------------------------------------------------
function   bit    intr_transaction::do_compare(uvm_object rhs, uvm_comparer comparer);

    intr_transaction that;

    if (!$cast(that, rhs)) begin
      return 0;
    end 

    return ((super.do_compare(rhs, comparer) &&
            (this.cq_occ_cq == that.cq_occ_cq)     &&  
            (this.cq_is_ldb == that.cq_is_ldb)  ));
endfunction
	    
`endif
