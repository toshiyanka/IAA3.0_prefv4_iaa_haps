// File output was printed on: Wednesday, March 20, 2013 9:00:22 AM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
//              TAP name,Opcode,   DR_length
`ifdef JTAG_BFM_TAPLINK_MODE
Create_Reg_Model (CLTAP,    12'h2,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is IDCODE [0x2]
Create_Reg_Model (CLTAP,    12'h1,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is SAMPLE_PRELOAD [0x1]
Create_Reg_Model (CLTAP,    12'h3,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is PRELOAD [0x3]
Create_Reg_Model (CLTAP,    12'h4,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is CLAMP [0x4]
Create_Reg_Model (CLTAP,    12'h6,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is INTEST [0x6]
Create_Reg_Model (CLTAP,    12'h8,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is HIGHZ [0x8]
Create_Reg_Model (CLTAP,    12'h9,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is EXTEST [0x9]
Create_Reg_Model (CLTAP,    12'hD,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is EXTEST_TOGGLE [0xD]
Create_Reg_Model (CLTAP,    12'hE,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is EXTEST_PULSE [0xE]
Create_Reg_Model (CLTAP,    12'hF,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is EXTEST_TRAIN [0xF]
Create_Reg_Model (CLTAP,    12'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is BYPASS [0xFF]
Create_Reg_Model (CLTAP,    12'h34,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is Opcode34_Width32 [0x34]
Create_Reg_Model (CLTAP,    12'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is OpcodeA0_WIdth32 [0xA0]
Create_Reg_Model (CLTAP,    12'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is CLTAPC_REMOVE [0x14]
Create_Reg_Model (CLTAP,    12'h5,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is USERCODE [0x5]
Create_Reg_Model (CLTAP,    12'h7,      'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is RUNBIST [0x7]
Create_Reg_Model (CLTAP,    12'h10,     'd6  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is CLTAPC_SEC_SEL [0x10]
Create_Reg_Model (CLTAP,    12'h11,     'd12 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is CLTAPC_SELECT [0x11]
Create_Reg_Model (CLTAP,    12'h12,     'd12 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif);   // opcode is CLTAPC_SELECT_OVR [0x12]
Create_Reg_Model (CLTAP,    12'h178,    'd0  `ifdef JTAG_BFM_TAPLINK_MODE ,     5,        8,            0 `endif);   // opcode is CLTAPC_SELECT_OVR [0x12]
Create_Reg_Model (CLTAP,    12'h179,    'd0  `ifdef JTAG_BFM_TAPLINK_MODE ,     6,        9,            0 `endif);   // opcode is CLTAPC_SELECT_OVR [0x12]

//
Create_Reg_Model (STAP0,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP0,    8'h50,     'd10 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode50_Width10 [0x50]
Create_Reg_Model (STAP0,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP0,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP1,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP1,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP1,    8'h51,     'd11 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode51_Width11 [0x51]
Create_Reg_Model (STAP1,    8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP1,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP1,    8'h10,     'd2  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP1,    8'h11,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP2,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP2,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP2,    8'h52,     'd12 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode52_Width12 [0x52]
Create_Reg_Model (STAP2,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP2,    8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP2,    8'h10,     'd3  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP2,    8'h11,     'd6  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP3,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP3,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP3,    8'h53,     'd13 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode53_Width13 [0x53]
Create_Reg_Model (STAP3,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP4,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP4,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP4,    8'h54,     'd14 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode54_Width14 [0x54]
Create_Reg_Model (STAP4,    8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP4,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP4,    8'h10,     'd2  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP4,    8'h11,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP5,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP5,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP5,    8'h55,     'd15 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode55_Width15 [0x55]
Create_Reg_Model (STAP5,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP6,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP6,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP6,    8'h56,     'd16 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode56_Width16 [0x56]
Create_Reg_Model (STAP6,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP7,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP7,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP7,    8'h57,     'd17 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode57_Width17 [0x57]
Create_Reg_Model (STAP7,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP8,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP8,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP8,    8'h58,     'd18 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode58_Width18 [0x58]
Create_Reg_Model (STAP8,    8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP8,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP8,    8'h10,     'd5  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP8,    8'h11,     'd10 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP9,    8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP9,    8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP9,    8'h59,     'd19 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode59_Width19 [0x59]
Create_Reg_Model (STAP9,    8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP10,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP10,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP10,   8'h60,     'd20 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode60_Width20 [0x60]
Create_Reg_Model (STAP10,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP11,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP11,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP11,   8'h61,     'd21 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode61_Width21 [0x61]
Create_Reg_Model (STAP11,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP12,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP12,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP12,   8'h62,     'd22 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode62_Width22 [0x62]
Create_Reg_Model (STAP12,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP13,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP13,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     2,        4,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP13,   8'h63,     'd23 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode63_Width23 [0x63]
Create_Reg_Model (STAP13,   8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP13,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP13,   8'h10,     'd2  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP13,   8'h11,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP14,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP14,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP14,   8'h64,     'd24 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode64_Width24 [0x64]
Create_Reg_Model (STAP14,   8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP14,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP14,   8'h10,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP14,   8'h11,     'd8  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP15,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP15,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP15,   8'h65,     'd25 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode65_Width25 [0x65]
Create_Reg_Model (STAP15,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP16,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP16,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP16,   8'h66,     'd26 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is Opcode66_Width26 [0x66]
Create_Reg_Model (STAP16,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0 `endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP17,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP17,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP17,   8'h67,     'd27 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode67_Width27 [0x67]
Create_Reg_Model (STAP17,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP18,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP18,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP18,   8'h68,     'd28 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode68_Width28 [0x68]
Create_Reg_Model (STAP18,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP19,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP19,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP19,   8'h69,     'd29 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode69_Width29 [0x69]
Create_Reg_Model (STAP19,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP20,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP20,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP20,   8'h70,     'd30 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode70_Width30 [0x70]
Create_Reg_Model (STAP20,   8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP20,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP20,   8'h10,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP20,   8'h11,     'd8  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP21,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP21,   8'h71,     'd31 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode71_Width31 [0x71]
Create_Reg_Model (STAP21,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP21,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP22,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP22,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP22,   8'h72,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode72_Width32 [0x72]
Create_Reg_Model (STAP22,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP23,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP23,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP23,   8'h73,     'd33 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode73_Width33 [0x73]
Create_Reg_Model (STAP23,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP24,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP24,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP24,   8'h74,     'd34 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode74_Width34 [0x74]
Create_Reg_Model (STAP24,   8'h14,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP24,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP24,   8'h10,     'd2  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP24,   8'h11,     'd4  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP25,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP25,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP25,   8'h75,     'd35 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode75_Width35 [0x75]
Create_Reg_Model (STAP25,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP26,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP26,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP26,   8'h76,     'd36 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode76_Width36 [0x76]
Create_Reg_Model (STAP26,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP27,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP27,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP27,   8'h77,     'd37 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode77_Width37 [0x77]
Create_Reg_Model (STAP27,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP28,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP28,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP28,   8'h78,     'd38 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode78_Width38 [0x78]
Create_Reg_Model (STAP28,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP29,   8'hFF,     'd1  `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP29,   8'hA0,     'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP29,   8'h79,     'd39 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is Opcode79_Width39 [0x79]
Create_Reg_Model (STAP29,   8'hC,      'd32 `ifdef JTAG_BFM_TAPLINK_MODE ,     0,        0,            0`endif     );   // opcode is IDCODE [0xC]
`else
Create_Reg_Model (CLTAP,    8'h2,      'd32     );   // opcode is IDCODE [0x2]
Create_Reg_Model (CLTAP,    8'h1,      'd1      );   // opcode is SAMPLE_PRELOAD [0x1]
Create_Reg_Model (CLTAP,    8'h3,      'd1      );   // opcode is PRELOAD [0x3]
Create_Reg_Model (CLTAP,    8'h4,      'd1      );   // opcode is CLAMP [0x4]
Create_Reg_Model (CLTAP,    8'h6,      'd1      );   // opcode is INTEST [0x6]
Create_Reg_Model (CLTAP,    8'h8,      'd1      );   // opcode is HIGHZ [0x8]
Create_Reg_Model (CLTAP,    8'h9,      'd1      );   // opcode is EXTEST [0x9]
Create_Reg_Model (CLTAP,    8'hD,      'd1      );   // opcode is EXTEST_TOGGLE [0xD]
Create_Reg_Model (CLTAP,    8'hE,      'd1      );   // opcode is EXTEST_PULSE [0xE]
Create_Reg_Model (CLTAP,    8'hF,      'd1      );   // opcode is EXTEST_TRAIN [0xF]
Create_Reg_Model (CLTAP,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (CLTAP,    8'h34,     'd32     );   // opcode is Opcode34_Width32 [0x34]
Create_Reg_Model (CLTAP,    8'hA0,     'd32     );   // opcode is OpcodeA0_WIdth32 [0xA0]
Create_Reg_Model (CLTAP,    8'h14,     'd1      );   // opcode is CLTAPC_REMOVE [0x14]
Create_Reg_Model (CLTAP,    8'h5,      'd1      );   // opcode is USERCODE [0x5]
Create_Reg_Model (CLTAP,    8'h7,      'd1      );   // opcode is RUNBIST [0x7]
Create_Reg_Model (CLTAP,    8'h10,     'd6      );   // opcode is CLTAPC_SEC_SEL [0x10]
Create_Reg_Model (CLTAP,    8'h11,     'd12     );   // opcode is CLTAPC_SELECT [0x11]
Create_Reg_Model (CLTAP,    8'h12,     'd12     );   // opcode is CLTAPC_SELECT_OVR [0x12]
//
Create_Reg_Model (STAP0,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP0,    8'h50,     'd10     );   // opcode is Opcode50_Width10 [0x50]
Create_Reg_Model (STAP0,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP0,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP1,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP1,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP1,    8'h51,     'd11     );   // opcode is Opcode51_Width11 [0x51]
Create_Reg_Model (STAP1,    8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP1,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP1,    8'h10,     'd2      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP1,    8'h11,     'd4      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP2,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP2,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP2,    8'h52,     'd12     );   // opcode is Opcode52_Width12 [0x52]
Create_Reg_Model (STAP2,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP2,    8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP2,    8'h10,     'd3      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP2,    8'h11,     'd6      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP3,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP3,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP3,    8'h53,     'd13     );   // opcode is Opcode53_Width13 [0x53]
Create_Reg_Model (STAP3,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP4,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP4,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP4,    8'h54,     'd14     );   // opcode is Opcode54_Width14 [0x54]
Create_Reg_Model (STAP4,    8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP4,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP4,    8'h10,     'd2      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP4,    8'h11,     'd4      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP5,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP5,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP5,    8'h55,     'd15     );   // opcode is Opcode55_Width15 [0x55]
Create_Reg_Model (STAP5,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP6,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP6,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP6,    8'h56,     'd16     );   // opcode is Opcode56_Width16 [0x56]
Create_Reg_Model (STAP6,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP7,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP7,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP7,    8'h57,     'd17     );   // opcode is Opcode57_Width17 [0x57]
Create_Reg_Model (STAP7,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP8,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP8,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP8,    8'h58,     'd18     );   // opcode is Opcode58_Width18 [0x58]
Create_Reg_Model (STAP8,    8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP8,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP8,    8'h10,     'd5      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP8,    8'h11,     'd10     );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP9,    8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP9,    8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP9,    8'h59,     'd19     );   // opcode is Opcode59_Width19 [0x59]
Create_Reg_Model (STAP9,    8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP10,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP10,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP10,   8'h60,     'd20     );   // opcode is Opcode60_Width20 [0x60]
Create_Reg_Model (STAP10,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP11,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP11,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP11,   8'h61,     'd21     );   // opcode is Opcode61_Width21 [0x61]
Create_Reg_Model (STAP11,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP12,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP12,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP12,   8'h62,     'd22     );   // opcode is Opcode62_Width22 [0x62]
Create_Reg_Model (STAP12,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP13,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP13,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP13,   8'h63,     'd23     );   // opcode is Opcode63_Width23 [0x63]
Create_Reg_Model (STAP13,   8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP13,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP13,   8'h10,     'd2      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP13,   8'h11,     'd4      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP14,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP14,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP14,   8'h64,     'd24     );   // opcode is Opcode64_Width24 [0x64]
Create_Reg_Model (STAP14,   8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP14,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP14,   8'h10,     'd4      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP14,   8'h11,     'd8      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP15,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP15,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP15,   8'h65,     'd25     );   // opcode is Opcode65_Width25 [0x65]
Create_Reg_Model (STAP15,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP16,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP16,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP16,   8'h66,     'd26     );   // opcode is Opcode66_Width26 [0x66]
Create_Reg_Model (STAP16,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP17,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP17,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP17,   8'h67,     'd27     );   // opcode is Opcode67_Width27 [0x67]
Create_Reg_Model (STAP17,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP18,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP18,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP18,   8'h68,     'd28     );   // opcode is Opcode68_Width28 [0x68]
Create_Reg_Model (STAP18,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP19,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP19,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP19,   8'h69,     'd29     );   // opcode is Opcode69_Width29 [0x69]
Create_Reg_Model (STAP19,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP20,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP20,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP20,   8'h70,     'd30     );   // opcode is Opcode70_Width30 [0x70]
Create_Reg_Model (STAP20,   8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP20,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP20,   8'h10,     'd4      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP20,   8'h11,     'd8      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP21,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP21,   8'h71,     'd31     );   // opcode is Opcode71_Width31 [0x71]
Create_Reg_Model (STAP21,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP21,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP22,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP22,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP22,   8'h72,     'd32     );   // opcode is Opcode72_Width32 [0x72]
Create_Reg_Model (STAP22,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP23,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP23,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP23,   8'h73,     'd33     );   // opcode is Opcode73_Width33 [0x73]
Create_Reg_Model (STAP23,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP24,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP24,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP24,   8'h74,     'd34     );   // opcode is Opcode74_Width34 [0x74]
Create_Reg_Model (STAP24,   8'h14,     'd1      );   // opcode is TAPC_REMOVE [0x14]
Create_Reg_Model (STAP24,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
Create_Reg_Model (STAP24,   8'h10,     'd2      );   // opcode is TAPC_SEC_SEL [0x10]
Create_Reg_Model (STAP24,   8'h11,     'd4      );   // opcode is TAPC_SELECT [0x11]
//
Create_Reg_Model (STAP25,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP25,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP25,   8'h75,     'd35     );   // opcode is Opcode75_Width35 [0x75]
Create_Reg_Model (STAP25,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP26,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP26,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP26,   8'h76,     'd36     );   // opcode is Opcode76_Width36 [0x76]
Create_Reg_Model (STAP26,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP27,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP27,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP27,   8'h77,     'd37     );   // opcode is Opcode77_Width37 [0x77]
Create_Reg_Model (STAP27,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP28,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP28,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP28,   8'h78,     'd38     );   // opcode is Opcode78_Width38 [0x78]
Create_Reg_Model (STAP28,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
Create_Reg_Model (STAP29,   8'hFF,     'd1      );   // opcode is BYPASS [0xFF]
Create_Reg_Model (STAP29,   8'hA0,     'd32     );   // opcode is OpcodeA0_Width32 [0xA0]
Create_Reg_Model (STAP29,   8'h79,     'd39     );   // opcode is Opcode79_Width39 [0x79]
Create_Reg_Model (STAP29,   8'hC,      'd32     );   // opcode is IDCODE [0xC]
//
`endif
