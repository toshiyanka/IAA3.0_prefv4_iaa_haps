`ifndef __VISA_IT__
`ifndef INTEL_GLOBAL_VISA_DISABLE

(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  0:  0] = visa_capture_reg_f.core_gated_rst_b             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  1:  1] = visa_capture_reg_f.constant_one                 ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  2:  2] = visa_capture_reg_f.rop_qed_force_clockon        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  3:  3] = visa_capture_reg_f.prim_clk_enable              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  4:  4] = visa_capture_reg_f.hqm_clk_enable               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  5:  5] = visa_capture_reg_f.hqm_clk_throttle             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  6:  6] = visa_capture_reg_f.hqm_gclock_enable            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  7:  7] = visa_capture_reg_f.hqm_cdc_clk_enable           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  8:  8] = visa_capture_reg_f.hqm_gated_local_override     ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[  9:  9] = visa_capture_reg_f.hqm_flr_prep                 ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 10: 10] = visa_capture_reg_f.pm_ip_clk_halt_b_2_rpt_0_iosf;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 11: 11] = visa_capture_reg_f.hqm_alarm_ready              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 12: 12] = visa_capture_reg_f.hqm_alarm_v                  ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 13: 13] = visa_capture_reg_f.hqm_unit_pipeidle            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 14: 14] = visa_capture_reg_f.hqm_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 15: 15] = visa_capture_reg_f.hqm_proc_reset_done          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 16: 16] = visa_capture_reg_f.sys_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 17: 17] = visa_capture_reg_f.sys_reset_done               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 18: 18] = visa_capture_reg_f.aqed_unit_pipeidle           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 19: 19] = visa_capture_reg_f.qed_unit_pipeidle            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 20: 20] = visa_capture_reg_f.dp_unit_pipeidle             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 21: 21] = visa_capture_reg_f.ap_unit_pipeidle             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 22: 22] = visa_capture_reg_f.nalb_unit_pipeidle           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 23: 23] = visa_capture_reg_f.lsp_unit_pipeidle            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 24: 24] = visa_capture_reg_f.rop_unit_pipeidle            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 25: 25] = visa_capture_reg_f.chp_unit_pipeidle            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 26: 26] = visa_capture_reg_f.aqed_unit_idle               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 27: 27] = visa_capture_reg_f.qed_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 28: 28] = visa_capture_reg_f.dp_unit_idle                 ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 29: 29] = visa_capture_reg_f.ap_unit_idle                 ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 30: 30] = visa_capture_reg_f.nalb_unit_idle               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 31: 31] = visa_capture_reg_f.lsp_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 32: 32] = visa_capture_reg_f.rop_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 33: 33] = visa_capture_reg_f.chp_unit_idle                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 34: 34] = visa_capture_reg_f.sys_hqm_proc_clk_en          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 35: 35] = visa_capture_reg_f.nalb_hqm_proc_clk_en         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 36: 36] = visa_capture_reg_f.dp_hqm_proc_clk_en           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 37: 37] = visa_capture_reg_f.qed_hqm_proc_clk_en          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 38: 38] = visa_capture_reg_f.lsp_hqm_proc_clk_en          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 39: 39] = visa_capture_reg_f.chp_hqm_proc_clk_en          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 40: 40] = visa_capture_reg_f.aqed_reset_done              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 41: 41] = visa_capture_reg_f.qed_reset_done               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 42: 42] = visa_capture_reg_f.dp_reset_done                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 43: 43] = visa_capture_reg_f.ap_reset_done                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 44: 44] = visa_capture_reg_f.nalb_reset_done              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 45: 45] = visa_capture_reg_f.lsp_reset_done               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 46: 46] = visa_capture_reg_f.rop_reset_done               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 47: 47] = visa_capture_reg_f.chp_reset_done               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 48: 48] = visa_capture_reg_f.cwdi_interrupt_w_req_ready   ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 49: 49] = visa_capture_reg_f.cwdi_interrupt_w_req_valid   ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 50: 50] = visa_capture_reg_f.interrupt_w_req_ready        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 51: 51] = visa_capture_reg_f.interrupt_w_req_valid        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 52: 52] = visa_capture_reg_f.aqed_chp_sch_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 53: 53] = visa_capture_reg_f.aqed_chp_sch_v               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 54: 54] = visa_capture_reg_f.aqed_ap_enq_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 55: 55] = visa_capture_reg_f.aqed_ap_enq_v                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 56: 56] = visa_capture_reg_f.aqed_lsp_sch_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 57: 57] = visa_capture_reg_f.aqed_lsp_sch_v               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 58: 58] = visa_capture_reg_f.qed_aqed_enq_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 59: 59] = visa_capture_reg_f.qed_aqed_enq_v               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 60: 60] = visa_capture_reg_f.qed_chp_sch_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 61: 61] = visa_capture_reg_f.qed_chp_sch_v                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 62: 62] = visa_capture_reg_f.ap_aqed_ready                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 63: 63] = visa_capture_reg_f.ap_aqed_v                    ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 64: 64] = visa_capture_reg_f.dp_lsp_enq_dir_ready         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 65: 65] = visa_capture_reg_f.dp_lsp_enq_dir_v             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 66: 66] = visa_capture_reg_f.nalb_lsp_enq_lb_ready        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 67: 67] = visa_capture_reg_f.nalb_lsp_enq_lb_v            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 68: 68] = visa_capture_reg_f.lsp_nalb_sch_atq_ready       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 69: 69] = visa_capture_reg_f.lsp_nalb_sch_atq_v           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 70: 70] = visa_capture_reg_f.lsp_dp_sch_rorply_ready      ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 71: 71] = visa_capture_reg_f.lsp_dp_sch_rorply_v          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 72: 72] = visa_capture_reg_f.lsp_nalb_sch_rorply_ready    ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 73: 73] = visa_capture_reg_f.lsp_nalb_sch_rorply_v        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 74: 74] = visa_capture_reg_f.lsp_dp_sch_dir_ready         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 75: 75] = visa_capture_reg_f.lsp_dp_sch_dir_v             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 76: 76] = visa_capture_reg_f.lsp_nalb_sch_unoord_ready    ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 77: 77] = visa_capture_reg_f.lsp_nalb_sch_unoord_v        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 78: 78] = visa_capture_reg_f.rop_dqed_enq_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 79: 79] = visa_capture_reg_f.rop_qed_enq_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 80: 80] = visa_capture_reg_f.rop_qed_dqed_enq_v           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 81: 81] = visa_capture_reg_f.rop_nalb_enq_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 82: 82] = visa_capture_reg_f.rop_nalb_enq_v               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 83: 83] = visa_capture_reg_f.rop_dp_enq_ready             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 84: 84] = visa_capture_reg_f.rop_dp_enq_v                 ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 85: 85] = visa_capture_reg_f.chp_lsp_token_ready          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 86: 86] = visa_capture_reg_f.chp_lsp_token_v              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 87: 87] = visa_capture_reg_f.chp_lsp_cmp_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 88: 88] = visa_capture_reg_f.chp_lsp_cmp_v                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 89: 89] = visa_capture_reg_f.chp_lsp_cmp_data             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 90: 90] = visa_capture_reg_f.chp_rop_hcw_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 91: 91] = visa_capture_reg_f.chp_rop_hcw_v                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 92: 92] = visa_capture_reg_f.hcw_enq_w_req_ready          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 93: 93] = visa_capture_reg_f.hcw_enq_w_req_valid          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 94: 94] = visa_capture_reg_f.hcw_sched_w_req_ready        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 95: 95] = visa_capture_reg_f.hcw_sched_w_req_valid        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 96: 96] = visa_capture_reg_f.rop_lsp_reordercmp_ready     ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 97: 97] = visa_capture_reg_f.rop_lsp_reordercmp_v         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 98: 98] = visa_capture_reg_f.dp_lsp_enq_rorply_ready      ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[ 99: 99] = visa_capture_reg_f.dp_lsp_enq_rorply_v          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[100:100] = visa_capture_reg_f.nalb_lsp_enq_rorply_ready    ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[101:101] = visa_capture_reg_f.nalb_lsp_enq_rorply_v        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[102:102] = visa_capture_reg_f.aqed_cfg_req_down_write      ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[103:103] = visa_capture_reg_f.aqed_cfg_req_down_read       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[105:104] = visa_capture_reg_f.aqed_cfg_req_down[1:0]       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[106:106] = visa_capture_reg_f.aqed_cfg_rsp_down_ack        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[108:107] = visa_capture_reg_f.aqed_cfg_rsp_down[1:0]       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[109:109] = visa_capture_reg_f.qed_cfg_req_down_write       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[110:110] = visa_capture_reg_f.qed_cfg_req_down_read        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[112:111] = visa_capture_reg_f.qed_cfg_req_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[113:113] = visa_capture_reg_f.qed_cfg_rsp_down_ack         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[115:114] = visa_capture_reg_f.qed_cfg_rsp_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[116:116] = visa_capture_reg_f.ap_cfg_req_down_write        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[117:117] = visa_capture_reg_f.ap_cfg_req_down_read         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[119:118] = visa_capture_reg_f.ap_cfg_req_down[1:0]         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[120:120] = visa_capture_reg_f.ap_cfg_rsp_down_ack          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[122:121] = visa_capture_reg_f.ap_cfg_rsp_down[1:0]         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[123:123] = visa_capture_reg_f.lsp_cfg_req_down_write       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[124:124] = visa_capture_reg_f.lsp_cfg_req_down_read        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[126:125] = visa_capture_reg_f.lsp_cfg_req_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[127:127] = visa_capture_reg_f.lsp_cfg_rsp_down_ack         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[129:128] = visa_capture_reg_f.lsp_cfg_rsp_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[130:130] = visa_capture_reg_f.rop_cfg_req_down_write       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[131:131] = visa_capture_reg_f.rop_cfg_req_down_read        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[133:132] = visa_capture_reg_f.rop_cfg_req_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[134:134] = visa_capture_reg_f.rop_cfg_rsp_down_ack         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[136:135] = visa_capture_reg_f.rop_cfg_rsp_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[137:137] = visa_capture_reg_f.chp_cfg_req_down_write       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[138:138] = visa_capture_reg_f.chp_cfg_req_down_read        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[140:139] = visa_capture_reg_f.chp_cfg_req_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[141:141] = visa_capture_reg_f.chp_cfg_rsp_down_ack         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[143:142] = visa_capture_reg_f.chp_cfg_rsp_down[1:0]        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[144:144] = visa_capture_reg_f.mstr_cfg_req_down_write      ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[145:145] = visa_capture_reg_f.mstr_cfg_req_down_read       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[147:146] = visa_capture_reg_f.mstr_cfg_req_down[1:0]       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[148:148] = visa_capture_reg_f.mstr_cfg_rsp_down_ack        ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[150:149] = visa_capture_reg_f.mstr_cfg_rsp_down[1:0]       ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[151:151] = visa_capture_reg_f.aqed_lsp_deq_v               ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[152:152] = visa_capture_reg_f.qed_lsp_deq_v                ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[153:153] = visa_capture_reg_f.rop_alarm_up_ready           ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[154:154] = visa_capture_reg_f.qed_alarm_down_v             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[155:155] = visa_capture_reg_f.ap_alarm_up_ready            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[156:156] = visa_capture_reg_f.aqed_alarm_down_v            ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[157:157] = visa_capture_reg_f.ap_alarm_down_ready          ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[158:158] = visa_capture_reg_f.ap_alarm_down_v              ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[159:159] = visa_capture_reg_f.lsp_alarm_down_ready         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[160:160] = visa_capture_reg_f.lsp_alarm_down_v             ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[161:161] = visa_capture_reg_f.rop_alarm_down_ready         ;
(* inserted_by="VISA IT" *) assign visaPrbsFrom_hqm_core_visa_block[162:162] = visa_capture_reg_f.rop_alarm_down_v             ;
(* inserted_by="VISA IT" *) assign visaRt_probe_from_i_hqm_core_visa_block   = visaPrbsFrom_hqm_core_visa_block                ;



`endif // INTEL_GLOBAL_VISA_DISABLE
`endif // __VISA_IT__
