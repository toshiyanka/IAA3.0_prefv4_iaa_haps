//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv0_sbr_cfg_1_ep_rtl/lv0_sbr_cfg_1_ep_rtl.csv rev -1.00
//
//------------------------------------------------------------------------------


//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------

module sbr
(
  // lintra push -80009, -80018, -70023
  // Synchronous Clock/Reset
          clk,
          rstb,

  // Power Well Isolation Input Signals
          pd1_pwrgd,

          p0_fab_init_idle_exit,
          p0_fab_init_idle_exit_ack,
          p1_fab_init_idle_exit,
          p1_fab_init_idle_exit_ack,
          p2_fab_init_idle_exit,
          p2_fab_init_idle_exit_ack,
          p3_fab_init_idle_exit,
          p3_fab_init_idle_exit_ack,
          p4_fab_init_idle_exit,
          p4_fab_init_idle_exit_ack,
          p5_fab_init_idle_exit,
          p5_fab_init_idle_exit_ack,
          p6_fab_init_idle_exit,
          p6_fab_init_idle_exit_ack,
          p7_fab_init_idle_exit,
          p7_fab_init_idle_exit_ack,
          sbr_idle,
  // VISA Debug Signal/Clock Outputs
 visa_arb_clk,
 visa_vp_clk,
 visa_p0_tier1_clk,
 visa_p0_tier2_clk,
 visa_p1_tier1_clk,
 visa_p1_tier2_clk,
 visa_p2_tier1_clk,
 visa_p2_tier2_clk,
 visa_p3_tier1_clk,
 visa_p3_tier2_clk,
 visa_p4_tier1_clk,
 visa_p4_tier2_clk,
 visa_p5_tier1_clk,
 visa_p5_tier2_clk,
 visa_p6_tier1_clk,
 visa_p6_tier2_clk,
 visa_p7_tier1_clk,
 visa_p7_tier2_clk,

  // DFx signals
          fscan_latchopen,
          fscan_latchclosed_b,
          fscan_clkungate,
          fscan_rstbypen,
          fscan_byprst_b,
  // Port 0 declarations
    ep0_sbr_side_ism_agent,
    sbr_ep0_side_ism_fabric,
          ep0_sbr_pccup,
          ep0_sbr_npcup,
          sbr_ep0_pcput,
          sbr_ep0_npput,
          sbr_ep0_eom,
    sbr_ep0_payload,
          sbr_ep0_pccup,
          sbr_ep0_npcup,
          ep0_sbr_pcput,
          ep0_sbr_npput,
          ep0_sbr_eom,
    ep0_sbr_payload,

  // Port 1 declarations
    ep1_sbr_side_ism_agent,
    sbr_ep1_side_ism_fabric,
          ep1_sbr_pccup,
          ep1_sbr_npcup,
          sbr_ep1_pcput,
          sbr_ep1_npput,
          sbr_ep1_eom,
    sbr_ep1_payload,
          sbr_ep1_pccup,
          sbr_ep1_npcup,
          ep1_sbr_pcput,
          ep1_sbr_npput,
          ep1_sbr_eom,
    ep1_sbr_payload,

  // Port 2 declarations
    ep2_sbr_side_ism_agent,
    sbr_ep2_side_ism_fabric,
          ep2_sbr_pccup,
          ep2_sbr_npcup,
          sbr_ep2_pcput,
          sbr_ep2_npput,
          sbr_ep2_eom,
    sbr_ep2_payload,
          sbr_ep2_pccup,
          sbr_ep2_npcup,
          ep2_sbr_pcput,
          ep2_sbr_npput,
          ep2_sbr_eom,
    ep2_sbr_payload,

  // Port 3 declarations
    ep3_sbr_side_ism_agent,
    sbr_ep3_side_ism_fabric,
          ep3_sbr_pccup,
          ep3_sbr_npcup,
          sbr_ep3_pcput,
          sbr_ep3_npput,
          sbr_ep3_eom,
    sbr_ep3_payload,
          sbr_ep3_pccup,
          sbr_ep3_npcup,
          ep3_sbr_pcput,
          ep3_sbr_npput,
          ep3_sbr_eom,
    ep3_sbr_payload,

  // Port 4 declarations
    ep4_sbr_side_ism_agent,
    sbr_ep4_side_ism_fabric,
          ep4_sbr_pccup,
          ep4_sbr_npcup,
          sbr_ep4_pcput,
          sbr_ep4_npput,
          sbr_ep4_eom,
    sbr_ep4_payload,
          sbr_ep4_pccup,
          sbr_ep4_npcup,
          ep4_sbr_pcput,
          ep4_sbr_npput,
          ep4_sbr_eom,
    ep4_sbr_payload,

  // Port 5 declarations
    ep5_sbr_side_ism_agent,
    sbr_ep5_side_ism_fabric,
          ep5_sbr_pccup,
          ep5_sbr_npcup,
          sbr_ep5_pcput,
          sbr_ep5_npput,
          sbr_ep5_eom,
    sbr_ep5_payload,
          sbr_ep5_pccup,
          sbr_ep5_npcup,
          ep5_sbr_pcput,
          ep5_sbr_npput,
          ep5_sbr_eom,
    ep5_sbr_payload,

  // Port 6 declarations
    ep6_sbr_side_ism_agent,
    sbr_ep6_side_ism_fabric,
          ep6_sbr_pccup,
          ep6_sbr_npcup,
          sbr_ep6_pcput,
          sbr_ep6_npput,
          sbr_ep6_eom,
    sbr_ep6_payload,
          sbr_ep6_pccup,
          sbr_ep6_npcup,
          ep6_sbr_pcput,
          ep6_sbr_npput,
          ep6_sbr_eom,
    ep6_sbr_payload,

  // Port 7 declarations
    ep7_sbr_side_ism_agent,
    sbr_ep7_side_ism_fabric,
          ep7_sbr_pccup,
          ep7_sbr_npcup,
          sbr_ep7_pcput,
          sbr_ep7_npput,
          sbr_ep7_eom,
    sbr_ep7_payload,
          sbr_ep7_pccup,
          sbr_ep7_npcup,
          ep7_sbr_pcput,
          ep7_sbr_npput,
          ep7_sbr_eom,
    ep7_sbr_payload
);

`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"
  
   // lintra push -80009, -80018, -70023
  // Synchronous Clock/Reset
  input  logic        clk;
  input  logic        rstb;

  // Power Well Isolation Input Signals
  input  logic        pd1_pwrgd;

  output logic        p0_fab_init_idle_exit;
  input  logic        p0_fab_init_idle_exit_ack;
  output logic        p1_fab_init_idle_exit;
  input  logic        p1_fab_init_idle_exit_ack;
  output logic        p2_fab_init_idle_exit;
  input  logic        p2_fab_init_idle_exit_ack;
  output logic        p3_fab_init_idle_exit;
  input  logic        p3_fab_init_idle_exit_ack;
  output logic        p4_fab_init_idle_exit;
  input  logic        p4_fab_init_idle_exit_ack;
  output logic        p5_fab_init_idle_exit;
  input  logic        p5_fab_init_idle_exit_ack;
  output logic        p6_fab_init_idle_exit;
  input  logic        p6_fab_init_idle_exit_ack;
  output logic        p7_fab_init_idle_exit;
  input  logic        p7_fab_init_idle_exit_ack;
  output logic        sbr_idle;
  // VISA Debug Signal/Clock Outputs
  output visa_arb visa_arb_clk;
  output visa_vp  visa_vp_clk;
  output visa_port_tier1 visa_p0_tier1_clk;
  output visa_port_tier2 visa_p0_tier2_clk;
  output visa_port_tier1 visa_p1_tier1_clk;
  output visa_port_tier2 visa_p1_tier2_clk;
  output visa_port_tier1 visa_p2_tier1_clk;
  output visa_port_tier2 visa_p2_tier2_clk;
  output visa_port_tier1 visa_p3_tier1_clk;
  output visa_port_tier2 visa_p3_tier2_clk;
  output visa_port_tier1 visa_p4_tier1_clk;
  output visa_port_tier2 visa_p4_tier2_clk;
  output visa_port_tier1 visa_p5_tier1_clk;
  output visa_port_tier2 visa_p5_tier2_clk;
  output visa_port_tier1 visa_p6_tier1_clk;
  output visa_port_tier2 visa_p6_tier2_clk;
  output visa_port_tier1 visa_p7_tier1_clk;
  output visa_port_tier2 visa_p7_tier2_clk;

  // DFx signals
  input  logic        fscan_latchopen;
  input  logic        fscan_latchclosed_b;
  input  logic        fscan_clkungate;
  input  logic        fscan_rstbypen;
  input  logic        fscan_byprst_b;
  // Port 0 declarations
  input  logic [ 2:0] ep0_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep0_side_ism_fabric;
  input  logic        ep0_sbr_pccup;
  input  logic        ep0_sbr_npcup;
  output logic        sbr_ep0_pcput;
  output logic        sbr_ep0_npput;
  output logic        sbr_ep0_eom;
  output logic [ 7:0] sbr_ep0_payload;
  output logic        sbr_ep0_pccup;
  output logic        sbr_ep0_npcup;
  input  logic        ep0_sbr_pcput;
  input  logic        ep0_sbr_npput;
  input  logic        ep0_sbr_eom;
  input  logic [ 7:0] ep0_sbr_payload;

  // Port 1 declarations
  input  logic [ 2:0] ep1_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep1_side_ism_fabric;
  input  logic        ep1_sbr_pccup;
  input  logic        ep1_sbr_npcup;
  output logic        sbr_ep1_pcput;
  output logic        sbr_ep1_npput;
  output logic        sbr_ep1_eom;
  output logic [ 7:0] sbr_ep1_payload;
  output logic        sbr_ep1_pccup;
  output logic        sbr_ep1_npcup;
  input  logic        ep1_sbr_pcput;
  input  logic        ep1_sbr_npput;
  input  logic        ep1_sbr_eom;
  input  logic [ 7:0] ep1_sbr_payload;

  // Port 2 declarations
  input  logic [ 2:0] ep2_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep2_side_ism_fabric;
  input  logic        ep2_sbr_pccup;
  input  logic        ep2_sbr_npcup;
  output logic        sbr_ep2_pcput;
  output logic        sbr_ep2_npput;
  output logic        sbr_ep2_eom;
  output logic [15:0] sbr_ep2_payload;
  output logic        sbr_ep2_pccup;
  output logic        sbr_ep2_npcup;
  input  logic        ep2_sbr_pcput;
  input  logic        ep2_sbr_npput;
  input  logic        ep2_sbr_eom;
  input  logic [15:0] ep2_sbr_payload;

  // Port 3 declarations
  input  logic [ 2:0] ep3_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep3_side_ism_fabric;
  input  logic        ep3_sbr_pccup;
  input  logic        ep3_sbr_npcup;
  output logic        sbr_ep3_pcput;
  output logic        sbr_ep3_npput;
  output logic        sbr_ep3_eom;
  output logic [15:0] sbr_ep3_payload;
  output logic        sbr_ep3_pccup;
  output logic        sbr_ep3_npcup;
  input  logic        ep3_sbr_pcput;
  input  logic        ep3_sbr_npput;
  input  logic        ep3_sbr_eom;
  input  logic [15:0] ep3_sbr_payload;

  // Port 4 declarations
  input  logic [ 2:0] ep4_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep4_side_ism_fabric;
  input  logic        ep4_sbr_pccup;
  input  logic        ep4_sbr_npcup;
  output logic        sbr_ep4_pcput;
  output logic        sbr_ep4_npput;
  output logic        sbr_ep4_eom;
  output logic [ 7:0] sbr_ep4_payload;
  output logic        sbr_ep4_pccup;
  output logic        sbr_ep4_npcup;
  input  logic        ep4_sbr_pcput;
  input  logic        ep4_sbr_npput;
  input  logic        ep4_sbr_eom;
  input  logic [ 7:0] ep4_sbr_payload;

  // Port 5 declarations
  input  logic [ 2:0] ep5_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep5_side_ism_fabric;
  input  logic        ep5_sbr_pccup;
  input  logic        ep5_sbr_npcup;
  output logic        sbr_ep5_pcput;
  output logic        sbr_ep5_npput;
  output logic        sbr_ep5_eom;
  output logic [ 7:0] sbr_ep5_payload;
  output logic        sbr_ep5_pccup;
  output logic        sbr_ep5_npcup;
  input  logic        ep5_sbr_pcput;
  input  logic        ep5_sbr_npput;
  input  logic        ep5_sbr_eom;
  input  logic [ 7:0] ep5_sbr_payload;

  // Port 6 declarations
  input  logic [ 2:0] ep6_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep6_side_ism_fabric;
  input  logic        ep6_sbr_pccup;
  input  logic        ep6_sbr_npcup;
  output logic        sbr_ep6_pcput;
  output logic        sbr_ep6_npput;
  output logic        sbr_ep6_eom;
  output logic [15:0] sbr_ep6_payload;
  output logic        sbr_ep6_pccup;
  output logic        sbr_ep6_npcup;
  input  logic        ep6_sbr_pcput;
  input  logic        ep6_sbr_npput;
  input  logic        ep6_sbr_eom;
  input  logic [15:0] ep6_sbr_payload;

  // Port 7 declarations
  input  logic [ 2:0] ep7_sbr_side_ism_agent;
  output logic [ 2:0] sbr_ep7_side_ism_fabric;
  input  logic        ep7_sbr_pccup;
  input  logic        ep7_sbr_npcup;
  output logic        sbr_ep7_pcput;
  output logic        sbr_ep7_npput;
  output logic        sbr_ep7_eom;
  output logic [15:0] sbr_ep7_payload;
  output logic        sbr_ep7_pccup;
  output logic        sbr_ep7_npcup;
  input  logic        ep7_sbr_pcput;
  input  logic        ep7_sbr_npput;
  input  logic        ep7_sbr_eom;
  input  logic [15:0] ep7_sbr_payload;
 
//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_sbcportmap;
always_comb sbr_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr (sbr)                                     SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  222 { 17'b0_0000_0000_0000_0000 }},   //   254: 33      SBCPORTMAPTABLE
               17'b1_0000_0000_0000_1111,      //    32          SBCPORTMAPTABLE
      {   18 { 17'b0_0000_0000_0000_0000 }},   //    31: 14      SBCPORTMAPTABLE
               17'b0_0000_0000_1000_0000,      //    13          SBCPORTMAPTABLE
               17'b0_0000_0000_0100_0000,      //    12          SBCPORTMAPTABLE
               17'b0_0000_0000_0010_0000,      //    11          SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //    10          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //     9          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //     8          SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0010 }},   //     7:  4      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }}    //     3:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  7;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;
logic                              p5_pcdstvld;
logic                              p6_pcdstvld;
logic                              p7_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic                              p5_npfence;
logic                              p6_npfence;
logic                              p7_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;
logic                              p5_npdstvld;
logic                              p6_npdstvld;
logic                              p7_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p1_ism_idle;
logic                              p2_ism_idle;
logic                              p3_ism_idle;
logic                              p4_ism_idle;
logic                              p5_ism_idle;
logic                              p6_ism_idle;
logic                              p7_ism_idle;
logic                              p0_cg_inprogress;
logic                              p1_cg_inprogress;
logic                              p2_cg_inprogress;
logic                              p3_cg_inprogress;
logic                              p4_cg_inprogress;
logic                              p5_cg_inprogress;
logic                              p6_cg_inprogress;
logic                              p7_cg_inprogress;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              pd1_pwrgd_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = '1;
always_comb cfg_clkgatedef    = '0;
always_comb cfg_idlecnt       = 8'h10;
always_comb jta_clkgate_ovrd  = '0;
always_comb jta_force_idle    = '0;
always_comb jta_force_notidle = '0;
always_comb jta_force_creditreq = '0;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( force_creditreq               )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_pd1_pwrgd (
  .d                   ( pd1_pwrgd                     ),
  .clr_b               ( rstb                          ),
  .clk                 ( clk                           ),
  .q                   ( pd1_pwrgd_ff2                 )
);


always_comb endpoint_pwrgd = { pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1,
                          pd1_pwrgd_ff2,
                          1'b1
                        };

logic p7_gated_clk;
sbc_clock_gate p7_pwr_clkgate  (
  .en ( endpoint_pwrgd[7] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk                           ),
  .enclk ( p7_gated_clk )
);

logic p5_gated_clk;
sbc_clock_gate p5_pwr_clkgate  (
  .en ( endpoint_pwrgd[5] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk                           ),
  .enclk ( p5_gated_clk )
);

logic p3_gated_clk;
sbc_clock_gate p3_pwr_clkgate  (
  .en ( endpoint_pwrgd[3] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk                           ),
  .enclk ( p3_gated_clk )
);

logic p1_gated_clk;
sbc_clock_gate p1_pwr_clkgate  (
  .en ( endpoint_pwrgd[1] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk                           ),
  .enclk ( p1_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p7_ism_idle | ~endpoint_pwrgd[7])
                  &  (p6_ism_idle | ~endpoint_pwrgd[6])
                  &  (p5_ism_idle | ~endpoint_pwrgd[5])
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
// SBR_IDLE signal for PMU
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle &
                  p2_ism_idle &
                  p3_ism_idle &
                  p4_ism_idle &
                  p5_ism_idle &
                  p6_ism_idle &
                  p7_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p7_npfence,
                 p6_npfence,
                 p5_npfence,
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p7_pcdstvld,
                 p6_pcdstvld,
                 p5_pcdstvld,
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p7_npdstvld,
                 p6_npdstvld,
                 p5_npdstvld,
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_clk = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk                           ),
  .side_rst_b          ( rstb                          ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_clk = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p0_fab_init_idle_exit <= '0;
    else
      p0_fab_init_idle_exit <= ~agent_idle[0] & (ep0_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p0_fab_init_idle_exit_ack & ~p0_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep0_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep0_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p0_side_clk_valid <= 1'b0;
        if ( p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack )
          p0_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_clk = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_clk = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport0 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( ep0_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep0_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .ism_idle            ( p0_ism_idle                   ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_ep0_pccup                 ),
  .tnpcup              ( sbr_ep0_npcup                 ),
  .tpcput              ( ep0_sbr_pcput                 ),
  .tnpput              ( ep0_sbr_npput                 ),
  .teom                ( ep0_sbr_eom                   ),
  .tpayload            ( ep0_sbr_payload               ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( ep0_sbr_pccup                 ),
  .mnpcup              ( ep0_sbr_npcup                 ),
  .mpcput              ( sbr_ep0_pcput                 ),
  .mnpput              ( sbr_ep0_npput                 ),
  .meom                ( sbr_ep0_eom                   ),
  .mpayload            ( sbr_ep0_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
logic p1_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p1_fab_init_idle_exit <= '0;
    else
      p1_fab_init_idle_exit <= ~agent_idle[1] & (ep1_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p1_fab_init_idle_exit_ack & ~p1_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep1_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep1_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p1_side_clk_valid <= 1'b0;
        if ( p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack )
          p1_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

  always_comb
    begin
      visa_p1_tier1_clk = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_clk = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport1 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( ep1_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep1_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .ism_idle            ( p1_ism_idle                   ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_ep1_pccup                 ),
  .tnpcup              ( sbr_ep1_npcup                 ),
  .tpcput              ( ep1_sbr_pcput                 ),
  .tnpput              ( ep1_sbr_npput                 ),
  .teom                ( ep1_sbr_eom                   ),
  .tpayload            ( ep1_sbr_payload               ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( ep1_sbr_pccup                 ),
  .mnpcup              ( ep1_sbr_npcup                 ),
  .mpcput              ( sbr_ep1_pcput                 ),
  .mnpput              ( sbr_ep1_npput                 ),
  .meom                ( sbr_ep1_eom                   ),
  .mpayload            ( sbr_ep1_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

// Port 2
logic p2_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p2_fab_init_idle_exit <= '0;
    else
      p2_fab_init_idle_exit <= ~agent_idle[2] & (ep2_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p2_fab_init_idle_exit_ack & ~p2_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep2_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep2_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p2_side_clk_valid <= 1'b0;
        if ( p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack )
          p2_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

  always_comb
    begin
      visa_p2_tier1_clk = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_clk = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport2 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( ep2_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep2_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .ism_idle            ( p2_ism_idle                   ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_ep2_pccup                 ),
  .tnpcup              ( sbr_ep2_npcup                 ),
  .tpcput              ( ep2_sbr_pcput                 ),
  .tnpput              ( ep2_sbr_npput                 ),
  .teom                ( ep2_sbr_eom                   ),
  .tpayload            ( ep2_sbr_payload               ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( ep2_sbr_pccup                 ),
  .mnpcup              ( ep2_sbr_npcup                 ),
  .mpcput              ( sbr_ep2_pcput                 ),
  .mnpput              ( sbr_ep2_npput                 ),
  .meom                ( sbr_ep2_eom                   ),
  .mpayload            ( sbr_ep2_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

// Port 3
logic p3_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p3_fab_init_idle_exit <= '0;
    else
      p3_fab_init_idle_exit <= ~agent_idle[3] & (ep3_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p3_fab_init_idle_exit_ack & ~p3_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep3_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep3_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p3_side_clk_valid <= 1'b0;
        if ( p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack )
          p3_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

  always_comb
    begin
      visa_p3_tier1_clk = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_clk = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport3 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p3_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( ep3_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep3_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .ism_idle            ( p3_ism_idle                   ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_ep3_pccup                 ),
  .tnpcup              ( sbr_ep3_npcup                 ),
  .tpcput              ( ep3_sbr_pcput                 ),
  .tnpput              ( ep3_sbr_npput                 ),
  .teom                ( ep3_sbr_eom                   ),
  .tpayload            ( ep3_sbr_payload               ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( ep3_sbr_pccup                 ),
  .mnpcup              ( ep3_sbr_npcup                 ),
  .mpcput              ( sbr_ep3_pcput                 ),
  .mnpput              ( sbr_ep3_npput                 ),
  .meom                ( sbr_ep3_eom                   ),
  .mpayload            ( sbr_ep3_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
logic p4_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p4_fab_init_idle_exit <= '0;
    else
      p4_fab_init_idle_exit <= ~agent_idle[4] & (ep4_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p4_fab_init_idle_exit_ack & ~p4_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep4_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep4_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p4_side_clk_valid <= 1'b0;
        if ( p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack )
          p4_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

  always_comb
    begin
      visa_p4_tier1_clk = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_clk = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport4 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( ep4_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep4_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .ism_idle            ( p4_ism_idle                   ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_ep4_pccup                 ),
  .tnpcup              ( sbr_ep4_npcup                 ),
  .tpcput              ( ep4_sbr_pcput                 ),
  .tnpput              ( ep4_sbr_npput                 ),
  .teom                ( ep4_sbr_eom                   ),
  .tpayload            ( ep4_sbr_payload               ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( ep4_sbr_pccup                 ),
  .mnpcup              ( ep4_sbr_npcup                 ),
  .mpcput              ( sbr_ep4_pcput                 ),
  .mnpput              ( sbr_ep4_npput                 ),
  .meom                ( sbr_ep4_eom                   ),
  .mpayload            ( sbr_ep4_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

// Port 5
logic p5_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p5_fab_init_idle_exit <= '0;
    else
      p5_fab_init_idle_exit <= ~agent_idle[5] & (ep5_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p5_fab_init_idle_exit_ack & ~p5_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p5_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep5_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep5_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p5_side_clk_valid <= 1'b0;
        if ( p5_fab_init_idle_exit & p5_fab_init_idle_exit_ack )
          p5_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p5_dbgbus;

  always_comb
    begin
      visa_p5_tier1_clk = { p5_dbgbus[31],
                            p5_dbgbus[27:24],
                            p5_dbgbus[21:19],
                            p5_dbgbus[15:12],
                            p5_dbgbus[7:4] };
      visa_p5_tier2_clk = { p5_dbgbus[30:28],
                            p5_dbgbus[23:22],
                            p5_dbgbus[18:16],
                            p5_dbgbus[11:8],
                            p5_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport5 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p5_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p5_side_clk_valid             ),
  .side_ism_in         ( ep5_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep5_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[5] ),
  .agent_idle          ( agent_idle[5]                 ),
  .port_idle           ( port_idle[5]                  ),
  .ism_idle            ( p5_ism_idle                   ),
  .cg_inprogress       ( p5_cg_inprogress              ),
  .tpccup              ( sbr_ep5_pccup                 ),
  .tnpcup              ( sbr_ep5_npcup                 ),
  .tpcput              ( ep5_sbr_pcput                 ),
  .tnpput              ( ep5_sbr_npput                 ),
  .teom                ( ep5_sbr_eom                   ),
  .tpayload            ( ep5_sbr_payload               ),
  .pctrdy              ( pctrdy[5]                     ),
  .pcirdy              ( pcirdy[5]                     ),
  .pcdata              ( pcdata[5]                     ),
  .pceom               ( pceom[5]                      ),
  .pcdstvld            ( p5_pcdstvld                   ),
  .nptrdy              ( nptrdy[5]                     ),
  .npirdy              ( npirdy[5]                     ),
  .npfence             ( p5_npfence                    ),
  .npdata              ( npdata[5]                     ),
  .npeom               ( npeom[5]                      ),
  .npdstvld            ( p5_npdstvld                   ),
  .mpccup              ( ep5_sbr_pccup                 ),
  .mnpcup              ( ep5_sbr_npcup                 ),
  .mpcput              ( sbr_ep5_pcput                 ),
  .mnpput              ( sbr_ep5_npput                 ),
  .meom                ( sbr_ep5_eom                   ),
  .mpayload            ( sbr_ep5_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[5]                    ),
  .enptrdy             ( enptrdy[5]                    ),
  .epcirdy             ( epcirdy[5]                    ),
  .enpirdy             ( enpirdy[5]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p5_dbgbus                     )
);

// Port 6
logic p6_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p6_fab_init_idle_exit <= '0;
    else
      p6_fab_init_idle_exit <= ~agent_idle[6] & (ep6_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p6_fab_init_idle_exit_ack & ~p6_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p6_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep6_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep6_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p6_side_clk_valid <= 1'b0;
        if ( p6_fab_init_idle_exit & p6_fab_init_idle_exit_ack )
          p6_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p6_dbgbus;

  always_comb
    begin
      visa_p6_tier1_clk = { p6_dbgbus[31],
                            p6_dbgbus[27:24],
                            p6_dbgbus[21:19],
                            p6_dbgbus[15:12],
                            p6_dbgbus[7:4] };
      visa_p6_tier2_clk = { p6_dbgbus[30:28],
                            p6_dbgbus[23:22],
                            p6_dbgbus[18:16],
                            p6_dbgbus[11:8],
                            p6_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport6 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p6_side_clk_valid             ),
  .side_ism_in         ( ep6_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep6_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[6] ),
  .agent_idle          ( agent_idle[6]                 ),
  .port_idle           ( port_idle[6]                  ),
  .ism_idle            ( p6_ism_idle                   ),
  .cg_inprogress       ( p6_cg_inprogress              ),
  .tpccup              ( sbr_ep6_pccup                 ),
  .tnpcup              ( sbr_ep6_npcup                 ),
  .tpcput              ( ep6_sbr_pcput                 ),
  .tnpput              ( ep6_sbr_npput                 ),
  .teom                ( ep6_sbr_eom                   ),
  .tpayload            ( ep6_sbr_payload               ),
  .pctrdy              ( pctrdy[6]                     ),
  .pcirdy              ( pcirdy[6]                     ),
  .pcdata              ( pcdata[6]                     ),
  .pceom               ( pceom[6]                      ),
  .pcdstvld            ( p6_pcdstvld                   ),
  .nptrdy              ( nptrdy[6]                     ),
  .npirdy              ( npirdy[6]                     ),
  .npfence             ( p6_npfence                    ),
  .npdata              ( npdata[6]                     ),
  .npeom               ( npeom[6]                      ),
  .npdstvld            ( p6_npdstvld                   ),
  .mpccup              ( ep6_sbr_pccup                 ),
  .mnpcup              ( ep6_sbr_npcup                 ),
  .mpcput              ( sbr_ep6_pcput                 ),
  .mnpput              ( sbr_ep6_npput                 ),
  .meom                ( sbr_ep6_eom                   ),
  .mpayload            ( sbr_ep6_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[6]                    ),
  .enptrdy             ( enptrdy[6]                    ),
  .epcirdy             ( epcirdy[6]                    ),
  .enpirdy             ( enpirdy[6]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p6_dbgbus                     )
);

// Port 7
logic p7_side_clk_valid;
  always_ff @(posedge clk or negedge rstb)
    if (~rstb)
      p7_fab_init_idle_exit <= '0;
    else
      p7_fab_init_idle_exit <= ~agent_idle[7] & (ep7_sbr_side_ism_agent == ISM_AGENT_IDLE) & ~p7_fab_init_idle_exit_ack & ~p7_side_clk_valid;

  always_ff @(posedge clk or negedge rstb)
    if ( ~rstb )
      p7_side_clk_valid <= 1'b0;
    else
      begin
        if ( ( ep7_sbr_side_ism_agent == ISM_AGENT_IDLEREQ ) & 
             ( sbr_ep7_side_ism_fabric == ISM_FABRIC_IDLE ) )
          p7_side_clk_valid <= 1'b0;
        if ( p7_fab_init_idle_exit & p7_fab_init_idle_exit_ack )
          p7_side_clk_valid <= 1'b1;
      end
//
// VISA tiered output assignments
//
logic [31:0] p7_dbgbus;

  always_comb
    begin
      visa_p7_tier1_clk = { p7_dbgbus[31],
                            p7_dbgbus[27:24],
                            p7_dbgbus[21:19],
                            p7_dbgbus[15:12],
                            p7_dbgbus[7:4] };
      visa_p7_tier2_clk = { p7_dbgbus[30:28],
                            p7_dbgbus[23:22],
                            p7_dbgbus[18:16],
                            p7_dbgbus[11:8],
                            p7_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        ( 15                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  1                            )
) sbcport7 (
  .side_clk            ( clk                           ),
  .gated_side_clk      ( p7_gated_clk                  ),
  .side_rst_b          ( rstb                          ),
  .side_clk_valid      ( p7_side_clk_valid             ),
  .side_ism_in         ( ep7_sbr_side_ism_agent        ),
  .side_ism_out        ( sbr_ep7_side_ism_fabric       ),
  .int_pok             ( endpoint_pwrgd[7] ),
  .agent_idle          ( agent_idle[7]                 ),
  .port_idle           ( port_idle[7]                  ),
  .ism_idle            ( p7_ism_idle                   ),
  .cg_inprogress       ( p7_cg_inprogress              ),
  .tpccup              ( sbr_ep7_pccup                 ),
  .tnpcup              ( sbr_ep7_npcup                 ),
  .tpcput              ( ep7_sbr_pcput                 ),
  .tnpput              ( ep7_sbr_npput                 ),
  .teom                ( ep7_sbr_eom                   ),
  .tpayload            ( ep7_sbr_payload               ),
  .pctrdy              ( pctrdy[7]                     ),
  .pcirdy              ( pcirdy[7]                     ),
  .pcdata              ( pcdata[7]                     ),
  .pceom               ( pceom[7]                      ),
  .pcdstvld            ( p7_pcdstvld                   ),
  .nptrdy              ( nptrdy[7]                     ),
  .npirdy              ( npirdy[7]                     ),
  .npfence             ( p7_npfence                    ),
  .npdata              ( npdata[7]                     ),
  .npeom               ( npeom[7]                      ),
  .npdstvld            ( p7_npdstvld                   ),
  .mpccup              ( ep7_sbr_pccup                 ),
  .mnpcup              ( ep7_sbr_npcup                 ),
  .mpcput              ( sbr_ep7_pcput                 ),
  .mnpput              ( sbr_ep7_npput                 ),
  .meom                ( sbr_ep7_eom                   ),
  .mpayload            ( sbr_ep7_payload               ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[7]                    ),
  .enptrdy             ( enptrdy[7]                    ),
  .epcirdy             ( epcirdy[7]                    ),
  .enpirdy             ( enpirdy[7]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p7_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

 // synopsys translate_off
    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk or negedge rstb)

      if (~rstb) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (~rstb)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk) disable iff (~rstb)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

 // synopsys translate_on
`endif
`endif

  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv0_sbr_cfg_1_ep_rtl/lv0_sbr_cfg_1_ep_rtl.csv
//
//------------------------------------------------------------------------------
/*
Endpoint, ep0,0, 1, 0, 1, 3, 3, 4, 0,1,2,3, 
Endpoint, ep1,1, 1, 0, 1, 3, 3, 4, 4,5,6,7, 
Endpoint, ep2,0, 2, 0, 1, 3, 3, 1, 8, 
Endpoint, ep3,1, 2, 0, 1, 3, 3, 1, 9, 
Endpoint, ep4,0, 1, 0, 1, 3, 3, 1, 10, 
Endpoint, ep5,1, 1, 0, 1, 3, 3, 1, 11, 
Endpoint, ep6,0, 2, 0, 1, 3, 3, 1, 12, 
Endpoint, ep7,1, 2, 0, 1, 3, 3, 1, 13, 
SyncRouter, sbr, sbr,0, 1, 0, 3, 4, 4, 0, 1, , , 0, 8, ep0, ep1, ep2, ep3, ep4, ep5, ep6, ep7, , , , , , , , , 
Multicast, 32, 4, 0,4,8,9
ClockReset, 0, clk, rstb, 0, , 1ns
PowerWell, 0, 
PowerWell, 1, pd1_pwrgd
*/
//------------------------------------------------------------------------------
