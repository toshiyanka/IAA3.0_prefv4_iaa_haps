`ifdef EP_CFG_GLS
`include "cfg_gls"
`endif
