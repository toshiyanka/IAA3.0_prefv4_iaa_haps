//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr_d : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr_d
(
  // Synchronous Clock/Reset
  clk_100,
  rst_b_100,

  // Asynchronous Clock/Reset(s)
  clk_200,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  p3_fab_init_idle_exit,
  p3_fab_init_idle_exit_ack,
  p4_fab_init_idle_exit,
  p4_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_clk_100,
  visa_vp_clk_100,
  visa_p0_tier1_clk_100,
  visa_p0_tier2_clk_100,
  visa_p1_tier1_clk_200,
  visa_p1_tier2_clk_200,
  visa_p1_ififo_tier1_clk_100,
  visa_p1_ififo_tier2_clk_100,
  visa_p1_efifo_tier1_clk_100,
  visa_p1_efifo_tier2_clk_100,
  visa_p2_tier1_clk_100,
  visa_p2_tier2_clk_100,
  visa_p3_tier1_clk_100,
  visa_p3_tier2_clk_100,
  visa_p4_tier1_clk_100,
  visa_p4_tier2_clk_100,


  // Register wires
  cfg_sbr_d_cgovrd,
  cfg_sbr_d_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  sbr_c_sbr_d_side_ism_agent,
  sbr_d_sbr_c_side_ism_fabric,
  sbr_c_sbr_d_pccup,
  sbr_c_sbr_d_npcup,
  sbr_d_sbr_c_pcput,
  sbr_d_sbr_c_npput,
  sbr_d_sbr_c_eom,
  sbr_d_sbr_c_payload,
  sbr_d_sbr_c_pccup,
  sbr_d_sbr_c_npcup,
  sbr_c_sbr_d_pcput,
  sbr_c_sbr_d_npput,
  sbr_c_sbr_d_eom,
  sbr_c_sbr_d_payload,

  // Port 1 declarations
  mcu_sbr_d_side_ism_agent,
  sbr_d_mcu_side_ism_fabric,
  mcu_sbr_d_pccup,
  mcu_sbr_d_npcup,
  sbr_d_mcu_pcput,
  sbr_d_mcu_npput,
  sbr_d_mcu_eom,
  sbr_d_mcu_payload,
  sbr_d_mcu_pccup,
  sbr_d_mcu_npcup,
  mcu_sbr_d_pcput,
  mcu_sbr_d_npput,
  mcu_sbr_d_eom,
  mcu_sbr_d_payload,

  // Port 2 declarations
  ddrio_sbr_d_side_ism_agent,
  sbr_d_ddrio_side_ism_fabric,
  ddrio_sbr_d_pccup,
  ddrio_sbr_d_npcup,
  sbr_d_ddrio_pcput,
  sbr_d_ddrio_npput,
  sbr_d_ddrio_eom,
  sbr_d_ddrio_payload,
  sbr_d_ddrio_pccup,
  sbr_d_ddrio_npcup,
  ddrio_sbr_d_pcput,
  ddrio_sbr_d_npput,
  ddrio_sbr_d_eom,
  ddrio_sbr_d_payload,

  // Port 3 declarations
  reut_0_sbr_d_side_ism_agent,
  sbr_d_reut_0_side_ism_fabric,
  reut_0_sbr_d_pccup,
  reut_0_sbr_d_npcup,
  sbr_d_reut_0_pcput,
  sbr_d_reut_0_npput,
  sbr_d_reut_0_eom,
  sbr_d_reut_0_payload,
  sbr_d_reut_0_pccup,
  sbr_d_reut_0_npcup,
  reut_0_sbr_d_pcput,
  reut_0_sbr_d_npput,
  reut_0_sbr_d_eom,
  reut_0_sbr_d_payload,

  // Port 4 declarations
  reut_1_sbr_d_side_ism_agent,
  sbr_d_reut_1_side_ism_fabric,
  reut_1_sbr_d_pccup,
  reut_1_sbr_d_npcup,
  sbr_d_reut_1_pcput,
  sbr_d_reut_1_npput,
  sbr_d_reut_1_eom,
  sbr_d_reut_1_payload,
  sbr_d_reut_1_pccup,
  sbr_d_reut_1_npcup,
  reut_1_sbr_d_pcput,
  reut_1_sbr_d_npput,
  reut_1_sbr_d_eom,
  reut_1_sbr_d_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic clk_100;
  input logic rst_b_100;

  // Asynchronous Clock/Reset(s)
  input logic clk_200;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic p3_fab_init_idle_exit;
  input logic p3_fab_init_idle_exit_ack;
  output logic p4_fab_init_idle_exit;
  input logic p4_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_clk_100;
  output visa_vp  visa_vp_clk_100;
  output visa_port_tier1 visa_p0_tier1_clk_100;
  output visa_port_tier2 visa_p0_tier2_clk_100;
  output visa_port_tier1 visa_p1_tier1_clk_200;
  output visa_port_tier2 visa_p1_tier2_clk_200;
  output visa_ififo_tier1 visa_p1_ififo_tier1_clk_100;
  output visa_ififo_tier2 visa_p1_ififo_tier2_clk_100;
  output visa_efifo_tier1 visa_p1_efifo_tier1_clk_100;
  output visa_efifo_tier2 visa_p1_efifo_tier2_clk_100;
  output visa_port_tier1 visa_p2_tier1_clk_100;
  output visa_port_tier2 visa_p2_tier2_clk_100;
  output visa_port_tier1 visa_p3_tier1_clk_100;
  output visa_port_tier2 visa_p3_tier2_clk_100;
  output visa_port_tier1 visa_p4_tier1_clk_100;
  output visa_port_tier2 visa_p4_tier2_clk_100;

  // Register wires
  input logic [4:0]  cfg_sbr_d_cgovrd;
  input logic [15:0] cfg_sbr_d_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic fscan_rstbypen;
  input logic fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] sbr_c_sbr_d_side_ism_agent;
  output logic [2:0] sbr_d_sbr_c_side_ism_fabric;
  input logic sbr_c_sbr_d_pccup;
  input logic sbr_c_sbr_d_npcup;
  output logic sbr_d_sbr_c_pcput;
  output logic sbr_d_sbr_c_npput;
  output logic sbr_d_sbr_c_eom;
  output logic [7:0] sbr_d_sbr_c_payload;
  output logic sbr_d_sbr_c_pccup;
  output logic sbr_d_sbr_c_npcup;
  input logic sbr_c_sbr_d_pcput;
  input logic sbr_c_sbr_d_npput;
  input logic sbr_c_sbr_d_eom;
  input logic [7:0] sbr_c_sbr_d_payload;

  // Port 1 declarations
  input logic [2:0] mcu_sbr_d_side_ism_agent;
  output logic [2:0] sbr_d_mcu_side_ism_fabric;
  input logic mcu_sbr_d_pccup;
  input logic mcu_sbr_d_npcup;
  output logic sbr_d_mcu_pcput;
  output logic sbr_d_mcu_npput;
  output logic sbr_d_mcu_eom;
  output logic [7:0] sbr_d_mcu_payload;
  output logic sbr_d_mcu_pccup;
  output logic sbr_d_mcu_npcup;
  input logic mcu_sbr_d_pcput;
  input logic mcu_sbr_d_npput;
  input logic mcu_sbr_d_eom;
  input logic [7:0] mcu_sbr_d_payload;

  // Port 2 declarations
  input logic [2:0] ddrio_sbr_d_side_ism_agent;
  output logic [2:0] sbr_d_ddrio_side_ism_fabric;
  input logic ddrio_sbr_d_pccup;
  input logic ddrio_sbr_d_npcup;
  output logic sbr_d_ddrio_pcput;
  output logic sbr_d_ddrio_npput;
  output logic sbr_d_ddrio_eom;
  output logic [7:0] sbr_d_ddrio_payload;
  output logic sbr_d_ddrio_pccup;
  output logic sbr_d_ddrio_npcup;
  input logic ddrio_sbr_d_pcput;
  input logic ddrio_sbr_d_npput;
  input logic ddrio_sbr_d_eom;
  input logic [7:0] ddrio_sbr_d_payload;

  // Port 3 declarations
  input logic [2:0] reut_0_sbr_d_side_ism_agent;
  output logic [2:0] sbr_d_reut_0_side_ism_fabric;
  input logic reut_0_sbr_d_pccup;
  input logic reut_0_sbr_d_npcup;
  output logic sbr_d_reut_0_pcput;
  output logic sbr_d_reut_0_npput;
  output logic sbr_d_reut_0_eom;
  output logic [7:0] sbr_d_reut_0_payload;
  output logic sbr_d_reut_0_pccup;
  output logic sbr_d_reut_0_npcup;
  input logic reut_0_sbr_d_pcput;
  input logic reut_0_sbr_d_npput;
  input logic reut_0_sbr_d_eom;
  input logic [7:0] reut_0_sbr_d_payload;

  // Port 4 declarations
  input logic [2:0] reut_1_sbr_d_side_ism_agent;
  output logic [2:0] sbr_d_reut_1_side_ism_fabric;
  input logic reut_1_sbr_d_pccup;
  input logic reut_1_sbr_d_npcup;
  output logic sbr_d_reut_1_pcput;
  output logic sbr_d_reut_1_npput;
  output logic sbr_d_reut_1_eom;
  output logic [7:0] sbr_d_reut_1_payload;
  output logic sbr_d_reut_1_pccup;
  output logic sbr_d_reut_1_npcup;
  input logic reut_1_sbr_d_pcput;
  input logic reut_1_sbr_d_npput;
  input logic reut_1_sbr_d_eom;
  input logic [7:0] reut_1_sbr_d_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr_d_sbcportmap;
always_comb sbr_d_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr_d (sbr_d)                                 SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {  107 { 17'b0_0000_0000_0000_0000 }},   //   254:148      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //   147          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   146          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //   145:144      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   143:140      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   139:136      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0000 }},   //   135:132      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //   131:128      SBCPORTMAPTABLE
      {   31 { 17'b0_0000_0000_0000_0000 }},   //   127: 97      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //    96          SBCPORTMAPTABLE
      {    6 { 17'b0_0000_0000_0000_0000 }},   //    95: 90      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    89: 88      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    87: 86      SBCPORTMAPTABLE
               17'b0_0000_0000_0001_0000,      //    85          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_1000,      //    84          SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0000 }},   //    83: 81      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //    80          SBCPORTMAPTABLE
      {   13 { 17'b0_0000_0000_0000_0000 }},   //    79: 67      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //    66: 64      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0000 }},   //    63: 59      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //    58: 56      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0000 }},   //    55: 53      SBCPORTMAPTABLE
      {    5 { 17'b0_0000_0000_0000_0001 }},   //    52: 48      SBCPORTMAPTABLE
      {    9 { 17'b0_0000_0000_0000_0000 }},   //    47: 39      SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_0000_0001 }},   //    38: 32      SBCPORTMAPTABLE
      {   14 { 17'b0_0000_0000_0000_0000 }},   //    31: 18      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //    17: 16      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //    15: 14      SBCPORTMAPTABLE
      {    4 { 17'b0_0000_0000_0000_0001 }},   //    13: 10      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     9:  8      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001,      //     7          SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0000 }},   //     6:  5      SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //     4:  2      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //     1          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0001       //     0          SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  4;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p2_pcdstvld;
logic                              p3_pcdstvld;
logic                              p4_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p2_npfence;
logic                              p3_npfence;
logic                              p4_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p2_npdstvld;
logic                              p3_npdstvld;
logic                              p4_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              p3_ism_idle;
logic                              p3_cg_inprogress;
logic                              p3_credit_reinit;
logic                              p4_ism_idle;
logic                              p4_cg_inprogress;
logic                              p4_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = cfg_sbr_d_cgctrl[15];
always_comb cfg_clkgatedef    = cfg_sbr_d_cgctrl[14];
always_comb cfg_idlecnt       = cfg_sbr_d_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = cfg_sbr_d_cgovrd[3];
always_comb jta_force_idle    = cfg_sbr_d_cgovrd[1];
always_comb jta_force_notidle = cfg_sbr_d_cgovrd[0];
always_comb jta_force_creditreq = cfg_sbr_d_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

// Asynchronous port signals
logic                              p1_clkgaten;
logic                              p1_clkgatedef;
logic                              p1_clkgate_ovrd;
logic                              p1_force_idle;
logic                              p1_force_notidle;
logic                              p1_force_creditreq;
logic                              p1_clken;
logic                              p1_gated_clk;
logic                              p1_agent_idle;
logic                              p1_eagent_idle;
logic                              p1_port_idle;
logic                              p1_ififo_idle;
logic                              p1_efifo_idle;
logic                              p1_pctrdy;
logic                              p1_pcirdy;
logic             [INTMAXPLDBIT:0] p1_pcdata;
logic                              p1_pceom;
logic                              p1_nptrdy;
logic                              p1_npirdy;
logic                              p1_npfence;
logic             [INTMAXPLDBIT:0] p1_npdata;
logic                              p1_npeom;
logic                              p1_enpstall;
logic                              p1_epctrdy;
logic                              p1_enptrdy;
logic                              p1_epcirdy;
logic                              p1_enpirdy;
logic                              p1_eom;
logic             [INTMAXPLDBIT:0] p1_data;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr_d_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr_d_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// Async clock reset synchronization
//
//------------------------------------------------------------------------------
logic clk_200_rst_b, clk_200_rst_b_pre;
sbc_doublesync sync_rst_clk_200 (
  .d     ( 1'b1 ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_200 ),
  .q     ( clk_200_rst_b_pre ));

always_comb clk_200_rst_b = fscan_rstbypen ? fscan_byprst_b : clk_200_rst_b_pre;


//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( rst_b_100                     ),
  .clk                 ( clk_100                       ),
  .q                   ( force_creditreq               )
);

sbc_doublesync sync_p1_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_force_idle                 )
);

sbc_doublesync sync_p1_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_force_notidle              )
);

sbc_doublesync sync_p1_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_force_creditreq            )
);

//------------------------------------------------------------------------------
//
// Asynchronous port local clock gating
//
//------------------------------------------------------------------------------
// Port 1
sbc_doublesync sync_p1_clkgaten (
  .d                   ( cfg_clkgaten                  ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_clkgaten                   )
);

sbc_doublesync sync_p1_clkgatedef (
  .d                   ( cfg_clkgatedef                ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_clkgatedef                 )
);

sbc_doublesync sync_p1_clkgate_ovrd (
  .d                   ( jta_clkgate_ovrd              ),
  .clr_b ( clk_200_rst_b ),
  .clk                 ( clk_200                       ),
  .q                   ( p1_clkgate_ovrd               )
);

always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if (~clk_200_rst_b)
    p1_clken <= '1;
  else
    p1_clken <= ~p1_clkgate_ovrd &
      (p1_clkgatedef | ~p1_clkgaten | ~p1_cg_inprogress |
       ((mcu_sbr_d_side_ism_agent == ISM_AGENT_ACTIVEREQ)  &
        (sbr_d_mcu_side_ism_fabric == ISM_FABRIC_ACTIVEREQ)) |
       (mcu_sbr_d_side_ism_agent == ISM_AGENT_ACTIVE)       |
       ((mcu_sbr_d_side_ism_agent == ISM_AGENT_IDLEREQ)    &
        (sbr_d_mcu_side_ism_fabric != ISM_FABRIC_IDLE)));

sbc_clock_gate p1_clkgate  (
  .en                  ( p1_clken                      ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( clk_200                       ),
  .enclk               ( p1_gated_clk                  )
);

always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          1'b1,
                          1'b1,
                          1'b1
                        };

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p4_ism_idle | ~endpoint_pwrgd[4])
                  &  (p3_ism_idle | ~endpoint_pwrgd[3])
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  &  p1_efifo_idle
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
logic p1_ism_idle_ff2, p1_ism_idle_pre;
always_ff @(posedge clk_200 or negedge clk_200_rst_b)
  if ( ~clk_200_rst_b)
    p1_ism_idle_pre <= '1;
  else
    p1_ism_idle_pre <= p1_ism_idle;

sbc_doublesync sync_idle_p1 (
  .d ( p1_ism_idle_pre ),
  .clr_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p1_ism_idle_ff2 ));

// SBR_IDLE signal for PMU
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle_ff2 &
                  p2_ism_idle &
                  p3_ism_idle &
                  p4_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p4_npfence,
                 p3_npfence,
                 p2_npfence,
                 1'b0,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p4_pcdstvld,
                 p3_pcdstvld,
                 p2_pcdstvld,
                 pcirdy[1],
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p4_npdstvld,
                 p3_npdstvld,
                 p2_npdstvld,
                 npirdy[1],
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_clk_100 = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( clk_100                       ),
  .side_rst_b          ( rst_b_100                     ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_clk_100 = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle & agent_idle[0] & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle & p0_side_clk_valid )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_clk_100 = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_clk_100 = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( sbr_c_sbr_d_side_ism_agent    ),
  .side_ism_out        ( sbr_d_sbr_c_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr_d_sbr_c_pccup             ),
  .tnpcup              ( sbr_d_sbr_c_npcup             ),
  .tpcput              ( sbr_c_sbr_d_pcput             ),
  .tnpput              ( sbr_c_sbr_d_npput             ),
  .teom                ( sbr_c_sbr_d_eom               ),
  .tpayload            ( sbr_c_sbr_d_payload           ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( sbr_c_sbr_d_pccup             ),
  .mnpcup              ( sbr_c_sbr_d_npcup             ),
  .mpcput              ( sbr_d_sbr_c_pcput             ),
  .mnpput              ( sbr_d_sbr_c_npput             ),
  .meom                ( sbr_d_sbr_c_eom               ),
  .mpayload            ( sbr_d_sbr_c_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1 (Asynchronous port)
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  logic p1_credit_reinit_ff2;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit_ff2 & p1_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & (~agent_idle[1] || ~p1_efifo_idle) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle_ff2 & agent_idle[1] & p1_efifo_idle & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle_ff2 & p1_side_clk_valid & ~p1_fab_init_idle_exit )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle_ff2 )
          p1_side_clk_valid <= '1;
      end

logic p1_side_clk_valid_ff2;
sbc_doublesync sync_p1_clk_valid (
  .d     ( p1_side_clk_valid ),
  .clr_b ( clk_200_rst_b ),
  .clk   ( clk_200 ),
  .q     ( p1_side_clk_valid_ff2 ));

sbc_doublesync_set sync_p1_credit_reinit (
  .d     ( p1_credit_reinit ),
  .set_b ( rst_b_100 ),
  .clk   ( clk_100 ),
  .q     ( p1_credit_reinit_ff2 ));

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

logic [15:0] p1_dbgbus_ing;
logic [15:0] p1_dbgbus_egr;
  always_comb
    begin
      visa_p1_tier1_clk_200 = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_clk_200 = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
      visa_p1_ififo_tier1_clk_100 = { p1_dbgbus_ing[15:14],
                             p1_dbgbus_ing[5:0]};
      visa_p1_ififo_tier2_clk_100 = { p1_dbgbus_ing[13:6] };
      visa_p1_efifo_tier1_clk_100 = { p1_dbgbus_egr[7:0] };
      visa_p1_efifo_tier2_clk_100 = { p1_dbgbus_egr[15:8] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( clk_200                       ),
  .gated_side_clk      ( p1_gated_clk                  ),
  .side_rst_b ( clk_200_rst_b ),
  .side_clk_valid      ( p1_side_clk_valid_ff2         ),
  .side_ism_in         ( mcu_sbr_d_side_ism_agent      ),
  .side_ism_out        ( sbr_d_mcu_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( p1_agent_idle                 ),
  .port_idle           ( p1_port_idle                  ),
  .idle_egress         (                               ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr_d_mcu_pccup               ),
  .tnpcup              ( sbr_d_mcu_npcup               ),
  .tpcput              ( mcu_sbr_d_pcput               ),
  .tnpput              ( mcu_sbr_d_npput               ),
  .teom                ( mcu_sbr_d_eom                 ),
  .tpayload            ( mcu_sbr_d_payload             ),
  .pctrdy              ( p1_pctrdy                     ),
  .pcirdy              ( p1_pcirdy                     ),
  .pcdata              ( p1_pcdata                     ),
  .pceom               ( p1_pceom                      ),
  .pcdstvld            (                               ),
  .nptrdy              ( p1_nptrdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( p1_npdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdstvld            (                               ),
  .mpccup              ( mcu_sbr_d_pccup               ),
  .mnpcup              ( mcu_sbr_d_npcup               ),
  .mpcput              ( sbr_d_mcu_pcput               ),
  .mnpput              ( sbr_d_mcu_npput               ),
  .meom                ( sbr_d_mcu_eom                 ),
  .mpayload            ( sbr_d_mcu_payload             ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .data                ( p1_data                       ),
  .eom                 ( p1_eom                        ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( p1_clkgaten                   ),
  .force_idle          ( p1_force_idle                 ),
  .force_notidle       ( p1_force_notidle              ),
  .force_creditreq     ( p1_force_creditreq            ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         ( 10                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  0                            ),
  .EGRSYNCROUTER       (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncingress1 (
  .ing_side_clk        ( p1_gated_clk                  ),
  .ing_side_rst_b ( clk_200_rst_b ),
  .port_idle           ( p1_port_idle                  ),
  .pcirdy              ( p1_pcirdy                     ),
  .npirdy              ( p1_npirdy                     ),
  .npfence             ( p1_npfence                    ),
  .pceom               ( p1_pceom                      ),
  .pcdata              ( p1_pcdata                     ),
  .npeom               ( p1_npeom                      ),
  .npdata              ( p1_npdata                     ),
  .pctrdy              ( p1_pctrdy                     ),
  .nptrdy              ( p1_nptrdy                     ),
  .npstall             (                               ),
  .fifo_idle           ( p1_ififo_idle                 ),
  .egr_side_clk        ( clk_100                       ),
  .gated_egr_side_clk  ( gated_side_clk                ),
  .egr_side_rst_b      ( rst_b_100                     ),
  .enpstall            ( 1'b0                          ),
  .epctrdy             ( pctrdy[1]                     ),
  .enptrdy             ( nptrdy[1]                     ),
  .epcirdy             ( pcirdy[1]                     ),
  .enpirdy             ( npirdy[1]                     ),
  .eom                 ( npeom[1]                      ),
  .data                ( npdata[1]                     ),
  .opceom              ( pceom[1]                      ),
  .opcdata             ( pcdata[1]                     ),
  .agent_idle          ( port_idle[1]                  ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           (                               ),
  .dbgbus_out          ( p1_dbgbus_ing                 )
);

sbcasyncfifo #(
  .ASYNCQDEPTH         (  4                            ),
  .MAXPLDBIT           ( INTMAXPLDBIT                  ),
  .INGSYNCROUTER       (  1                            ),
  .EGRSYNCROUTER       (  0                            ),
  .LATCHQUEUES         (  0                            )
) sbcasyncegress1 (
  .ing_side_clk        ( clk_100                       ),
  .ing_side_rst_b      ( rst_b_100                     ),
  .port_idle           ( agent_idle[1]                 ),
  .pcirdy              ( epcirdy[1]                    ),
  .npirdy              ( enpirdy[1]                    ),
  .npfence             ( 1'b0                          ),
  .pceom               ( eom                           ),
  .pcdata              ( data                          ),
  .npeom               ( eom                           ),
  .npdata              ( data                          ),
  .pctrdy              ( epctrdy[1]                    ),
  .nptrdy              ( enptrdy[1]                    ),
  .npstall             (                               ),
  .fifo_idle           ( p1_efifo_idle                 ),
  .egr_side_clk        ( clk_200                       ),
  .gated_egr_side_clk  ( p1_gated_clk                  ),
  .egr_side_rst_b ( clk_200_rst_b ),
  .enpstall            ( p1_enpstall                   ),
  .epctrdy             ( p1_epctrdy                    ),
  .enptrdy             ( p1_enptrdy                    ),
  .epcirdy             ( p1_epcirdy                    ),
  .enpirdy             ( p1_enpirdy                    ),
  .eom                 ( p1_eom                        ),
  .data                ( p1_data                       ),
  .opceom              (                               ),
  .opcdata             (                               ),
  .agent_idle          ( p1_eagent_idle                ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus_in           ( p1_dbgbus_egr                 ),
  .dbgbus_out          (                               )
);

always_comb p1_agent_idle  = p1_eagent_idle & p1_ififo_idle;

// Port 2
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit & p2_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle & (~agent_idle[2] || ~p2_idle_egress) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle & agent_idle[2] & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle & p2_side_clk_valid )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle )
          p2_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

  always_comb
    begin
      visa_p2_tier1_clk_100 = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_clk_100 = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( ddrio_sbr_d_side_ism_agent    ),
  .side_ism_out        ( sbr_d_ddrio_side_ism_fabric   ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .idle_egress         ( p2_idle_egress                ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr_d_ddrio_pccup             ),
  .tnpcup              ( sbr_d_ddrio_npcup             ),
  .tpcput              ( ddrio_sbr_d_pcput             ),
  .tnpput              ( ddrio_sbr_d_npput             ),
  .teom                ( ddrio_sbr_d_eom               ),
  .tpayload            ( ddrio_sbr_d_payload           ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( ddrio_sbr_d_pccup             ),
  .mnpcup              ( ddrio_sbr_d_npcup             ),
  .mpcput              ( sbr_d_ddrio_pcput             ),
  .mnpput              ( sbr_d_ddrio_npput             ),
  .meom                ( sbr_d_ddrio_eom               ),
  .mpayload            ( sbr_d_ddrio_payload           ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

// Port 3
logic p3_side_clk_valid, p3_idle_egress, p3_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_rst_suppress <= 1'b1;
    else
      p3_rst_suppress <= p3_credit_reinit & p3_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p3_fab_init_idle_exit <= '1;
    else
      if ( ~p3_rst_suppress & (p3_ism_idle & (~agent_idle[3] || ~p3_idle_egress) & ~p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '1;
      else if ( ~p3_rst_suppress & (p3_ism_idle & agent_idle[3] & p3_fab_init_idle_exit_ack ))
        p3_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p3_side_clk_valid <= 1'b0;
    else
      begin
        if ( p3_ism_idle & p3_side_clk_valid )
          p3_side_clk_valid <= '0;
        else if ( (p3_fab_init_idle_exit & p3_fab_init_idle_exit_ack) || ~p3_ism_idle )
          p3_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p3_dbgbus;

  always_comb
    begin
      visa_p3_tier1_clk_100 = { p3_dbgbus[31],
                            p3_dbgbus[27:24],
                            p3_dbgbus[21:19],
                            p3_dbgbus[15:12],
                            p3_dbgbus[7:4] };
      visa_p3_tier2_clk_100 = { p3_dbgbus[30:28],
                            p3_dbgbus[23:22],
                            p3_dbgbus[18:16],
                            p3_dbgbus[11:8],
                            p3_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport3 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p3_side_clk_valid             ),
  .side_ism_in         ( reut_0_sbr_d_side_ism_agent   ),
  .side_ism_out        ( sbr_d_reut_0_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[3] ),
  .agent_idle          ( agent_idle[3]                 ),
  .port_idle           ( port_idle[3]                  ),
  .idle_egress         ( p3_idle_egress                ),
  .ism_idle            ( p3_ism_idle                   ),
  .credit_reinit       ( p3_credit_reinit              ),
  .cg_inprogress       ( p3_cg_inprogress              ),
  .tpccup              ( sbr_d_reut_0_pccup            ),
  .tnpcup              ( sbr_d_reut_0_npcup            ),
  .tpcput              ( reut_0_sbr_d_pcput            ),
  .tnpput              ( reut_0_sbr_d_npput            ),
  .teom                ( reut_0_sbr_d_eom              ),
  .tpayload            ( reut_0_sbr_d_payload          ),
  .pctrdy              ( pctrdy[3]                     ),
  .pcirdy              ( pcirdy[3]                     ),
  .pcdata              ( pcdata[3]                     ),
  .pceom               ( pceom[3]                      ),
  .pcdstvld            ( p3_pcdstvld                   ),
  .nptrdy              ( nptrdy[3]                     ),
  .npirdy              ( npirdy[3]                     ),
  .npfence             ( p3_npfence                    ),
  .npdata              ( npdata[3]                     ),
  .npeom               ( npeom[3]                      ),
  .npdstvld            ( p3_npdstvld                   ),
  .mpccup              ( reut_0_sbr_d_pccup            ),
  .mnpcup              ( reut_0_sbr_d_npcup            ),
  .mpcput              ( sbr_d_reut_0_pcput            ),
  .mnpput              ( sbr_d_reut_0_npput            ),
  .meom                ( sbr_d_reut_0_eom              ),
  .mpayload            ( sbr_d_reut_0_payload          ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[3]                    ),
  .enptrdy             ( enptrdy[3]                    ),
  .epcirdy             ( epcirdy[3]                    ),
  .enpirdy             ( enpirdy[3]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p3_dbgbus                     )
);

// Port 4
logic p4_side_clk_valid, p4_idle_egress, p4_rst_suppress;
  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_rst_suppress <= 1'b1;
    else
      p4_rst_suppress <= p4_credit_reinit & p4_rst_suppress;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if (~rst_b_100)
      p4_fab_init_idle_exit <= '1;
    else
      if ( ~p4_rst_suppress & (p4_ism_idle & (~agent_idle[4] || ~p4_idle_egress) & ~p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '1;
      else if ( ~p4_rst_suppress & (p4_ism_idle & agent_idle[4] & p4_fab_init_idle_exit_ack ))
        p4_fab_init_idle_exit <= '0;

  always_ff @(posedge clk_100 or negedge rst_b_100)
    if ( ~rst_b_100 )
      p4_side_clk_valid <= 1'b0;
    else
      begin
        if ( p4_ism_idle & p4_side_clk_valid )
          p4_side_clk_valid <= '0;
        else if ( (p4_fab_init_idle_exit & p4_fab_init_idle_exit_ack) || ~p4_ism_idle )
          p4_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p4_dbgbus;

  always_comb
    begin
      visa_p4_tier1_clk_100 = { p4_dbgbus[31],
                            p4_dbgbus[27:24],
                            p4_dbgbus[21:19],
                            p4_dbgbus[15:12],
                            p4_dbgbus[7:4] };
      visa_p4_tier2_clk_100 = { p4_dbgbus[30:28],
                            p4_dbgbus[23:22],
                            p4_dbgbus[18:16],
                            p4_dbgbus[11:8],
                            p4_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport4 (
  .side_clk            ( clk_100                       ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( rst_b_100                     ),
  .side_clk_valid      ( p4_side_clk_valid             ),
  .side_ism_in         ( reut_1_sbr_d_side_ism_agent   ),
  .side_ism_out        ( sbr_d_reut_1_side_ism_fabric  ),
  .int_pok             ( endpoint_pwrgd[4] ),
  .agent_idle          ( agent_idle[4]                 ),
  .port_idle           ( port_idle[4]                  ),
  .idle_egress         ( p4_idle_egress                ),
  .ism_idle            ( p4_ism_idle                   ),
  .credit_reinit       ( p4_credit_reinit              ),
  .cg_inprogress       ( p4_cg_inprogress              ),
  .tpccup              ( sbr_d_reut_1_pccup            ),
  .tnpcup              ( sbr_d_reut_1_npcup            ),
  .tpcput              ( reut_1_sbr_d_pcput            ),
  .tnpput              ( reut_1_sbr_d_npput            ),
  .teom                ( reut_1_sbr_d_eom              ),
  .tpayload            ( reut_1_sbr_d_payload          ),
  .pctrdy              ( pctrdy[4]                     ),
  .pcirdy              ( pcirdy[4]                     ),
  .pcdata              ( pcdata[4]                     ),
  .pceom               ( pceom[4]                      ),
  .pcdstvld            ( p4_pcdstvld                   ),
  .nptrdy              ( nptrdy[4]                     ),
  .npirdy              ( npirdy[4]                     ),
  .npfence             ( p4_npfence                    ),
  .npdata              ( npdata[4]                     ),
  .npeom               ( npeom[4]                      ),
  .npdstvld            ( p4_npdstvld                   ),
  .mpccup              ( reut_1_sbr_d_pccup            ),
  .mnpcup              ( reut_1_sbr_d_npcup            ),
  .mpcput              ( sbr_d_reut_1_pcput            ),
  .mnpput              ( sbr_d_reut_1_npput            ),
  .meom                ( sbr_d_reut_1_eom              ),
  .mpayload            ( sbr_d_reut_1_payload          ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[4]                    ),
  .enptrdy             ( enptrdy[4]                    ),
  .epcirdy             ( epcirdy[4]                    ),
  .enpirdy             ( enpirdy[4]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p4_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr_d_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr_d_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge clk_100 or negedge rst_b_100)

      if (~rst_b_100) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge clk_100) disable iff (rst_b_100 !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_9_BVL/lv2_sbn_cfg_9_BVL.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 1, clk_100, rst_b_100, 0, , 5ns
ClockReset, 0, clk_200, rst_b_200, 0, , 2.5ns
ClockReset, 2, clk_27, rst_b_27, 0, , 18.5ns
Endpoint, SAPms,3, 1, 1, 0, 3, 3, 1, 65, 2, 2, 
Endpoint, adac,0, 1, 1, 0, 3, 3, 1, 129, 2, 2, 
Endpoint, apll,0, 1, 2, 0, 3, 3, 1, 139, 2, 2, 
Endpoint, bunit,2, 1, 0, 0, 3, 3, 1, 03, 2, 2, 
Endpoint, cpunit,2, 1, 1, 0, 3, 3, 1, 10, 2, 2, 
Endpoint, cunit,2, 1, 0, 0, 3, 3, 1, 07, 2, 2, 
Endpoint, ddrio,2, 1, 1, 0, 3, 3, 1, 80, 2, 2, 
Endpoint, dfx_jtag,2, 1, 1, 0, 3, 3, 1, 58, 2, 2, 
Endpoint, dfx_lakemore,2, 1, 1, 0, 3, 3, 1, 56, 2, 2, 
Endpoint, dfx_omar,2, 1, 1, 0, 3, 3, 1, 57, 2, 2, 
Endpoint, dpll,0, 1, 2, 0, 3, 3, 1, 138, 2, 2, 
Endpoint, fpll,0, 1, 2, 0, 3, 3, 1, 136, 2, 2, 
Endpoint, hdmi_rx,0, 1, 1, 0, 3, 3, 1, 131, 2, 2, 
Endpoint, hdmi_tx,0, 1, 1, 0, 3, 3, 1, 130, 2, 2, 
Endpoint, hpll,0, 1, 2, 0, 3, 3, 1, 137, 2, 2, 
Endpoint, hunit,2, 1, 0, 0, 3, 3, 1, 02, 2, 2, 
Endpoint, itunit,2, 1, 1, 0, 3, 3, 1, 64, 2, 2, 
Endpoint, itunit2,2, 1, 1, 0, 3, 3, 1, 66, 2, 2, 
Endpoint, legacy,2, 1, 1, 0, 3, 3, 10, 11,12,13,32,33,34,35,36,37,38, 2, 2, 
Endpoint, mcu,2, 1, 0, 0, 3, 3, 1, 01, 2, 2, 
Endpoint, pcie_afe,4, 1, 1, 0, 3, 3, 1, 17, 2, 2, 
Endpoint, pcie_ctrl,4, 1, 1, 0, 3, 3, 1, 16, 2, 2, 
Endpoint, psf_0_north,4, 1, 0, 0, 3, 3, 1, 50, 2, 2, 
Endpoint, psf_0_south,4, 1, 1, 0, 3, 3, 1, 144, 2, 2, 
Endpoint, psf_1,4, 1, 0, 0, 3, 3, 1, 145, 2, 2, 
Endpoint, psf_3,2, 1, 0, 0, 3, 3, 1, 147, 2, 2, 
Endpoint, punit,1, 1, 2, 0, 3, 3, 1, 04, 2, 2, 
Endpoint, reut_0,2, 1, 1, 0, 3, 3, 1, 84, 2, 2, 
Endpoint, reut_1,2, 1, 1, 0, 3, 3, 1, 85, 2, 2, 
Endpoint, sata_afe,4, 1, 1, 0, 3, 3, 1, 89, 2, 2, 
Endpoint, sata_ctrl,4, 1, 1, 0, 3, 3, 1, 88, 2, 2, 
SyncRouter, sbr_a, sbr_a,1, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 2, 8, sbr_e, sbr_b, sbr_c, dpll, apll, hpll, fpll, punit, , , , , , , , , 
RouterAgentPort, sbr_a, 0
RouterAgentPort, sbr_a, 1
RouterAgentPort, sbr_a, 2
RouterRange, sbr_a, 0, 48,49
SyncRouter, sbr_b, sbr_b,4, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 9, sbr_a, pcie_afe, sata_afe, usb_afe, sata_ctrl, pcie_ctrl, psf_1, psf_0_south, psf_0_north, , , , , , , , 
RouterRange, sbr_b, 0, 51,51
SyncRouter, sbr_c, sbr_c,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 15, sbr_a, sbr_d, vtunit, hunit, bunit, cunit, cpunit, legacy, dfx_lakemore, dfx_omar, dfx_jtag, itunit, psf_3, SAPms, itunit2, , 
RouterAgentPort, sbr_c, 1
RouterRange, sbr_c, 0, 52,52
SyncRouter, sbr_d, sbr_d,2, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_c, mcu, ddrio, reut_0, reut_1, , , , , , , , , , , , 
RouterRange, sbr_d, 0, 54,55
SyncRouter, sbr_e, sbr_e,5, 0, 0, 3, 4, 1, 0, 1, visa, cfg, 1, 5, sbr_a, vdac, adac, hdmi_tx, hdmi_rx, , , , , , , , , , , , 
Endpoint, usb_afe,4, 1, 1, 0, 3, 3, 1, 96, 2, 2, 
Endpoint, vdac,0, 1, 1, 0, 3, 3, 1, 128, 2, 2, 
Endpoint, vtunit,2, 1, 0, 0, 3, 3, 1, 00, 2, 2, 
AsyncPort, sbr_a, 0, 10, 4, 0, 
AsyncPort, sbr_a, 1, 10, 4, 0, 
AsyncPort, sbr_a, 2, 10, 4, 0, 
AsyncPort, sbr_b, 6, 4, 2, 0, 
AsyncPort, sbr_b, 8, 4, 2, 0, 
AsyncPort, sbr_c, 12, 4, 2, 0, 
AsyncPort, sbr_c, 2, 10, 4, 0, 
AsyncPort, sbr_c, 3, 10, 4, 0, 
AsyncPort, sbr_c, 4, 10, 4, 0, 
AsyncPort, sbr_c, 5, 10, 4, 0, 
AsyncPort, sbr_d, 1, 10, 4, 0, 
PowerWell, 0, 
PowerWell, 1, island0_pok
PowerWell, 2, island1_pok
PowerWell, 3, island2_pok
PowerWell, 4, island3_pok
PowerWell, 5, island8_pok
*/
//------------------------------------------------------------------------------
