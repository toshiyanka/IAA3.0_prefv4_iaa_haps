typedef enum int {
	   cltap           =  'd0,
      dfx_aggregator           = 'd1,
      stap0           = 'd2,
      stap1           = 'd3,
      stap3           = 'd4,
      stap4           = 'd5,
      stap5           = 'd6,
      stap6           = 'd7,
      stap7           = 'd8,
      stap8           = 'd9,
      stap_extr           = 'd10,
      stap_extr3           = 'd11,
      stap_extr4           = 'd12,
      stap_extr1           = 'd13,
      stap_extr2           = 'd14,
      NOTAP           = 'hFFFF_FFFF
} Tap_t;
