VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf132b032e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  FOREIGN arf132b032e1r1w0cbbehbaa4acw ;
  ORIGIN 0 0 ;
  SIZE 19.8 BY 29.76 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 16.68 10.928 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.184 14.76 8.228 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 16.68 11.828 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 16.68 6.772 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 16.68 7.028 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 16.68 7.116 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.284 16.68 7.328 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 16.68 11.016 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 16.68 11.272 17.88 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 16.68 11.528 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 16.68 11.616 17.88 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 14.76 9.728 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 14.76 9.816 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 14.76 10.028 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 14.76 10.628 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 14.76 10.716 15.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.272 14.76 8.316 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 14.76 8.828 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 0.24 8.916 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 22.56 8.828 23.76 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 22.56 8.916 23.76 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 22.56 10.628 23.76 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 22.56 10.028 23.76 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 23.28 8.572 24.48 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 23.28 9.128 24.48 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 23.28 10.116 24.48 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 23.28 10.372 24.48 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 24 9.216 25.2 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 24 9.472 25.2 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 1.68 10.628 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 24 9.728 25.2 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 24 9.816 25.2 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 24.72 8.828 25.92 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 24.72 8.916 25.92 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 24.72 10.628 25.92 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 24.72 10.028 25.92 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 25.44 8.572 26.64 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 25.44 9.128 26.64 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 25.44 10.116 26.64 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 25.44 10.372 26.64 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 1.68 10.028 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 26.16 9.216 27.36 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 26.16 9.472 27.36 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 26.16 9.728 27.36 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 26.16 9.816 27.36 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 26.88 8.828 28.08 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 26.88 8.916 28.08 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 26.88 10.628 28.08 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 26.88 10.028 28.08 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 27.6 8.572 28.8 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 27.6 9.128 28.8 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 2.4 8.572 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 27.6 10.116 28.8 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 27.6 10.372 28.8 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 28.32 9.216 29.52 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 28.32 9.472 29.52 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 28.32 9.728 29.52 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 28.32 9.816 29.52 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 2.4 9.128 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 2.4 10.116 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 2.4 10.372 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 3.12 9.216 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 3.12 9.472 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 3.12 9.728 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 3.12 9.816 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 0.24 9.128 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 3.84 8.828 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 3.84 8.916 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 3.84 10.628 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 3.84 10.028 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 4.56 8.572 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 4.56 9.128 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 4.56 10.116 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 4.56 10.372 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 5.28 9.216 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 5.28 9.472 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.24 10.372 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 5.28 9.728 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 5.28 9.816 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 6 8.828 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 6 8.916 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 6 10.628 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 6 10.028 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 6.72 8.572 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 6.72 9.128 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 6.72 10.116 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 6.72 10.372 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 0.24 10.628 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 7.44 9.216 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 7.44 9.472 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 7.44 9.728 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 7.44 9.816 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 8.16 8.828 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 8.16 8.916 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 8.16 10.628 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 8.16 10.028 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 8.88 8.572 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 8.88 9.128 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 0.96 9.216 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 8.88 10.116 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 8.88 10.372 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 9.6 9.216 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 9.6 9.472 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 9.6 9.728 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 9.6 9.816 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 10.32 8.828 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 10.32 8.916 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 10.32 10.628 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 10.32 10.028 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 0.96 9.472 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 11.04 8.572 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 11.04 9.128 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 11.04 10.116 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 11.04 10.372 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 11.76 9.216 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 11.76 9.472 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 11.76 9.728 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 11.76 9.816 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 12.48 8.828 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 12.48 8.916 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 0.96 9.728 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 12.48 10.628 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 12.48 10.028 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 13.2 8.572 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 13.2 9.128 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 13.2 10.116 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 13.2 10.372 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 18.24 8.916 19.44 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 18.24 9.128 19.44 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 18.24 10.372 19.44 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 18.24 10.628 19.44 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 0.96 9.816 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 18.96 8.572 20.16 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 18.96 8.828 20.16 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 18.96 10.028 20.16 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 18.96 10.116 20.16 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 19.68 9.216 20.88 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 19.68 9.472 20.88 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 19.68 9.728 20.88 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 19.68 9.816 20.88 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 20.4 8.828 21.6 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 20.4 8.916 21.6 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.784 1.68 8.828 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 20.4 10.628 21.6 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 20.4 10.028 21.6 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.528 21.12 8.572 22.32 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.084 21.12 9.128 22.32 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 21.12 10.116 22.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 21.12 10.372 22.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 21.84 9.216 23.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 21.84 9.472 23.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.684 21.84 9.728 23.04 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.772 21.84 9.816 23.04 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 1.68 8.916 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.172 14.76 9.216 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.428 14.76 9.472 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 8.872 14.76 8.916 15.96 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 0.24 6.772 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 22.56 7.928 23.76 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 22.56 7.116 23.76 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 22.56 11.016 23.76 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 22.56 11.616 23.76 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 23.28 7.416 24.48 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 23.28 7.672 24.48 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 23.28 11.916 24.48 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 23.28 12.172 24.48 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 24 6.772 25.2 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 24 7.028 25.2 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 1.68 11.016 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 24 11.272 25.2 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 24 11.528 25.2 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 24.72 7.928 25.92 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 24.72 7.116 25.92 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 24.72 11.016 25.92 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 24.72 11.616 25.92 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 25.44 7.416 26.64 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 25.44 7.672 26.64 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 25.44 11.916 26.64 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 25.44 12.172 26.64 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 1.68 11.616 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 26.16 6.772 27.36 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 26.16 7.028 27.36 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 26.16 11.272 27.36 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 26.16 11.528 27.36 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 26.88 7.928 28.08 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 26.88 7.116 28.08 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 26.88 11.016 28.08 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 26.88 11.616 28.08 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 27.6 7.416 28.8 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 27.6 7.672 28.8 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 2.4 7.416 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 27.6 11.916 28.8 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 27.6 12.172 28.8 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 28.32 6.772 29.52 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 28.32 7.028 29.52 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 28.32 11.272 29.52 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 28.32 11.528 29.52 ;
    END
  END rddatap0[135]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 2.4 7.672 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 2.4 11.916 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 2.4 12.172 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 3.12 6.772 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 3.12 7.028 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 3.12 11.272 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 3.12 11.528 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 0.24 7.028 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 3.84 7.928 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 3.84 7.116 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 3.84 11.016 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 3.84 11.616 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 4.56 7.416 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 4.56 7.672 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 4.56 11.916 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 4.56 12.172 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 5.28 6.772 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 5.28 7.028 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 0.24 11.916 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 5.28 11.272 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 5.28 11.528 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 6 7.928 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 6 7.116 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 6 11.016 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 6 11.616 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 6.72 7.416 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 6.72 7.672 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 6.72 11.916 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 6.72 12.172 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 0.24 12.172 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 7.44 6.772 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 7.44 7.028 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 7.44 11.272 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 7.44 11.528 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 8.16 7.928 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 8.16 7.116 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 8.16 11.016 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 8.16 11.616 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 8.88 7.416 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 8.88 7.672 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 0.96 7.116 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 8.88 11.916 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 8.88 12.172 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 9.6 6.772 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 9.6 7.028 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 9.6 11.272 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 9.6 11.528 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 10.32 7.928 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 10.32 7.116 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 10.32 11.016 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 10.32 11.616 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.284 0.96 7.328 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 11.04 7.416 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 11.04 7.672 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 11.04 11.916 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 11.04 12.172 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 11.76 6.772 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 11.76 7.028 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 11.76 11.272 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 11.76 11.528 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 12.48 7.928 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 12.48 7.116 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 0.96 11.272 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 12.48 11.016 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 12.48 11.616 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 13.2 7.416 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 13.2 7.672 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 13.2 11.916 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 13.2 12.172 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 18.24 7.416 19.44 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 18.24 7.672 19.44 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 18.24 11.916 19.44 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 18.24 12.172 19.44 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 0.96 11.528 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 18.96 7.116 20.16 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.284 18.96 7.328 20.16 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 18.96 11.616 20.16 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 18.96 11.828 20.16 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 19.68 6.772 20.88 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 19.68 7.028 20.88 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 19.68 11.272 20.88 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 19.68 11.528 20.88 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 20.4 7.928 21.6 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.072 20.4 7.116 21.6 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.884 1.68 7.928 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 20.4 11.016 21.6 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 20.4 11.616 21.6 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.372 21.12 7.416 22.32 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 7.628 21.12 7.672 22.32 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 21.12 11.916 22.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 21.12 12.172 22.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 21.84 6.772 23.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 21.84 7.028 23.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 21.84 11.272 23.04 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 21.84 11.528 23.04 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 1.68 6.772 2.88 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 29.7 ;
        RECT 2.662 0.06 2.738 29.7 ;
        RECT 4.462 0.06 4.538 29.7 ;
        RECT 6.262 0.06 6.338 29.7 ;
        RECT 8.062 0.06 8.138 29.7 ;
        RECT 9.862 0.06 9.938 29.7 ;
        RECT 11.662 0.06 11.738 29.7 ;
        RECT 13.462 0.06 13.538 29.7 ;
        RECT 15.262 0.06 15.338 29.7 ;
        RECT 17.062 0.06 17.138 29.7 ;
        RECT 18.862 0.06 18.938 29.7 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 29.7 ;
        RECT 3.562 0.06 3.638 29.7 ;
        RECT 5.362 0.06 5.438 29.7 ;
        RECT 7.162 0.06 7.238 29.7 ;
        RECT 8.962 0.06 9.038 29.7 ;
        RECT 10.762 0.06 10.838 29.7 ;
        RECT 12.562 0.06 12.638 29.7 ;
        RECT 14.362 0.06 14.438 29.7 ;
        RECT 16.162 0.06 16.238 29.7 ;
        RECT 17.962 0.06 18.038 29.7 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 19.816 29.774 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 19.82 29.78 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 19.8705 29.798 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 19.835 29.83 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 19.87 29.798 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 19.859 29.85 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 19.89 29.822 ;
    LAYER m7 SPACING 0 ;
      RECT 18.938 29.82 19.84 29.88 ;
      RECT 18.938 -0.06 19.892 29.82 ;
      RECT 18.938 -0.12 19.84 -0.06 ;
      RECT 18.038 -0.12 18.862 29.88 ;
      RECT 17.138 -0.12 17.962 29.88 ;
      RECT 16.238 -0.12 17.062 29.88 ;
      RECT 15.338 -0.12 16.162 29.88 ;
      RECT 14.438 -0.12 15.262 29.88 ;
      RECT 13.538 -0.12 14.362 29.88 ;
      RECT 12.638 -0.12 13.462 29.88 ;
      RECT 11.738 28.8 12.562 29.88 ;
      RECT 11.738 27.6 11.872 28.8 ;
      RECT 11.916 27.6 12.128 28.8 ;
      RECT 12.172 27.6 12.562 28.8 ;
      RECT 11.738 26.64 12.562 27.6 ;
      RECT 11.738 25.44 11.872 26.64 ;
      RECT 11.916 25.44 12.128 26.64 ;
      RECT 12.172 25.44 12.562 26.64 ;
      RECT 11.738 24.48 12.562 25.44 ;
      RECT 11.738 23.28 11.872 24.48 ;
      RECT 11.916 23.28 12.128 24.48 ;
      RECT 12.172 23.28 12.562 24.48 ;
      RECT 11.738 22.32 12.562 23.28 ;
      RECT 11.738 21.12 11.872 22.32 ;
      RECT 11.916 21.12 12.128 22.32 ;
      RECT 12.172 21.12 12.562 22.32 ;
      RECT 11.738 20.16 12.562 21.12 ;
      RECT 11.828 19.44 12.562 20.16 ;
      RECT 11.738 18.96 11.784 20.16 ;
      RECT 11.828 18.96 11.872 19.44 ;
      RECT 11.916 18.24 12.128 19.44 ;
      RECT 12.172 18.24 12.562 19.44 ;
      RECT 11.738 18.24 11.872 18.96 ;
      RECT 11.738 17.88 12.562 18.24 ;
      RECT 11.738 16.68 11.784 17.88 ;
      RECT 11.828 16.68 12.562 17.88 ;
      RECT 11.738 14.4 12.562 16.68 ;
      RECT 11.738 13.2 11.872 14.4 ;
      RECT 11.916 13.2 12.128 14.4 ;
      RECT 12.172 13.2 12.562 14.4 ;
      RECT 11.738 12.24 12.562 13.2 ;
      RECT 11.738 11.04 11.872 12.24 ;
      RECT 11.916 11.04 12.128 12.24 ;
      RECT 12.172 11.04 12.562 12.24 ;
      RECT 11.738 10.08 12.562 11.04 ;
      RECT 11.738 8.88 11.872 10.08 ;
      RECT 11.916 8.88 12.128 10.08 ;
      RECT 12.172 8.88 12.562 10.08 ;
      RECT 11.738 7.92 12.562 8.88 ;
      RECT 11.738 6.72 11.872 7.92 ;
      RECT 11.916 6.72 12.128 7.92 ;
      RECT 12.172 6.72 12.562 7.92 ;
      RECT 11.738 5.76 12.562 6.72 ;
      RECT 11.738 4.56 11.872 5.76 ;
      RECT 11.916 4.56 12.128 5.76 ;
      RECT 12.172 4.56 12.562 5.76 ;
      RECT 11.738 3.6 12.562 4.56 ;
      RECT 11.738 2.4 11.872 3.6 ;
      RECT 11.916 2.4 12.128 3.6 ;
      RECT 12.172 2.4 12.562 3.6 ;
      RECT 11.738 1.44 12.562 2.4 ;
      RECT 11.738 0.24 11.872 1.44 ;
      RECT 11.916 0.24 12.128 1.44 ;
      RECT 12.172 0.24 12.562 1.44 ;
      RECT 11.738 -0.12 12.562 0.24 ;
      RECT 10.838 29.52 11.662 29.88 ;
      RECT 10.838 28.32 11.228 29.52 ;
      RECT 11.272 28.32 11.484 29.52 ;
      RECT 11.528 28.32 11.662 29.52 ;
      RECT 10.838 28.08 11.662 28.32 ;
      RECT 11.016 27.36 11.572 28.08 ;
      RECT 10.838 26.88 10.972 28.08 ;
      RECT 11.616 26.88 11.662 28.08 ;
      RECT 11.016 26.88 11.228 27.36 ;
      RECT 11.528 26.88 11.572 27.36 ;
      RECT 11.272 26.16 11.484 27.36 ;
      RECT 10.838 26.16 11.228 26.88 ;
      RECT 11.528 26.16 11.662 26.88 ;
      RECT 10.838 25.92 11.662 26.16 ;
      RECT 11.016 25.2 11.572 25.92 ;
      RECT 10.838 24.72 10.972 25.92 ;
      RECT 11.616 24.72 11.662 25.92 ;
      RECT 11.016 24.72 11.228 25.2 ;
      RECT 11.528 24.72 11.572 25.2 ;
      RECT 11.272 24 11.484 25.2 ;
      RECT 10.838 24 11.228 24.72 ;
      RECT 11.528 24 11.662 24.72 ;
      RECT 10.838 23.76 11.662 24 ;
      RECT 11.016 23.04 11.572 23.76 ;
      RECT 10.838 22.56 10.972 23.76 ;
      RECT 11.616 22.56 11.662 23.76 ;
      RECT 11.016 22.56 11.228 23.04 ;
      RECT 11.528 22.56 11.572 23.04 ;
      RECT 11.272 21.84 11.484 23.04 ;
      RECT 10.838 21.84 11.228 22.56 ;
      RECT 11.528 21.84 11.662 22.56 ;
      RECT 10.838 21.6 11.662 21.84 ;
      RECT 11.016 20.88 11.572 21.6 ;
      RECT 10.838 20.4 10.972 21.6 ;
      RECT 11.616 20.4 11.662 21.6 ;
      RECT 11.016 20.4 11.228 20.88 ;
      RECT 11.528 20.4 11.572 20.88 ;
      RECT 11.528 20.16 11.662 20.4 ;
      RECT 11.272 19.68 11.484 20.88 ;
      RECT 10.838 19.68 11.228 20.4 ;
      RECT 11.528 19.68 11.572 20.16 ;
      RECT 11.616 18.96 11.662 20.16 ;
      RECT 10.838 18.96 11.572 19.68 ;
      RECT 10.838 17.88 11.662 18.96 ;
      RECT 10.838 16.68 10.884 17.88 ;
      RECT 10.928 16.68 10.972 17.88 ;
      RECT 11.016 16.68 11.228 17.88 ;
      RECT 11.272 16.68 11.484 17.88 ;
      RECT 11.528 16.68 11.572 17.88 ;
      RECT 11.616 16.68 11.662 17.88 ;
      RECT 10.838 13.68 11.662 16.68 ;
      RECT 11.016 12.96 11.572 13.68 ;
      RECT 10.838 12.48 10.972 13.68 ;
      RECT 11.616 12.48 11.662 13.68 ;
      RECT 11.016 12.48 11.228 12.96 ;
      RECT 11.528 12.48 11.572 12.96 ;
      RECT 11.272 11.76 11.484 12.96 ;
      RECT 10.838 11.76 11.228 12.48 ;
      RECT 11.528 11.76 11.662 12.48 ;
      RECT 10.838 11.52 11.662 11.76 ;
      RECT 11.016 10.8 11.572 11.52 ;
      RECT 10.838 10.32 10.972 11.52 ;
      RECT 11.616 10.32 11.662 11.52 ;
      RECT 11.016 10.32 11.228 10.8 ;
      RECT 11.528 10.32 11.572 10.8 ;
      RECT 11.272 9.6 11.484 10.8 ;
      RECT 10.838 9.6 11.228 10.32 ;
      RECT 11.528 9.6 11.662 10.32 ;
      RECT 10.838 9.36 11.662 9.6 ;
      RECT 11.016 8.64 11.572 9.36 ;
      RECT 10.838 8.16 10.972 9.36 ;
      RECT 11.616 8.16 11.662 9.36 ;
      RECT 11.016 8.16 11.228 8.64 ;
      RECT 11.528 8.16 11.572 8.64 ;
      RECT 11.272 7.44 11.484 8.64 ;
      RECT 10.838 7.44 11.228 8.16 ;
      RECT 11.528 7.44 11.662 8.16 ;
      RECT 10.838 7.2 11.662 7.44 ;
      RECT 11.016 6.48 11.572 7.2 ;
      RECT 10.838 6 10.972 7.2 ;
      RECT 11.616 6 11.662 7.2 ;
      RECT 11.016 6 11.228 6.48 ;
      RECT 11.528 6 11.572 6.48 ;
      RECT 11.272 5.28 11.484 6.48 ;
      RECT 10.838 5.28 11.228 6 ;
      RECT 11.528 5.28 11.662 6 ;
      RECT 10.838 5.04 11.662 5.28 ;
      RECT 11.016 4.32 11.572 5.04 ;
      RECT 10.838 3.84 10.972 5.04 ;
      RECT 11.616 3.84 11.662 5.04 ;
      RECT 11.016 3.84 11.228 4.32 ;
      RECT 11.528 3.84 11.572 4.32 ;
      RECT 11.272 3.12 11.484 4.32 ;
      RECT 10.838 3.12 11.228 3.84 ;
      RECT 11.528 3.12 11.662 3.84 ;
      RECT 10.838 2.88 11.662 3.12 ;
      RECT 11.016 2.16 11.572 2.88 ;
      RECT 10.838 1.68 10.972 2.88 ;
      RECT 11.616 1.68 11.662 2.88 ;
      RECT 11.016 1.68 11.228 2.16 ;
      RECT 11.528 1.68 11.572 2.16 ;
      RECT 11.272 0.96 11.484 2.16 ;
      RECT 10.838 0.96 11.228 1.68 ;
      RECT 11.528 0.96 11.662 1.68 ;
      RECT 10.838 -0.12 11.662 0.96 ;
      RECT 9.938 28.8 10.762 29.88 ;
      RECT 9.938 28.08 10.072 28.8 ;
      RECT 10.372 28.08 10.762 28.8 ;
      RECT 10.116 27.6 10.328 28.8 ;
      RECT 10.028 27.6 10.072 28.08 ;
      RECT 10.372 27.6 10.584 28.08 ;
      RECT 9.938 26.88 9.984 28.08 ;
      RECT 10.628 26.88 10.762 28.08 ;
      RECT 10.028 26.88 10.584 27.6 ;
      RECT 9.938 26.64 10.762 26.88 ;
      RECT 9.938 25.92 10.072 26.64 ;
      RECT 10.372 25.92 10.762 26.64 ;
      RECT 10.116 25.44 10.328 26.64 ;
      RECT 10.028 25.44 10.072 25.92 ;
      RECT 10.372 25.44 10.584 25.92 ;
      RECT 9.938 24.72 9.984 25.92 ;
      RECT 10.628 24.72 10.762 25.92 ;
      RECT 10.028 24.72 10.584 25.44 ;
      RECT 9.938 24.48 10.762 24.72 ;
      RECT 9.938 23.76 10.072 24.48 ;
      RECT 10.372 23.76 10.762 24.48 ;
      RECT 10.116 23.28 10.328 24.48 ;
      RECT 10.028 23.28 10.072 23.76 ;
      RECT 10.372 23.28 10.584 23.76 ;
      RECT 9.938 22.56 9.984 23.76 ;
      RECT 10.628 22.56 10.762 23.76 ;
      RECT 10.028 22.56 10.584 23.28 ;
      RECT 9.938 22.32 10.762 22.56 ;
      RECT 9.938 21.6 10.072 22.32 ;
      RECT 10.372 21.6 10.762 22.32 ;
      RECT 10.116 21.12 10.328 22.32 ;
      RECT 10.028 21.12 10.072 21.6 ;
      RECT 10.372 21.12 10.584 21.6 ;
      RECT 9.938 20.4 9.984 21.6 ;
      RECT 10.628 20.4 10.762 21.6 ;
      RECT 10.028 20.4 10.584 21.12 ;
      RECT 9.938 20.16 10.762 20.4 ;
      RECT 10.116 19.44 10.762 20.16 ;
      RECT 9.938 18.96 9.984 20.16 ;
      RECT 10.028 18.96 10.072 20.16 ;
      RECT 10.116 18.96 10.328 19.44 ;
      RECT 10.372 18.24 10.584 19.44 ;
      RECT 10.628 18.24 10.762 19.44 ;
      RECT 9.938 18.24 10.328 18.96 ;
      RECT 9.938 15.96 10.762 18.24 ;
      RECT 9.938 14.76 9.984 15.96 ;
      RECT 10.028 14.76 10.584 15.96 ;
      RECT 10.628 14.76 10.672 15.96 ;
      RECT 10.716 14.76 10.762 15.96 ;
      RECT 9.938 14.4 10.762 14.76 ;
      RECT 9.938 13.68 10.072 14.4 ;
      RECT 10.372 13.68 10.762 14.4 ;
      RECT 10.116 13.2 10.328 14.4 ;
      RECT 10.028 13.2 10.072 13.68 ;
      RECT 10.372 13.2 10.584 13.68 ;
      RECT 9.938 12.48 9.984 13.68 ;
      RECT 10.628 12.48 10.762 13.68 ;
      RECT 10.028 12.48 10.584 13.2 ;
      RECT 9.938 12.24 10.762 12.48 ;
      RECT 9.938 11.52 10.072 12.24 ;
      RECT 10.372 11.52 10.762 12.24 ;
      RECT 10.116 11.04 10.328 12.24 ;
      RECT 10.028 11.04 10.072 11.52 ;
      RECT 10.372 11.04 10.584 11.52 ;
      RECT 9.938 10.32 9.984 11.52 ;
      RECT 10.628 10.32 10.762 11.52 ;
      RECT 10.028 10.32 10.584 11.04 ;
      RECT 9.938 10.08 10.762 10.32 ;
      RECT 9.938 9.36 10.072 10.08 ;
      RECT 10.372 9.36 10.762 10.08 ;
      RECT 10.116 8.88 10.328 10.08 ;
      RECT 10.028 8.88 10.072 9.36 ;
      RECT 10.372 8.88 10.584 9.36 ;
      RECT 9.938 8.16 9.984 9.36 ;
      RECT 10.628 8.16 10.762 9.36 ;
      RECT 10.028 8.16 10.584 8.88 ;
      RECT 9.938 7.92 10.762 8.16 ;
      RECT 9.938 7.2 10.072 7.92 ;
      RECT 10.372 7.2 10.762 7.92 ;
      RECT 10.116 6.72 10.328 7.92 ;
      RECT 10.028 6.72 10.072 7.2 ;
      RECT 10.372 6.72 10.584 7.2 ;
      RECT 9.938 6 9.984 7.2 ;
      RECT 10.628 6 10.762 7.2 ;
      RECT 10.028 6 10.584 6.72 ;
      RECT 9.938 5.76 10.762 6 ;
      RECT 9.938 5.04 10.072 5.76 ;
      RECT 10.372 5.04 10.762 5.76 ;
      RECT 10.116 4.56 10.328 5.76 ;
      RECT 10.028 4.56 10.072 5.04 ;
      RECT 10.372 4.56 10.584 5.04 ;
      RECT 9.938 3.84 9.984 5.04 ;
      RECT 10.628 3.84 10.762 5.04 ;
      RECT 10.028 3.84 10.584 4.56 ;
      RECT 9.938 3.6 10.762 3.84 ;
      RECT 9.938 2.88 10.072 3.6 ;
      RECT 10.372 2.88 10.762 3.6 ;
      RECT 10.116 2.4 10.328 3.6 ;
      RECT 10.028 2.4 10.072 2.88 ;
      RECT 10.372 2.4 10.584 2.88 ;
      RECT 9.938 1.68 9.984 2.88 ;
      RECT 10.628 1.68 10.762 2.88 ;
      RECT 10.028 1.68 10.584 2.4 ;
      RECT 9.938 1.44 10.762 1.68 ;
      RECT 9.938 0.24 10.328 1.44 ;
      RECT 10.372 0.24 10.584 1.44 ;
      RECT 10.628 0.24 10.762 1.44 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 29.52 9.862 29.88 ;
      RECT 9.038 28.8 9.172 29.52 ;
      RECT 9.216 28.32 9.428 29.52 ;
      RECT 9.472 28.32 9.684 29.52 ;
      RECT 9.728 28.32 9.772 29.52 ;
      RECT 9.816 28.32 9.862 29.52 ;
      RECT 9.128 28.32 9.172 28.8 ;
      RECT 9.038 27.6 9.084 28.8 ;
      RECT 9.128 27.6 9.862 28.32 ;
      RECT 9.038 27.36 9.862 27.6 ;
      RECT 9.038 26.64 9.172 27.36 ;
      RECT 9.216 26.16 9.428 27.36 ;
      RECT 9.472 26.16 9.684 27.36 ;
      RECT 9.728 26.16 9.772 27.36 ;
      RECT 9.816 26.16 9.862 27.36 ;
      RECT 9.128 26.16 9.172 26.64 ;
      RECT 9.038 25.44 9.084 26.64 ;
      RECT 9.128 25.44 9.862 26.16 ;
      RECT 9.038 25.2 9.862 25.44 ;
      RECT 9.038 24.48 9.172 25.2 ;
      RECT 9.216 24 9.428 25.2 ;
      RECT 9.472 24 9.684 25.2 ;
      RECT 9.728 24 9.772 25.2 ;
      RECT 9.816 24 9.862 25.2 ;
      RECT 9.128 24 9.172 24.48 ;
      RECT 9.038 23.28 9.084 24.48 ;
      RECT 9.128 23.28 9.862 24 ;
      RECT 9.038 23.04 9.862 23.28 ;
      RECT 9.038 22.32 9.172 23.04 ;
      RECT 9.216 21.84 9.428 23.04 ;
      RECT 9.472 21.84 9.684 23.04 ;
      RECT 9.728 21.84 9.772 23.04 ;
      RECT 9.816 21.84 9.862 23.04 ;
      RECT 9.128 21.84 9.172 22.32 ;
      RECT 9.038 21.12 9.084 22.32 ;
      RECT 9.128 21.12 9.862 21.84 ;
      RECT 9.038 20.88 9.862 21.12 ;
      RECT 9.038 19.68 9.172 20.88 ;
      RECT 9.216 19.68 9.428 20.88 ;
      RECT 9.472 19.68 9.684 20.88 ;
      RECT 9.728 19.68 9.772 20.88 ;
      RECT 9.816 19.68 9.862 20.88 ;
      RECT 9.038 19.44 9.862 19.68 ;
      RECT 9.038 18.24 9.084 19.44 ;
      RECT 9.128 18.24 9.862 19.44 ;
      RECT 9.038 15.96 9.862 18.24 ;
      RECT 9.038 14.76 9.172 15.96 ;
      RECT 9.216 14.76 9.428 15.96 ;
      RECT 9.472 14.76 9.684 15.96 ;
      RECT 9.728 14.76 9.772 15.96 ;
      RECT 9.816 14.76 9.862 15.96 ;
      RECT 9.038 14.4 9.862 14.76 ;
      RECT 9.038 13.2 9.084 14.4 ;
      RECT 9.128 13.2 9.862 14.4 ;
      RECT 9.038 12.96 9.862 13.2 ;
      RECT 9.038 12.24 9.172 12.96 ;
      RECT 9.216 11.76 9.428 12.96 ;
      RECT 9.472 11.76 9.684 12.96 ;
      RECT 9.728 11.76 9.772 12.96 ;
      RECT 9.816 11.76 9.862 12.96 ;
      RECT 9.128 11.76 9.172 12.24 ;
      RECT 9.038 11.04 9.084 12.24 ;
      RECT 9.128 11.04 9.862 11.76 ;
      RECT 9.038 10.8 9.862 11.04 ;
      RECT 9.038 10.08 9.172 10.8 ;
      RECT 9.216 9.6 9.428 10.8 ;
      RECT 9.472 9.6 9.684 10.8 ;
      RECT 9.728 9.6 9.772 10.8 ;
      RECT 9.816 9.6 9.862 10.8 ;
      RECT 9.128 9.6 9.172 10.08 ;
      RECT 9.038 8.88 9.084 10.08 ;
      RECT 9.128 8.88 9.862 9.6 ;
      RECT 9.038 8.64 9.862 8.88 ;
      RECT 9.038 7.92 9.172 8.64 ;
      RECT 9.216 7.44 9.428 8.64 ;
      RECT 9.472 7.44 9.684 8.64 ;
      RECT 9.728 7.44 9.772 8.64 ;
      RECT 9.816 7.44 9.862 8.64 ;
      RECT 9.128 7.44 9.172 7.92 ;
      RECT 9.038 6.72 9.084 7.92 ;
      RECT 9.128 6.72 9.862 7.44 ;
      RECT 9.038 6.48 9.862 6.72 ;
      RECT 9.038 5.76 9.172 6.48 ;
      RECT 9.216 5.28 9.428 6.48 ;
      RECT 9.472 5.28 9.684 6.48 ;
      RECT 9.728 5.28 9.772 6.48 ;
      RECT 9.816 5.28 9.862 6.48 ;
      RECT 9.128 5.28 9.172 5.76 ;
      RECT 9.038 4.56 9.084 5.76 ;
      RECT 9.128 4.56 9.862 5.28 ;
      RECT 9.038 4.32 9.862 4.56 ;
      RECT 9.038 3.6 9.172 4.32 ;
      RECT 9.216 3.12 9.428 4.32 ;
      RECT 9.472 3.12 9.684 4.32 ;
      RECT 9.728 3.12 9.772 4.32 ;
      RECT 9.816 3.12 9.862 4.32 ;
      RECT 9.128 3.12 9.172 3.6 ;
      RECT 9.038 2.4 9.084 3.6 ;
      RECT 9.128 2.4 9.862 3.12 ;
      RECT 9.038 2.16 9.862 2.4 ;
      RECT 9.038 1.44 9.172 2.16 ;
      RECT 9.216 0.96 9.428 2.16 ;
      RECT 9.472 0.96 9.684 2.16 ;
      RECT 9.728 0.96 9.772 2.16 ;
      RECT 9.816 0.96 9.862 2.16 ;
      RECT 9.128 0.96 9.172 1.44 ;
      RECT 9.038 0.24 9.084 1.44 ;
      RECT 9.128 0.24 9.862 0.96 ;
      RECT 9.038 -0.12 9.862 0.24 ;
      RECT 8.138 28.8 8.962 29.88 ;
      RECT 8.572 28.08 8.962 28.8 ;
      RECT 8.138 27.6 8.528 28.8 ;
      RECT 8.572 27.6 8.784 28.08 ;
      RECT 8.828 26.88 8.872 28.08 ;
      RECT 8.916 26.88 8.962 28.08 ;
      RECT 8.138 26.88 8.784 27.6 ;
      RECT 8.138 26.64 8.962 26.88 ;
      RECT 8.572 25.92 8.962 26.64 ;
      RECT 8.138 25.44 8.528 26.64 ;
      RECT 8.572 25.44 8.784 25.92 ;
      RECT 8.828 24.72 8.872 25.92 ;
      RECT 8.916 24.72 8.962 25.92 ;
      RECT 8.138 24.72 8.784 25.44 ;
      RECT 8.138 24.48 8.962 24.72 ;
      RECT 8.572 23.76 8.962 24.48 ;
      RECT 8.138 23.28 8.528 24.48 ;
      RECT 8.572 23.28 8.784 23.76 ;
      RECT 8.828 22.56 8.872 23.76 ;
      RECT 8.916 22.56 8.962 23.76 ;
      RECT 8.138 22.56 8.784 23.28 ;
      RECT 8.138 22.32 8.962 22.56 ;
      RECT 8.572 21.6 8.962 22.32 ;
      RECT 8.138 21.12 8.528 22.32 ;
      RECT 8.572 21.12 8.784 21.6 ;
      RECT 8.828 20.4 8.872 21.6 ;
      RECT 8.916 20.4 8.962 21.6 ;
      RECT 8.138 20.4 8.784 21.12 ;
      RECT 8.138 20.16 8.962 20.4 ;
      RECT 8.828 19.44 8.962 20.16 ;
      RECT 8.138 18.96 8.528 20.16 ;
      RECT 8.572 18.96 8.784 20.16 ;
      RECT 8.828 18.96 8.872 19.44 ;
      RECT 8.916 18.24 8.962 19.44 ;
      RECT 8.138 18.24 8.872 18.96 ;
      RECT 8.138 15.96 8.962 18.24 ;
      RECT 8.138 14.76 8.184 15.96 ;
      RECT 8.228 14.76 8.272 15.96 ;
      RECT 8.316 14.76 8.784 15.96 ;
      RECT 8.828 14.76 8.872 15.96 ;
      RECT 8.916 14.76 8.962 15.96 ;
      RECT 8.138 14.4 8.962 14.76 ;
      RECT 8.572 13.68 8.962 14.4 ;
      RECT 8.138 13.2 8.528 14.4 ;
      RECT 8.572 13.2 8.784 13.68 ;
      RECT 8.828 12.48 8.872 13.68 ;
      RECT 8.916 12.48 8.962 13.68 ;
      RECT 8.138 12.48 8.784 13.2 ;
      RECT 8.138 12.24 8.962 12.48 ;
      RECT 8.572 11.52 8.962 12.24 ;
      RECT 8.138 11.04 8.528 12.24 ;
      RECT 8.572 11.04 8.784 11.52 ;
      RECT 8.828 10.32 8.872 11.52 ;
      RECT 8.916 10.32 8.962 11.52 ;
      RECT 8.138 10.32 8.784 11.04 ;
      RECT 8.138 10.08 8.962 10.32 ;
      RECT 8.572 9.36 8.962 10.08 ;
      RECT 8.138 8.88 8.528 10.08 ;
      RECT 8.572 8.88 8.784 9.36 ;
      RECT 8.828 8.16 8.872 9.36 ;
      RECT 8.916 8.16 8.962 9.36 ;
      RECT 8.138 8.16 8.784 8.88 ;
      RECT 8.138 7.92 8.962 8.16 ;
      RECT 8.572 7.2 8.962 7.92 ;
      RECT 8.138 6.72 8.528 7.92 ;
      RECT 8.572 6.72 8.784 7.2 ;
      RECT 8.828 6 8.872 7.2 ;
      RECT 8.916 6 8.962 7.2 ;
      RECT 8.138 6 8.784 6.72 ;
      RECT 8.138 5.76 8.962 6 ;
      RECT 8.572 5.04 8.962 5.76 ;
      RECT 8.138 4.56 8.528 5.76 ;
      RECT 8.572 4.56 8.784 5.04 ;
      RECT 8.828 3.84 8.872 5.04 ;
      RECT 8.916 3.84 8.962 5.04 ;
      RECT 8.138 3.84 8.784 4.56 ;
      RECT 8.138 3.6 8.962 3.84 ;
      RECT 8.572 2.88 8.962 3.6 ;
      RECT 8.138 2.4 8.528 3.6 ;
      RECT 8.572 2.4 8.784 2.88 ;
      RECT 8.828 1.68 8.872 2.88 ;
      RECT 8.916 1.68 8.962 2.88 ;
      RECT 8.138 1.68 8.784 2.4 ;
      RECT 8.138 1.44 8.962 1.68 ;
      RECT 8.138 0.24 8.872 1.44 ;
      RECT 8.916 0.24 8.962 1.44 ;
      RECT 8.138 -0.12 8.962 0.24 ;
      RECT 7.238 28.8 8.062 29.88 ;
      RECT 7.672 28.08 8.062 28.8 ;
      RECT 7.238 27.6 7.372 28.8 ;
      RECT 7.416 27.6 7.628 28.8 ;
      RECT 7.672 27.6 7.884 28.08 ;
      RECT 7.928 26.88 8.062 28.08 ;
      RECT 7.238 26.88 7.884 27.6 ;
      RECT 7.238 26.64 8.062 26.88 ;
      RECT 7.672 25.92 8.062 26.64 ;
      RECT 7.238 25.44 7.372 26.64 ;
      RECT 7.416 25.44 7.628 26.64 ;
      RECT 7.672 25.44 7.884 25.92 ;
      RECT 7.928 24.72 8.062 25.92 ;
      RECT 7.238 24.72 7.884 25.44 ;
      RECT 7.238 24.48 8.062 24.72 ;
      RECT 7.672 23.76 8.062 24.48 ;
      RECT 7.238 23.28 7.372 24.48 ;
      RECT 7.416 23.28 7.628 24.48 ;
      RECT 7.672 23.28 7.884 23.76 ;
      RECT 7.928 22.56 8.062 23.76 ;
      RECT 7.238 22.56 7.884 23.28 ;
      RECT 7.238 22.32 8.062 22.56 ;
      RECT 7.672 21.6 8.062 22.32 ;
      RECT 7.238 21.12 7.372 22.32 ;
      RECT 7.416 21.12 7.628 22.32 ;
      RECT 7.672 21.12 7.884 21.6 ;
      RECT 7.928 20.4 8.062 21.6 ;
      RECT 7.238 20.4 7.884 21.12 ;
      RECT 7.238 20.16 8.062 20.4 ;
      RECT 7.328 19.44 8.062 20.16 ;
      RECT 7.238 18.96 7.284 20.16 ;
      RECT 7.328 18.96 7.372 19.44 ;
      RECT 7.416 18.24 7.628 19.44 ;
      RECT 7.672 18.24 8.062 19.44 ;
      RECT 7.238 18.24 7.372 18.96 ;
      RECT 7.238 17.88 8.062 18.24 ;
      RECT 7.238 16.68 7.284 17.88 ;
      RECT 7.328 16.68 8.062 17.88 ;
      RECT 7.238 14.4 8.062 16.68 ;
      RECT 7.672 13.68 8.062 14.4 ;
      RECT 7.238 13.2 7.372 14.4 ;
      RECT 7.416 13.2 7.628 14.4 ;
      RECT 7.672 13.2 7.884 13.68 ;
      RECT 7.928 12.48 8.062 13.68 ;
      RECT 7.238 12.48 7.884 13.2 ;
      RECT 7.238 12.24 8.062 12.48 ;
      RECT 7.672 11.52 8.062 12.24 ;
      RECT 7.238 11.04 7.372 12.24 ;
      RECT 7.416 11.04 7.628 12.24 ;
      RECT 7.672 11.04 7.884 11.52 ;
      RECT 7.928 10.32 8.062 11.52 ;
      RECT 7.238 10.32 7.884 11.04 ;
      RECT 7.238 10.08 8.062 10.32 ;
      RECT 7.672 9.36 8.062 10.08 ;
      RECT 7.238 8.88 7.372 10.08 ;
      RECT 7.416 8.88 7.628 10.08 ;
      RECT 7.672 8.88 7.884 9.36 ;
      RECT 7.928 8.16 8.062 9.36 ;
      RECT 7.238 8.16 7.884 8.88 ;
      RECT 7.238 7.92 8.062 8.16 ;
      RECT 7.672 7.2 8.062 7.92 ;
      RECT 7.238 6.72 7.372 7.92 ;
      RECT 7.416 6.72 7.628 7.92 ;
      RECT 7.672 6.72 7.884 7.2 ;
      RECT 7.928 6 8.062 7.2 ;
      RECT 7.238 6 7.884 6.72 ;
      RECT 7.238 5.76 8.062 6 ;
      RECT 7.672 5.04 8.062 5.76 ;
      RECT 7.238 4.56 7.372 5.76 ;
      RECT 7.416 4.56 7.628 5.76 ;
      RECT 7.672 4.56 7.884 5.04 ;
      RECT 7.928 3.84 8.062 5.04 ;
      RECT 7.238 3.84 7.884 4.56 ;
      RECT 7.238 3.6 8.062 3.84 ;
      RECT 7.672 2.88 8.062 3.6 ;
      RECT 7.238 2.4 7.372 3.6 ;
      RECT 7.416 2.4 7.628 3.6 ;
      RECT 7.672 2.4 7.884 2.88 ;
      RECT 7.238 2.16 7.884 2.4 ;
      RECT 7.928 1.68 8.062 2.88 ;
      RECT 7.328 1.68 7.884 2.16 ;
      RECT 7.238 0.96 7.284 2.16 ;
      RECT 7.328 0.96 8.062 1.68 ;
      RECT 7.238 -0.12 8.062 0.96 ;
      RECT 6.338 29.52 7.162 29.88 ;
      RECT 6.338 28.32 6.728 29.52 ;
      RECT 6.772 28.32 6.984 29.52 ;
      RECT 7.028 28.32 7.162 29.52 ;
      RECT 6.338 28.08 7.162 28.32 ;
      RECT 6.338 27.36 7.072 28.08 ;
      RECT 7.116 26.88 7.162 28.08 ;
      RECT 7.028 26.88 7.072 27.36 ;
      RECT 6.338 26.16 6.728 27.36 ;
      RECT 6.772 26.16 6.984 27.36 ;
      RECT 7.028 26.16 7.162 26.88 ;
      RECT 6.338 25.92 7.162 26.16 ;
      RECT 6.338 25.2 7.072 25.92 ;
      RECT 7.116 24.72 7.162 25.92 ;
      RECT 7.028 24.72 7.072 25.2 ;
      RECT 6.338 24 6.728 25.2 ;
      RECT 6.772 24 6.984 25.2 ;
      RECT 7.028 24 7.162 24.72 ;
      RECT 6.338 23.76 7.162 24 ;
      RECT 6.338 23.04 7.072 23.76 ;
      RECT 7.116 22.56 7.162 23.76 ;
      RECT 7.028 22.56 7.072 23.04 ;
      RECT 6.338 21.84 6.728 23.04 ;
      RECT 6.772 21.84 6.984 23.04 ;
      RECT 7.028 21.84 7.162 22.56 ;
      RECT 6.338 21.6 7.162 21.84 ;
      RECT 6.338 20.88 7.072 21.6 ;
      RECT 7.116 20.4 7.162 21.6 ;
      RECT 7.028 20.4 7.072 20.88 ;
      RECT 7.028 20.16 7.162 20.4 ;
      RECT 6.338 19.68 6.728 20.88 ;
      RECT 6.772 19.68 6.984 20.88 ;
      RECT 7.028 19.68 7.072 20.16 ;
      RECT 7.116 18.96 7.162 20.16 ;
      RECT 6.338 18.96 7.072 19.68 ;
      RECT 6.338 17.88 7.162 18.96 ;
      RECT 6.338 16.68 6.728 17.88 ;
      RECT 6.772 16.68 6.984 17.88 ;
      RECT 7.028 16.68 7.072 17.88 ;
      RECT 7.116 16.68 7.162 17.88 ;
      RECT 6.338 13.68 7.162 16.68 ;
      RECT 6.338 12.96 7.072 13.68 ;
      RECT 7.116 12.48 7.162 13.68 ;
      RECT 7.028 12.48 7.072 12.96 ;
      RECT 6.338 11.76 6.728 12.96 ;
      RECT 6.772 11.76 6.984 12.96 ;
      RECT 7.028 11.76 7.162 12.48 ;
      RECT 6.338 11.52 7.162 11.76 ;
      RECT 6.338 10.8 7.072 11.52 ;
      RECT 7.116 10.32 7.162 11.52 ;
      RECT 7.028 10.32 7.072 10.8 ;
      RECT 6.338 9.6 6.728 10.8 ;
      RECT 6.772 9.6 6.984 10.8 ;
      RECT 7.028 9.6 7.162 10.32 ;
      RECT 6.338 9.36 7.162 9.6 ;
      RECT 6.338 8.64 7.072 9.36 ;
      RECT 7.116 8.16 7.162 9.36 ;
      RECT 7.028 8.16 7.072 8.64 ;
      RECT 6.338 7.44 6.728 8.64 ;
      RECT 6.772 7.44 6.984 8.64 ;
      RECT 7.028 7.44 7.162 8.16 ;
      RECT 6.338 7.2 7.162 7.44 ;
      RECT 6.338 6.48 7.072 7.2 ;
      RECT 7.116 6 7.162 7.2 ;
      RECT 7.028 6 7.072 6.48 ;
      RECT 6.338 5.28 6.728 6.48 ;
      RECT 6.772 5.28 6.984 6.48 ;
      RECT 7.028 5.28 7.162 6 ;
      RECT 6.338 5.04 7.162 5.28 ;
      RECT 6.338 4.32 7.072 5.04 ;
      RECT 7.116 3.84 7.162 5.04 ;
      RECT 7.028 3.84 7.072 4.32 ;
      RECT 6.338 3.12 6.728 4.32 ;
      RECT 6.772 3.12 6.984 4.32 ;
      RECT 7.028 3.12 7.162 3.84 ;
      RECT 6.338 2.88 7.162 3.12 ;
      RECT 6.772 2.16 7.162 2.88 ;
      RECT 6.338 1.68 6.728 2.88 ;
      RECT 6.772 1.68 7.072 2.16 ;
      RECT 6.338 1.44 7.072 1.68 ;
      RECT 7.116 0.96 7.162 2.16 ;
      RECT 7.028 0.96 7.072 1.44 ;
      RECT 6.338 0.24 6.728 1.44 ;
      RECT 6.772 0.24 6.984 1.44 ;
      RECT 7.028 0.24 7.162 0.96 ;
      RECT 6.338 -0.12 7.162 0.24 ;
      RECT 5.438 -0.12 6.262 29.88 ;
      RECT 4.538 -0.12 5.362 29.88 ;
      RECT 3.638 -0.12 4.462 29.88 ;
      RECT 2.738 -0.12 3.562 29.88 ;
      RECT 1.838 -0.12 2.662 29.88 ;
      RECT 0.938 -0.12 1.762 29.88 ;
      RECT -0.04 29.82 0.862 29.88 ;
      RECT -0.092 -0.06 0.862 29.82 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 19.058 0 19.72 29.76 ;
      RECT 18.158 0 18.742 29.76 ;
      RECT 17.258 0 17.842 29.76 ;
      RECT 16.358 0 16.942 29.76 ;
      RECT 15.458 0 16.042 29.76 ;
      RECT 14.558 0 15.142 29.76 ;
      RECT 13.658 0 14.242 29.76 ;
      RECT 12.758 0 13.342 29.76 ;
      RECT 11.858 28.92 12.442 29.76 ;
      RECT 12.292 27.48 12.442 28.92 ;
      RECT 11.858 26.76 12.442 27.48 ;
      RECT 12.292 25.32 12.442 26.76 ;
      RECT 11.858 24.6 12.442 25.32 ;
      RECT 12.292 23.16 12.442 24.6 ;
      RECT 11.858 22.44 12.442 23.16 ;
      RECT 12.292 21 12.442 22.44 ;
      RECT 11.858 20.28 12.442 21 ;
      RECT 11.948 19.56 12.442 20.28 ;
      RECT 12.292 18.12 12.442 19.56 ;
      RECT 11.858 18 12.442 18.12 ;
      RECT 11.948 16.56 12.442 18 ;
      RECT 11.858 14.52 12.442 16.56 ;
      RECT 12.292 13.08 12.442 14.52 ;
      RECT 11.858 12.36 12.442 13.08 ;
      RECT 12.292 10.92 12.442 12.36 ;
      RECT 11.858 10.2 12.442 10.92 ;
      RECT 12.292 8.76 12.442 10.2 ;
      RECT 11.858 8.04 12.442 8.76 ;
      RECT 12.292 6.6 12.442 8.04 ;
      RECT 11.858 5.88 12.442 6.6 ;
      RECT 12.292 4.44 12.442 5.88 ;
      RECT 11.858 3.72 12.442 4.44 ;
      RECT 12.292 2.28 12.442 3.72 ;
      RECT 11.858 1.56 12.442 2.28 ;
      RECT 12.292 0.12 12.442 1.56 ;
      RECT 11.858 0 12.442 0.12 ;
      RECT 10.958 29.64 11.542 29.76 ;
      RECT 10.958 28.2 11.108 29.64 ;
      RECT 10.058 28.92 10.642 29.76 ;
      RECT 10.492 28.2 10.642 28.92 ;
      RECT 9.158 29.64 9.742 29.76 ;
      RECT 8.258 28.92 8.842 29.76 ;
      RECT 8.692 28.2 8.842 28.92 ;
      RECT 8.258 27.48 8.408 28.92 ;
      RECT 8.258 26.76 8.664 27.48 ;
      RECT 8.258 25.32 8.408 26.76 ;
      RECT 8.258 24.6 8.664 25.32 ;
      RECT 8.258 23.16 8.408 24.6 ;
      RECT 8.258 22.44 8.664 23.16 ;
      RECT 8.258 21 8.408 22.44 ;
      RECT 8.258 20.28 8.664 21 ;
      RECT 8.258 18.84 8.408 20.28 ;
      RECT 8.258 18.12 8.752 18.84 ;
      RECT 8.258 16.08 8.842 18.12 ;
      RECT 8.436 14.64 8.664 16.08 ;
      RECT 8.258 14.52 8.842 14.64 ;
      RECT 8.692 13.8 8.842 14.52 ;
      RECT 8.258 13.08 8.408 14.52 ;
      RECT 8.258 12.36 8.664 13.08 ;
      RECT 8.258 10.92 8.408 12.36 ;
      RECT 8.258 10.2 8.664 10.92 ;
      RECT 8.258 8.76 8.408 10.2 ;
      RECT 8.258 8.04 8.664 8.76 ;
      RECT 8.258 6.6 8.408 8.04 ;
      RECT 8.258 5.88 8.664 6.6 ;
      RECT 8.258 4.44 8.408 5.88 ;
      RECT 8.258 3.72 8.664 4.44 ;
      RECT 8.258 2.28 8.408 3.72 ;
      RECT 8.258 1.56 8.664 2.28 ;
      RECT 8.258 0.12 8.752 1.56 ;
      RECT 8.258 0 8.842 0.12 ;
      RECT 7.358 28.92 7.942 29.76 ;
      RECT 7.792 28.2 7.942 28.92 ;
      RECT 6.458 29.64 7.042 29.76 ;
      RECT 6.458 28.2 6.608 29.64 ;
      RECT 6.458 27.48 6.952 28.2 ;
      RECT 6.458 26.04 6.608 27.48 ;
      RECT 6.458 25.32 6.952 26.04 ;
      RECT 6.458 23.88 6.608 25.32 ;
      RECT 6.458 23.16 6.952 23.88 ;
      RECT 6.458 21.72 6.608 23.16 ;
      RECT 6.458 21 6.952 21.72 ;
      RECT 6.458 19.56 6.608 21 ;
      RECT 6.458 18.84 6.952 19.56 ;
      RECT 6.458 18 7.042 18.84 ;
      RECT 6.458 16.56 6.608 18 ;
      RECT 6.458 13.8 7.042 16.56 ;
      RECT 6.458 13.08 6.952 13.8 ;
      RECT 6.458 11.64 6.608 13.08 ;
      RECT 6.458 10.92 6.952 11.64 ;
      RECT 6.458 9.48 6.608 10.92 ;
      RECT 6.458 8.76 6.952 9.48 ;
      RECT 6.458 7.32 6.608 8.76 ;
      RECT 6.458 6.6 6.952 7.32 ;
      RECT 6.458 5.16 6.608 6.6 ;
      RECT 6.458 4.44 6.952 5.16 ;
      RECT 6.458 0.12 6.608 4.44 ;
      RECT 6.458 0 7.042 0.12 ;
      RECT 5.558 0 6.142 29.76 ;
      RECT 4.658 0 5.242 29.76 ;
      RECT 3.758 0 4.342 29.76 ;
      RECT 2.858 0 3.442 29.76 ;
      RECT 1.958 0 2.542 29.76 ;
      RECT 1.058 0 1.642 29.76 ;
      RECT 0.08 0 0.742 29.76 ;
      RECT 11.136 27.48 11.452 28.2 ;
      RECT 9.248 27.48 9.742 28.2 ;
      RECT 10.148 26.76 10.464 27.48 ;
      RECT 7.358 26.76 7.764 27.48 ;
      RECT 10.958 26.04 11.108 26.76 ;
      RECT 10.492 26.04 10.642 26.76 ;
      RECT 8.692 26.04 8.842 26.76 ;
      RECT 7.792 26.04 7.942 26.76 ;
      RECT 11.136 25.32 11.452 26.04 ;
      RECT 9.248 25.32 9.742 26.04 ;
      RECT 10.148 24.6 10.464 25.32 ;
      RECT 7.358 24.6 7.764 25.32 ;
      RECT 10.958 23.88 11.108 24.6 ;
      RECT 10.492 23.88 10.642 24.6 ;
      RECT 8.692 23.88 8.842 24.6 ;
      RECT 7.792 23.88 7.942 24.6 ;
      RECT 11.136 23.16 11.452 23.88 ;
      RECT 9.248 23.16 9.742 23.88 ;
      RECT 10.148 22.44 10.464 23.16 ;
      RECT 7.358 22.44 7.764 23.16 ;
      RECT 10.958 21.72 11.108 22.44 ;
      RECT 10.492 21.72 10.642 22.44 ;
      RECT 8.692 21.72 8.842 22.44 ;
      RECT 7.792 21.72 7.942 22.44 ;
      RECT 11.136 21 11.452 21.72 ;
      RECT 9.248 21 9.742 21.72 ;
      RECT 10.148 20.28 10.464 21 ;
      RECT 10.236 19.56 10.642 20.28 ;
      RECT 7.358 20.28 7.764 21 ;
      RECT 7.448 19.56 7.942 20.28 ;
      RECT 7.792 18.12 7.942 19.56 ;
      RECT 7.358 18 7.942 18.12 ;
      RECT 7.448 16.56 7.942 18 ;
      RECT 7.358 14.52 7.942 16.56 ;
      RECT 7.792 13.8 7.942 14.52 ;
      RECT 10.958 19.56 11.108 20.28 ;
      RECT 10.958 18.84 11.452 19.56 ;
      RECT 10.958 18 11.542 18.84 ;
      RECT 9.248 18.12 9.742 19.56 ;
      RECT 9.158 16.08 9.742 18.12 ;
      RECT 10.058 18.12 10.208 18.84 ;
      RECT 10.058 16.08 10.642 18.12 ;
      RECT 10.148 14.64 10.464 16.08 ;
      RECT 10.058 14.52 10.642 14.64 ;
      RECT 10.492 13.8 10.642 14.52 ;
      RECT 10.958 13.8 11.542 16.56 ;
      RECT 11.136 13.08 11.452 13.8 ;
      RECT 9.158 14.52 9.742 14.64 ;
      RECT 9.248 13.08 9.742 14.52 ;
      RECT 10.148 12.36 10.464 13.08 ;
      RECT 7.358 12.36 7.764 13.08 ;
      RECT 10.958 11.64 11.108 12.36 ;
      RECT 10.492 11.64 10.642 12.36 ;
      RECT 8.692 11.64 8.842 12.36 ;
      RECT 7.792 11.64 7.942 12.36 ;
      RECT 11.136 10.92 11.452 11.64 ;
      RECT 9.248 10.92 9.742 11.64 ;
      RECT 10.148 10.2 10.464 10.92 ;
      RECT 7.358 10.2 7.764 10.92 ;
      RECT 10.958 9.48 11.108 10.2 ;
      RECT 10.492 9.48 10.642 10.2 ;
      RECT 8.692 9.48 8.842 10.2 ;
      RECT 7.792 9.48 7.942 10.2 ;
      RECT 11.136 8.76 11.452 9.48 ;
      RECT 9.248 8.76 9.742 9.48 ;
      RECT 10.148 8.04 10.464 8.76 ;
      RECT 7.358 8.04 7.764 8.76 ;
      RECT 10.958 7.32 11.108 8.04 ;
      RECT 10.492 7.32 10.642 8.04 ;
      RECT 8.692 7.32 8.842 8.04 ;
      RECT 7.792 7.32 7.942 8.04 ;
      RECT 11.136 6.6 11.452 7.32 ;
      RECT 9.248 6.6 9.742 7.32 ;
      RECT 10.148 5.88 10.464 6.6 ;
      RECT 7.358 5.88 7.764 6.6 ;
      RECT 10.958 5.16 11.108 5.88 ;
      RECT 10.492 5.16 10.642 5.88 ;
      RECT 8.692 5.16 8.842 5.88 ;
      RECT 7.792 5.16 7.942 5.88 ;
      RECT 11.136 4.44 11.452 5.16 ;
      RECT 9.248 4.44 9.742 5.16 ;
      RECT 10.148 3.72 10.464 4.44 ;
      RECT 7.358 3.72 7.764 4.44 ;
      RECT 10.958 3 11.108 3.72 ;
      RECT 10.492 3 10.642 3.72 ;
      RECT 8.692 3 8.842 3.72 ;
      RECT 7.792 3 7.942 3.72 ;
      RECT 11.136 2.28 11.452 3 ;
      RECT 9.248 2.28 9.742 3 ;
      RECT 6.892 2.28 7.042 3 ;
      RECT 6.892 1.56 6.952 2.28 ;
      RECT 10.148 1.56 10.464 2.28 ;
      RECT 10.058 0.12 10.208 1.56 ;
      RECT 10.058 0 10.642 0.12 ;
      RECT 7.448 1.56 7.764 2.28 ;
      RECT 7.448 0.84 7.942 1.56 ;
      RECT 7.358 0 7.942 0.84 ;
      RECT 10.958 0.84 11.108 1.56 ;
      RECT 10.958 0 11.542 0.84 ;
      RECT 9.248 0.12 9.742 0.84 ;
      RECT 9.158 0 9.742 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 19.8 29.758 ;
    LAYER m1 ;
      RECT 0 0 19.8 29.76 ;
    LAYER m2 ;
      RECT 0 0.015 19.8 29.745 ;
    LAYER m3 ;
      RECT 0.015 0 19.785 29.76 ;
    LAYER m4 ;
      RECT 0 0.02 19.8 29.74 ;
    LAYER m5 ;
      RECT 0.012 0 19.788 29.76 ;
    LAYER m6 ;
      RECT 0 0.012 19.8 29.748 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf132b032e1r1w0cbbehbaa4acw

END LIBRARY
