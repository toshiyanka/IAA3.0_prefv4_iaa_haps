VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf192b080e1r1w0cbbehbaa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf192b080e1r1w0cbbehbaa4acw 0 0 ;
  SIZE 34.2 BY 41.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 21.48 18.128 22.68 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 19.56 15.128 20.76 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 21.48 13.628 22.68 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 21.48 13.716 22.68 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 21.48 13.972 22.68 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 21.48 14.228 22.68 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 21.48 14.316 22.68 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 21.48 14.528 22.68 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.084 21.48 15.128 22.68 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 21.48 18.216 22.68 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.428 21.48 18.472 22.68 ;
    END
  END rdaddrp0_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 0.24 13.628 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 23.28 14.616 24.48 ;
    END
  END rddatap0[100]
  PIN rddatap0[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 23.28 14.872 24.48 ;
    END
  END rddatap0[101]
  PIN rddatap0[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.784 23.28 17.828 24.48 ;
    END
  END rddatap0[102]
  PIN rddatap0[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 23.28 17.916 24.48 ;
    END
  END rddatap0[103]
  PIN rddatap0[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 24 13.972 25.2 ;
    END
  END rddatap0[104]
  PIN rddatap0[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 24 14.228 25.2 ;
    END
  END rddatap0[105]
  PIN rddatap0[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 24 18.728 25.2 ;
    END
  END rddatap0[106]
  PIN rddatap0[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 24 18.816 25.2 ;
    END
  END rddatap0[107]
  PIN rddatap0[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 24.72 14.872 25.92 ;
    END
  END rddatap0[108]
  PIN rddatap0[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 24.72 13.628 25.92 ;
    END
  END rddatap0[109]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 1.68 18.816 2.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 24.72 17.916 25.92 ;
    END
  END rddatap0[110]
  PIN rddatap0[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 24.72 18.128 25.92 ;
    END
  END rddatap0[111]
  PIN rddatap0[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 25.44 14.316 26.64 ;
    END
  END rddatap0[112]
  PIN rddatap0[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 25.44 14.528 26.64 ;
    END
  END rddatap0[113]
  PIN rddatap0[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 25.44 18.816 26.64 ;
    END
  END rddatap0[114]
  PIN rddatap0[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 25.44 19.028 26.64 ;
    END
  END rddatap0[115]
  PIN rddatap0[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 26.16 13.628 27.36 ;
    END
  END rddatap0[116]
  PIN rddatap0[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 26.16 13.716 27.36 ;
    END
  END rddatap0[117]
  PIN rddatap0[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 26.16 18.128 27.36 ;
    END
  END rddatap0[118]
  PIN rddatap0[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 26.16 18.216 27.36 ;
    END
  END rddatap0[119]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 1.68 19.028 2.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 26.88 14.616 28.08 ;
    END
  END rddatap0[120]
  PIN rddatap0[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 26.88 14.872 28.08 ;
    END
  END rddatap0[121]
  PIN rddatap0[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 26.88 18.816 28.08 ;
    END
  END rddatap0[122]
  PIN rddatap0[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 26.88 19.028 28.08 ;
    END
  END rddatap0[123]
  PIN rddatap0[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 27.6 13.628 28.8 ;
    END
  END rddatap0[124]
  PIN rddatap0[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 27.6 13.716 28.8 ;
    END
  END rddatap0[125]
  PIN rddatap0[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 27.6 18.128 28.8 ;
    END
  END rddatap0[126]
  PIN rddatap0[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 27.6 18.216 28.8 ;
    END
  END rddatap0[127]
  PIN rddatap0[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 28.32 14.616 29.52 ;
    END
  END rddatap0[128]
  PIN rddatap0[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 28.32 14.872 29.52 ;
    END
  END rddatap0[129]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 2.4 13.628 3.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 28.32 18.816 29.52 ;
    END
  END rddatap0[130]
  PIN rddatap0[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 28.32 19.028 29.52 ;
    END
  END rddatap0[131]
  PIN rddatap0[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 29.04 13.628 30.24 ;
    END
  END rddatap0[132]
  PIN rddatap0[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 29.04 13.716 30.24 ;
    END
  END rddatap0[133]
  PIN rddatap0[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 29.04 18.128 30.24 ;
    END
  END rddatap0[134]
  PIN rddatap0[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 29.04 18.216 30.24 ;
    END
  END rddatap0[135]
  PIN rddatap0[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 29.76 14.616 30.96 ;
    END
  END rddatap0[136]
  PIN rddatap0[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 29.76 14.872 30.96 ;
    END
  END rddatap0[137]
  PIN rddatap0[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 29.76 18.816 30.96 ;
    END
  END rddatap0[138]
  PIN rddatap0[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 29.76 19.028 30.96 ;
    END
  END rddatap0[139]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 2.4 13.716 3.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 30.48 13.628 31.68 ;
    END
  END rddatap0[140]
  PIN rddatap0[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 30.48 13.716 31.68 ;
    END
  END rddatap0[141]
  PIN rddatap0[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 30.48 18.128 31.68 ;
    END
  END rddatap0[142]
  PIN rddatap0[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 30.48 18.216 31.68 ;
    END
  END rddatap0[143]
  PIN rddatap0[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 31.2 14.616 32.4 ;
    END
  END rddatap0[144]
  PIN rddatap0[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 31.2 14.872 32.4 ;
    END
  END rddatap0[145]
  PIN rddatap0[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 31.2 18.816 32.4 ;
    END
  END rddatap0[146]
  PIN rddatap0[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 31.2 19.028 32.4 ;
    END
  END rddatap0[147]
  PIN rddatap0[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 31.92 13.628 33.12 ;
    END
  END rddatap0[148]
  PIN rddatap0[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 31.92 13.716 33.12 ;
    END
  END rddatap0[149]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 2.4 18.128 3.6 ;
    END
  END rddatap0[14]
  PIN rddatap0[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 31.92 18.128 33.12 ;
    END
  END rddatap0[150]
  PIN rddatap0[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 31.92 18.216 33.12 ;
    END
  END rddatap0[151]
  PIN rddatap0[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 32.64 14.616 33.84 ;
    END
  END rddatap0[152]
  PIN rddatap0[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 32.64 14.872 33.84 ;
    END
  END rddatap0[153]
  PIN rddatap0[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 32.64 18.816 33.84 ;
    END
  END rddatap0[154]
  PIN rddatap0[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 32.64 19.028 33.84 ;
    END
  END rddatap0[155]
  PIN rddatap0[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 33.36 13.628 34.56 ;
    END
  END rddatap0[156]
  PIN rddatap0[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 33.36 13.716 34.56 ;
    END
  END rddatap0[157]
  PIN rddatap0[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 33.36 18.128 34.56 ;
    END
  END rddatap0[158]
  PIN rddatap0[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 33.36 18.216 34.56 ;
    END
  END rddatap0[159]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 2.4 18.216 3.6 ;
    END
  END rddatap0[15]
  PIN rddatap0[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 34.08 14.616 35.28 ;
    END
  END rddatap0[160]
  PIN rddatap0[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 34.08 14.872 35.28 ;
    END
  END rddatap0[161]
  PIN rddatap0[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 34.08 18.816 35.28 ;
    END
  END rddatap0[162]
  PIN rddatap0[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 34.08 19.028 35.28 ;
    END
  END rddatap0[163]
  PIN rddatap0[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 34.8 13.628 36 ;
    END
  END rddatap0[164]
  PIN rddatap0[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 34.8 13.716 36 ;
    END
  END rddatap0[165]
  PIN rddatap0[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 34.8 18.128 36 ;
    END
  END rddatap0[166]
  PIN rddatap0[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 34.8 18.216 36 ;
    END
  END rddatap0[167]
  PIN rddatap0[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 35.52 14.616 36.72 ;
    END
  END rddatap0[168]
  PIN rddatap0[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 35.52 14.872 36.72 ;
    END
  END rddatap0[169]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 3.12 14.616 4.32 ;
    END
  END rddatap0[16]
  PIN rddatap0[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 35.52 18.816 36.72 ;
    END
  END rddatap0[170]
  PIN rddatap0[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 35.52 19.028 36.72 ;
    END
  END rddatap0[171]
  PIN rddatap0[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 36.24 13.628 37.44 ;
    END
  END rddatap0[172]
  PIN rddatap0[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 36.24 13.716 37.44 ;
    END
  END rddatap0[173]
  PIN rddatap0[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 36.24 18.128 37.44 ;
    END
  END rddatap0[174]
  PIN rddatap0[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 36.24 18.216 37.44 ;
    END
  END rddatap0[175]
  PIN rddatap0[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 36.96 14.616 38.16 ;
    END
  END rddatap0[176]
  PIN rddatap0[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 36.96 14.872 38.16 ;
    END
  END rddatap0[177]
  PIN rddatap0[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 36.96 18.816 38.16 ;
    END
  END rddatap0[178]
  PIN rddatap0[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 36.96 19.028 38.16 ;
    END
  END rddatap0[179]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 3.12 14.872 4.32 ;
    END
  END rddatap0[17]
  PIN rddatap0[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 37.68 13.628 38.88 ;
    END
  END rddatap0[180]
  PIN rddatap0[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 37.68 13.716 38.88 ;
    END
  END rddatap0[181]
  PIN rddatap0[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 37.68 18.128 38.88 ;
    END
  END rddatap0[182]
  PIN rddatap0[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 37.68 18.216 38.88 ;
    END
  END rddatap0[183]
  PIN rddatap0[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 38.4 14.616 39.6 ;
    END
  END rddatap0[184]
  PIN rddatap0[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 38.4 14.872 39.6 ;
    END
  END rddatap0[185]
  PIN rddatap0[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 38.4 18.816 39.6 ;
    END
  END rddatap0[186]
  PIN rddatap0[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 38.4 19.028 39.6 ;
    END
  END rddatap0[187]
  PIN rddatap0[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 39.12 13.628 40.32 ;
    END
  END rddatap0[188]
  PIN rddatap0[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 39.12 13.716 40.32 ;
    END
  END rddatap0[189]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 3.12 18.816 4.32 ;
    END
  END rddatap0[18]
  PIN rddatap0[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 39.12 18.128 40.32 ;
    END
  END rddatap0[190]
  PIN rddatap0[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 39.12 18.216 40.32 ;
    END
  END rddatap0[191]
  PIN rddatap0[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 39.84 14.616 41.04 ;
    END
  END rddatap0[192]
  PIN rddatap0[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 39.84 14.872 41.04 ;
    END
  END rddatap0[193]
  PIN rddatap0[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 39.84 18.816 41.04 ;
    END
  END rddatap0[194]
  PIN rddatap0[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 39.84 19.028 41.04 ;
    END
  END rddatap0[195]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 3.12 19.028 4.32 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 0.24 13.716 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 3.84 13.628 5.04 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 3.84 13.716 5.04 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 3.84 18.128 5.04 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 3.84 18.216 5.04 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 4.56 14.616 5.76 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 4.56 14.872 5.76 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 4.56 18.816 5.76 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 4.56 19.028 5.76 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 5.28 13.628 6.48 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 5.28 13.716 6.48 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 0.24 18.816 1.44 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 5.28 18.128 6.48 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 5.28 18.216 6.48 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6 14.616 7.2 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 6 14.872 7.2 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 6 18.816 7.2 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 6 19.028 7.2 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 6.72 13.628 7.92 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 6.72 13.716 7.92 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 6.72 18.128 7.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 6.72 18.216 7.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 0.24 19.028 1.44 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 7.44 14.616 8.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 7.44 14.872 8.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 7.44 18.816 8.64 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 7.44 19.028 8.64 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 8.16 13.628 9.36 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 8.16 13.716 9.36 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 8.16 18.128 9.36 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 8.16 18.216 9.36 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 8.88 14.616 10.08 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 8.88 14.872 10.08 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 0.96 13.972 2.16 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 8.88 18.816 10.08 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 8.88 19.028 10.08 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 9.6 13.628 10.8 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 9.6 13.716 10.8 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 9.6 18.128 10.8 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 9.6 18.216 10.8 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 10.32 14.616 11.52 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 10.32 14.872 11.52 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 10.32 18.816 11.52 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 10.32 19.028 11.52 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 0.96 14.228 2.16 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 11.04 13.628 12.24 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 11.04 13.716 12.24 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 11.04 18.128 12.24 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 11.04 18.216 12.24 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 11.76 14.616 12.96 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 11.76 14.872 12.96 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 11.76 18.816 12.96 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 11.76 19.028 12.96 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 12.48 13.628 13.68 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 12.48 13.716 13.68 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 0.96 18.128 2.16 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 12.48 18.128 13.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 12.48 18.216 13.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 13.2 14.616 14.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 13.2 14.872 14.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 13.2 18.816 14.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 13.2 19.028 14.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 13.92 13.628 15.12 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 13.92 13.716 15.12 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 13.92 18.128 15.12 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 13.92 18.216 15.12 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 0.96 18.216 2.16 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 14.64 14.616 15.84 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 14.64 14.872 15.84 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 14.64 18.816 15.84 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 14.64 19.028 15.84 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 15.36 13.628 16.56 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 15.36 13.716 16.56 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 15.36 18.128 16.56 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 15.36 18.216 16.56 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 16.08 14.616 17.28 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 16.08 14.872 17.28 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 1.68 14.616 2.88 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 16.08 18.816 17.28 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 16.08 19.028 17.28 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 16.8 13.628 18 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 16.8 13.716 18 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.084 16.8 18.128 18 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.172 16.8 18.216 18 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 17.52 14.616 18.72 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 17.52 14.872 18.72 ;
    END
  END rddatap0[97]
  PIN rddatap0[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.772 17.52 18.816 18.72 ;
    END
  END rddatap0[98]
  PIN rddatap0[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.984 17.52 19.028 18.72 ;
    END
  END rddatap0[99]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.828 1.68 14.872 2.88 ;
    END
  END rddatap0[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 18.684 21.48 18.728 22.68 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 19.072 21.48 19.116 22.68 ;
    END
  END sdl_initp0
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 33.262 0.06 33.338 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.462 0.06 31.538 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.662 0.06 29.738 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 27.862 0.06 27.938 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.062 0.06 26.138 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.262 0.06 24.338 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 22.462 0.06 22.538 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.662 0.06 20.738 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.862 0.06 18.938 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.062 0.06 17.138 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.262 0.06 15.338 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 41.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 32.362 0.06 32.438 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.562 0.06 30.638 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 28.762 0.06 28.838 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.962 0.06 27.038 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.162 0.06 25.238 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.362 0.06 23.438 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 21.562 0.06 21.638 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 19.762 0.06 19.838 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.962 0.06 18.038 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 16.162 0.06 16.238 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.362 0.06 14.438 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 41.22 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 41.22 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 19.56 16.416 20.76 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 19.56 16.672 20.76 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 19.56 16.928 20.76 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 19.56 17.016 20.76 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 19.56 17.228 20.76 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.784 19.56 17.828 20.76 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.872 19.56 17.916 20.76 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.172 19.56 15.216 20.76 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 19.56 15.772 20.76 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 0.24 15.772 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 23.28 15.772 24.48 ;
    END
  END wrdatap0[100]
  PIN wrdatap0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 23.28 16.028 24.48 ;
    END
  END wrdatap0[101]
  PIN wrdatap0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 23.28 17.316 24.48 ;
    END
  END wrdatap0[102]
  PIN wrdatap0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 23.28 17.572 24.48 ;
    END
  END wrdatap0[103]
  PIN wrdatap0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.372 24 16.416 25.2 ;
    END
  END wrdatap0[104]
  PIN wrdatap0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 24 15.428 25.2 ;
    END
  END wrdatap0[105]
  PIN wrdatap0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 24 16.928 25.2 ;
    END
  END wrdatap0[106]
  PIN wrdatap0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.972 24 17.016 25.2 ;
    END
  END wrdatap0[107]
  PIN wrdatap0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.728 24.72 15.772 25.92 ;
    END
  END wrdatap0[108]
  PIN wrdatap0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 24.72 16.028 25.92 ;
    END
  END wrdatap0[109]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 1.68 17.316 2.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 24.72 17.572 25.92 ;
    END
  END wrdatap0[110]
  PIN wrdatap0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 24.72 16.672 25.92 ;
    END
  END wrdatap0[111]
  PIN wrdatap0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 25.44 15.428 26.64 ;
    END
  END wrdatap0[112]
  PIN wrdatap0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 25.44 15.516 26.64 ;
    END
  END wrdatap0[113]
  PIN wrdatap0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.184 25.44 17.228 26.64 ;
    END
  END wrdatap0[114]
  PIN wrdatap0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 25.44 17.316 26.64 ;
    END
  END wrdatap0[115]
  PIN wrdatap0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 26.16 16.116 27.36 ;
    END
  END wrdatap0[116]
  PIN wrdatap0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 26.16 16.328 27.36 ;
    END
  END wrdatap0[117]
  PIN wrdatap0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 26.16 16.672 27.36 ;
    END
  END wrdatap0[118]
  PIN wrdatap0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 26.16 16.928 27.36 ;
    END
  END wrdatap0[119]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 1.68 17.572 2.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 26.88 15.428 28.08 ;
    END
  END wrdatap0[120]
  PIN wrdatap0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 26.88 15.516 28.08 ;
    END
  END wrdatap0[121]
  PIN wrdatap0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 26.88 17.316 28.08 ;
    END
  END wrdatap0[122]
  PIN wrdatap0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 26.88 17.572 28.08 ;
    END
  END wrdatap0[123]
  PIN wrdatap0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 27.6 16.116 28.8 ;
    END
  END wrdatap0[124]
  PIN wrdatap0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 27.6 16.328 28.8 ;
    END
  END wrdatap0[125]
  PIN wrdatap0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 27.6 16.672 28.8 ;
    END
  END wrdatap0[126]
  PIN wrdatap0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 27.6 16.928 28.8 ;
    END
  END wrdatap0[127]
  PIN wrdatap0[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 28.32 15.428 29.52 ;
    END
  END wrdatap0[128]
  PIN wrdatap0[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 28.32 15.516 29.52 ;
    END
  END wrdatap0[129]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 2.4 16.116 3.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 28.32 17.316 29.52 ;
    END
  END wrdatap0[130]
  PIN wrdatap0[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 28.32 17.572 29.52 ;
    END
  END wrdatap0[131]
  PIN wrdatap0[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 29.04 16.116 30.24 ;
    END
  END wrdatap0[132]
  PIN wrdatap0[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 29.04 16.328 30.24 ;
    END
  END wrdatap0[133]
  PIN wrdatap0[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 29.04 16.672 30.24 ;
    END
  END wrdatap0[134]
  PIN wrdatap0[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 29.04 16.928 30.24 ;
    END
  END wrdatap0[135]
  PIN wrdatap0[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 29.76 15.428 30.96 ;
    END
  END wrdatap0[136]
  PIN wrdatap0[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 29.76 15.516 30.96 ;
    END
  END wrdatap0[137]
  PIN wrdatap0[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 29.76 17.316 30.96 ;
    END
  END wrdatap0[138]
  PIN wrdatap0[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 29.76 17.572 30.96 ;
    END
  END wrdatap0[139]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 2.4 16.328 3.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 30.48 16.116 31.68 ;
    END
  END wrdatap0[140]
  PIN wrdatap0[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 30.48 16.328 31.68 ;
    END
  END wrdatap0[141]
  PIN wrdatap0[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 30.48 16.672 31.68 ;
    END
  END wrdatap0[142]
  PIN wrdatap0[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 30.48 16.928 31.68 ;
    END
  END wrdatap0[143]
  PIN wrdatap0[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 31.2 15.428 32.4 ;
    END
  END wrdatap0[144]
  PIN wrdatap0[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 31.2 15.516 32.4 ;
    END
  END wrdatap0[145]
  PIN wrdatap0[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 31.2 17.316 32.4 ;
    END
  END wrdatap0[146]
  PIN wrdatap0[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 31.2 17.572 32.4 ;
    END
  END wrdatap0[147]
  PIN wrdatap0[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 31.92 16.116 33.12 ;
    END
  END wrdatap0[148]
  PIN wrdatap0[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 31.92 16.328 33.12 ;
    END
  END wrdatap0[149]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 2.4 16.672 3.6 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 31.92 16.672 33.12 ;
    END
  END wrdatap0[150]
  PIN wrdatap0[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 31.92 16.928 33.12 ;
    END
  END wrdatap0[151]
  PIN wrdatap0[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 32.64 15.428 33.84 ;
    END
  END wrdatap0[152]
  PIN wrdatap0[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 32.64 15.516 33.84 ;
    END
  END wrdatap0[153]
  PIN wrdatap0[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 32.64 17.316 33.84 ;
    END
  END wrdatap0[154]
  PIN wrdatap0[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 32.64 17.572 33.84 ;
    END
  END wrdatap0[155]
  PIN wrdatap0[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 33.36 16.116 34.56 ;
    END
  END wrdatap0[156]
  PIN wrdatap0[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 33.36 16.328 34.56 ;
    END
  END wrdatap0[157]
  PIN wrdatap0[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 33.36 16.672 34.56 ;
    END
  END wrdatap0[158]
  PIN wrdatap0[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 33.36 16.928 34.56 ;
    END
  END wrdatap0[159]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 2.4 16.928 3.6 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 34.08 15.428 35.28 ;
    END
  END wrdatap0[160]
  PIN wrdatap0[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 34.08 15.516 35.28 ;
    END
  END wrdatap0[161]
  PIN wrdatap0[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 34.08 17.316 35.28 ;
    END
  END wrdatap0[162]
  PIN wrdatap0[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 34.08 17.572 35.28 ;
    END
  END wrdatap0[163]
  PIN wrdatap0[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 34.8 16.116 36 ;
    END
  END wrdatap0[164]
  PIN wrdatap0[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 34.8 16.328 36 ;
    END
  END wrdatap0[165]
  PIN wrdatap0[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 34.8 16.672 36 ;
    END
  END wrdatap0[166]
  PIN wrdatap0[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 34.8 16.928 36 ;
    END
  END wrdatap0[167]
  PIN wrdatap0[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 35.52 15.428 36.72 ;
    END
  END wrdatap0[168]
  PIN wrdatap0[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 35.52 15.516 36.72 ;
    END
  END wrdatap0[169]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 3.12 15.428 4.32 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 35.52 17.316 36.72 ;
    END
  END wrdatap0[170]
  PIN wrdatap0[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 35.52 17.572 36.72 ;
    END
  END wrdatap0[171]
  PIN wrdatap0[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 36.24 16.116 37.44 ;
    END
  END wrdatap0[172]
  PIN wrdatap0[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 36.24 16.328 37.44 ;
    END
  END wrdatap0[173]
  PIN wrdatap0[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 36.24 16.672 37.44 ;
    END
  END wrdatap0[174]
  PIN wrdatap0[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 36.24 16.928 37.44 ;
    END
  END wrdatap0[175]
  PIN wrdatap0[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 36.96 15.428 38.16 ;
    END
  END wrdatap0[176]
  PIN wrdatap0[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 36.96 15.516 38.16 ;
    END
  END wrdatap0[177]
  PIN wrdatap0[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 36.96 17.316 38.16 ;
    END
  END wrdatap0[178]
  PIN wrdatap0[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 36.96 17.572 38.16 ;
    END
  END wrdatap0[179]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 3.12 15.516 4.32 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 37.68 16.116 38.88 ;
    END
  END wrdatap0[180]
  PIN wrdatap0[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 37.68 16.328 38.88 ;
    END
  END wrdatap0[181]
  PIN wrdatap0[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 37.68 16.672 38.88 ;
    END
  END wrdatap0[182]
  PIN wrdatap0[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 37.68 16.928 38.88 ;
    END
  END wrdatap0[183]
  PIN wrdatap0[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 38.4 15.428 39.6 ;
    END
  END wrdatap0[184]
  PIN wrdatap0[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 38.4 15.516 39.6 ;
    END
  END wrdatap0[185]
  PIN wrdatap0[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 38.4 17.316 39.6 ;
    END
  END wrdatap0[186]
  PIN wrdatap0[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 38.4 17.572 39.6 ;
    END
  END wrdatap0[187]
  PIN wrdatap0[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 39.12 16.116 40.32 ;
    END
  END wrdatap0[188]
  PIN wrdatap0[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 39.12 16.328 40.32 ;
    END
  END wrdatap0[189]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 3.12 17.316 4.32 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 39.12 16.672 40.32 ;
    END
  END wrdatap0[190]
  PIN wrdatap0[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 39.12 16.928 40.32 ;
    END
  END wrdatap0[191]
  PIN wrdatap0[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 39.84 15.428 41.04 ;
    END
  END wrdatap0[192]
  PIN wrdatap0[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 39.84 15.516 41.04 ;
    END
  END wrdatap0[193]
  PIN wrdatap0[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 39.84 17.316 41.04 ;
    END
  END wrdatap0[194]
  PIN wrdatap0[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 39.84 17.572 41.04 ;
    END
  END wrdatap0[195]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 3.12 17.572 4.32 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 0.24 16.028 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 3.84 16.116 5.04 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 3.84 16.328 5.04 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 3.84 16.672 5.04 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 3.84 16.928 5.04 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 4.56 15.428 5.76 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 4.56 15.516 5.76 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 4.56 17.316 5.76 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 4.56 17.572 5.76 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 5.28 16.116 6.48 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 5.28 16.328 6.48 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 0.24 17.316 1.44 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 5.28 16.672 6.48 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 5.28 16.928 6.48 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 6 15.428 7.2 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 6 15.516 7.2 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 6 17.316 7.2 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 6 17.572 7.2 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 6.72 16.116 7.92 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 6.72 16.328 7.92 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 6.72 16.672 7.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 6.72 16.928 7.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 0.24 17.572 1.44 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 7.44 15.428 8.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 7.44 15.516 8.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 7.44 17.316 8.64 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 7.44 17.572 8.64 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 8.16 16.116 9.36 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 8.16 16.328 9.36 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 8.16 16.672 9.36 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 8.16 16.928 9.36 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 8.88 15.428 10.08 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 8.88 15.516 10.08 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 0.96 16.116 2.16 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 8.88 17.316 10.08 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 8.88 17.572 10.08 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 9.6 16.116 10.8 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 9.6 16.328 10.8 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 9.6 16.672 10.8 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 9.6 16.928 10.8 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 10.32 15.428 11.52 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 10.32 15.516 11.52 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 10.32 17.316 11.52 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 10.32 17.572 11.52 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 0.96 16.328 2.16 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 11.04 16.116 12.24 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 11.04 16.328 12.24 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 11.04 16.672 12.24 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 11.04 16.928 12.24 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 11.76 15.428 12.96 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 11.76 15.516 12.96 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 11.76 17.316 12.96 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 11.76 17.572 12.96 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 12.48 16.116 13.68 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 12.48 16.328 13.68 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 0.96 16.672 2.16 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 12.48 16.672 13.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 12.48 16.928 13.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 13.2 15.428 14.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 13.2 15.516 14.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 13.2 17.316 14.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 13.2 17.572 14.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 13.92 16.116 15.12 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 13.92 16.328 15.12 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 13.92 16.672 15.12 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 13.92 16.928 15.12 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 0.96 16.928 2.16 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 14.64 15.428 15.84 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 14.64 15.516 15.84 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 14.64 17.316 15.84 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 14.64 17.572 15.84 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 15.36 16.116 16.56 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 15.36 16.328 16.56 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 15.36 16.672 16.56 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 15.36 16.928 16.56 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 16.08 15.428 17.28 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 16.08 15.516 17.28 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 1.68 15.428 2.88 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 16.08 17.316 17.28 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 16.08 17.572 17.28 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 16.8 16.116 18 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 16.8 16.328 18 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.628 16.8 16.672 18 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.884 16.8 16.928 18 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.384 17.52 15.428 18.72 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 17.52 15.516 18.72 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.272 17.52 17.316 18.72 ;
    END
  END wrdatap0[98]
  PIN wrdatap0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 17.528 17.52 17.572 18.72 ;
    END
  END wrdatap0[99]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.472 1.68 15.516 2.88 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.072 19.56 16.116 20.76 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 16.284 19.56 16.328 20.76 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 15.984 19.56 16.028 20.76 ;
    END
  END wrenp0
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 34.2 41.28 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 34.2 41.28 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 34.2705 41.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 34.235 41.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 34.27 41.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 34.259 41.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 34.29 41.342 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 34.292 41.34 ;
  END
END arf192b080e1r1w0cbbehbaa4acw
END LIBRARY
