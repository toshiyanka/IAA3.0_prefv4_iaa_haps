VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

MACRO arf074b064e1r1w0cbbehsaa4acw
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN arf074b064e1r1w0cbbehsaa4acw 0 0 ;
  SIZE 14.4 BY 32.64 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 16.68 3.172 17.88 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 14.76 0.728 15.96 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 16.68 0.472 17.88 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 16.68 0.728 17.88 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 16.68 0.816 17.88 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 16.68 1.028 17.88 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 16.68 1.116 17.88 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 16.68 1.372 17.88 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.68 3.516 17.88 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 16.68 3.728 17.88 ;
    END
  END rdaddrp0_rd
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 0.24 3.516 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.84 3.516 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.84 3.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.56 3.428 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 4.56 3.816 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 5.28 3.172 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.28 3.516 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6 4.328 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6 3.428 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 6.72 3.816 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.72 4.072 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.24 3.728 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.44 3.516 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 7.44 3.728 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 8.16 3.428 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 8.16 3.816 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 8.88 3.172 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.88 3.516 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.6 4.328 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9.6 3.428 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 10.32 3.816 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 10.32 4.072 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.96 3.428 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.04 3.516 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 11.04 3.728 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 11.76 3.428 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 11.76 3.816 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 12.48 3.172 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.48 3.516 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 13.2 4.328 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 13.2 3.428 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 18.24 4.328 19.44 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 18.24 3.428 19.44 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 0.96 3.816 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 18.96 3.816 20.16 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 18.96 4.072 20.16 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.68 3.516 20.88 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 19.68 3.728 20.88 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.4 3.428 21.6 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 20.4 3.816 21.6 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 21.12 3.172 22.32 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 21.12 3.516 22.32 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 21.84 4.328 23.04 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 21.84 3.428 23.04 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 1.68 3.172 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 22.56 3.816 23.76 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 22.56 4.072 23.76 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 23.28 3.516 24.48 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 23.28 3.728 24.48 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 24 3.428 25.2 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 24 3.816 25.2 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 24.72 3.172 25.92 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 24.72 3.516 25.92 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 25.44 4.328 26.64 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 25.44 3.428 26.64 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 1.68 3.516 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 26.16 3.816 27.36 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 26.16 4.072 27.36 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 26.88 3.516 28.08 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 26.88 3.728 28.08 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 27.6 3.428 28.8 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 27.6 3.816 28.8 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 28.32 3.172 29.52 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 28.32 3.516 29.52 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 29.04 4.328 30.24 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 29.04 3.428 30.24 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 2.4 4.328 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 29.76 3.816 30.96 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 29.76 4.072 30.96 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 30.48 3.516 31.68 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 30.48 3.728 31.68 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 31.2 3.428 32.4 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 31.2 3.816 32.4 ;
    END
  END rddatap0[75]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.4 3.428 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 3.12 3.816 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 3.12 4.072 4.32 ;
    END
  END rddatap0[9]
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 16.68 3.816 17.88 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.68 4.072 17.88 ;
    END
  END sdl_initp0
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 13.462 0.06 13.538 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.662 0.06 11.738 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.862 0.06 9.938 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.062 0.06 8.138 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.262 0.06 6.338 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.462 0.06 4.538 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.662 0.06 2.738 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 32.58 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 12.562 0.06 12.638 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.762 0.06 10.838 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.962 0.06 9.038 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.162 0.06 7.238 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.362 0.06 5.438 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.562 0.06 3.638 32.58 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 32.58 ;
    END
  END vss
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 14.76 1.716 15.96 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 14.76 1.928 15.96 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 14.76 2.016 15.96 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.76 2.616 15.96 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 14.76 2.828 15.96 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 14.76 2.916 15.96 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 14.76 0.816 15.96 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 14.76 1.028 15.96 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.24 1.928 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 3.84 1.928 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 3.84 2.272 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 4.56 2.916 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 4.56 2.016 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.28 2.616 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.28 2.828 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 6 2.272 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6 2.528 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 6.72 2.016 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 6.72 2.616 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 0.24 2.016 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 7.44 1.928 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 7.44 2.272 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 8.16 2.916 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 8.16 2.016 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 8.88 2.616 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 8.88 2.828 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 9.6 2.272 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 9.6 2.528 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 10.32 2.016 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 10.32 2.616 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.96 2.916 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 11.04 1.928 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 11.04 2.272 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 11.76 2.916 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 11.76 2.016 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 12.48 2.616 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12.48 2.828 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 13.2 2.272 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 13.2 2.528 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 18.24 2.916 19.44 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 18.24 1.928 19.44 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.96 2.272 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 18.96 2.272 20.16 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 18.96 2.528 20.16 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 19.68 1.928 20.88 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 19.68 2.016 20.88 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 20.4 2.916 21.6 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 20.4 2.272 21.6 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 21.12 2.616 22.32 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 21.12 2.828 22.32 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 21.84 2.272 23.04 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 21.84 2.528 23.04 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 1.68 2.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 22.56 2.016 23.76 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 22.56 2.616 23.76 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 23.28 1.928 24.48 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 23.28 2.272 24.48 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 24 2.916 25.2 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 24 2.016 25.2 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 24.72 2.616 25.92 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 24.72 2.828 25.92 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 25.44 2.272 26.64 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 25.44 2.528 26.64 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 1.68 2.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 26.16 2.016 27.36 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 26.16 2.616 27.36 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 26.88 1.928 28.08 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 26.88 2.272 28.08 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 27.6 2.916 28.8 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 27.6 2.016 28.8 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 28.32 2.616 29.52 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 28.32 2.828 29.52 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 29.04 2.272 30.24 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 29.04 2.528 30.24 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 2.4 2.272 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 29.76 2.016 30.96 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 29.76 2.616 30.96 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 30.48 1.928 31.68 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 30.48 2.272 31.68 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 31.2 2.916 32.4 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 31.2 2.016 32.4 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.4 2.528 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 3.12 2.016 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.12 2.616 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 14.76 1.372 15.96 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 14.76 1.628 15.96 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 14.76 1.116 15.96 ;
    END
  END wrenp0
  OBS
    LAYER m0 SPACING 0 ;
      RECT 0 0 14.4 32.64 ;
    LAYER m1 SPACING 0 ;
      RECT 0 0 14.4 32.64 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 14.4705 32.678 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 14.435 32.71 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 14.47 32.678 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 14.459 32.73 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 14.49 32.702 ;
    LAYER m7 SPACING 0 ;
      RECT -0.092 -0.06 14.492 32.7 ;
  END
END arf074b064e1r1w0cbbehsaa4acw
END LIBRARY
