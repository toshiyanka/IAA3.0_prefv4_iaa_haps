//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2021 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//  
//  Collateral Description:
//  IOSF - Sideband Channel IP
//  
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//  
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//  
//  Revision:
//  2021WW02_PICr35
//  
//  Module sbr2 : 
//
//         This is a project specific RTL wrapper for the IOSF sideband
//         channel synchronous N-Port router.
//
//  This RTL file generated by: ../../unsupported/gen/sbccfg rev 0.61
//  Fabric configuration file:  ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv rev -1.00
//
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
// The Router Module
//
//------------------------------------------------------------------------------
  // lintra push -80099, -80009, -80018, -70023

module sbr2
(
  // Synchronous Clock/Reset
  iosf_swf_side_clk,
  iosf_swf_side_rst_b,

  // Power Well Isolation Input Signals
  eva_present,

  p0_fab_init_idle_exit,
  p0_fab_init_idle_exit_ack,
  p1_fab_init_idle_exit,
  p1_fab_init_idle_exit_ack,
  p2_fab_init_idle_exit,
  p2_fab_init_idle_exit_ack,
  sbr_idle,

  // VISA Debug Interface IO
  visa_all_disable,
  visa_customer_disable,
  avisa_data_out,
  avisa_clk_out,
  visa_ser_cfg_in,
  visa_arb_iosf_swf_side_clk,
  visa_vp_iosf_swf_side_clk,
  visa_p0_tier1_iosf_swf_side_clk,
  visa_p0_tier2_iosf_swf_side_clk,
  visa_p1_tier1_iosf_swf_side_clk,
  visa_p1_tier2_iosf_swf_side_clk,
  visa_p2_tier1_iosf_swf_side_clk,
  visa_p2_tier2_iosf_swf_side_clk,


  // Register wires
  dfxa_sbr2_cgovrd,
  dfxa_sbr2_cgctrl,

  fscan_mode,
  fscan_clkungate,
  fscan_clkungate_syn,
  fscan_rstbypen,
  fscan_byprst_b,
  // Port 0 declarations
  sbr1_sbr2_side_ism_agent,
  sbr2_sbr1_side_ism_fabric,
  sbr1_sbr2_pccup,
  sbr1_sbr2_npcup,
  sbr2_sbr1_pcput,
  sbr2_sbr1_npput,
  sbr2_sbr1_eom,
  sbr2_sbr1_payload,
  sbr2_sbr1_pccup,
  sbr2_sbr1_npcup,
  sbr1_sbr2_pcput,
  sbr1_sbr2_npput,
  sbr1_sbr2_eom,
  sbr1_sbr2_payload,

  // Port 1 declarations
  xut_sbr2_side_ism_agent,
  sbr2_xut_side_ism_fabric,
  xut_sbr2_pccup,
  xut_sbr2_npcup,
  sbr2_xut_pcput,
  sbr2_xut_npput,
  sbr2_xut_eom,
  sbr2_xut_payload,
  sbr2_xut_pccup,
  sbr2_xut_npcup,
  xut_sbr2_pcput,
  xut_sbr2_npput,
  xut_sbr2_eom,
  xut_sbr2_payload,

  // Port 2 declarations
  swf_sbr2_side_ism_agent,
  sbr2_swf_side_ism_fabric,
  swf_sbr2_pccup,
  swf_sbr2_npcup,
  sbr2_swf_pcput,
  sbr2_swf_npput,
  sbr2_swf_eom,
  sbr2_swf_payload,
  sbr2_swf_pccup,
  sbr2_swf_npcup,
  swf_sbr2_pcput,
  swf_sbr2_npput,
  swf_sbr2_eom,
  swf_sbr2_payload);


`include "sbcglobal_params.vm"
`include "sbcstruct_local.vm"

  parameter SBR_VISA_ID_PARAM = 11;
  parameter NUMBER_OF_BITS_PER_LANE = 8;
  parameter NUMBER_OF_VISAMUX_MODULES = 1;
  parameter NUMBER_OF_OUTPUT_LANES = (NUMBER_OF_VISAMUX_MODULES == 1)? 2 : NUMBER_OF_VISAMUX_MODULES;

  input logic iosf_swf_side_clk;
  input logic iosf_swf_side_rst_b;

  // Power Well Isolation Input Signals
  input logic eva_present;

  output logic p0_fab_init_idle_exit;
  input logic p0_fab_init_idle_exit_ack;
  output logic p1_fab_init_idle_exit;
  input logic p1_fab_init_idle_exit_ack;
  output logic p2_fab_init_idle_exit;
  input logic p2_fab_init_idle_exit_ack;
  output logic sbr_idle;

  // VISA Debug Interface IO
  input logic visa_all_disable;
  input logic visa_customer_disable;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0][(NUMBER_OF_BITS_PER_LANE-1):0] avisa_data_out;
  output logic [(NUMBER_OF_OUTPUT_LANES-1):0] avisa_clk_out;
  input logic [2:0] visa_ser_cfg_in;

  // VISA Debug Signal/Clock Structs
  output visa_arb visa_arb_iosf_swf_side_clk;
  output visa_vp  visa_vp_iosf_swf_side_clk;
  output visa_port_tier1 visa_p0_tier1_iosf_swf_side_clk;
  output visa_port_tier2 visa_p0_tier2_iosf_swf_side_clk;
  output visa_port_tier1 visa_p1_tier1_iosf_swf_side_clk;
  output visa_port_tier2 visa_p1_tier2_iosf_swf_side_clk;
  output visa_port_tier1 visa_p2_tier1_iosf_swf_side_clk;
  output visa_port_tier2 visa_p2_tier2_iosf_swf_side_clk;

  // Register wires
  input logic [4:0]  dfxa_sbr2_cgovrd;
  input logic [15:0] dfxa_sbr2_cgctrl;

  input logic fscan_mode;
  input logic fscan_clkungate;
  input logic fscan_clkungate_syn;
  input logic fscan_rstbypen;
  input logic fscan_byprst_b;
  // Port 0 declarations
  input logic [2:0] sbr1_sbr2_side_ism_agent;
  output logic [2:0] sbr2_sbr1_side_ism_fabric;
  input logic sbr1_sbr2_pccup;
  input logic sbr1_sbr2_npcup;
  output logic sbr2_sbr1_pcput;
  output logic sbr2_sbr1_npput;
  output logic sbr2_sbr1_eom;
  output logic [7:0] sbr2_sbr1_payload;
  output logic sbr2_sbr1_pccup;
  output logic sbr2_sbr1_npcup;
  input logic sbr1_sbr2_pcput;
  input logic sbr1_sbr2_npput;
  input logic sbr1_sbr2_eom;
  input logic [7:0] sbr1_sbr2_payload;

  // Port 1 declarations
  input logic [2:0] xut_sbr2_side_ism_agent;
  output logic [2:0] sbr2_xut_side_ism_fabric;
  input logic xut_sbr2_pccup;
  input logic xut_sbr2_npcup;
  output logic sbr2_xut_pcput;
  output logic sbr2_xut_npput;
  output logic sbr2_xut_eom;
  output logic [7:0] sbr2_xut_payload;
  output logic sbr2_xut_pccup;
  output logic sbr2_xut_npcup;
  input logic xut_sbr2_pcput;
  input logic xut_sbr2_npput;
  input logic xut_sbr2_eom;
  input logic [7:0] xut_sbr2_payload;

  // Port 2 declarations
  input logic [2:0] swf_sbr2_side_ism_agent;
  output logic [2:0] sbr2_swf_side_ism_fabric;
  input logic swf_sbr2_pccup;
  input logic swf_sbr2_npcup;
  output logic sbr2_swf_pcput;
  output logic sbr2_swf_npput;
  output logic sbr2_swf_eom;
  output logic [7:0] sbr2_swf_payload;
  output logic sbr2_swf_pccup;
  output logic sbr2_swf_npcup;
  input logic swf_sbr2_pcput;
  input logic swf_sbr2_npput;
  input logic swf_sbr2_eom;
  input logic [7:0] swf_sbr2_payload;



//------------------------------------------------------------------------------
//
// Router Port Map Table
//
//------------------------------------------------------------------------------
logic [255:0][16:0] sbr2_sbcportmap;
always_comb sbr2_sbcportmap = {

      //-----------------------------------------------------    SBCPORTMAPTABLE
      //  Module:  sbr2 (sbr2)                                   SBCPORTMAPTABLE
      //  Ports:   M 1111 11                                     SBCPORTMAPTABLE
      //           C 5432 1098 7654 3210           Port ID       SBCPORTMAPTABLE
      //---------------------------------------//                SBCPORTMAPTABLE
               17'b1_1111_1111_1111_1111,      //   255          SBCPORTMAPTABLE
      {   15 { 17'b0_0000_0000_0000_0000 }},   //   254:240      SBCPORTMAPTABLE
      {    2 { 17'b0_0000_0000_0000_0001 }},   //   239:238      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //   237          SBCPORTMAPTABLE
      {    3 { 17'b0_0000_0000_0000_0001 }},   //   236:234      SBCPORTMAPTABLE
      {  224 { 17'b0_0000_0000_0000_0000 }},   //   233: 10      SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0100,      //     9          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0010,      //     8          SBCPORTMAPTABLE
               17'b0_0000_0000_0000_0000,      //     7          SBCPORTMAPTABLE
      {    7 { 17'b0_0000_0000_0000_0001 }}    //     6:  0      SBCPORTMAPTABLE
    };

//------------------------------------------------------------------------------
//
// Local Parameters
//
//------------------------------------------------------------------------------
localparam MAXPORT      =  2;
localparam INTMAXPLDBIT = 31;

//------------------------------------------------------------------------------
//
// Signal declarations
//
//------------------------------------------------------------------------------

// Router Port Arrays
logic [MAXPORT:0]                  agent_idle;
logic [MAXPORT:0]                  port_idle;
logic [MAXPORT:0]                  pctrdy;
logic [MAXPORT:0]                  pcirdy;
logic [MAXPORT:0]                  pceom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] pcdata;
logic [MAXPORT:0]                  pcdstvld;
logic                              p0_pcdstvld;
logic                              p1_pcdstvld;
logic                              p2_pcdstvld;

logic [MAXPORT:0]                  nptrdy;
logic [MAXPORT:0]                  npirdy;
logic [MAXPORT:0]                  npfence;
logic                              p0_npfence;
logic                              p1_npfence;
logic                              p2_npfence;
logic [MAXPORT:0]                  npeom;
logic [MAXPORT:0] [INTMAXPLDBIT:0] npdata;
logic [MAXPORT:0]                  npdstvld;
logic                              p0_npdstvld;
logic                              p1_npdstvld;
logic                              p2_npdstvld;

logic [MAXPORT:0]                  epctrdy;
logic [MAXPORT:0]                  enptrdy;
logic [MAXPORT:0]                  epcirdy;
logic [MAXPORT:0]                  enpirdy;

// Datapath
logic [MAXPORT:0]                  portmapgnt;
logic [MAXPORT:0]                  pcportmapdone;
logic [MAXPORT:0]                  npportmapdone;
logic                              destnp;
logic                              eom;
logic             [INTMAXPLDBIT:0] data;

// Virtual Port Signals
logic                              pctrdy_vp;
logic                              pcirdy_vp;
logic                              pceom_vp;
logic             [INTMAXPLDBIT:0] pcdata_vp;
logic [MAXPORT:0]                  pcdstvec_vp;
logic                              enptrdy_vp;
logic                              epcirdy_vp;
logic                              enpirdy_vp;
logic [MAXPORT:0]                  enpirdy_pwrdn;

// Port Mapping Signals
logic                       [ 7:0] destportid;
logic [MAXPORT:0]                  destvector;
logic                              multicast;
logic                              dest0xFE;

logic [MAXPORT:0]                  endpoint_pwrgd ;
logic                              p0_ism_idle;
logic                              p0_cg_inprogress;
logic                              p0_credit_reinit;
logic                              p1_ism_idle;
logic                              p1_cg_inprogress;
logic                              p1_credit_reinit;
logic                              p2_ism_idle;
logic                              p2_cg_inprogress;
logic                              p2_credit_reinit;
logic                              all_idle;
logic                              arbiter_idle;
logic                              gated_side_clk;
logic                       [31:0] dbgbus_arb;
logic                       [31:0] dbgbus_vp;
logic                              eva_present_ff2;

logic                              cfg_clkgaten;
logic                              cfg_clkgatedef;
logic                        [7:0] cfg_idlecnt;
logic                              jta_clkgate_ovrd;
logic                              jta_force_idle;
logic                              jta_force_notidle;
logic                              jta_force_creditreq;
logic                              force_idle;
logic                              force_notidle;
logic                              force_creditreq;

always_comb cfg_clkgaten      = dfxa_sbr2_cgctrl[15];
always_comb cfg_clkgatedef    = dfxa_sbr2_cgctrl[14];
always_comb cfg_idlecnt       = dfxa_sbr2_cgctrl[7:0];
always_comb jta_clkgate_ovrd  = dfxa_sbr2_cgovrd[3];
always_comb jta_force_idle    = dfxa_sbr2_cgovrd[1];
always_comb jta_force_notidle = dfxa_sbr2_cgovrd[0];
always_comb jta_force_creditreq = dfxa_sbr2_cgovrd[4];

logic                              fscan_latchopen;
logic                              fscan_latchclosed_b;

always_comb fscan_latchopen     = '0;
always_comb fscan_latchclosed_b = '1;

//------------------------------------------------------------------------------
//
// Destination Port ID to Egress Vector Mapping
//
//------------------------------------------------------------------------------
always_comb destvector = sbr2_sbcportmap[destportid][MAXPORT:0];
always_comb multicast  = sbr2_sbcportmap[destportid][16];

//------------------------------------------------------------------------------
//
// DFx clock syncs
//
//------------------------------------------------------------------------------
sbc_doublesync sync_force_idle (
  .d                   ( jta_force_idle                ),
  .clr_b               ( iosf_swf_side_rst_b           ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( force_idle                    )
);

sbc_doublesync sync_force_notidle (
  .d                   ( jta_force_notidle             ),
  .clr_b               ( iosf_swf_side_rst_b           ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( force_notidle                 )
);

sbc_doublesync sync_force_creditreq (
  .d                   ( jta_force_creditreq           ),
  .clr_b               ( iosf_swf_side_rst_b           ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( force_creditreq               )
);

//------------------------------------------------------------------------------
//
// Power well isolation signal synchronizers
//
//------------------------------------------------------------------------------
sbc_doublesync sync_eva_present (
  .d                   ( eva_present                   ),
  .clr_b               ( iosf_swf_side_rst_b           ),
  .clk                 ( iosf_swf_side_clk             ),
  .q                   ( eva_present_ff2               )
);


always_comb endpoint_pwrgd = { 1'b1,
                          1'b1,
                          eva_present_ff2
                        };

logic p0_gated_clk;
sbc_clock_gate p0_pwr_clkgate  (
  .en ( endpoint_pwrgd[0] ),
  .te                  ( fscan_clkungate               ),
  .clk                 ( gated_side_clk                ),
  .enclk ( p0_gated_clk )
);

//------------------------------------------------------------------------------
//
// ISM idle signal for all synchronous port ISMs
//
//------------------------------------------------------------------------------
always_comb all_idle =   &(port_idle | ~endpoint_pwrgd)
                  &  (p2_ism_idle | ~endpoint_pwrgd[2])
                  &  (p1_ism_idle | ~endpoint_pwrgd[1])
                  &  (p0_ism_idle | ~endpoint_pwrgd[0]);

// ISM IDLE cross into router clock domain
// SBR_IDLE signal for PMU
  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if (~iosf_swf_side_rst_b)
      sbr_idle <= '0;
    else
      sbr_idle <= arbiter_idle & all_idle &
                  p0_ism_idle &
                  p1_ism_idle &
                  p2_ism_idle;

//------------------------------------------------------------------------------
//
// The router datapath and destination port ID selection
//
//------------------------------------------------------------------------------
always_comb begin : sbcrouterdp
  destportid = '0;
  destnp     = '0;
  eom        = pctrdy_vp ? pceom_vp  : '0;
  data       = pctrdy_vp ? pcdata_vp : '0;
  for (int i=0; i<=MAXPORT; i++) begin
    if (portmapgnt[i]) begin
      destportid |= npdstvld[i] & ~npportmapdone[i] & ~npfence[i]
                    ? npdata[i][7:0]
                    : pcdstvld[i] & ~pcportmapdone[i]
                      ? pcdata[i][7:0] : npdata[i][7:0];
      destnp |= npdstvld[i] & ~npportmapdone[i] &
                (~npfence[i] | ~pcdstvld[i] | pcportmapdone[i]);
    end
    if (pctrdy[i]) begin
      eom  |= pceom[i];
      data |= pcdata[i];
    end
    if (nptrdy[i]) begin
      eom  |= npeom[i];
      data |= npdata[i];
    end
  end
end

always_comb dest0xFE = destportid == 8'hFE;

always_comb
  begin
    npfence = { 
                 p2_npfence,
                 p1_npfence,
                 p0_npfence
               };
  end

always_comb
  begin
    pcdstvld = { 
                 p2_pcdstvld,
                 p1_pcdstvld,
                 p0_pcdstvld
               };
  end

always_comb
  begin
    npdstvld = { 
                 p2_npdstvld,
                 p1_npdstvld,
                 p0_npdstvld
               };
  end

//------------------------------------------------------------------------------
//
// The arbiter instantiation
//
//------------------------------------------------------------------------------

logic [MAXPORT:0] rsp_scbd;

always_comb visa_arb_iosf_swf_side_clk = dbgbus_arb;
sbcarbiter #(
  .MAXPORT             ( MAXPORT                       ),
  .FASTPEND2IP         (  0                            ),
  .PIPELINE            (  1                            )
) sbcarbiter (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( iosf_swf_side_clk             ),
  .side_rst_b          ( iosf_swf_side_rst_b           ),
  .endpoint_pwrgd      ( endpoint_pwrgd                ),
  .all_idle            ( all_idle                      ),
  .agent_idle          ( agent_idle                    ),
  .gated_side_clk      ( gated_side_clk                ),
  .arbiter_idle        ( arbiter_idle                  ),
  .jta_clkgate_ovrd    ( jta_clkgate_ovrd              ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .cfg_clkgatedef      ( cfg_clkgatedef                ),
  .cfg_idlecnt         ( cfg_idlecnt                   ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .pcdstvld            ( pcdstvld                      ),
  .npdstvld            ( npdstvld                      ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcirdy              ( pcirdy                        ),
  .npirdy              ( npirdy                        ),
  .npfence             ( npfence                       ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .portmapgnt          ( portmapgnt                    ),
  .pcportmapdone       ( pcportmapdone                 ),
  .npportmapdone       ( npportmapdone                 ),
  .multicast           ( multicast                     ),
  .destvector          ( destvector                    ),
  .destnp              ( destnp                        ),
  .dest0xFE            ( dest0xFE                      ),
  .eom                 ( eom                           ),
  .epctrdy             ( epctrdy                       ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .enptrdy             ( enptrdy                       ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .epcirdy             ( epcirdy                       ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .su_local_ugt        ( fscan_clkungate               ),
  .dbgbus              ( dbgbus_arb                    )
);

//------------------------------------------------------------------------------
//
// The virtual port instantiation
//
//------------------------------------------------------------------------------
always_comb visa_vp_iosf_swf_side_clk = dbgbus_vp;
sbcvirtport #(
  .MAXPORT             ( MAXPORT                       ),
  .INTMAXPLDBIT        ( INTMAXPLDBIT                  )
) sbcvirtport (
  .rsp_scbd            ( rsp_scbd                      ),
  .side_clk            ( gated_side_clk                ),
  .side_rst_b          ( iosf_swf_side_rst_b           ),
  .pctrdy_vp           ( pctrdy_vp                     ),
  .pcirdy_vp           ( pcirdy_vp                     ),
  .pcdata_vp           ( pcdata_vp                     ),
  .pceom_vp            ( pceom_vp                      ),
  .pcdstvec_vp         ( pcdstvec_vp                   ),
  .eom                 ( eom                           ),
  .data                ( data                          ),
  .enptrdy_vp          ( enptrdy_vp                    ),
  .epcirdy_vp          ( epcirdy_vp                    ),
  .enpirdy_vp          ( enpirdy_vp                    ),
  .enpirdy             ( enpirdy                       ),
  .enpirdy_pwrdn       ( enpirdy_pwrdn                 ),
  .pctrdy              ( pctrdy                        ),
  .nptrdy              ( nptrdy                        ),
  .dbgbus              ( dbgbus_vp                     )
);

//------------------------------------------------------------------------------
//
// Instantiation of the sideband port (fabric ISMs, ingress/egress port)
//
//------------------------------------------------------------------------------

// Port 0
logic p0_side_clk_valid, p0_idle_egress, p0_rst_suppress;
  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p0_rst_suppress <= 1'b1;
    else
      p0_rst_suppress <= p0_credit_reinit & p0_rst_suppress;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if (~iosf_swf_side_rst_b)
      p0_fab_init_idle_exit <= '1;
    else
      if ( ~p0_rst_suppress & (p0_ism_idle & (~agent_idle[0] || ~p0_idle_egress) & ~p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '1;
      else if ( ~p0_rst_suppress & (p0_ism_idle & agent_idle[0] & p0_fab_init_idle_exit_ack ))
        p0_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p0_side_clk_valid <= 1'b0;
    else
      begin
        if ( p0_ism_idle & p0_side_clk_valid )
          p0_side_clk_valid <= '0;
        else if ( (p0_fab_init_idle_exit & p0_fab_init_idle_exit_ack) || ~p0_ism_idle )
          p0_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p0_dbgbus;

  always_comb
    begin
      visa_p0_tier1_iosf_swf_side_clk = { p0_dbgbus[31],
                            p0_dbgbus[27:24],
                            p0_dbgbus[21:19],
                            p0_dbgbus[15:12],
                            p0_dbgbus[7:4] };
      visa_p0_tier2_iosf_swf_side_clk = { p0_dbgbus[30:28],
                            p0_dbgbus[23:22],
                            p0_dbgbus[18:16],
                            p0_dbgbus[11:8],
                            p0_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport0 (
  .side_clk            ( iosf_swf_side_clk             ),
  .gated_side_clk      ( p0_gated_clk                  ),
  .side_rst_b          ( iosf_swf_side_rst_b           ),
  .side_clk_valid      ( p0_side_clk_valid             ),
  .side_ism_in         ( sbr1_sbr2_side_ism_agent      ),
  .side_ism_out        ( sbr2_sbr1_side_ism_fabric     ),
  .int_pok             ( endpoint_pwrgd[0] ),
  .agent_idle          ( agent_idle[0]                 ),
  .port_idle           ( port_idle[0]                  ),
  .idle_egress         ( p0_idle_egress                ),
  .ism_idle            ( p0_ism_idle                   ),
  .credit_reinit       ( p0_credit_reinit              ),
  .cg_inprogress       ( p0_cg_inprogress              ),
  .tpccup              ( sbr2_sbr1_pccup               ),
  .tnpcup              ( sbr2_sbr1_npcup               ),
  .tpcput              ( sbr1_sbr2_pcput               ),
  .tnpput              ( sbr1_sbr2_npput               ),
  .teom                ( sbr1_sbr2_eom                 ),
  .tpayload            ( sbr1_sbr2_payload             ),
  .pctrdy              ( pctrdy[0]                     ),
  .pcirdy              ( pcirdy[0]                     ),
  .pcdata              ( pcdata[0]                     ),
  .pceom               ( pceom[0]                      ),
  .pcdstvld            ( p0_pcdstvld                   ),
  .nptrdy              ( nptrdy[0]                     ),
  .npirdy              ( npirdy[0]                     ),
  .npfence             ( p0_npfence                    ),
  .npdata              ( npdata[0]                     ),
  .npeom               ( npeom[0]                      ),
  .npdstvld            ( p0_npdstvld                   ),
  .mpccup              ( sbr1_sbr2_pccup               ),
  .mnpcup              ( sbr1_sbr2_npcup               ),
  .mpcput              ( sbr2_sbr1_pcput               ),
  .mnpput              ( sbr2_sbr1_npput               ),
  .meom                ( sbr2_sbr1_eom                 ),
  .mpayload            ( sbr2_sbr1_payload             ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[0]                    ),
  .enptrdy             ( enptrdy[0]                    ),
  .epcirdy             ( epcirdy[0]                    ),
  .enpirdy             ( enpirdy[0]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p0_dbgbus                     )
);

// Port 1
logic p1_side_clk_valid, p1_idle_egress, p1_rst_suppress;
  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p1_rst_suppress <= 1'b1;
    else
      p1_rst_suppress <= p1_credit_reinit & p1_rst_suppress;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if (~iosf_swf_side_rst_b)
      p1_fab_init_idle_exit <= '1;
    else
      if ( ~p1_rst_suppress & (p1_ism_idle & (~agent_idle[1] || ~p1_idle_egress) & ~p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '1;
      else if ( ~p1_rst_suppress & (p1_ism_idle & agent_idle[1] & p1_fab_init_idle_exit_ack ))
        p1_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p1_side_clk_valid <= 1'b0;
    else
      begin
        if ( p1_ism_idle & p1_side_clk_valid )
          p1_side_clk_valid <= '0;
        else if ( (p1_fab_init_idle_exit & p1_fab_init_idle_exit_ack) || ~p1_ism_idle )
          p1_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p1_dbgbus;

  always_comb
    begin
      visa_p1_tier1_iosf_swf_side_clk = { p1_dbgbus[31],
                            p1_dbgbus[27:24],
                            p1_dbgbus[21:19],
                            p1_dbgbus[15:12],
                            p1_dbgbus[7:4] };
      visa_p1_tier2_iosf_swf_side_clk = { p1_dbgbus[30:28],
                            p1_dbgbus[23:22],
                            p1_dbgbus[18:16],
                            p1_dbgbus[11:8],
                            p1_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport1 (
  .side_clk            ( iosf_swf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_swf_side_rst_b           ),
  .side_clk_valid      ( p1_side_clk_valid             ),
  .side_ism_in         ( xut_sbr2_side_ism_agent       ),
  .side_ism_out        ( sbr2_xut_side_ism_fabric      ),
  .int_pok             ( endpoint_pwrgd[1] ),
  .agent_idle          ( agent_idle[1]                 ),
  .port_idle           ( port_idle[1]                  ),
  .idle_egress         ( p1_idle_egress                ),
  .ism_idle            ( p1_ism_idle                   ),
  .credit_reinit       ( p1_credit_reinit              ),
  .cg_inprogress       ( p1_cg_inprogress              ),
  .tpccup              ( sbr2_xut_pccup                ),
  .tnpcup              ( sbr2_xut_npcup                ),
  .tpcput              ( xut_sbr2_pcput                ),
  .tnpput              ( xut_sbr2_npput                ),
  .teom                ( xut_sbr2_eom                  ),
  .tpayload            ( xut_sbr2_payload              ),
  .pctrdy              ( pctrdy[1]                     ),
  .pcirdy              ( pcirdy[1]                     ),
  .pcdata              ( pcdata[1]                     ),
  .pceom               ( pceom[1]                      ),
  .pcdstvld            ( p1_pcdstvld                   ),
  .nptrdy              ( nptrdy[1]                     ),
  .npirdy              ( npirdy[1]                     ),
  .npfence             ( p1_npfence                    ),
  .npdata              ( npdata[1]                     ),
  .npeom               ( npeom[1]                      ),
  .npdstvld            ( p1_npdstvld                   ),
  .mpccup              ( xut_sbr2_pccup                ),
  .mnpcup              ( xut_sbr2_npcup                ),
  .mpcput              ( sbr2_xut_pcput                ),
  .mnpput              ( sbr2_xut_npput                ),
  .meom                ( sbr2_xut_eom                  ),
  .mpayload            ( sbr2_xut_payload              ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[1]                    ),
  .enptrdy             ( enptrdy[1]                    ),
  .epcirdy             ( epcirdy[1]                    ),
  .enpirdy             ( enpirdy[1]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p1_dbgbus                     )
);

// Port 2
logic p2_side_clk_valid, p2_idle_egress, p2_rst_suppress;
  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p2_rst_suppress <= 1'b1;
    else
      p2_rst_suppress <= p2_credit_reinit & p2_rst_suppress;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if (~iosf_swf_side_rst_b)
      p2_fab_init_idle_exit <= '1;
    else
      if ( ~p2_rst_suppress & (p2_ism_idle & (~agent_idle[2] || ~p2_idle_egress) & ~p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '1;
      else if ( ~p2_rst_suppress & (p2_ism_idle & agent_idle[2] & p2_fab_init_idle_exit_ack ))
        p2_fab_init_idle_exit <= '0;

  always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)
    if ( ~iosf_swf_side_rst_b )
      p2_side_clk_valid <= 1'b0;
    else
      begin
        if ( p2_ism_idle & p2_side_clk_valid )
          p2_side_clk_valid <= '0;
        else if ( (p2_fab_init_idle_exit & p2_fab_init_idle_exit_ack) || ~p2_ism_idle )
          p2_side_clk_valid <= '1;
      end

//
// VISA tiered output assignments
//
logic [31:0] p2_dbgbus;

  always_comb
    begin
      visa_p2_tier1_iosf_swf_side_clk = { p2_dbgbus[31],
                            p2_dbgbus[27:24],
                            p2_dbgbus[21:19],
                            p2_dbgbus[15:12],
                            p2_dbgbus[7:4] };
      visa_p2_tier2_iosf_swf_side_clk = { p2_dbgbus[30:28],
                            p2_dbgbus[23:22],
                            p2_dbgbus[18:16],
                            p2_dbgbus[11:8],
                            p2_dbgbus[3:0] };
    end

sbcport #(
  .EXTMAXPLDBIT        (  7                            ),
  .INGMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .EGRMAXPLDBIT        ( INTMAXPLDBIT                  ),
  .CUP2PUT1CYC         (  0                            ),
  .NPQUEUEDEPTH        (  3                            ),
  .PCQUEUEDEPTH        (  3                            ),
  .SBCISMISAGENT       (  0                            ),
  .SYNCROUTER          (  1                            ),
  .LATCHQUEUES         (  0                            )
) sbcport2 (
  .side_clk            ( iosf_swf_side_clk             ),
  .gated_side_clk      ( gated_side_clk                ),
  .side_rst_b          ( iosf_swf_side_rst_b           ),
  .side_clk_valid      ( p2_side_clk_valid             ),
  .side_ism_in         ( swf_sbr2_side_ism_agent       ),
  .side_ism_out        ( sbr2_swf_side_ism_fabric      ),
  .int_pok             ( endpoint_pwrgd[2] ),
  .agent_idle          ( agent_idle[2]                 ),
  .port_idle           ( port_idle[2]                  ),
  .idle_egress         ( p2_idle_egress                ),
  .ism_idle            ( p2_ism_idle                   ),
  .credit_reinit       ( p2_credit_reinit              ),
  .cg_inprogress       ( p2_cg_inprogress              ),
  .tpccup              ( sbr2_swf_pccup                ),
  .tnpcup              ( sbr2_swf_npcup                ),
  .tpcput              ( swf_sbr2_pcput                ),
  .tnpput              ( swf_sbr2_npput                ),
  .teom                ( swf_sbr2_eom                  ),
  .tpayload            ( swf_sbr2_payload              ),
  .pctrdy              ( pctrdy[2]                     ),
  .pcirdy              ( pcirdy[2]                     ),
  .pcdata              ( pcdata[2]                     ),
  .pceom               ( pceom[2]                      ),
  .pcdstvld            ( p2_pcdstvld                   ),
  .nptrdy              ( nptrdy[2]                     ),
  .npirdy              ( npirdy[2]                     ),
  .npfence             ( p2_npfence                    ),
  .npdata              ( npdata[2]                     ),
  .npeom               ( npeom[2]                      ),
  .npdstvld            ( p2_npdstvld                   ),
  .mpccup              ( swf_sbr2_pccup                ),
  .mnpcup              ( swf_sbr2_npcup                ),
  .mpcput              ( sbr2_swf_pcput                ),
  .mnpput              ( sbr2_swf_npput                ),
  .meom                ( sbr2_swf_eom                  ),
  .mpayload            ( sbr2_swf_payload              ),
  .enpstall            (                               ),
  .epctrdy             ( epctrdy[2]                    ),
  .enptrdy             ( enptrdy[2]                    ),
  .epcirdy             ( epcirdy[2]                    ),
  .enpirdy             ( enpirdy[2]                    ),
  .data                ( data                          ),
  .eom                 ( eom                           ),
  .cfg_idlecnt         ( 8'h10                         ),
  .cfg_clkgaten        ( cfg_clkgaten                  ),
  .force_idle          ( force_idle                    ),
  .force_notidle       ( force_notidle                 ),
  .force_creditreq     ( force_creditreq               ),
  .dt_latchopen        ( fscan_latchopen               ),
  .dt_latchclosed_b    ( fscan_latchclosed_b           ),
  .dbgbus              ( p2_dbgbus                     )
);

//------------------------------------------------------------------------------
//
// SV Assertions
//
//------------------------------------------------------------------------------
 // synopsys translate_off

`ifndef INTEL_SVA_OFF
`ifndef IOSF_SB_ASSERT_OFF

    localparam SRCBIT = 8;

    logic [MAXPORT:0] pcwait4src;
    logic [MAXPORT:0] pcwait4eom;
    logic [MAXPORT:0] npwait4src;
    logic [MAXPORT:0] npwait4eom;
    logic [MAXPORT:0] eomvec;
    logic [MAXPORT:0] srcvec;
    logic [MAXPORT:0] mcastsrc;

    always_comb begin
      eomvec   = {MAXPORT+1{eom}};
      mcastsrc = {MAXPORT+1{ (data[SRCBIT+7:SRCBIT] == 8'hfe) |
                             sbr2_sbcportmap[data[SRCBIT+7:SRCBIT]][16] }};
      srcvec   = sbr2_sbcportmap[data[SRCBIT+7:SRCBIT]][MAXPORT:0];
      pcwait4src = ~pcwait4eom;
      npwait4src = ~npwait4eom;
    end

    always_ff @(posedge iosf_swf_side_clk or negedge iosf_swf_side_rst_b)

      if (~iosf_swf_side_rst_b) begin
        pcwait4eom <= '0;
        npwait4eom <= '0;
      end else begin
        pcwait4eom <= (pcwait4eom & ~(pcirdy & pctrdy & eomvec)) |
                      (pcwait4src & ~pcwait4eom & pcirdy & pctrdy & ~eomvec);
        npwait4eom <= (npwait4eom & ~(npirdy & nptrdy & eomvec)) |
                      (npwait4src & ~npwait4eom & npirdy & nptrdy & ~eomvec);
      end

    pc_source_port_id_check: //samassert
    assert property (@(posedge iosf_swf_side_clk) disable iff (iosf_swf_side_rst_b !== 1'b1)
        ~(pcwait4src & pcirdy & pctrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband pc message recieved on wrong ingress port", $time);

    np_source_port_id_check: //samassert
    assert property (@(posedge iosf_swf_side_clk) disable iff (iosf_swf_side_rst_b !== 1'b1)
        ~(npwait4src & npirdy & nptrdy & ~mcastsrc & ~srcvec) ) else
        $display("%0t: %m: ERROR: Sideband np message recieved on wrong ingress port", $time);

`endif
`endif

 // synopsys translate_on
  // lintra pop
endmodule

//------------------------------------------------------------------------------
//
// Fabric configuration file: ../tb/top_tb/lv2_sbn_cfg_8_pbg/lv2_sbn_cfg_8_pbg.csv
//
//------------------------------------------------------------------------------
/*
ClockReset, 0, bb_cclk, bb_rst_b, 0, , 4ns
ClockReset, 3, iosf_fust_side_clk, iosf_fust_side_rst_b, 0, , 2ns
ClockReset, 4, iosf_idf_side_clk, iosf_idf_side_rst_b, 0, cgc0, 2ns
ClockReset, 5, iosf_swf_side_clk, iosf_swf_side_rst_b, 0, cgc1, 2ns
ClockReset, 1, sosc_125_clk_core, sbi_rst_125_core_b, 0, , 4ns
ClockReset, 2, sosc_25_clk_core, sbi_rst_25_core_b, 0, , 40ns
SyncRouter, ccsb, ccsb,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 2, sbra, sbr1, , , , , , , , , , , , , , , 
RouterAgentPort, ccsb, 0
RouterAgentPort, ccsb, 1
Endpoint, dfxa,1, 1, 4, 0, 3, 3, 1, 2, 3, 3, 
Endpoint, fust,1, 1, 3, 0, 3, 3, 1, 0, 3, 3, 
Endpoint, idf,1, 1, 4, 0, 3, 3, 1, 5, 3, 3, 
Endpoint, io_dmi,0, 1, 2, 0, 1, 1, 1, 235, 3, 3, 
Endpoint, io_pxp,0, 1, 2, 0, 1, 1, 1, 236, 3, 3, 
Endpoint, io_st,0, 1, 2, 0, 1, 1, 1, 234, 3, 3, 
Endpoint, isa,1, 1, 4, 0, 3, 3, 1, 1, 3, 3, 
Endpoint, npsb,0, 1, 0, 0, 1, 1, 1, 239, 3, 3, 
Endpoint, rsp,1, 1, 4, 0, 3, 3, 1, 6, 3, 3, 
SyncRouter, sbr1, sbr1,1, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 4, 9, ccsb, fust, sbr2, isa, dfxa, scu0, scu1, idf, rsp, , , , , , , , 
RouterAgentPort, sbr1, 2
SyncRouter, sbr2, sbr2,2, 0, 0, 3, 4, 1, 0, 1, noa, dfxa, 5, 3, sbr1, xut, swf, , , , , , , , , , , , , , 
SyncRouter, sbra, sbra,0, 0, 0, 1, 4, 1, 0, 1, noa, dfxa, 2, 6, npsb, xpsb, ccsb, io_pxp, io_dmi, io_st, , , , , , , , , , , 
Endpoint, scu0,1, 1, 4, 0, 3, 3, 1, 3, 3, 3, 
Endpoint, scu1,3, 1, 4, 0, 3, 3, 1, 4, 3, 3, 
Endpoint, swf,2, 1, 5, 0, 3, 3, 1, 9, 3, 3, 
Endpoint, xpsb,0, 1, 1, 0, 1, 1, 1, 238, 3, 3, 
Endpoint, xut,2, 1, 5, 0, 3, 3, 1, 8, 3, 3, 
AsyncPort, ccsb, 0, 4, 4, 0, 
AsyncPort, sbr1, 1, 4, 4, 0, 
AsyncPort, sbr1, 2, 4, 4, 0, 
AsyncPort, sbra, 0, 2, 2, 0, 
AsyncPort, sbra, 1, 2, 2, 0, 
PowerWell, 0, 
PowerWell, 1, eva_present
PowerWell, 2, crp_sbr1_xu_en
PowerWell, 3, crp_sbr1_scu1_en
*/
//------------------------------------------------------------------------------
