module ctech_lib_firewall_and (a, en, o);
     input a, en;
     output o;
     d04swa00ld0b0 ctech_lib_dcszo (.a(a),.en(en),.o(o));
endmodule
