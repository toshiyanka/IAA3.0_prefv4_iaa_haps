//------------------------------------------------------------------------------
//  INTEL CONFIDENTIAL
//
//  Copyright 2016 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//
//  Collateral Description:
//  %header_collateral%
//
//  Source organization:
//  %header_organization%
//
//  Support Information:
//  %header_support%
//
//  Revision:
//  %header_tag%
//
//  Module <module name> :  < put your functional description here in plain text >
//
//------------------------------------------------------------------------------

//----------------------------------------------------------------------
// Intel Proprietary -- Copyright 2016 Intel -- All rights reserved
//----------------------------------------------------------------------
// NOTE: Log history is at end of file.
//----------------------------------------------------------------------
//
//    FILENAME    : DfxSecurePlugin_ClkGen.sv
//    CREATED BY  : Sudheer V Bandana
//    PROJECT     : DfxSecurePlugin
//    PURPOSE     : Clock Generation for the ENV
//    DESCRIPTION : This module is generic Clock Generator for
//                  the DfxSecurePlugin Environment.
//    PARAMETERS  :
//    TB_CLK_PERIOD
//                  This value is the peroid of the clock at which
//                  we want to run the environment.
//----------------------------------------------------------------------

module DfxSecurePlugin_ClkGen #(parameter TB_CLK_PERIOD = 10ns)(output logic DfxSecurePlugin_tb_clk);

    initial begin
        DfxSecurePlugin_tb_clk = 1'b0;
    end

    // 100 MHz always on TB Clock
    always begin
        #(TB_CLK_PERIOD/2) DfxSecurePlugin_tb_clk = ~(DfxSecurePlugin_tb_clk);
    end

endmodule

