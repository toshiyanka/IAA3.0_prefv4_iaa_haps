class hqm_ral_base_seq extends hqm_sla_pcie_base_seq;

   `ovm_sequence_utils(hqm_ral_base_seq, sla_sequencer)

   int                   registers_per_seg;
   int                   segment_number;

   sla_ral_access_path_t backdoor_id, ral_access_path;
   sla_ral_reg           reg_list[$];
   sla_ral_reg           reconfig_registers[$];
   sla_ral_reg           pf_cfg_reg_list[$];
   sla_ral_reg           list_sel_pipe_reg_list[$];
   sla_ral_reg           dir_pipe_reg_list[$];
   sla_ral_reg           qed_pipe_reg_list[$];
   sla_ral_reg           nalb_pipe_reg_list[$];
   sla_ral_reg           atm_pipe_reg_list[$];
   sla_ral_reg           aqed_pipe_reg_list[$];
   sla_ral_reg           reorder_pipe_reg_list[$];
   sla_ral_reg           credit_hist_pipe_reg_list[$];
   sla_ral_reg           config_master_reg_list[$];
   sla_ral_reg           system_csr_reg_list[$];
   sla_ral_reg           sif_csr_reg_list[$];
   sla_ral_reg           msix_mem_reg_list[$];
   static int            modified_reg[string];
   int                   exclude_reg[string];
   int                   reconfig_reg[string];
   int                   regs_read_via_backdoor;
   bit                   read_counter;
   bit [7:0]             legal_sai;
   string                log = "";
   string                reg_name = "";
   int                   register_wr_index;
   string                updated_register = "";
   int                   regs_written;
   logic [31:0]          mask = 32'hffff_ffff;
   sla_status_t          status;
   sla_ral_addr_t        reg_addr;
   logic [31:0]          comp_val; 

function new(string name = "hqm_ral_base_seq");

   super.new(name);

   pf_cfg_regs.get_regs(pf_cfg_reg_list);   
   list_sel_pipe_regs.get_regs(list_sel_pipe_reg_list);   
   dp_regs.get_regs(dir_pipe_reg_list);   
   qed_regs.get_regs(qed_pipe_reg_list);   
   nalb_regs.get_regs(nalb_pipe_reg_list);
   atm_pipe_regs.get_regs(atm_pipe_reg_list);
   aqed_pipe_regs.get_regs(aqed_pipe_reg_list);
   rop_regs.get_regs(reorder_pipe_reg_list);
   credit_hist_pipe_regs.get_regs(credit_hist_pipe_reg_list);
   master_regs.get_regs(config_master_reg_list);
   hqm_system_csr_regs.get_regs(system_csr_reg_list);
   hqm_sif_csr_regs.get_regs(sif_csr_reg_list);
   hqm_msix_mem_regs.get_regs(msix_mem_reg_list);

   reg_list = {pf_cfg_reg_list, list_sel_pipe_reg_list, dir_pipe_reg_list, qed_pipe_reg_list, nalb_pipe_reg_list, atm_pipe_reg_list, aqed_pipe_reg_list, reorder_pipe_reg_list, credit_hist_pipe_reg_list, config_master_reg_list, system_csr_reg_list, sif_csr_reg_list, msix_mem_reg_list};

   `ovm_info(get_full_name(),$psprintf("reg_list size is %d", reg_list.size()),OVM_LOW); 

endfunction   

//Contains the list of registers which have been modifed
//either in config sequence or in current sequence

virtual function modified_reg_list();

   modified_reg["DEVICE_COMMAND"         ] = 0;
   modified_reg["CSR_BAR_U"              ] = 1;
   modified_reg["CSR_BAR_L"              ] = 2; 
   modified_reg["FUNC_BAR_L"             ] = 3;
   modified_reg["FUNC_BAR_U"             ] = 4; 
   modified_reg["HQM_CSR_RAC_LO"         ] = 5;
   modified_reg["HQM_CSR_RAC_HI"         ] = 6;    
   modified_reg["HQM_CSR_WAC_LO"         ] = 7;    
   modified_reg["HQM_CSR_WAC_HI"         ] = 8;    
   modified_reg["HQM_CSR_CP_LO"          ] = 9;    
   modified_reg["HQM_CSR_CP_HI"          ] = 10;   
   modified_reg["PCIE_CAP_DEVICE_CONTROL"] = 11;
   modified_reg["PCIE_CAP_DEVICE_CONTROL_2"] = 12;
endfunction   
   
//Contains the list of registers which should be 
//excluded from being written. The list is generally set 
//of registers which trigger other HQM registers

virtual function excluded_reg_list();  

   exclude_reg["DEVICE_COMMAND"         ] = 0;
   exclude_reg["CSR_BAR_U"              ] = 1;
   exclude_reg["CSR_BAR_L"              ] = 2; 
   exclude_reg["FUNC_BAR_L"             ] = 3;
   exclude_reg["FUNC_BAR_U"             ] = 4; 
   exclude_reg["HQM_CSR_RAC_LO"         ] = 5;
   exclude_reg["HQM_CSR_RAC_HI"         ] = 6;    
   exclude_reg["HQM_CSR_WAC_LO"         ] = 7;    
   exclude_reg["HQM_CSR_WAC_HI"         ] = 8;    
   exclude_reg["HQM_CSR_CP_LO"          ] = 9;    
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[0]"]     = 10 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[1]"]     = 11 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[2]"]     = 12 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[3]"]     = 13 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[4]"]     = 14 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[5]"]     = 15 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[6]"]     = 16 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[7]"]     = 17 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[8]"]     = 18 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[9]"]     = 19 ;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[10]"]    = 20;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[11]"]    = 21;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[12]"]    = 22;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[13]"]    = 23;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[14]"]    = 24;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[15]"]    = 25;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[16]"]    = 26;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[17]"]    = 27;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[18]"]    = 28;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[19]"]    = 29;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[20]"]    = 30;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[21]"]    = 31;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[22]"]    = 32;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[23]"]    = 33;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[24]"]    = 34;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[25]"]    = 35;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[26]"]    = 36;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[27]"]    = 37;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[28]"]    = 38;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[29]"]    = 39;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[30]"]    = 40;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[31]"]    = 41;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[32]"]    = 42;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[33]"]    = 43;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[34]"]    = 44;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[35]"]    = 45;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[36]"]    = 46;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[37]"]    = 47;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[38]"]    = 48;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[39]"]    = 49;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[40]"]    = 50;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[41]"]    = 51;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[42]"]    = 52;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[43]"]    = 53;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[44]"]    = 54;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[45]"]    = 55;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[46]"]    = 56;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[47]"]    = 57;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[48]"]    = 58;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[49]"]    = 59;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[50]"]    = 60;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[51]"]    = 61;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[52]"]    = 62;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[53]"]    = 63;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[54]"]    = 64;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[55]"]    = 65;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[56]"]    = 66;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[57]"]    = 67;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[58]"]    = 68;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[59]"]    = 69;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[60]"]    = 70;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[61]"]    = 71;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[62]"]    = 72;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[63]"]    = 73;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[64]"]    = 74;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[65]"]    = 75;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[66]"]    = 76;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[67]"]    = 77;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[68]"]    = 78;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[69]"]    = 79;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[70]"]    = 70;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[71]"]    = 71;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[72]"]    = 72;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[73]"]    = 73;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[74]"]    = 74;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[75]"]    = 75;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[76]"]    = 76;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[77]"]    = 77;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[78]"]    = 78;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[79]"]    = 79;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[80]"]    = 80;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[81]"]    = 81;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[82]"]    = 82;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[83]"]    = 83;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[84]"]    = 84;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[85]"]    = 85;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[86]"]    = 86;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[87]"]    = 87;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[88]"]    = 88;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[89]"]    = 89;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[90]"]    = 90;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[91]"]    = 91;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[92]"]    = 92;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[93]"]    = 93;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[94]"]    = 94;
   exclude_reg["CFG_CQ_DIR_TOKEN_COUNT[95]"]    = 95;
   exclude_reg["HQM_CSR_CP_HI"          ] = 96;   
   exclude_reg["PCIE_CAP_DEVICE_CONTROL"] = 97;
   exclude_reg["CFG_PM_PMCSR_DISABLE   "] = 98;
   exclude_reg["PCIE_CAP_DEVICE_CONTROL_2"] = 99;
   exclude_reg["CFG_ERROR_INJECT"]            = 113;
   exclude_reg["CFG_DIAGNOSTIC_STATUS_1"]     = 114;
   exclude_reg["CFG_CONTROL_GENERAL"]         = 115;
   exclude_reg["CFG_CONTROL_GENERAL_01"]      = 117;
   exclude_reg["CFG_CONTROL_GENERAL_02"]      = 118;
   exclude_reg["CFG_LDB_SCHED_CONTROL"]      = 203;
   exclude_reg["ECC_CTL"]                    = 204;
   exclude_reg["AL_SIF_ALARM_AFULL_AGITATE_CONTROL"] = 205;
   exclude_reg["AL_HQM_ALARM_DB_AGITATE_CONTROL"] = 206;
   exclude_reg["AL_CWD_ALARM_DB_AGITATE_CONTROL"] = 207;
   ////HQMV30  exclude_reg["AL_MSI_MSIX_DB_AGITATE_CONTROL"] = 208;
   exclude_reg["EG_HCW_SCHED_DB_AGITATE_CONTROL"] = 208; //--reuse EG_HCW_SCHED_DB_AGITATE_CONTROL to replace AL_MSI_MSIX_DB_AGITATE_CONTROL
   exclude_reg["EG_HCW_SCHED_DB_AGITATE_CONTROL"] = 209;
   exclude_reg["IG_HCW_ENQ_W_DB_AGITATE_CONTROL"] = 210;
   exclude_reg["IG_HCW_ENQ_AFULL_AGITATE_CONTROL"] = 211;
   exclude_reg["WB_SCH_OUT_AFULL_AGITATE_CONTROL"] = 212;
   exclude_reg["PARITY_CTL"] = 213;
   exclude_reg["SIF_ALARM_FIFO_STATUS"] = 214;
   exclude_reg["HQM_ALARM_RX_FIFO_STATUS"] = 215;
   exclude_reg["CWDI_RX_FIFO_STATUS"] = 216;
   exclude_reg["CFG_RX_FIFO_STATUS"] = 217;
   exclude_reg["SCH_OUT_FIFO_STATUS"] = 218;
   exclude_reg["HCW_SCH_FIFO_STATUS"] = 219;
   exclude_reg["HCW_ENQ_FIFO_STATUS"] = 220;
   exclude_reg["PRIM_CDC_CTL"]        = 221;
   exclude_reg["INT_SIG_NUM_FIFO_STATUS"] = 222;
   exclude_reg["IOSFS_CGCTL"] = 223;
   exclude_reg["IOSFP_CGCTL"] = 224;
   exclude_reg["SIF_ALARM_ERR"] = 225;
   exclude_reg["RI_PARITY_ERR"] = 226;
   exclude_reg["TI_PARITY_ERR"] = 227;
   exclude_reg["SIF_PARITY_ERR"] = 228;
   exclude_reg["CFG_HQM_CDC_CONTROL"] = 229;
   exclude_reg["ALARM_ERR"] = 230;
   exclude_reg["EGRESS_LUT_ERR"] = 231;
   exclude_reg["ALARM_LUT_PERR"] = 232;
   exclude_reg["INGRESS_LUT_ERR"] = 233;
   exclude_reg["ALARM_MB_ECC_ERR"] = 234;
   exclude_reg["ALARM_SB_ECC_ERR"] = 235;
   exclude_reg["CFG_HQM_PGCB_CONTROL"] = 236; //FIXME
   exclude_reg["SIDE_CDC_CTL"]        = 237;
   exclude_reg["HQM_SIF_CNT_CTL"]= 238;
   exclude_reg["CFG_PATCH_CONTROL"]= 239;
   exclude_reg["PASID_CONTROL"]= 240;
   exclude_reg["AW_SMON_CONFIGURATION0[0]"]= 241;
   exclude_reg["AW_SMON_CONFIGURATION0[1]"]= 242;
   exclude_reg["PERF_SMON_CONFIGURATION0"]= 243;
   exclude_reg["MSIX_CAP_CONTROL"]= 244;
   exclude_reg["PM_CAP_CONTROL_STATUS"] = 245;
   exclude_reg["CFG_MASTER_CTL"] = 246;

endfunction

virtual function reconfig_excluded_reg_list();
   reconfig_reg["CFG_CONTROL_GENERAL_00"]        = 4;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[0]"]=   10;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[1]"]=   11;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[2]"]=   12;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[3]"]=   13;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[4]"]=   14;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[5]"]=   15;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[6]"]=   16;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[7]"]=   17;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[8]"]=   18;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[9]"]=   19;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[10]"]= 20;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[11]"]= 21;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[12]"]= 22;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[13]"]= 23;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[14]"]= 24;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[15]"]= 25;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[16]"]= 26;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[17]"]= 27;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[18]"]= 28;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[19]"]= 29;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[20]"]= 30;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[21]"]= 31;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[22]"]= 32;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[23]"]= 33;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[24]"]= 34;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[25]"]= 35;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[26]"]= 36;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[27]"]= 37;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[28]"]= 38;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[29]"]= 39;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[30]"]= 40;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[31]"]= 41;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[32]"]= 42;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[33]"]= 43;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[34]"]= 44;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[35]"]= 45;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[36]"]= 46;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[37]"]= 47;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[38]"]= 48;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[39]"]= 49;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[40]"]= 50;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[41]"]= 51;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[42]"]= 52;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[43]"]= 53;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[44]"]= 54;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[45]"]= 55;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[46]"]= 56;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[47]"]= 57;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[48]"]= 58;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[49]"]= 59;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[50]"]= 60;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[51]"]= 61;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[52]"]= 62;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[53]"]= 63;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[54]"]= 64;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[55]"]= 65;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[56]"]= 66;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[57]"]= 67;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[58]"]= 68;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[59]"]= 69;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[60]"]= 70;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[61]"]= 71;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[62]"]= 72;
   reconfig_reg["CFG_HIST_LIST_POP_PTR[63]"]= 73;
   reconfig_reg["CFG_DIR_CQ_DEPTH[0]"]= 74;
   reconfig_reg["CFG_DIR_CQ_DEPTH[1]"]= 75;
   reconfig_reg["CFG_DIR_CQ_DEPTH[2]"]= 76;
   reconfig_reg["CFG_DIR_CQ_DEPTH[3]"]= 77;
   reconfig_reg["CFG_DIR_CQ_DEPTH[4]"]= 78;
   reconfig_reg["CFG_DIR_CQ_DEPTH[5]"]= 79;
   reconfig_reg["CFG_DIR_CQ_DEPTH[6]"]= 80;
   reconfig_reg["CFG_DIR_CQ_DEPTH[7]"]= 81;
   reconfig_reg["CFG_DIR_CQ_DEPTH[8]"]= 82;
   reconfig_reg["CFG_DIR_CQ_DEPTH[9]"]= 83;
   reconfig_reg["CFG_DIR_CQ_DEPTH[10]"]= 84;
   reconfig_reg["CFG_DIR_CQ_DEPTH[11]"]= 85;
   reconfig_reg["CFG_DIR_CQ_DEPTH[12]"]= 86;
   reconfig_reg["CFG_DIR_CQ_DEPTH[13]"]= 88;
   reconfig_reg["CFG_DIR_CQ_DEPTH[14]"]= 89;
   reconfig_reg["CFG_DIR_CQ_DEPTH[15]"]= 90;
   reconfig_reg["CFG_DIR_CQ_DEPTH[16]"]= 91;
   reconfig_reg["CFG_DIR_CQ_DEPTH[17]"]= 92;
   reconfig_reg["CFG_DIR_CQ_DEPTH[18]"]= 93;
   reconfig_reg["CFG_DIR_CQ_DEPTH[19]"]= 94;
   reconfig_reg["CFG_DIR_CQ_DEPTH[20]"]= 95;
   reconfig_reg["CFG_DIR_CQ_DEPTH[21]"]= 96;
   reconfig_reg["CFG_DIR_CQ_DEPTH[22]"]= 97;
   reconfig_reg["CFG_DIR_CQ_DEPTH[23]"]= 98;
   reconfig_reg["CFG_DIR_CQ_DEPTH[24]"]= 99;
   reconfig_reg["CFG_DIR_CQ_DEPTH[25]"]= 100;
   reconfig_reg["CFG_DIR_CQ_DEPTH[26]"]= 101;
   reconfig_reg["CFG_DIR_CQ_DEPTH[27]"]= 102;
   reconfig_reg["CFG_DIR_CQ_DEPTH[28]"]= 103;
   reconfig_reg["CFG_DIR_CQ_DEPTH[29]"]= 104;
   reconfig_reg["CFG_DIR_CQ_DEPTH[30]"]= 105;
   reconfig_reg["CFG_DIR_CQ_DEPTH[31]"]= 106;
   reconfig_reg["CFG_DIR_CQ_DEPTH[32]"]= 107;
   reconfig_reg["CFG_DIR_CQ_DEPTH[33]"]= 108;
   reconfig_reg["CFG_DIR_CQ_DEPTH[34]"]= 109;
   reconfig_reg["CFG_DIR_CQ_DEPTH[35]"]= 200;
   reconfig_reg["CFG_DIR_CQ_DEPTH[36]"]= 201;
   reconfig_reg["CFG_DIR_CQ_DEPTH[37]"]= 202;
   reconfig_reg["CFG_DIR_CQ_DEPTH[38]"]= 203;
   reconfig_reg["CFG_DIR_CQ_DEPTH[39]"]= 204;
   reconfig_reg["CFG_DIR_CQ_DEPTH[40]"]= 205;
   reconfig_reg["CFG_DIR_CQ_DEPTH[41]"]= 206;
   reconfig_reg["CFG_DIR_CQ_DEPTH[42]"]= 207;
   reconfig_reg["CFG_DIR_CQ_DEPTH[43]"]= 208;
   reconfig_reg["CFG_DIR_CQ_DEPTH[44]"]= 209;
   reconfig_reg["CFG_DIR_CQ_DEPTH[45]"]= 210;
   reconfig_reg["CFG_DIR_CQ_DEPTH[46]"]= 211;
   reconfig_reg["CFG_DIR_CQ_DEPTH[47]"]= 212;
   reconfig_reg["CFG_DIR_CQ_DEPTH[48]"]= 213;
   reconfig_reg["CFG_DIR_CQ_DEPTH[49]"]= 214;
   reconfig_reg["CFG_DIR_CQ_DEPTH[50]"]= 215;
   reconfig_reg["CFG_DIR_CQ_DEPTH[51]"]= 216;
   reconfig_reg["CFG_DIR_CQ_DEPTH[52]"]= 217;
   reconfig_reg["CFG_DIR_CQ_DEPTH[53]"]= 218;
   reconfig_reg["CFG_DIR_CQ_DEPTH[54]"]= 219;
   reconfig_reg["CFG_DIR_CQ_DEPTH[55]"]= 220;
   reconfig_reg["CFG_DIR_CQ_DEPTH[56]"]= 221;
   reconfig_reg["CFG_DIR_CQ_DEPTH[57]"]= 222;
   reconfig_reg["CFG_DIR_CQ_DEPTH[58]"]= 223;
   reconfig_reg["CFG_DIR_CQ_DEPTH[59]"]= 224;
   reconfig_reg["CFG_DIR_CQ_DEPTH[60]"]= 225;
   reconfig_reg["CFG_DIR_CQ_DEPTH[61]"]= 226;
   reconfig_reg["CFG_DIR_CQ_DEPTH[62]"]= 227;
   reconfig_reg["CFG_DIR_CQ_DEPTH[63]"]= 228;
   reconfig_reg["CFG_DIR_CQ_DEPTH[64]"]= 229;
   reconfig_reg["CFG_DIR_CQ_DEPTH[65]"]= 230;
   reconfig_reg["CFG_DIR_CQ_DEPTH[66]"]= 231;
   reconfig_reg["CFG_DIR_CQ_DEPTH[67]"]= 232;
   reconfig_reg["CFG_DIR_CQ_DEPTH[68]"]= 233;
   reconfig_reg["CFG_DIR_CQ_DEPTH[69]"]= 234;
   reconfig_reg["CFG_DIR_CQ_DEPTH[70]"]= 235;
   reconfig_reg["CFG_DIR_CQ_DEPTH[71]"]= 236;
   reconfig_reg["CFG_DIR_CQ_DEPTH[72]"]= 237;
   reconfig_reg["CFG_DIR_CQ_DEPTH[73]"]= 238;
   reconfig_reg["CFG_DIR_CQ_DEPTH[74]"]= 239;
   reconfig_reg["CFG_DIR_CQ_DEPTH[75]"]= 240;
   reconfig_reg["CFG_DIR_CQ_DEPTH[76]"]= 241;
   reconfig_reg["CFG_DIR_CQ_DEPTH[77]"]= 242;
   reconfig_reg["CFG_DIR_CQ_DEPTH[78]"]= 243;
   reconfig_reg["CFG_DIR_CQ_DEPTH[79]"]= 244;
   reconfig_reg["CFG_DIR_CQ_DEPTH[80]"]= 245;
   reconfig_reg["CFG_DIR_CQ_DEPTH[81]"]= 246;
   reconfig_reg["CFG_DIR_CQ_DEPTH[82]"]= 247;
   reconfig_reg["CFG_DIR_CQ_DEPTH[83]"]= 248;
   reconfig_reg["CFG_DIR_CQ_DEPTH[84]"]= 249;
   reconfig_reg["CFG_DIR_CQ_DEPTH[85]"]= 250;
   reconfig_reg["CFG_DIR_CQ_DEPTH[86]"]= 251;
   reconfig_reg["CFG_DIR_CQ_DEPTH[87]"]= 252;
   reconfig_reg["CFG_DIR_CQ_DEPTH[88]"]= 253;
   reconfig_reg["CFG_DIR_CQ_DEPTH[89]"]= 254;
   reconfig_reg["CFG_DIR_CQ_DEPTH[90]"]= 255;
   reconfig_reg["CFG_DIR_CQ_DEPTH[91]"]= 256;
   reconfig_reg["CFG_DIR_CQ_DEPTH[92]"]= 257;
   reconfig_reg["CFG_DIR_CQ_DEPTH[93]"]= 258;
   reconfig_reg["CFG_DIR_CQ_DEPTH[94]"]= 259;
   reconfig_reg["CFG_DIR_CQ_DEPTH[95]"]= 260;
   reconfig_reg["CFG_LDB_CQ_DEPTH[0]"]= 261;
   reconfig_reg["CFG_LDB_CQ_DEPTH[1]"]= 262;
   reconfig_reg["CFG_LDB_CQ_DEPTH[2]"]= 263;
   reconfig_reg["CFG_LDB_CQ_DEPTH[3]"]= 264;
   reconfig_reg["CFG_LDB_CQ_DEPTH[4]"]= 265;
   reconfig_reg["CFG_LDB_CQ_DEPTH[5]"]= 266;
   reconfig_reg["CFG_LDB_CQ_DEPTH[6]"]= 267;
   reconfig_reg["CFG_LDB_CQ_DEPTH[7]"]= 268;
   reconfig_reg["CFG_LDB_CQ_DEPTH[8]"]= 269;
   reconfig_reg["CFG_LDB_CQ_DEPTH[9]"]= 270;
   reconfig_reg["CFG_LDB_CQ_DEPTH[10]"]= 271;
   reconfig_reg["CFG_LDB_CQ_DEPTH[11]"]= 272;
   reconfig_reg["CFG_LDB_CQ_DEPTH[12]"]= 273;
   reconfig_reg["CFG_LDB_CQ_DEPTH[13]"]= 274;
   reconfig_reg["CFG_LDB_CQ_DEPTH[14]"]= 275;
   reconfig_reg["CFG_LDB_CQ_DEPTH[15]"]= 276;
   reconfig_reg["CFG_LDB_CQ_DEPTH[16]"]= 277;
   reconfig_reg["CFG_LDB_CQ_DEPTH[17]"]= 278;
   reconfig_reg["CFG_LDB_CQ_DEPTH[18]"]= 279;
   reconfig_reg["CFG_LDB_CQ_DEPTH[19]"]= 280;
   reconfig_reg["CFG_LDB_CQ_DEPTH[20]"]= 281;
   reconfig_reg["CFG_LDB_CQ_DEPTH[21]"]= 282;
   reconfig_reg["CFG_LDB_CQ_DEPTH[22]"]= 283;
   reconfig_reg["CFG_LDB_CQ_DEPTH[23]"]= 284;
   reconfig_reg["CFG_LDB_CQ_DEPTH[24]"]= 285;
   reconfig_reg["CFG_LDB_CQ_DEPTH[25]"]= 286;
   reconfig_reg["CFG_LDB_CQ_DEPTH[26]"]= 287;
   reconfig_reg["CFG_LDB_CQ_DEPTH[27]"]= 288;
   reconfig_reg["CFG_LDB_CQ_DEPTH[28]"]= 289;
   reconfig_reg["CFG_LDB_CQ_DEPTH[29]"]= 290;
   reconfig_reg["CFG_LDB_CQ_DEPTH[30]"]= 291;
   reconfig_reg["CFG_LDB_CQ_DEPTH[31]"]= 292;
   reconfig_reg["CFG_LDB_CQ_DEPTH[32]"]= 293;
   reconfig_reg["CFG_LDB_CQ_DEPTH[33]"]= 294;
   reconfig_reg["CFG_LDB_CQ_DEPTH[34]"]= 295;
   reconfig_reg["CFG_LDB_CQ_DEPTH[35]"]= 296;
   reconfig_reg["CFG_LDB_CQ_DEPTH[36]"]= 297;
   reconfig_reg["CFG_LDB_CQ_DEPTH[37]"]= 298;
   reconfig_reg["CFG_LDB_CQ_DEPTH[38]"]= 299;
   reconfig_reg["CFG_LDB_CQ_DEPTH[39]"]= 300;
   reconfig_reg["CFG_LDB_CQ_DEPTH[40]"]= 301;
   reconfig_reg["CFG_LDB_CQ_DEPTH[41]"]= 302;
   reconfig_reg["CFG_LDB_CQ_DEPTH[42]"]= 303;
   reconfig_reg["CFG_LDB_CQ_DEPTH[43]"]= 304;
   reconfig_reg["CFG_LDB_CQ_DEPTH[44]"]= 305;
   reconfig_reg["CFG_LDB_CQ_DEPTH[45]"]= 306;
   reconfig_reg["CFG_LDB_CQ_DEPTH[46]"]= 307;
   reconfig_reg["CFG_LDB_CQ_DEPTH[47]"]= 308;
   reconfig_reg["CFG_LDB_CQ_DEPTH[48]"]= 309;
   reconfig_reg["CFG_LDB_CQ_DEPTH[49]"]= 340;
   reconfig_reg["CFG_LDB_CQ_DEPTH[50]"]= 341;
   reconfig_reg["CFG_LDB_CQ_DEPTH[51]"]= 342;
   reconfig_reg["CFG_LDB_CQ_DEPTH[52]"]= 343;
   reconfig_reg["CFG_LDB_CQ_DEPTH[53]"]= 344;
   reconfig_reg["CFG_LDB_CQ_DEPTH[54]"]= 345;
   reconfig_reg["CFG_LDB_CQ_DEPTH[55]"]= 346;
   reconfig_reg["CFG_LDB_CQ_DEPTH[56]"]= 347;
   reconfig_reg["CFG_LDB_CQ_DEPTH[57]"]= 348;
   reconfig_reg["CFG_LDB_CQ_DEPTH[58]"]= 349;
   reconfig_reg["CFG_LDB_CQ_DEPTH[59]"]= 350;
   reconfig_reg["CFG_LDB_CQ_DEPTH[60]"]= 351;
   reconfig_reg["CFG_LDB_CQ_DEPTH[61]"]= 352;
   reconfig_reg["CFG_LDB_CQ_DEPTH[62]"]= 353;
   reconfig_reg["CFG_LDB_CQ_DEPTH[63]"]= 354;
   reconfig_reg["LDB_PP_CQ_CFG[0]"]=   355 ;
   reconfig_reg["LDB_PP_CQ_CFG[1]"]=   356 ;
   reconfig_reg["LDB_PP_CQ_CFG[2]"]=   357 ;
   reconfig_reg["LDB_PP_CQ_CFG[3]"]=   358 ;
   reconfig_reg["LDB_PP_CQ_CFG[4]"]=   359 ;
   reconfig_reg["LDB_PP_CQ_CFG[5]"]=   360 ;
   reconfig_reg["LDB_PP_CQ_CFG[6]"]=   361 ;
   reconfig_reg["LDB_PP_CQ_CFG[7]"]=   362 ;
   reconfig_reg["LDB_PP_CQ_CFG[8]"]=   363 ;
   reconfig_reg["LDB_PP_CQ_CFG[9]"]=   364 ;
   reconfig_reg["LDB_PP_CQ_CFG[10]"]=  365  ;
   reconfig_reg["LDB_PP_CQ_CFG[11]"]=  366  ;
   reconfig_reg["LDB_PP_CQ_CFG[12]"]=  367  ;
   reconfig_reg["LDB_PP_CQ_CFG[13]"]=  368  ;
   reconfig_reg["LDB_PP_CQ_CFG[14]"]=  369  ;
   reconfig_reg["LDB_PP_CQ_CFG[15]"]=  370  ;
   reconfig_reg["LDB_PP_CQ_CFG[16]"]=  371  ;
   reconfig_reg["LDB_PP_CQ_CFG[17]"]=  372  ;
   reconfig_reg["LDB_PP_CQ_CFG[18]"]=  373  ;
   reconfig_reg["LDB_PP_CQ_CFG[19]"]=  374  ;
   reconfig_reg["LDB_PP_CQ_CFG[20]"]=  375  ;
   reconfig_reg["LDB_PP_CQ_CFG[21]"]=  376  ;
   reconfig_reg["LDB_PP_CQ_CFG[22]"]=  377  ;
   reconfig_reg["LDB_PP_CQ_CFG[23]"]=  378  ;
   reconfig_reg["LDB_PP_CQ_CFG[24]"]=  379  ;
   reconfig_reg["LDB_PP_CQ_CFG[25]"]=  380  ;
   reconfig_reg["LDB_PP_CQ_CFG[26]"]=  381  ;
   reconfig_reg["LDB_PP_CQ_CFG[27]"]=  382  ;
   reconfig_reg["LDB_PP_CQ_CFG[28]"]=  383  ;
   reconfig_reg["LDB_PP_CQ_CFG[29]"]=  384  ;
   reconfig_reg["LDB_PP_CQ_CFG[30]"]=  385  ;
   reconfig_reg["LDB_PP_CQ_CFG[31]"]=  386  ;
   reconfig_reg["LDB_PP_CQ_CFG[32]"]=  387 ;
   reconfig_reg["LDB_PP_CQ_CFG[33]"]=  388  ;
   reconfig_reg["LDB_PP_CQ_CFG[34]"]=  389  ;
   reconfig_reg["LDB_PP_CQ_CFG[35]"]=  390  ;
   reconfig_reg["LDB_PP_CQ_CFG[36]"]=  391  ;
   reconfig_reg["LDB_PP_CQ_CFG[37]"]=  392  ;
   reconfig_reg["LDB_PP_CQ_CFG[38]"]=  393  ;
   reconfig_reg["LDB_PP_CQ_CFG[39]"]=  394  ;
   reconfig_reg["LDB_PP_CQ_CFG[40]"]=  395  ;
   reconfig_reg["LDB_PP_CQ_CFG[41]"]=  396  ;
   reconfig_reg["LDB_PP_CQ_CFG[42]"]=  397  ;
   reconfig_reg["LDB_PP_CQ_CFG[43]"]=  398  ;
   reconfig_reg["LDB_PP_CQ_CFG[44]"]=  399  ;
   reconfig_reg["LDB_PP_CQ_CFG[45]"]=  400  ;
   reconfig_reg["LDB_PP_CQ_CFG[46]"]=  401  ;
   reconfig_reg["LDB_PP_CQ_CFG[47]"]=  402  ;
   reconfig_reg["LDB_PP_CQ_CFG[48]"]=  403  ;
   reconfig_reg["LDB_PP_CQ_CFG[49]"]=  404  ;
   reconfig_reg["LDB_PP_CQ_CFG[50]"]=  405  ;
   reconfig_reg["LDB_PP_CQ_CFG[51]"]=  406  ;
   reconfig_reg["LDB_PP_CQ_CFG[52]"]=  407  ;
   reconfig_reg["LDB_PP_CQ_CFG[53]"]=  408  ;
   reconfig_reg["LDB_PP_CQ_CFG[54]"]=  409  ;
   reconfig_reg["LDB_PP_CQ_CFG[55]"]=  410  ;
   reconfig_reg["LDB_PP_CQ_CFG[56]"]=  411  ;
   reconfig_reg["LDB_PP_CQ_CFG[57]"]=  412  ;
   reconfig_reg["LDB_PP_CQ_CFG[58]"]=  413  ;
   reconfig_reg["LDB_PP_CQ_CFG[59]"]=  414  ;
   reconfig_reg["LDB_PP_CQ_CFG[60]"]=  415  ;
   reconfig_reg["LDB_PP_CQ_CFG[61]"]=  416  ;
   reconfig_reg["LDB_PP_CQ_CFG[62]"]=  417  ;
   reconfig_reg["LDB_PP_CQ_CFG[63]"]=  418  ;

   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[9]"]=   419;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[10]"]= 420;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[11]"]= 421;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[12]"]= 422;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[13]"]= 423;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[14]"]= 424;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[15]"]= 425;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[16]"]= 426;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[17]"]= 427;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[18]"]= 428;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[19]"]= 429;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[20]"]= 430;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[21]"]= 431;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[22]"]= 432;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[23]"]= 433;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[24]"]= 434;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[25]"]= 435;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[26]"]= 436;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[27]"]= 437;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[28]"]= 438;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[29]"]= 439;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[30]"]= 440;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[31]"]= 441;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[32]"]= 442;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[33]"]= 443;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[34]"]= 444;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[35]"]= 445;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[36]"]= 446;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[37]"]= 447;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[38]"]= 448;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[39]"]= 449;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[40]"]= 450;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[41]"]= 451;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[42]"]= 452;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[43]"]= 453;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[44]"]= 454;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[45]"]= 455;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[46]"]= 456;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[47]"]= 457;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[48]"]= 458;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[49]"]= 459;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[50]"]= 460;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[51]"]= 461;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[52]"]= 462;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[53]"]= 463;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[54]"]= 464;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[55]"]= 465;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[56]"]= 466;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[57]"]= 467;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[58]"]= 468;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[59]"]= 469;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[60]"]= 470;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[61]"]= 471;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[62]"]= 472;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[63]"]= 473;  
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[0]"]=  474;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[1]"]=  475;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[2]"]=  476;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[3]"]=  477;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[4]"]=  478;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[5]"]=  478;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[6]"]=  479;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[7]"]=  480;
   reconfig_reg["CFG_HIST_LIST_PUSH_PTR[8]"]=  481;

endfunction


endclass
