### Tool : gds2def
### Version 14.1     Linux64
### Vendor : Apache Design, Inc. A Subsidiary of ANSYS, Inc. 
### Date : Jun 19 2014 02:20:56 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO c73p4hdxrom_iopwrcell
 CLASS CORE ;
 ORIGIN -0.224 -0.042 ;
 SIZE 2.912 BY 1.197 ;
 PIN vccd_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 2.912 0.042 2.968 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.744 0.042 2.8 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.408 0.042 2.464 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.576 0.042 2.632 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.24 0.042 2.296 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.072 0.042 2.128 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.736 0.042 1.792 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.904 0.042 1.96 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.08 0.042 3.136 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.4 0.042 1.456 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.98 0.21 1.036 1.223 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.812 0.209 0.868 1.222 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.224 0.042 0.28 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.568 0.042 1.624 1.236 ;
  END
 END vccd_1p0
 PIN vccdgt_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 2.996 0.042 3.052 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.66 0.042 2.716 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.652 0.9 1.708 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.988 0.042 2.044 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.324 0.042 2.38 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.652 0.042 1.708 0.858 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.316 0.042 1.372 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.484 0.042 1.54 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.064 0.042 1.12 1.236 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.728 0.042 0.784 1.236 ;
  END
 END vccdgt_1p0
 PIN vss
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER m1 ;
   RECT 1.148 0.474 1.204 1.16 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.392 0.609 0.448 0.912 ;
  END
 END vss
 PIN pwren_in
  DIRECTION INPUT ;
  USE SIGNAL ;
 END pwren_in
END c73p4hdxrom_iopwrcell

MACRO c73p4hdxrom_x4pwrcell
 CLASS CORE ;
 ORIGIN -0.001 -1.097 ;
 SIZE 0.728 BY 0.898 ;
 PIN vccd_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 0.673 1.582 0.729 1.65 ;
   LAYER m1 ;
   RECT 0.673 1.097 0.729 1.582 ;
   LAYER m1 ;
   RECT 0.673 1.582 0.729 1.767 ;
   LAYER m1 ;
   RECT 0.673 1.65 0.729 1.767 ;
   LAYER m1 ;
   RECT 0.673 1.097 0.729 1.582 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.169 1.778 0.225 1.848 ;
   LAYER m1 ;
   RECT 0.169 1.133 0.225 1.872 ;
   LAYER m1 ;
   RECT 0.169 1.31 0.225 1.378 ;
   LAYER m1 ;
   RECT 0.169 1.133 0.225 1.872 ;
   LAYER m1 ;
   RECT 0.169 1.442 0.225 1.512 ;
   LAYER m1 ;
   RECT 0.169 1.65 0.225 1.71 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.001 1.442 0.057 1.512 ;
   LAYER m1 ;
   RECT 0.001 1.133 0.057 1.767 ;
   LAYER m1 ;
   RECT 0.001 1.582 0.057 1.65 ;
   LAYER m1 ;
   RECT 0.001 1.133 0.057 1.767 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.337 1.31 0.393 1.378 ;
   LAYER m1 ;
   RECT 0.337 1.133 0.393 1.872 ;
   LAYER m1 ;
   RECT 0.337 1.582 0.393 1.65 ;
   LAYER m1 ;
   RECT 0.337 1.133 0.393 1.872 ;
   LAYER m1 ;
   RECT 0.337 1.442 0.393 1.512 ;
   LAYER m1 ;
   RECT 0.337 1.778 0.393 1.848 ;
  END
 END vccd_1p0
 PIN vccdgt_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 0.589 1.71 0.645 1.778 ;
   LAYER m1 ;
   RECT 0.589 1.133 0.645 1.995 ;
   LAYER m1 ;
   RECT 0.589 1.848 0.645 1.918 ;
   LAYER m1 ;
   RECT 0.589 1.106 0.645 1.995 ;
   LAYER m1 ;
   RECT 0.589 1.392 0.645 1.428 ;
   LAYER m1 ;
   RECT 0.589 1.512 0.645 1.582 ;
   LAYER m1 ;
   RECT 0.589 1.106 0.645 1.176 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.421 1.71 0.477 1.778 ;
   LAYER m1 ;
   RECT 0.421 1.133 0.477 1.995 ;
   LAYER m1 ;
   RECT 0.421 1.392 0.477 1.428 ;
   LAYER m1 ;
   RECT 0.421 1.133 0.477 1.995 ;
   LAYER m1 ;
   RECT 0.421 1.512 0.477 1.582 ;
   LAYER m1 ;
   RECT 0.421 1.26 0.477 1.296 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.253 1.848 0.309 1.918 ;
   LAYER m1 ;
   RECT 0.253 1.133 0.309 1.995 ;
   LAYER m1 ;
   RECT 0.253 1.106 0.309 1.176 ;
   LAYER m1 ;
   RECT 0.253 1.106 0.309 1.995 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.085 1.71 0.141 1.778 ;
   LAYER m1 ;
   RECT 0.085 1.133 0.141 1.995 ;
   LAYER m1 ;
   RECT 0.085 1.26 0.141 1.296 ;
   LAYER m1 ;
   RECT 0.085 1.133 0.141 1.995 ;
  END
 END vccdgt_1p0
 PIN pwren_in
  DIRECTION INPUT ;
  USE SIGNAL ;
 END pwren_in
END c73p4hdxrom_x4pwrcell

MACRO c73p4hdxrom_wldrvgappwrcell
 CLASS CORE ;
 ORIGIN -0.14 -0.034 ;
 SIZE 5.348 BY 1.958 ;
 PIN vccd_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 5.432 1.778 5.488 1.848 ;
   LAYER m1 ;
   RECT 5.432 0.034 5.488 1.932 ;
   LAYER m1 ;
   RECT 5.432 1.442 5.488 1.512 ;
   LAYER m1 ;
   RECT 5.432 0.034 5.488 1.932 ;
   LAYER m1 ;
   RECT 5.432 1.31 5.488 1.378 ;
   LAYER m1 ;
   RECT 5.432 1.038 5.488 1.106 ;
   LAYER m1 ;
   RECT 5.432 1.176 5.488 1.246 ;
   LAYER m1 ;
   RECT 5.432 0.048 5.488 0.084 ;
   LAYER m1 ;
   RECT 5.432 0.91 5.488 0.978 ;
   LAYER m1 ;
   RECT 5.432 0.306 5.488 0.366 ;
   LAYER m1 ;
   RECT 5.432 0.588 5.488 0.624 ;
   LAYER m1 ;
   RECT 5.432 0.434 5.488 0.504 ;
   LAYER m1 ;
   RECT 5.432 0.77 5.488 0.84 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.76 1.778 4.816 1.848 ;
   LAYER m1 ;
   RECT 4.76 0.034 4.816 1.932 ;
   LAYER m1 ;
   RECT 4.76 1.442 4.816 1.512 ;
   LAYER m1 ;
   RECT 4.76 0.034 4.816 1.932 ;
   LAYER m1 ;
   RECT 4.76 1.038 4.816 1.106 ;
   LAYER m1 ;
   RECT 4.76 1.176 4.816 1.246 ;
   LAYER m1 ;
   RECT 4.76 1.31 4.816 1.378 ;
   LAYER m1 ;
   RECT 4.76 1.65 4.816 1.71 ;
   LAYER m1 ;
   RECT 4.76 0.91 4.816 0.978 ;
   LAYER m1 ;
   RECT 4.76 0.588 4.816 0.624 ;
   LAYER m1 ;
   RECT 4.76 0.434 4.816 0.504 ;
   LAYER m1 ;
   RECT 4.76 0.77 4.816 0.84 ;
   LAYER m1 ;
   RECT 4.76 0.048 4.816 0.084 ;
   LAYER m1 ;
   RECT 4.76 0.306 4.816 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.928 1.778 4.984 1.848 ;
   LAYER m1 ;
   RECT 4.928 0.034 4.984 1.932 ;
   LAYER m1 ;
   RECT 4.928 1.038 4.984 1.106 ;
   LAYER m1 ;
   RECT 4.928 0.034 4.984 1.932 ;
   LAYER m1 ;
   RECT 4.928 1.176 4.984 1.246 ;
   LAYER m1 ;
   RECT 4.928 1.31 4.984 1.378 ;
   LAYER m1 ;
   RECT 4.928 1.442 4.984 1.512 ;
   LAYER m1 ;
   RECT 4.928 1.65 4.984 1.71 ;
   LAYER m1 ;
   RECT 4.928 0.91 4.984 0.978 ;
   LAYER m1 ;
   RECT 4.928 0.72 4.984 0.756 ;
   LAYER m1 ;
   RECT 4.928 0.434 4.984 0.504 ;
   LAYER m1 ;
   RECT 4.928 0.588 4.984 0.624 ;
   LAYER m1 ;
   RECT 4.928 0.048 4.984 0.084 ;
   LAYER m1 ;
   RECT 4.928 0.306 4.984 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 5.096 1.778 5.152 1.848 ;
   LAYER m1 ;
   RECT 5.096 0.034 5.152 1.932 ;
   LAYER m1 ;
   RECT 5.096 1.038 5.152 1.106 ;
   LAYER m1 ;
   RECT 5.096 0.034 5.152 1.932 ;
   LAYER m1 ;
   RECT 5.096 1.176 5.152 1.246 ;
   LAYER m1 ;
   RECT 5.096 1.31 5.152 1.378 ;
   LAYER m1 ;
   RECT 5.096 1.442 5.152 1.512 ;
   LAYER m1 ;
   RECT 5.096 1.65 5.152 1.71 ;
   LAYER m1 ;
   RECT 5.096 0.91 5.152 0.978 ;
   LAYER m1 ;
   RECT 5.096 0.72 5.152 0.756 ;
   LAYER m1 ;
   RECT 5.096 0.588 5.152 0.624 ;
   LAYER m1 ;
   RECT 5.096 0.434 5.152 0.504 ;
   LAYER m1 ;
   RECT 5.096 0.048 5.152 0.084 ;
   LAYER m1 ;
   RECT 5.096 0.306 5.152 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 5.264 1.778 5.32 1.848 ;
   LAYER m1 ;
   RECT 5.264 0.034 5.32 1.932 ;
   LAYER m1 ;
   RECT 5.264 1.038 5.32 1.106 ;
   LAYER m1 ;
   RECT 5.264 0.034 5.32 1.932 ;
   LAYER m1 ;
   RECT 5.264 1.176 5.32 1.246 ;
   LAYER m1 ;
   RECT 5.264 1.31 5.32 1.378 ;
   LAYER m1 ;
   RECT 5.264 1.442 5.32 1.512 ;
   LAYER m1 ;
   RECT 5.264 1.65 5.32 1.71 ;
   LAYER m1 ;
   RECT 5.264 0.91 5.32 0.978 ;
   LAYER m1 ;
   RECT 5.264 0.434 5.32 0.504 ;
   LAYER m1 ;
   RECT 5.264 0.77 5.32 0.84 ;
   LAYER m1 ;
   RECT 5.264 0.588 5.32 0.624 ;
   LAYER m1 ;
   RECT 5.264 0.048 5.32 0.084 ;
   LAYER m1 ;
   RECT 5.264 0.306 5.32 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.248 0.034 3.304 1.991 ;
   LAYER m1 ;
   RECT 3.248 1.038 3.304 1.106 ;
   LAYER m1 ;
   RECT 3.248 0.034 3.304 1.991 ;
   LAYER m1 ;
   RECT 3.248 1.65 3.304 1.71 ;
   LAYER m1 ;
   RECT 3.248 0.91 3.304 0.978 ;
   LAYER m1 ;
   RECT 3.248 0.434 3.304 0.504 ;
   LAYER m1 ;
   RECT 3.248 0.77 3.304 0.84 ;
   LAYER m1 ;
   RECT 3.248 0.588 3.304 0.624 ;
   LAYER m1 ;
   RECT 3.248 0.048 3.304 0.084 ;
   LAYER m1 ;
   RECT 3.248 0.306 3.304 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.08 1.932 3.136 1.968 ;
   LAYER m1 ;
   RECT 3.08 0.034 3.136 1.991 ;
   LAYER m1 ;
   RECT 3.08 1.038 3.136 1.106 ;
   LAYER m1 ;
   RECT 3.08 0.034 3.136 1.991 ;
   LAYER m1 ;
   RECT 3.08 1.65 3.136 1.71 ;
   LAYER m1 ;
   RECT 3.08 0.91 3.136 0.978 ;
   LAYER m1 ;
   RECT 3.08 0.72 3.136 0.756 ;
   LAYER m1 ;
   RECT 3.08 0.434 3.136 0.504 ;
   LAYER m1 ;
   RECT 3.08 0.588 3.136 0.624 ;
   LAYER m1 ;
   RECT 3.08 0.048 3.136 0.084 ;
   LAYER m1 ;
   RECT 3.08 0.306 3.136 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.744 0.034 2.8 1.991 ;
   LAYER m1 ;
   RECT 2.744 1.038 2.8 1.106 ;
   LAYER m1 ;
   RECT 2.744 0.034 2.8 1.991 ;
   LAYER m1 ;
   RECT 2.744 1.65 2.8 1.71 ;
   LAYER m1 ;
   RECT 2.744 0.72 2.8 0.756 ;
   LAYER m1 ;
   RECT 2.744 0.91 2.8 0.978 ;
   LAYER m1 ;
   RECT 2.744 0.434 2.8 0.504 ;
   LAYER m1 ;
   RECT 2.744 0.588 2.8 0.624 ;
   LAYER m1 ;
   RECT 2.744 0.048 2.8 0.084 ;
   LAYER m1 ;
   RECT 2.744 0.306 2.8 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.576 1.932 2.632 1.968 ;
   LAYER m1 ;
   RECT 2.576 0.034 2.632 1.991 ;
   LAYER m1 ;
   RECT 2.576 1.038 2.632 1.106 ;
   LAYER m1 ;
   RECT 2.576 0.034 2.632 1.991 ;
   LAYER m1 ;
   RECT 2.576 1.65 2.632 1.71 ;
   LAYER m1 ;
   RECT 2.576 0.91 2.632 0.978 ;
   LAYER m1 ;
   RECT 2.576 0.434 2.632 0.504 ;
   LAYER m1 ;
   RECT 2.576 0.77 2.632 0.84 ;
   LAYER m1 ;
   RECT 2.576 0.588 2.632 0.624 ;
   LAYER m1 ;
   RECT 2.576 0.048 2.632 0.084 ;
   LAYER m1 ;
   RECT 2.576 0.306 2.632 0.366 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.408 0.034 2.464 1.991 ;
   LAYER m1 ;
   RECT 2.408 1.31 2.464 1.378 ;
   LAYER m1 ;
   RECT 2.408 0.034 2.464 1.991 ;
   LAYER m1 ;
   RECT 2.408 1.038 2.464 1.106 ;
   LAYER m1 ;
   RECT 2.408 1.442 2.464 1.512 ;
   LAYER m1 ;
   RECT 2.408 1.65 2.464 1.71 ;
   LAYER m1 ;
   RECT 2.408 0.91 2.464 0.978 ;
   LAYER m1 ;
   RECT 2.408 0.72 2.464 0.756 ;
   LAYER m1 ;
   RECT 2.408 0.588 2.464 0.624 ;
   LAYER m1 ;
   RECT 2.408 0.434 2.464 0.504 ;
   LAYER m1 ;
   RECT 2.408 0.048 2.464 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.24 0.034 2.296 1.991 ;
   LAYER m1 ;
   RECT 2.24 1.65 2.296 1.71 ;
   LAYER m1 ;
   RECT 2.24 0.034 2.296 1.991 ;
   LAYER m1 ;
   RECT 2.24 0.91 2.296 0.978 ;
   LAYER m1 ;
   RECT 2.24 0.77 2.296 0.84 ;
   LAYER m1 ;
   RECT 2.24 0.588 2.296 0.624 ;
   LAYER m1 ;
   RECT 2.24 0.048 2.296 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.568 1.932 1.624 1.968 ;
   LAYER m1 ;
   RECT 1.568 0.034 1.624 1.991 ;
   LAYER m1 ;
   RECT 1.568 1.038 1.624 1.106 ;
   LAYER m1 ;
   RECT 1.568 0.034 1.624 1.991 ;
   LAYER m1 ;
   RECT 1.568 1.442 1.624 1.512 ;
   LAYER m1 ;
   RECT 1.568 1.65 1.624 1.71 ;
   LAYER m1 ;
   RECT 1.568 0.91 1.624 0.978 ;
   LAYER m1 ;
   RECT 1.568 0.72 1.624 0.756 ;
   LAYER m1 ;
   RECT 1.568 0.048 1.624 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.4 1.932 1.456 1.968 ;
   LAYER m1 ;
   RECT 1.4 0.034 1.456 1.991 ;
   LAYER m1 ;
   RECT 1.4 1.778 1.456 1.848 ;
   LAYER m1 ;
   RECT 1.4 0.034 1.456 1.991 ;
   LAYER m1 ;
   RECT 1.4 1.038 1.456 1.106 ;
   LAYER m1 ;
   RECT 1.4 1.442 1.456 1.512 ;
   LAYER m1 ;
   RECT 1.4 1.65 1.456 1.71 ;
   LAYER m1 ;
   RECT 1.4 0.91 1.456 0.978 ;
   LAYER m1 ;
   RECT 1.4 0.72 1.456 0.756 ;
   LAYER m1 ;
   RECT 1.4 0.048 1.456 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.736 0.034 1.792 1.991 ;
   LAYER m1 ;
   RECT 1.736 1.038 1.792 1.106 ;
   LAYER m1 ;
   RECT 1.736 0.034 1.792 1.991 ;
   LAYER m1 ;
   RECT 1.736 1.442 1.792 1.512 ;
   LAYER m1 ;
   RECT 1.736 1.65 1.792 1.71 ;
   LAYER m1 ;
   RECT 1.736 0.91 1.792 0.978 ;
   LAYER m1 ;
   RECT 1.736 0.72 1.792 0.756 ;
   LAYER m1 ;
   RECT 1.736 0.048 1.792 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.904 0.034 1.96 1.991 ;
   LAYER m1 ;
   RECT 1.904 1.038 1.96 1.106 ;
   LAYER m1 ;
   RECT 1.904 0.034 1.96 1.991 ;
   LAYER m1 ;
   RECT 1.904 1.65 1.96 1.71 ;
   LAYER m1 ;
   RECT 1.904 0.91 1.96 0.978 ;
   LAYER m1 ;
   RECT 1.904 0.72 1.96 0.756 ;
   LAYER m1 ;
   RECT 1.904 0.048 1.96 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.072 0.034 2.128 1.991 ;
   LAYER m1 ;
   RECT 2.072 1.932 2.128 1.968 ;
   LAYER m1 ;
   RECT 2.072 0.034 2.128 1.991 ;
   LAYER m1 ;
   RECT 2.072 1.65 2.128 1.71 ;
   LAYER m1 ;
   RECT 2.072 0.91 2.128 0.978 ;
   LAYER m1 ;
   RECT 2.072 0.72 2.128 0.756 ;
   LAYER m1 ;
   RECT 2.072 0.048 2.128 0.084 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.896 1.442 0.952 1.512 ;
   LAYER m1 ;
   RECT 0.896 0.085 0.952 1.528 ;
   LAYER m1 ;
   RECT 0.896 0.91 0.952 0.978 ;
   LAYER m1 ;
   RECT 0.896 0.91 0.952 0.978 ;
   LAYER m1 ;
   RECT 0.896 0.085 0.952 1.528 ;
   LAYER m1 ;
   RECT 0.896 0.306 0.952 0.366 ;
   LAYER m1 ;
   RECT 0.896 0.306 0.952 0.366 ;
   LAYER m1 ;
   RECT 0.896 1.442 0.952 1.512 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.392 1.778 0.448 1.848 ;
   LAYER m1 ;
   RECT 0.392 0.074 0.448 1.932 ;
   LAYER m1 ;
   RECT 0.392 1.442 0.448 1.512 ;
   LAYER m1 ;
   RECT 0.392 0.074 0.448 1.932 ;
   LAYER m1 ;
   RECT 0.392 1.31 0.448 1.378 ;
   LAYER m1 ;
   RECT 0.392 1.038 0.448 1.106 ;
   LAYER m1 ;
   RECT 0.392 0.72 0.448 0.756 ;
   LAYER m1 ;
   RECT 0.392 0.306 0.448 0.366 ;
   LAYER m1 ;
   RECT 0.392 0.91 0.448 0.978 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.224 1.778 0.28 1.848 ;
   LAYER m1 ;
   RECT 0.224 0.074 0.28 1.932 ;
   LAYER m1 ;
   RECT 0.224 1.31 0.28 1.378 ;
   LAYER m1 ;
   RECT 0.224 0.074 0.28 1.932 ;
   LAYER m1 ;
   RECT 0.224 1.65 0.28 1.71 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.912 0.034 2.968 1.991 ;
   LAYER m1 ;
   RECT 2.912 0.91 2.968 0.978 ;
   LAYER m1 ;
   RECT 2.912 0.034 2.968 1.991 ;
   LAYER m1 ;
   RECT 2.912 0.048 2.968 0.084 ;
   LAYER m1 ;
   RECT 2.912 0.306 2.968 0.366 ;
   LAYER m1 ;
   RECT 2.912 0.588 2.968 0.624 ;
   LAYER m1 ;
   RECT 2.912 0.72 2.968 0.756 ;
   LAYER m1 ;
   RECT 2.912 0.434 2.968 0.504 ;
   LAYER m1 ;
   RECT 2.912 1.038 2.968 1.106 ;
   LAYER m1 ;
   RECT 2.912 1.65 2.968 1.71 ;
   LAYER m1 ;
   RECT 2.912 1.778 2.968 1.848 ;
   LAYER m1 ;
   RECT 2.912 1.932 2.968 1.968 ;
  END
 END vccd_1p0
 PIN vccdgt_1p0
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER m1 ;
   RECT 4.844 1.848 4.9 1.918 ;
   LAYER m1 ;
   RECT 4.844 0.034 4.9 1.932 ;
   LAYER m1 ;
   RECT 4.844 1.512 4.9 1.582 ;
   LAYER m1 ;
   RECT 4.844 0.034 4.9 1.932 ;
   LAYER m1 ;
   RECT 4.844 0.238 4.9 0.306 ;
   LAYER m1 ;
   RECT 4.844 0.098 4.9 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 5.012 1.848 5.068 1.918 ;
   LAYER m1 ;
   RECT 5.012 0.034 5.068 1.932 ;
   LAYER m1 ;
   RECT 5.012 1.512 5.068 1.582 ;
   LAYER m1 ;
   RECT 5.012 0.034 5.068 1.932 ;
   LAYER m1 ;
   RECT 5.012 0.84 5.068 0.91 ;
   LAYER m1 ;
   RECT 5.012 0.238 5.068 0.306 ;
   LAYER m1 ;
   RECT 5.012 0.098 5.068 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 5.18 1.848 5.236 1.918 ;
   LAYER m1 ;
   RECT 5.18 0.034 5.236 1.932 ;
   LAYER m1 ;
   RECT 5.18 1.512 5.236 1.582 ;
   LAYER m1 ;
   RECT 5.18 0.034 5.236 1.932 ;
   LAYER m1 ;
   RECT 5.18 0.238 5.236 0.306 ;
   LAYER m1 ;
   RECT 5.18 0.098 5.236 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.676 1.512 4.732 1.582 ;
   LAYER m1 ;
   RECT 4.676 0.034 4.732 1.813 ;
   LAYER m1 ;
   RECT 4.676 0.638 4.732 0.706 ;
   LAYER m1 ;
   RECT 4.676 0.034 4.732 1.813 ;
   LAYER m1 ;
   RECT 4.676 0.098 4.732 0.168 ;
   LAYER m1 ;
   RECT 4.676 0.238 4.732 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 5.348 1.512 5.404 1.582 ;
   LAYER m1 ;
   RECT 5.348 0.034 5.404 1.932 ;
   LAYER m1 ;
   RECT 5.348 1.848 5.404 1.918 ;
   LAYER m1 ;
   RECT 5.348 0.034 5.404 1.932 ;
   LAYER m1 ;
   RECT 5.348 0.238 5.404 0.306 ;
   LAYER m1 ;
   RECT 5.348 0.098 5.404 0.168 ;
   LAYER m1 ;
   RECT 5.348 0.638 5.404 0.706 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.836 0.034 3.892 1.991 ;
   LAYER m1 ;
   RECT 3.836 1.512 3.892 1.582 ;
   LAYER m1 ;
   RECT 3.836 0.034 3.892 1.991 ;
   LAYER m1 ;
   RECT 3.836 1.392 3.892 1.428 ;
   LAYER m1 ;
   RECT 3.836 1.26 3.892 1.296 ;
   LAYER m1 ;
   RECT 3.836 0.098 3.892 0.168 ;
   LAYER m1 ;
   RECT 3.836 0.238 3.892 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.172 0.034 4.228 1.991 ;
   LAYER m1 ;
   RECT 4.172 1.512 4.228 1.582 ;
   LAYER m1 ;
   RECT 4.172 0.034 4.228 1.991 ;
   LAYER m1 ;
   RECT 4.172 0.638 4.228 0.706 ;
   LAYER m1 ;
   RECT 4.172 0.098 4.228 0.168 ;
   LAYER m1 ;
   RECT 4.172 0.238 4.228 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.34 0.034 4.396 1.991 ;
   LAYER m1 ;
   RECT 4.34 1.512 4.396 1.582 ;
   LAYER m1 ;
   RECT 4.34 0.034 4.396 1.991 ;
   LAYER m1 ;
   RECT 4.34 0.638 4.396 0.706 ;
   LAYER m1 ;
   RECT 4.34 0.238 4.396 0.306 ;
   LAYER m1 ;
   RECT 4.34 0.098 4.396 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.004 0.034 4.06 1.991 ;
   LAYER m1 ;
   RECT 4.004 0.638 4.06 0.706 ;
   LAYER m1 ;
   RECT 4.004 0.034 4.06 1.991 ;
   LAYER m1 ;
   RECT 4.004 0.098 4.06 0.168 ;
   LAYER m1 ;
   RECT 4.004 0.238 4.06 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.164 0.034 3.22 1.991 ;
   LAYER m1 ;
   RECT 3.164 1.106 3.22 1.176 ;
   LAYER m1 ;
   RECT 3.164 0.034 3.22 1.991 ;
   LAYER m1 ;
   RECT 3.164 1.26 3.22 1.296 ;
   LAYER m1 ;
   RECT 3.164 1.512 3.22 1.582 ;
   LAYER m1 ;
   RECT 3.164 1.392 3.22 1.428 ;
   LAYER m1 ;
   RECT 3.164 0.098 3.22 0.168 ;
   LAYER m1 ;
   RECT 3.164 0.238 3.22 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.332 0.034 3.388 1.991 ;
   LAYER m1 ;
   RECT 3.332 1.106 3.388 1.176 ;
   LAYER m1 ;
   RECT 3.332 0.034 3.388 1.991 ;
   LAYER m1 ;
   RECT 3.332 1.26 3.388 1.296 ;
   LAYER m1 ;
   RECT 3.332 1.512 3.388 1.582 ;
   LAYER m1 ;
   RECT 3.332 0.098 3.388 0.168 ;
   LAYER m1 ;
   RECT 3.332 0.238 3.388 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.668 0.034 3.724 1.991 ;
   LAYER m1 ;
   RECT 3.668 1.106 3.724 1.176 ;
   LAYER m1 ;
   RECT 3.668 0.034 3.724 1.991 ;
   LAYER m1 ;
   RECT 3.668 1.26 3.724 1.296 ;
   LAYER m1 ;
   RECT 3.668 1.392 3.724 1.428 ;
   LAYER m1 ;
   RECT 3.668 0.84 3.724 0.91 ;
   LAYER m1 ;
   RECT 3.668 0.098 3.724 0.168 ;
   LAYER m1 ;
   RECT 3.668 0.238 3.724 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 3.5 0.034 3.556 1.991 ;
   LAYER m1 ;
   RECT 3.5 1.26 3.556 1.296 ;
   LAYER m1 ;
   RECT 3.5 0.034 3.556 1.991 ;
   LAYER m1 ;
   RECT 3.5 1.512 3.556 1.582 ;
   LAYER m1 ;
   RECT 3.5 0.84 3.556 0.91 ;
   LAYER m1 ;
   RECT 3.5 0.098 3.556 0.168 ;
   LAYER m1 ;
   RECT 3.5 0.238 3.556 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.996 0.034 3.052 1.991 ;
   LAYER m1 ;
   RECT 2.996 1.26 3.052 1.296 ;
   LAYER m1 ;
   RECT 2.996 0.034 3.052 1.991 ;
   LAYER m1 ;
   RECT 2.996 1.512 3.052 1.582 ;
   LAYER m1 ;
   RECT 2.996 1.392 3.052 1.428 ;
   LAYER m1 ;
   RECT 2.996 0.84 3.052 0.91 ;
   LAYER m1 ;
   RECT 2.996 0.098 3.052 0.168 ;
   LAYER m1 ;
   RECT 2.996 0.238 3.052 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 4.508 0.034 4.564 1.991 ;
   LAYER m1 ;
   RECT 4.508 1.512 4.564 1.582 ;
   LAYER m1 ;
   RECT 4.508 0.034 4.564 1.991 ;
   LAYER m1 ;
   RECT 4.508 0.238 4.564 0.306 ;
   LAYER m1 ;
   RECT 4.508 0.098 4.564 0.168 ;
   LAYER m1 ;
   RECT 4.508 0.638 4.564 0.706 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.66 0.034 2.716 1.991 ;
   LAYER m1 ;
   RECT 2.66 1.106 2.716 1.176 ;
   LAYER m1 ;
   RECT 2.66 0.034 2.716 1.991 ;
   LAYER m1 ;
   RECT 2.66 1.26 2.716 1.296 ;
   LAYER m1 ;
   RECT 2.66 1.392 2.716 1.428 ;
   LAYER m1 ;
   RECT 2.66 1.512 2.716 1.582 ;
   LAYER m1 ;
   RECT 2.66 0.098 2.716 0.168 ;
   LAYER m1 ;
   RECT 2.66 0.238 2.716 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.156 0.034 2.212 1.991 ;
   LAYER m1 ;
   RECT 2.156 1.71 2.212 1.77 ;
   LAYER m1 ;
   RECT 2.156 0.034 2.212 1.991 ;
   LAYER m1 ;
   RECT 2.156 1.106 2.212 1.176 ;
   LAYER m1 ;
   RECT 2.156 1.26 2.212 1.296 ;
   LAYER m1 ;
   RECT 2.156 1.392 2.212 1.428 ;
   LAYER m1 ;
   RECT 2.156 1.512 2.212 1.582 ;
   LAYER m1 ;
   RECT 2.156 0.366 2.212 0.434 ;
   LAYER m1 ;
   RECT 2.156 0.504 2.212 0.574 ;
   LAYER m1 ;
   RECT 2.156 0.638 2.212 0.706 ;
   LAYER m1 ;
   RECT 2.156 0.098 2.212 0.168 ;
   LAYER m1 ;
   RECT 2.156 0.238 2.212 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.324 0.034 2.38 1.991 ;
   LAYER m1 ;
   RECT 2.324 1.106 2.38 1.176 ;
   LAYER m1 ;
   RECT 2.324 0.034 2.38 1.991 ;
   LAYER m1 ;
   RECT 2.324 1.26 2.38 1.296 ;
   LAYER m1 ;
   RECT 2.324 1.512 2.38 1.582 ;
   LAYER m1 ;
   RECT 2.324 0.366 2.38 0.434 ;
   LAYER m1 ;
   RECT 2.324 0.098 2.38 0.168 ;
   LAYER m1 ;
   RECT 2.324 0.238 2.38 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.492 0.034 2.548 1.991 ;
   LAYER m1 ;
   RECT 2.492 1.106 2.548 1.176 ;
   LAYER m1 ;
   RECT 2.492 0.034 2.548 1.991 ;
   LAYER m1 ;
   RECT 2.492 1.26 2.548 1.296 ;
   LAYER m1 ;
   RECT 2.492 1.512 2.548 1.582 ;
   LAYER m1 ;
   RECT 2.492 0.098 2.548 0.168 ;
   LAYER m1 ;
   RECT 2.492 0.238 2.548 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 2.828 0.034 2.884 1.991 ;
   LAYER m1 ;
   RECT 2.828 1.26 2.884 1.296 ;
   LAYER m1 ;
   RECT 2.828 0.034 2.884 1.991 ;
   LAYER m1 ;
   RECT 2.828 1.512 2.884 1.582 ;
   LAYER m1 ;
   RECT 2.828 1.392 2.884 1.428 ;
   LAYER m1 ;
   RECT 2.828 0.84 2.884 0.91 ;
   LAYER m1 ;
   RECT 2.828 0.098 2.884 0.168 ;
   LAYER m1 ;
   RECT 2.828 0.238 2.884 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.652 0.034 1.708 1.991 ;
   LAYER m1 ;
   RECT 1.652 1.106 1.708 1.176 ;
   LAYER m1 ;
   RECT 1.652 0.034 1.708 1.991 ;
   LAYER m1 ;
   RECT 1.652 1.26 1.708 1.296 ;
   LAYER m1 ;
   RECT 1.652 1.512 1.708 1.582 ;
   LAYER m1 ;
   RECT 1.652 0.638 1.708 0.706 ;
   LAYER m1 ;
   RECT 1.652 0.84 1.708 0.91 ;
   LAYER m1 ;
   RECT 1.652 0.504 1.708 0.574 ;
   LAYER m1 ;
   RECT 1.652 0.366 1.708 0.434 ;
   LAYER m1 ;
   RECT 1.652 0.098 1.708 0.168 ;
   LAYER m1 ;
   RECT 1.652 0.238 1.708 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.82 0.034 1.876 1.991 ;
   LAYER m1 ;
   RECT 1.82 1.106 1.876 1.176 ;
   LAYER m1 ;
   RECT 1.82 0.034 1.876 1.991 ;
   LAYER m1 ;
   RECT 1.82 1.26 1.876 1.296 ;
   LAYER m1 ;
   RECT 1.82 1.512 1.876 1.582 ;
   LAYER m1 ;
   RECT 1.82 0.638 1.876 0.706 ;
   LAYER m1 ;
   RECT 1.82 0.84 1.876 0.91 ;
   LAYER m1 ;
   RECT 1.82 0.366 1.876 0.434 ;
   LAYER m1 ;
   RECT 1.82 0.504 1.876 0.574 ;
   LAYER m1 ;
   RECT 1.82 0.238 1.876 0.306 ;
   LAYER m1 ;
   RECT 1.82 0.098 1.876 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.988 0.034 2.044 1.991 ;
   LAYER m1 ;
   RECT 1.988 1.26 2.044 1.296 ;
   LAYER m1 ;
   RECT 1.988 0.034 2.044 1.991 ;
   LAYER m1 ;
   RECT 1.988 1.512 2.044 1.582 ;
   LAYER m1 ;
   RECT 1.988 1.392 2.044 1.428 ;
   LAYER m1 ;
   RECT 1.988 0.638 2.044 0.706 ;
   LAYER m1 ;
   RECT 1.988 0.84 2.044 0.91 ;
   LAYER m1 ;
   RECT 1.988 0.366 2.044 0.434 ;
   LAYER m1 ;
   RECT 1.988 0.504 2.044 0.574 ;
   LAYER m1 ;
   RECT 1.988 0.238 2.044 0.306 ;
   LAYER m1 ;
   RECT 1.988 0.098 2.044 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.484 0.034 1.54 1.991 ;
   LAYER m1 ;
   RECT 1.484 1.26 1.54 1.296 ;
   LAYER m1 ;
   RECT 1.484 0.034 1.54 1.991 ;
   LAYER m1 ;
   RECT 1.484 1.392 1.54 1.428 ;
   LAYER m1 ;
   RECT 1.484 0.638 1.54 0.706 ;
   LAYER m1 ;
   RECT 1.484 0.84 1.54 0.91 ;
   LAYER m1 ;
   RECT 1.484 0.366 1.54 0.434 ;
   LAYER m1 ;
   RECT 1.484 0.504 1.54 0.574 ;
   LAYER m1 ;
   RECT 1.484 0.098 1.54 0.168 ;
   LAYER m1 ;
   RECT 1.484 0.238 1.54 0.306 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.308 1.848 0.364 1.918 ;
   LAYER m1 ;
   RECT 0.308 0.074 0.364 1.932 ;
   LAYER m1 ;
   RECT 0.308 1.512 0.364 1.582 ;
   LAYER m1 ;
   RECT 0.308 0.074 0.364 1.932 ;
   LAYER m1 ;
   RECT 0.308 0.238 0.364 0.306 ;
   LAYER m1 ;
   RECT 0.308 0.098 0.364 0.168 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.14 1.106 0.196 1.176 ;
   LAYER m1 ;
   RECT 0.14 0.074 0.196 1.932 ;
   LAYER m1 ;
   RECT 0.14 1.512 0.196 1.582 ;
   LAYER m1 ;
   RECT 0.14 0.074 0.196 1.932 ;
   LAYER m1 ;
   RECT 0.14 1.392 0.196 1.428 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.476 1.106 0.532 1.176 ;
   LAYER m1 ;
   RECT 0.476 0.074 0.532 1.932 ;
   LAYER m1 ;
   RECT 0.476 1.392 0.532 1.428 ;
   LAYER m1 ;
   RECT 0.476 0.074 0.532 1.932 ;
   LAYER m1 ;
   RECT 0.476 0.238 0.532 0.306 ;
   LAYER m1 ;
   RECT 0.476 0.111 0.532 0.167 ;
   LAYER m1 ;
   RECT 0.476 0.84 0.532 0.91 ;
   LAYER m1 ;
   RECT 0.476 0.978 0.532 1.038 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.316 0.034 1.372 1.991 ;
   LAYER m1 ;
   RECT 1.316 1.26 1.372 1.296 ;
   LAYER m1 ;
   RECT 1.316 0.034 1.372 1.991 ;
   LAYER m1 ;
   RECT 1.316 1.392 1.372 1.428 ;
   LAYER m1 ;
   RECT 1.316 0.366 1.372 0.434 ;
   LAYER m1 ;
   RECT 1.316 0.112 1.372 0.154 ;
   LAYER m1 ;
   RECT 1.316 0.238 1.372 0.306 ;
   LAYER m1 ;
   RECT 1.316 0.504 1.372 0.574 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.98 0.098 1.036 0.168 ;
   LAYER m1 ;
   RECT 0.98 0.063 1.036 0.519 ;
   LAYER m1 ;
   RECT 0.98 0.238 1.036 0.306 ;
   LAYER m1 ;
   RECT 0.98 0.063 1.036 0.519 ;
  END
 END vccdgt_1p0
 PIN vss
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER m1 ;
   RECT 4.676 1.855 4.732 1.992 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.896 1.778 0.952 1.848 ;
   LAYER m1 ;
   RECT 0.896 1.57 0.952 1.915 ;
   LAYER m1 ;
   RECT 0.896 1.582 0.952 1.65 ;
   LAYER m1 ;
   RECT 0.896 1.57 0.952 1.915 ;
  END
  PORT
   LAYER m1 ;
   RECT 1.064 1.778 1.12 1.848 ;
   LAYER m1 ;
   RECT 1.064 0.352 1.12 1.915 ;
   LAYER m1 ;
   RECT 1.064 1.582 1.12 1.65 ;
   LAYER m1 ;
   RECT 1.064 0.352 1.12 1.915 ;
   LAYER m1 ;
   RECT 1.064 0.77 1.12 0.84 ;
   LAYER m1 ;
   RECT 1.064 0.366 1.12 0.434 ;
   LAYER m1 ;
   RECT 1.064 0.588 1.12 0.624 ;
  END
  PORT
   LAYER m1 ;
   RECT 0.812 0.366 0.868 0.434 ;
   LAYER m1 ;
   RECT 0.812 0.085 0.868 0.802 ;
   LAYER m1 ;
   RECT 0.812 0.77 0.868 0.84 ;
   LAYER m1 ;
   RECT 0.812 0.085 0.868 0.802 ;
   LAYER m1 ;
   RECT 0.812 0.588 0.868 0.624 ;
   LAYER m1 ;
   RECT 0.812 0.085 0.868 0.802 ;
   LAYER m1 ;
   RECT 0.812 0.168 0.868 0.238 ;
   LAYER m1 ;
   RECT 0.812 0.366 0.868 0.434 ;
  END
 END vss
 PIN pwren_in
  DIRECTION INPUT ;
  USE SIGNAL ;
 END pwren_in
END c73p4hdxrom_wldrvgappwrcell


END LIBRARY
