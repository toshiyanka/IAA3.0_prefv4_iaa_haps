// File output was printed on: Thursday, March 21, 2013 4:21:02 PM
// Chassis TAP Tool version: 0.6.1.2
// ---------------------------------------------------- 
case (Node)
   'd0 : begin
            Tap_Info_Int.Next_Tap[0] = NOTAP;
        end
endcase


