//-----------------------------------------------------------------
// Intel Proprietary -- Copyright 2013 Intel -- All rights reserved 
//-----------------------------------------------------------------
// Author       : Chris Sadler
// Date Created : 01-2014
//-----------------------------------------------------------------
// Description:
// Systeminit socket picker - this picker should generate the knobs
// that SocketShrTbCfg reads
// except for sim_type, which is generated by topo_base_picker.sv
//------------------------------------------------------------------

// Define & register this picker
`picker_class_begin(socket_picker, base_socket_picker)
//`add_knob_enum("mem_usage", mem_usage, mem_usage_t)
//`add_knob_string("rtl_path", rtl_path)

//`include "socket_picker_cms_knobs.sv"
//constraint mem_usage_c {
//   soft mem_usage == mu_flat_1lm;
//}
  
//  rand pm_integ_socket_picker pm_integ_picker;
//  function void init();
//    super.init();
//    pm_integ_picker = pm_integ_socket_picker::type_id::create("pm_integ_socket_picker", this);
//  endfunction: init;
 
function void pre_randomizes();
   super.pre_randomize();
endfunction: pre_randomizes;

function void post_randomizes();
   super.pre_randomize();
   //set_config_int("*.mc0", "dir_enable", dir_enable);
endfunction: post_randomizes;
  
function void build();
   //topo_base_picker mc_pickers[$];
   //mc_picker my_mc_picker;
   //int size_mb;
   //`ovm_info(get_name(), "build()", OVM_NONE)
   //   size_mb = 0;
   //get_pickers_of_type("MC",mc_pickers);
   //foreach(mc_pickers[i]) begin
   //   //$display("%p", mc_pickers[i]);
   //   $cast(my_mc_picker,mc_pickers[i]);
   //   size_mb = size_mb + my_mc_picker.total_mb_mem;
   //end
   //$display("S0 Size MB %d\n", size_mb);
   //total_mb_mem = size_mb;

   super.build();
endfunction: build;

function void connect();
   topo_base_picker sapma_pickers[$];
 //  sapma_picker my_sapma_picker;

   //topo_base_picker mcddr_pll_pickers[$];
   //mcddr_pll_picker my_mcddr_pll_picker;

   //topo_base_picker mcddr_mee_pickers[$];
   //base_mcddr_mee_chassis_picker my_mcddr_mee_picker;

   //topo_base_picker domain_pickers[$];
   //domain_picker my_domain_picker;

 //  get_pickers_of_type("SAPMA",sapma_pickers);
   //get_pickers_of_type("MCDDR_PLL",mcddr_pll_pickers);
   //get_pickers_of_type("MCDDR_MEE_CHASSIS",mcddr_mee_pickers);
   
  // foreach(sapma_pickers[i]) begin
  //    $cast(my_sapma_picker,sapma_pickers[i]);
      //if ( !$cast(my_mcddr_pll_picker,mcddr_pll_pickers[i]) )`ovm_fatal( "socket_picker", "cast failed to my_mcddr_pll_picker" )	
      //$cast(my_mcddr_mee_picker,mcddr_mee_pickers[i]);
      	
  //    `override_cfg_val(my_sapma_picker.domains[0].pll_ratio, socket_clocks.pll_pickers[5].multiplier); 
      //`override_cfg_val(my_sapma_picker.domains[0].pll_ratio,my_mcddr_pll_picker.mltiplier);  
      //`override_cfg_val(my_sapma_picker.domains[0].pll_ratio,my_mcddr_mee_picker.pll_ratio);	
  // end

   super.connect();
endfunction: connect

`picker_class_end
