`iosf_sb_port_agent_inst(8,0,1,4,1,0,0)
