
///
///  INTEL CONFIDENTIAL
///
///  Copyright 2015 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

 module hqm_rcfwl_gclk_psocclkdist 
 #(
	NUM_OF_OUTPUTS    = 'd1
    
    )
 (
  input  logic			        clk_in,
  output logic  [NUM_OF_OUTPUTS-1:0]	clk_out
   
);


 generate
genvar i;

  for( i=0;i<NUM_OF_OUTPUTS ; i=i+1)
   begin: gen_clkdist_rptrs
    assign clk_out[i] = clk_in; 
    end
endgenerate
   
 
 endmodule
 
 

 
