// RTL Generated using Collage

module hqm_sip_gated_wrap (
    output          ap_alarm_down_v,
    output          ap_alarm_up_ready,
    output          ap_aqed_ready,
    output          ap_aqed_v,
    output          ap_cfg_req_down_read,
    output          ap_cfg_req_down_write,
    output          ap_cfg_rsp_down_ack,
    output          aqed_alarm_down_v,
    output          aqed_ap_enq_ready,
    output          aqed_ap_enq_v,
    output          aqed_chp_sch_ready,
    output          aqed_chp_sch_v,
    output          aqed_lsp_sch_ready,
    output          aqed_lsp_sch_v,
    output          aqed_unit_idle,
    output          chp_alarm_up_ready,
    output          chp_cfg_req_down_read,
    output          chp_cfg_req_down_write,
    output          chp_cfg_rsp_down_ack,
    output          chp_lsp_cmp_ready,
    output          chp_lsp_cmp_v,
    output          chp_lsp_token_ready,
    output          chp_lsp_token_v,
    output          chp_rop_hcw_ready,
    output          chp_rop_hcw_v,
    output          cwdi_interrupt_w_req_ready,
    output          cwdi_interrupt_w_req_valid,
    output          dp_lsp_enq_dir_ready,
    output          dp_lsp_enq_dir_v,
    output          dp_lsp_enq_rorply_ready,
    output          dp_lsp_enq_rorply_v,
    output          hcw_enq_w_req_ready,
    output          hcw_enq_w_req_valid,
    output          hcw_sched_w_req_ready,
    output          hcw_sched_w_req_valid,
    output          hqm_alarm_ready,
    output          hqm_alarm_v,
    output          hqm_proc_clk_en_chp,
    output          hqm_proc_clk_en_dir,
    output          hqm_proc_clk_en_lsp,
    output          hqm_proc_clk_en_nalb,
    output          hqm_proc_clk_en_sys,
    output          interrupt_w_req_ready,
    output          interrupt_w_req_valid,
    output          lsp_alarm_down_v,
    output          lsp_alarm_up_ready,
    output          lsp_cfg_req_down_read,
    output          lsp_cfg_req_down_write,
    output          lsp_cfg_rsp_down_ack,
    output          lsp_dp_sch_dir_ready,
    output          lsp_dp_sch_dir_v,
    output          lsp_dp_sch_rorply_ready,
    output          lsp_dp_sch_rorply_v,
    output          lsp_nalb_sch_atq_ready,
    output          lsp_nalb_sch_atq_v,
    output          lsp_nalb_sch_rorply_ready,
    output          lsp_nalb_sch_rorply_v,
    output          lsp_nalb_sch_unoord_ready,
    output          lsp_nalb_sch_unoord_v,
    output          nalb_lsp_enq_lb_ready,
    output          nalb_lsp_enq_lb_v,
    output          nalb_lsp_enq_rorply_ready,
    output          nalb_lsp_enq_rorply_v,
    output          qed_alarm_down_v,
    output          qed_alarm_up_ready,
    output          qed_aqed_enq_ready,
    output          qed_aqed_enq_v,
    output          qed_cfg_req_down_read,
    output          qed_cfg_req_down_write,
    output          qed_cfg_rsp_down_ack,
    output          qed_chp_sch_ready,
    output          qed_chp_sch_v,
    output          rop_alarm_down_v,
    output          rop_alarm_up_ready,
    output          rop_cfg_req_down_read,
    output          rop_cfg_req_down_write,
    output          rop_cfg_rsp_down_ack,
    output          rop_dp_enq_ready,
    output          rop_dp_enq_v,
    output          rop_dqed_enq_ready,
    output          rop_lsp_reordercmp_ready,
    output          rop_lsp_reordercmp_v,
    output          rop_nalb_enq_ready,
    output          rop_nalb_enq_v,
    output          rop_qed_dqed_enq_v,
    output          rop_qed_enq_ready,
    output          rop_qed_force_clockon,
    output          rop_unit_idle,
    output          system_cfg_req_down_read,
    output          system_cfg_req_down_write,
    output          system_cfg_rsp_down_ack,
    // Ports for Manually exported pins
    input           fscan_byprst_b,
    input           fscan_clkungate,
    input           fscan_rstbypen,
    input   [160:0] hcw_enq_in_data,
    input           hcw_enq_in_v,
    input           hqm_clk_enable,
    input           hqm_clk_rptr_rst_b,
    input           hqm_clk_trunk,
    input           hqm_clk_ungate,
    input           hqm_flr_prep,
    input           hqm_gated_local_override,
    input           hqm_gated_rst_b,
    input           hqm_proc_reset_done_sync_hqm,
    input   [2047:0] i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cmatch,
    input   [207:0] i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_rdata,
    input   [16:0]  i_hqm_aqed_pipe_rf_aqed_fid_cnt_rdata,
    input   [44:0]  i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rdata,
    input   [23:0]  i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rdata,
    input   [179:0] i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rdata,
    input   [31:0]  i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rdata,
    input   [34:0]  i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rdata,
    input   [152:0] i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rdata,
    input   [154:0] i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rdata,
    input   [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rdata,
    input   [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rdata,
    input   [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rdata,
    input   [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rdata,
    input   [14:0]  i_hqm_aqed_pipe_rf_aqed_qid_cnt_rdata,
    input   [13:0]  i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rdata,
    input   [138:0] i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rdata,
    input   [15:0]  i_hqm_aqed_pipe_sr_aqed_freelist_rdata,
    input   [15:0]  i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_rdata,
    input   [138:0] i_hqm_aqed_pipe_sr_aqed_rdata,
    input   [178:0] i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rdata,
    input   [200:0] i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rdata,
    input   [73:0]  i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rdata,
    input   [28:0]  i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rdata,
    input   [199:0] i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rdata,
    input   [1:0]   i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rdata,
    input   [9:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rdata,
    input   [9:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rdata,
    input   [12:0]  i_hqm_credit_hist_pipe_rf_dir_cq_depth_rdata,
    input   [14:0]  i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rdata,
    input   [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rdata,
    input   [12:0]  i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rdata,
    input   [159:0] i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rdata,
    input   [29:0]  i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rdata,
    input   [31:0]  i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rdata,
    input   [29:0]  i_hqm_credit_hist_pipe_rf_hist_list_minmax_rdata,
    input   [31:0]  i_hqm_credit_hist_pipe_rf_hist_list_ptr_rdata,
    input   [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rdata,
    input   [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rdata,
    input   [31:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rdata,
    input   [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rdata,
    input   [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rdata,
    input   [11:0]  i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rdata,
    input   [11:0]  i_hqm_credit_hist_pipe_rf_ord_qid_sn_rdata,
    input   [159:0] i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rdata,
    input   [25:0]  i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rdata,
    input   [176:0] i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rdata,
    input   [196:0] i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rdata,
    input   [13:0]  i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rdata,
    input   [13:0]  i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_0_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_1_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_2_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_3_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_4_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_5_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_6_rdata,
    input   [15:0]  i_hqm_credit_hist_pipe_sr_freelist_7_rdata,
    input   [65:0]  i_hqm_credit_hist_pipe_sr_hist_list_a_rdata,
    input   [65:0]  i_hqm_credit_hist_pipe_sr_hist_list_rdata,
    input   [8:0]   i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rdata,
    input   [527:0] i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rdata,
    input   [54:0]  i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rdata,
    input   [44:0]  i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rdata,
    input   [23:0]  i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rdata,
    input   [32:0]  i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rdata,
    input   [32:0]  i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rdata,
    input   [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rdata,
    input   [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rdata,
    input   [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rdata,
    input   [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rdata,
    input   [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rdata,
    input   [12:0]  i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rdata,
    input   [12:0]  i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rdata,
    input   [527:0] i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rdata,
    input   [527:0] i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rdata,
    input   [72:0]  i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata,
    input   [24:0]  i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rdata,
    input   [95:0]  i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rdata,
    input   [65:0]  i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rdata,
    input   [14:0]  i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rdata,
    input   [12:0]  i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rdata,
    input   [65:0]  i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rdata,
    input   [18:0]  i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rdata,
    input   [95:0]  i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rdata,
    input   [12:0]  i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rdata,
    input   [7:0]   i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rdata,
    input   [7:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata,
    input   [22:0]  i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata,
    input   [9:0]   i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rdata,
    input   [11:0]  i_hqm_list_sel_pipe_rf_fid2cqqidix_rdata,
    input   [24:0]  i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rdata,
    input   [55:0]  i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rdata,
    input   [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rdata,
    input   [59:0]  i_hqm_list_sel_pipe_rf_ll_slst_cnt_rdata,
    input   [17:0]  i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rdata,
    input   [9:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata,
    input   [26:0]  i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata,
    input   [26:0]  i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rdata,
    input   [8:0]   i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rdata,
    input   [65:0]  i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rdata,
    input   [14:0]  i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rdata,
    input   [65:0]  i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rdata,
    input   [13:0]  i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rdata,
    input   [14:0]  i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rdata,
    input   [65:0]  i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rdata,
    input   [5:0]   i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rdata,
    input   [16:0]  i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata,
    input   [34:0]  i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rdata,
    input   [19:0]  i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rdata,
    input   [67:0]  i_hqm_qed_pipe_rf_atq_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_atq_hp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_atq_tp_rdata,
    input   [67:0]  i_hqm_qed_pipe_rf_dir_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_hp_rdata,
    input   [67:0]  i_hqm_qed_pipe_rf_dir_replay_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_replay_hp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_replay_tp_rdata,
    input   [16:0]  i_hqm_qed_pipe_rf_dir_rofrag_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_rofrag_hp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_rofrag_tp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_dir_tp_rdata,
    input   [44:0]  i_hqm_qed_pipe_rf_dp_dqed_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rdata,
    input   [22:0]  i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rdata,
    input   [26:0]  i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rdata,
    input   [26:0]  i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rdata,
    input   [67:0]  i_hqm_qed_pipe_rf_nalb_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_hp_rdata,
    input   [26:0]  i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rdata,
    input   [9:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rdata,
    input   [44:0]  i_hqm_qed_pipe_rf_nalb_qed_rdata,
    input   [67:0]  i_hqm_qed_pipe_rf_nalb_replay_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_replay_hp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_replay_tp_rdata,
    input   [16:0]  i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_rofrag_hp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_rofrag_tp_rdata,
    input   [14:0]  i_hqm_qed_pipe_rf_nalb_tp_rdata,
    input   [176:0] i_hqm_qed_pipe_rf_qed_chp_sch_data_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rop_dp_enq_dir_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rop_dp_enq_ro_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rdata,
    input   [44:0]  i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rdata,
    input   [26:0]  i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rdata,
    input   [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rdata,
    input   [26:0]  i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rdata,
    input   [44:0]  i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rdata,
    input   [99:0]  i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rdata,
    input   [156:0] i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rdata,
    input   [20:0]  i_hqm_qed_pipe_sr_dir_nxthp_rdata,
    input   [20:0]  i_hqm_qed_pipe_sr_nalb_nxthp_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_0_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_1_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_2_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_3_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_4_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_5_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_6_rdata,
    input   [138:0] i_hqm_qed_pipe_sr_qed_7_rdata,
    input   [59:0]  i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rdata,
    input   [59:0]  i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rdata,
    input   [18:0]  i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rdata,
    input   [15:0]  i_hqm_reorder_pipe_rf_reord_cnt_mem_rdata,
    input   [16:0]  i_hqm_reorder_pipe_rf_reord_dirhp_mem_rdata,
    input   [16:0]  i_hqm_reorder_pipe_rf_reord_dirtp_mem_rdata,
    input   [16:0]  i_hqm_reorder_pipe_rf_reord_lbhp_mem_rdata,
    input   [16:0]  i_hqm_reorder_pipe_rf_reord_lbtp_mem_rdata,
    input   [24:0]  i_hqm_reorder_pipe_rf_reord_st_mem_rdata,
    input   [203:0] i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rdata,
    input   [11:0]  i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rdata,
    input   [11:0]  i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rdata,
    input   [20:0]  i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rdata,
    input   [12:0]  i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rdata,
    input   [29:0]  i_hqm_system_rf_alarm_vf_synd0_rdata,
    input   [31:0]  i_hqm_system_rf_alarm_vf_synd1_rdata,
    input   [31:0]  i_hqm_system_rf_alarm_vf_synd2_rdata,
    input   [143:0] i_hqm_system_rf_dir_wb0_rdata,
    input   [143:0] i_hqm_system_rf_dir_wb1_rdata,
    input   [143:0] i_hqm_system_rf_dir_wb2_rdata,
    input   [166:0] i_hqm_system_rf_hcw_enq_fifo_rdata,
    input   [143:0] i_hqm_system_rf_ldb_wb0_rdata,
    input   [143:0] i_hqm_system_rf_ldb_wb1_rdata,
    input   [143:0] i_hqm_system_rf_ldb_wb2_rdata,
    input   [12:0]  i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rdata,
    input   [26:0]  i_hqm_system_rf_lut_dir_cq_addr_l_rdata,
    input   [32:0]  i_hqm_system_rf_lut_dir_cq_addr_u_rdata,
    input   [30:0]  i_hqm_system_rf_lut_dir_cq_ai_addr_l_rdata,
    input   [32:0]  i_hqm_system_rf_lut_dir_cq_ai_addr_u_rdata,
    input   [32:0]  i_hqm_system_rf_lut_dir_cq_ai_data_rdata,
    input   [12:0]  i_hqm_system_rf_lut_dir_cq_isr_rdata,
    input   [23:0]  i_hqm_system_rf_lut_dir_cq_pasid_rdata,
    input   [10:0]  i_hqm_system_rf_lut_dir_pp2vas_rdata,
    input   [16:0]  i_hqm_system_rf_lut_dir_pp_v_rdata,
    input   [32:0]  i_hqm_system_rf_lut_dir_vasqid_v_rdata,
    input   [12:0]  i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rdata,
    input   [26:0]  i_hqm_system_rf_lut_ldb_cq_addr_l_rdata,
    input   [32:0]  i_hqm_system_rf_lut_ldb_cq_addr_u_rdata,
    input   [30:0]  i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rdata,
    input   [32:0]  i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rdata,
    input   [32:0]  i_hqm_system_rf_lut_ldb_cq_ai_data_rdata,
    input   [12:0]  i_hqm_system_rf_lut_ldb_cq_isr_rdata,
    input   [23:0]  i_hqm_system_rf_lut_ldb_cq_pasid_rdata,
    input   [10:0]  i_hqm_system_rf_lut_ldb_pp2vas_rdata,
    input   [20:0]  i_hqm_system_rf_lut_ldb_qid2vqid_rdata,
    input   [16:0]  i_hqm_system_rf_lut_ldb_vasqid_v_rdata,
    input   [30:0]  i_hqm_system_rf_lut_vf_dir_vpp2pp_rdata,
    input   [16:0]  i_hqm_system_rf_lut_vf_dir_vpp_v_rdata,
    input   [30:0]  i_hqm_system_rf_lut_vf_dir_vqid2qid_rdata,
    input   [16:0]  i_hqm_system_rf_lut_vf_dir_vqid_v_rdata,
    input   [24:0]  i_hqm_system_rf_lut_vf_ldb_vpp2pp_rdata,
    input   [16:0]  i_hqm_system_rf_lut_vf_ldb_vpp_v_rdata,
    input   [26:0]  i_hqm_system_rf_lut_vf_ldb_vqid2qid_rdata,
    input   [16:0]  i_hqm_system_rf_lut_vf_ldb_vqid_v_rdata,
    input   [32:0]  i_hqm_system_rf_msix_tbl_word0_rdata,
    input   [32:0]  i_hqm_system_rf_msix_tbl_word1_rdata,
    input   [32:0]  i_hqm_system_rf_msix_tbl_word2_rdata,
    input   [269:0] i_hqm_system_rf_sch_out_fifo_rdata,
    input           i_hqm_system_side_rst_sync_prim_n_rst_n,
    input   [155:0] i_hqm_system_sr_rob_mem_rdata,
    input   [15:0]  master_chp_timestamp,
    input   [92:0]  mstr_cfg_req_down,
    input           mstr_cfg_req_down_read,
    input           mstr_cfg_req_down_write,
    input           pci_cfg_pmsixctl_fm,
    input           pci_cfg_pmsixctl_msie,
    input           pci_cfg_sciov_en,
    input           pgcb_clk,
    input           prim_clk,
    input           prim_clk_enable,
    input           prim_clk_ungate,
    input   [24:0]  sif_alarm_data,
    input           sif_alarm_v,
    input           write_buffer_mstr_ready,
    output          ap_reset_done,
    output          ap_unit_idle,
    output          ap_unit_pipeidle,
    output  [92:0]  aqed_cfg_req_down,
    output          aqed_cfg_req_down_read,
    output          aqed_cfg_req_down_write,
    output  [38:0]  aqed_cfg_rsp_down,
    output          aqed_cfg_rsp_down_ack,
    output          aqed_reset_done,
    output          aqed_unit_pipeidle,
    output          chp_reset_done,
    output          chp_unit_idle,
    output          chp_unit_pipeidle,
    output          dp_reset_done,
    output          dp_unit_idle,
    output          dp_unit_pipeidle,
    output          hcw_enq_in_ready,
    output          hqm_proc_clk_en_qed,
    output  [29:0]  hqm_system_visa_str,
    output          i_hqm_aqed_pipe_aqed_lsp_deq_v,
    output          i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cclk,
    output  [207:0] i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cdata,
    output  [7:0]   i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_ce,
    output          i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_dfx_clk,
    output  [7:0]   i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_raddr,
    output          i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_rclk,
    output          i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_re,
    output  [63:0]  i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_waddr,
    output          i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_wclk,
    output  [207:0] i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_wdata,
    output  [7:0]   i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_fid_cnt_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_fid_cnt_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_wclk_rst_n,
    output  [16:0]  i_hqm_aqed_pipe_rf_aqed_fid_cnt_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fid_cnt_we,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_re,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wclk_rst_n,
    output  [44:0]  i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_we,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_re,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wclk_rst_n,
    output  [23:0]  i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_we,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_re,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wclk_rst_n,
    output  [179:0] i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_we,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_re,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wclk_rst_n,
    output  [31:0]  i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_we,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_re,
    output  [3:0]   i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wclk_rst_n,
    output  [34:0]  i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_we,
    output  [2:0]   i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_re,
    output  [2:0]   i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wclk_rst_n,
    output  [152:0] i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_we,
    output  [1:0]   i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_re,
    output  [1:0]   i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wclk_rst_n,
    output  [154:0] i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wclk_rst_n,
    output  [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wclk_rst_n,
    output  [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wclk_rst_n,
    output  [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wclk_rst_n,
    output  [15:0]  i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_we,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_re,
    output  [10:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_we,
    output  [4:0]   i_hqm_aqed_pipe_rf_aqed_qid_cnt_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_re,
    output  [4:0]   i_hqm_aqed_pipe_rf_aqed_qid_cnt_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_wclk_rst_n,
    output  [14:0]  i_hqm_aqed_pipe_rf_aqed_qid_cnt_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_qid_cnt_we,
    output  [4:0]   i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_raddr,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rclk,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_re,
    output  [4:0]   i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_waddr,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wclk,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wclk_rst_n,
    output  [13:0]  i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wdata,
    output          i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_we,
    output  [1:0]   i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_raddr,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rclk,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rclk_rst_n,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_re,
    output  [1:0]   i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_waddr,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wclk,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wclk_rst_n,
    output  [138:0] i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wdata,
    output          i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_we,
    output  [10:0]  i_hqm_aqed_pipe_sr_aqed_addr,
    output          i_hqm_aqed_pipe_sr_aqed_clk,
    output          i_hqm_aqed_pipe_sr_aqed_clk_rst_n,
    output  [10:0]  i_hqm_aqed_pipe_sr_aqed_freelist_addr,
    output          i_hqm_aqed_pipe_sr_aqed_freelist_clk,
    output          i_hqm_aqed_pipe_sr_aqed_freelist_clk_rst_n,
    output          i_hqm_aqed_pipe_sr_aqed_freelist_re,
    output  [15:0]  i_hqm_aqed_pipe_sr_aqed_freelist_wdata,
    output          i_hqm_aqed_pipe_sr_aqed_freelist_we,
    output  [10:0]  i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_addr,
    output          i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_clk,
    output          i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_clk_rst_n,
    output          i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_re,
    output  [15:0]  i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_wdata,
    output          i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_we,
    output          i_hqm_aqed_pipe_sr_aqed_re,
    output  [138:0] i_hqm_aqed_pipe_sr_aqed_wdata,
    output          i_hqm_aqed_pipe_sr_aqed_we,
    output  [1:0]   i_hqm_credit_hist_pipe_chp_cfg_req_down_1_0,
    output  [1:0]   i_hqm_credit_hist_pipe_chp_cfg_rsp_down_5_4,
    output  [1:0]   i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_re,
    output  [1:0]   i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wclk_rst_n,
    output  [178:0] i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_we,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_re,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wclk_rst_n,
    output  [200:0] i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_we,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_re,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wclk_rst_n,
    output  [73:0]  i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_we,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_re,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wclk_rst_n,
    output  [28:0]  i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_we,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_re,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wclk_rst_n,
    output  [199:0] i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wclk_rst_n,
    output  [1:0]   i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wclk_rst_n,
    output  [15:0]  i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wclk_rst_n,
    output  [15:0]  i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wclk_rst_n,
    output  [9:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wclk_rst_n,
    output  [9:0]   i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_depth_raddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_rclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_depth_waddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_wclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_wclk_rst_n,
    output  [12:0]  i_hqm_credit_hist_pipe_rf_dir_cq_depth_wdata,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_depth_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_raddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_waddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wclk_rst_n,
    output  [14:0]  i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wdata,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_raddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_waddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wclk_rst_n,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wdata,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_wptr_raddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_dir_cq_wptr_waddr,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wclk,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wclk_rst_n,
    output  [12:0]  i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wdata,
    output          i_hqm_credit_hist_pipe_rf_dir_cq_wptr_we,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_re,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wclk_rst_n,
    output  [159:0] i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_raddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_waddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wclk_rst_n,
    output  [29:0]  i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wdata,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_raddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_waddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wclk_rst_n,
    output  [31:0]  i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wdata,
    output          i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_minmax_raddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_rclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_minmax_waddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_wclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_wclk_rst_n,
    output  [29:0]  i_hqm_credit_hist_pipe_rf_hist_list_minmax_wdata,
    output          i_hqm_credit_hist_pipe_rf_hist_list_minmax_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_ptr_raddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_rclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_hist_list_ptr_waddr,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_wclk,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_wclk_rst_n,
    output  [31:0]  i_hqm_credit_hist_pipe_rf_hist_list_ptr_wdata,
    output          i_hqm_credit_hist_pipe_rf_hist_list_ptr_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_depth_raddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_depth_waddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wclk_rst_n,
    output  [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wdata,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_depth_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_raddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_waddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wclk_rst_n,
    output  [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wdata,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_raddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_waddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wclk_rst_n,
    output  [31:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wdata,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_raddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_waddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wclk_rst_n,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wdata,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_raddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_waddr,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wclk,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wclk_rst_n,
    output  [12:0]  i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wdata,
    output          i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_we,
    output  [4:0]   i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_raddr,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rclk,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_re,
    output  [4:0]   i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_waddr,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wclk,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wclk_rst_n,
    output  [11:0]  i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wdata,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_we,
    output  [4:0]   i_hqm_credit_hist_pipe_rf_ord_qid_sn_raddr,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_rclk,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_re,
    output  [4:0]   i_hqm_credit_hist_pipe_rf_ord_qid_sn_waddr,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_wclk,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_wclk_rst_n,
    output  [11:0]  i_hqm_credit_hist_pipe_rf_ord_qid_sn_wdata,
    output          i_hqm_credit_hist_pipe_rf_ord_qid_sn_we,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_re,
    output  [3:0]   i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wclk_rst_n,
    output  [159:0] i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_we,
    output  [1:0]   i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_re,
    output  [1:0]   i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk_rst_n,
    output  [25:0]  i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_we,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_re,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wclk_rst_n,
    output  [176:0] i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_we,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_re,
    output  [2:0]   i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wclk_rst_n,
    output  [196:0] i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wclk_rst_n,
    output  [13:0]  i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_we,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_raddr,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rclk,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rclk_rst_n,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_re,
    output  [5:0]   i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_waddr,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wclk,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wclk_rst_n,
    output  [13:0]  i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wdata,
    output          i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_0_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_0_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_0_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_0_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_0_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_0_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_1_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_1_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_1_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_1_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_1_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_1_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_2_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_2_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_2_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_2_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_2_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_2_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_3_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_3_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_3_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_3_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_3_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_3_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_4_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_4_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_4_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_4_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_4_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_4_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_5_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_5_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_5_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_5_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_5_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_5_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_6_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_6_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_6_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_6_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_6_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_6_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_freelist_7_addr,
    output          i_hqm_credit_hist_pipe_sr_freelist_7_clk,
    output          i_hqm_credit_hist_pipe_sr_freelist_7_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_freelist_7_re,
    output  [15:0]  i_hqm_credit_hist_pipe_sr_freelist_7_wdata,
    output          i_hqm_credit_hist_pipe_sr_freelist_7_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_hist_list_a_addr,
    output          i_hqm_credit_hist_pipe_sr_hist_list_a_clk,
    output          i_hqm_credit_hist_pipe_sr_hist_list_a_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_hist_list_a_re,
    output  [65:0]  i_hqm_credit_hist_pipe_sr_hist_list_a_wdata,
    output          i_hqm_credit_hist_pipe_sr_hist_list_a_we,
    output  [10:0]  i_hqm_credit_hist_pipe_sr_hist_list_addr,
    output          i_hqm_credit_hist_pipe_sr_hist_list_clk,
    output          i_hqm_credit_hist_pipe_sr_hist_list_clk_rst_n,
    output          i_hqm_credit_hist_pipe_sr_hist_list_re,
    output  [65:0]  i_hqm_credit_hist_pipe_sr_hist_list_wdata,
    output          i_hqm_credit_hist_pipe_sr_hist_list_we,
    output  [1:0]   i_hqm_list_sel_pipe_ap_cfg_req_down_1_0,
    output  [1:0]   i_hqm_list_sel_pipe_ap_cfg_rsp_down_5_4,
    output  [1:0]   i_hqm_list_sel_pipe_lsp_cfg_req_down_1_0,
    output  [1:0]   i_hqm_list_sel_pipe_lsp_cfg_rsp_down_5_4,
    output  [4:0]   i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wclk_rst_n,
    output  [8:0]   i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_raddr,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rclk,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_waddr,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wclk,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wclk_rst_n,
    output  [527:0] i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wdata,
    output          i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_we,
    output  [2:0]   i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_re,
    output  [2:0]   i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wclk_rst_n,
    output  [54:0]  i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_we,
    output  [3:0]   i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_raddr,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rclk,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_re,
    output  [3:0]   i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_waddr,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wclk,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wclk_rst_n,
    output  [44:0]  i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wdata,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_raddr,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rclk,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_waddr,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wclk,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wclk_rst_n,
    output  [23:0]  i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wdata,
    output          i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wclk_rst_n,
    output  [32:0]  i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wclk_rst_n,
    output  [32:0]  i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wclk_rst_n,
    output  [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wclk_rst_n,
    output  [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wclk_rst_n,
    output  [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wclk_rst_n,
    output  [28:0]  i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n,
    output  [12:0]  i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n,
    output  [12:0]  i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n,
    output  [527:0] i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n,
    output  [527:0] i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n,
    output  [72:0]  i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n,
    output  [24:0]  i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wclk_rst_n,
    output  [95:0]  i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n,
    output  [65:0]  i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wclk_rst_n,
    output  [14:0]  i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wclk_rst_n,
    output  [12:0]  i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n,
    output  [65:0]  i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wclk_rst_n,
    output  [18:0]  i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wclk_rst_n,
    output  [95:0]  i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wclk_rst_n,
    output  [12:0]  i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wclk_rst_n,
    output  [7:0]   i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n,
    output  [7:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n,
    output  [22:0]  i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wclk_rst_n,
    output  [9:0]   i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_fid2cqqidix_raddr,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_rclk,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_fid2cqqidix_waddr,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_wclk,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_wclk_rst_n,
    output  [11:0]  i_hqm_list_sel_pipe_rf_fid2cqqidix_wdata,
    output          i_hqm_list_sel_pipe_rf_fid2cqqidix_we,
    output  [2:0]   i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_re,
    output  [2:0]   i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wclk_rst_n,
    output  [24:0]  i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rlst_cnt_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_ll_rlst_cnt_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wclk_rst_n,
    output  [55:0]  i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_rlst_cnt_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_we,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_re,
    output  [10:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wclk_rst_n,
    output  [15:0]  i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_we,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_slst_cnt_raddr,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_rclk,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_re,
    output  [8:0]   i_hqm_list_sel_pipe_rf_ll_slst_cnt_waddr,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_wclk,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_wclk_rst_n,
    output  [59:0]  i_hqm_list_sel_pipe_rf_ll_slst_cnt_wdata,
    output          i_hqm_list_sel_pipe_rf_ll_slst_cnt_we,
    output  [2:0]   i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_re,
    output  [2:0]   i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wclk_rst_n,
    output  [17:0]  i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n,
    output  [9:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n,
    output  [26:0]  i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we,
    output  [3:0]   i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_re,
    output  [3:0]   i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wclk_rst_n,
    output  [26:0]  i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wclk_rst_n,
    output  [8:0]   i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atm_active_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atm_active_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_atm_active_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n,
    output  [65:0]  i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wclk_rst_n,
    output  [14:0]  i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_we,
    output  [5:0]   i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_re,
    output  [5:0]   i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n,
    output  [65:0]  i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wclk_rst_n,
    output  [13:0]  i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wclk_rst_n,
    output  [14:0]  i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n,
    output  [65:0]  i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_we,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_raddr,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rclk,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_re,
    output  [4:0]   i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_waddr,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wclk,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wclk_rst_n,
    output  [5:0]   i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wdata,
    output          i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_we,
    output  [2:0]   i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re,
    output  [2:0]   i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n,
    output  [16:0]  i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we,
    output  [1:0]   i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_re,
    output  [1:0]   i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n,
    output  [34:0]  i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_we,
    output  [2:0]   i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_raddr,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rclk,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rclk_rst_n,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_re,
    output  [2:0]   i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_waddr,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wclk,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wclk_rst_n,
    output  [19:0]  i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wdata,
    output          i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_we,
    output  [1:0]   i_hqm_qed_pipe_qed_cfg_req_down_1_0,
    output  [1:0]   i_hqm_qed_pipe_qed_cfg_rsp_down_5_4,
    output          i_hqm_qed_pipe_qed_lsp_deq_v,
    output  [4:0]   i_hqm_qed_pipe_rf_atq_cnt_raddr,
    output          i_hqm_qed_pipe_rf_atq_cnt_rclk,
    output          i_hqm_qed_pipe_rf_atq_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_atq_cnt_re,
    output  [4:0]   i_hqm_qed_pipe_rf_atq_cnt_waddr,
    output          i_hqm_qed_pipe_rf_atq_cnt_wclk,
    output          i_hqm_qed_pipe_rf_atq_cnt_wclk_rst_n,
    output  [67:0]  i_hqm_qed_pipe_rf_atq_cnt_wdata,
    output          i_hqm_qed_pipe_rf_atq_cnt_we,
    output  [6:0]   i_hqm_qed_pipe_rf_atq_hp_raddr,
    output          i_hqm_qed_pipe_rf_atq_hp_rclk,
    output          i_hqm_qed_pipe_rf_atq_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_atq_hp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_atq_hp_waddr,
    output          i_hqm_qed_pipe_rf_atq_hp_wclk,
    output          i_hqm_qed_pipe_rf_atq_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_atq_hp_wdata,
    output          i_hqm_qed_pipe_rf_atq_hp_we,
    output  [6:0]   i_hqm_qed_pipe_rf_atq_tp_raddr,
    output          i_hqm_qed_pipe_rf_atq_tp_rclk,
    output          i_hqm_qed_pipe_rf_atq_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_atq_tp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_atq_tp_waddr,
    output          i_hqm_qed_pipe_rf_atq_tp_wclk,
    output          i_hqm_qed_pipe_rf_atq_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_atq_tp_wdata,
    output          i_hqm_qed_pipe_rf_atq_tp_we,
    output  [5:0]   i_hqm_qed_pipe_rf_dir_cnt_raddr,
    output          i_hqm_qed_pipe_rf_dir_cnt_rclk,
    output          i_hqm_qed_pipe_rf_dir_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_cnt_re,
    output  [5:0]   i_hqm_qed_pipe_rf_dir_cnt_waddr,
    output          i_hqm_qed_pipe_rf_dir_cnt_wclk,
    output          i_hqm_qed_pipe_rf_dir_cnt_wclk_rst_n,
    output  [67:0]  i_hqm_qed_pipe_rf_dir_cnt_wdata,
    output          i_hqm_qed_pipe_rf_dir_cnt_we,
    output  [7:0]   i_hqm_qed_pipe_rf_dir_hp_raddr,
    output          i_hqm_qed_pipe_rf_dir_hp_rclk,
    output          i_hqm_qed_pipe_rf_dir_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_hp_re,
    output  [7:0]   i_hqm_qed_pipe_rf_dir_hp_waddr,
    output          i_hqm_qed_pipe_rf_dir_hp_wclk,
    output          i_hqm_qed_pipe_rf_dir_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_hp_wdata,
    output          i_hqm_qed_pipe_rf_dir_hp_we,
    output  [4:0]   i_hqm_qed_pipe_rf_dir_replay_cnt_raddr,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_rclk,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_re,
    output  [4:0]   i_hqm_qed_pipe_rf_dir_replay_cnt_waddr,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_wclk,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_wclk_rst_n,
    output  [67:0]  i_hqm_qed_pipe_rf_dir_replay_cnt_wdata,
    output          i_hqm_qed_pipe_rf_dir_replay_cnt_we,
    output  [6:0]   i_hqm_qed_pipe_rf_dir_replay_hp_raddr,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_rclk,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_dir_replay_hp_waddr,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_wclk,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_replay_hp_wdata,
    output          i_hqm_qed_pipe_rf_dir_replay_hp_we,
    output  [6:0]   i_hqm_qed_pipe_rf_dir_replay_tp_raddr,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_rclk,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_dir_replay_tp_waddr,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_wclk,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_replay_tp_wdata,
    output          i_hqm_qed_pipe_rf_dir_replay_tp_we,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_cnt_raddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_rclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_re,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_cnt_waddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_wclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_wclk_rst_n,
    output  [16:0]  i_hqm_qed_pipe_rf_dir_rofrag_cnt_wdata,
    output          i_hqm_qed_pipe_rf_dir_rofrag_cnt_we,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_hp_raddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_rclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_re,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_hp_waddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_wclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_rofrag_hp_wdata,
    output          i_hqm_qed_pipe_rf_dir_rofrag_hp_we,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_tp_raddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_rclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_re,
    output  [8:0]   i_hqm_qed_pipe_rf_dir_rofrag_tp_waddr,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_wclk,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_rofrag_tp_wdata,
    output          i_hqm_qed_pipe_rf_dir_rofrag_tp_we,
    output  [7:0]   i_hqm_qed_pipe_rf_dir_tp_raddr,
    output          i_hqm_qed_pipe_rf_dir_tp_rclk,
    output          i_hqm_qed_pipe_rf_dir_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dir_tp_re,
    output  [7:0]   i_hqm_qed_pipe_rf_dir_tp_waddr,
    output          i_hqm_qed_pipe_rf_dir_tp_wclk,
    output          i_hqm_qed_pipe_rf_dir_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_dir_tp_wdata,
    output          i_hqm_qed_pipe_rf_dir_tp_we,
    output  [4:0]   i_hqm_qed_pipe_rf_dp_dqed_raddr,
    output          i_hqm_qed_pipe_rf_dp_dqed_rclk,
    output          i_hqm_qed_pipe_rf_dp_dqed_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dp_dqed_re,
    output  [4:0]   i_hqm_qed_pipe_rf_dp_dqed_waddr,
    output          i_hqm_qed_pipe_rf_dp_dqed_wclk,
    output          i_hqm_qed_pipe_rf_dp_dqed_wclk_rst_n,
    output  [44:0]  i_hqm_qed_pipe_rf_dp_dqed_wdata,
    output          i_hqm_qed_pipe_rf_dp_dqed_we,
    output  [3:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_dir_raddr,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rclk,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_re,
    output  [3:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_dir_waddr,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wclk,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wdata,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_dir_we,
    output  [3:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_raddr,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rclk,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_re,
    output  [3:0]   i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_waddr,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wclk,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wclk_rst_n,
    output  [22:0]  i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wdata,
    output          i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_we,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_dir_raddr,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rclk,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_re,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_dir_waddr,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wclk,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wclk_rst_n,
    output  [26:0]  i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wdata,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_dir_we,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_raddr,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rclk,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_re,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_waddr,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wclk,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wdata,
    output          i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_we,
    output  [4:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_raddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_re,
    output  [4:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_waddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wdata,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_we,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_raddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_re,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_waddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wdata,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_we,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_raddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_re,
    output  [1:0]   i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_waddr,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wclk,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wclk_rst_n,
    output  [26:0]  i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wdata,
    output          i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_we,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_cnt_raddr,
    output          i_hqm_qed_pipe_rf_nalb_cnt_rclk,
    output          i_hqm_qed_pipe_rf_nalb_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_cnt_re,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_cnt_waddr,
    output          i_hqm_qed_pipe_rf_nalb_cnt_wclk,
    output          i_hqm_qed_pipe_rf_nalb_cnt_wclk_rst_n,
    output  [67:0]  i_hqm_qed_pipe_rf_nalb_cnt_wdata,
    output          i_hqm_qed_pipe_rf_nalb_cnt_we,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_hp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_hp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_hp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_hp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_hp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_hp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_hp_we,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_raddr,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rclk,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_re,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_waddr,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wclk,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wclk_rst_n,
    output  [26:0]  i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wdata,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_we,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_raddr,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rclk,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_re,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_waddr,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wclk,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wclk_rst_n,
    output  [9:0]   i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wdata,
    output          i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_we,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_qed_raddr,
    output          i_hqm_qed_pipe_rf_nalb_qed_rclk,
    output          i_hqm_qed_pipe_rf_nalb_qed_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_qed_re,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_qed_waddr,
    output          i_hqm_qed_pipe_rf_nalb_qed_wclk,
    output          i_hqm_qed_pipe_rf_nalb_qed_wclk_rst_n,
    output  [44:0]  i_hqm_qed_pipe_rf_nalb_qed_wdata,
    output          i_hqm_qed_pipe_rf_nalb_qed_we,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_replay_cnt_raddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_rclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_re,
    output  [4:0]   i_hqm_qed_pipe_rf_nalb_replay_cnt_waddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_wclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_wclk_rst_n,
    output  [67:0]  i_hqm_qed_pipe_rf_nalb_replay_cnt_wdata,
    output          i_hqm_qed_pipe_rf_nalb_replay_cnt_we,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_replay_hp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_replay_hp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_replay_hp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_replay_hp_we,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_replay_tp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_replay_tp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_replay_tp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_replay_tp_we,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_cnt_raddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_re,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_cnt_waddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wclk_rst_n,
    output  [16:0]  i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wdata,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_cnt_we,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_hp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_re,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_hp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_rofrag_hp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_hp_we,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_tp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_re,
    output  [8:0]   i_hqm_qed_pipe_rf_nalb_rofrag_tp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_rofrag_tp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_rofrag_tp_we,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_tp_raddr,
    output          i_hqm_qed_pipe_rf_nalb_tp_rclk,
    output          i_hqm_qed_pipe_rf_nalb_tp_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_nalb_tp_re,
    output  [6:0]   i_hqm_qed_pipe_rf_nalb_tp_waddr,
    output          i_hqm_qed_pipe_rf_nalb_tp_wclk,
    output          i_hqm_qed_pipe_rf_nalb_tp_wclk_rst_n,
    output  [14:0]  i_hqm_qed_pipe_rf_nalb_tp_wdata,
    output          i_hqm_qed_pipe_rf_nalb_tp_we,
    output  [2:0]   i_hqm_qed_pipe_rf_qed_chp_sch_data_raddr,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_rclk,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_re,
    output  [2:0]   i_hqm_qed_pipe_rf_qed_chp_sch_data_waddr,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_wclk,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_wclk_rst_n,
    output  [176:0] i_hqm_qed_pipe_rf_qed_chp_sch_data_wdata,
    output          i_hqm_qed_pipe_rf_qed_chp_sch_data_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_dp_enq_dir_raddr,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_rclk,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_dp_enq_dir_waddr,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_wclk,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rop_dp_enq_dir_wdata,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_dir_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_dp_enq_ro_raddr,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_rclk,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_dp_enq_ro_waddr,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_wclk,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rop_dp_enq_ro_wdata,
    output          i_hqm_qed_pipe_rf_rop_dp_enq_ro_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_nalb_enq_ro_raddr,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rclk,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_nalb_enq_ro_waddr,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wclk,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wdata,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_ro_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_raddr,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rclk,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_waddr,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wclk,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wdata,
    output          i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wclk_rst_n,
    output  [44:0]  i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wclk_rst_n,
    output  [26:0]  i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wclk_rst_n,
    output  [7:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wclk_rst_n,
    output  [26:0]  i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wclk_rst_n,
    output  [44:0]  i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wclk_rst_n,
    output  [99:0]  i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_we,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_raddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rclk_rst_n,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_re,
    output  [1:0]   i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_waddr,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wclk,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wclk_rst_n,
    output  [156:0] i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wdata,
    output          i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_we,
    output  [13:0]  i_hqm_qed_pipe_sr_dir_nxthp_addr,
    output          i_hqm_qed_pipe_sr_dir_nxthp_clk,
    output          i_hqm_qed_pipe_sr_dir_nxthp_clk_rst_n,
    output          i_hqm_qed_pipe_sr_dir_nxthp_re,
    output  [20:0]  i_hqm_qed_pipe_sr_dir_nxthp_wdata,
    output          i_hqm_qed_pipe_sr_dir_nxthp_we,
    output  [13:0]  i_hqm_qed_pipe_sr_nalb_nxthp_addr,
    output          i_hqm_qed_pipe_sr_nalb_nxthp_clk,
    output          i_hqm_qed_pipe_sr_nalb_nxthp_clk_rst_n,
    output          i_hqm_qed_pipe_sr_nalb_nxthp_re,
    output  [20:0]  i_hqm_qed_pipe_sr_nalb_nxthp_wdata,
    output          i_hqm_qed_pipe_sr_nalb_nxthp_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_0_addr,
    output          i_hqm_qed_pipe_sr_qed_0_clk,
    output          i_hqm_qed_pipe_sr_qed_0_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_0_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_0_wdata,
    output          i_hqm_qed_pipe_sr_qed_0_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_1_addr,
    output          i_hqm_qed_pipe_sr_qed_1_clk,
    output          i_hqm_qed_pipe_sr_qed_1_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_1_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_1_wdata,
    output          i_hqm_qed_pipe_sr_qed_1_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_2_addr,
    output          i_hqm_qed_pipe_sr_qed_2_clk,
    output          i_hqm_qed_pipe_sr_qed_2_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_2_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_2_wdata,
    output          i_hqm_qed_pipe_sr_qed_2_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_3_addr,
    output          i_hqm_qed_pipe_sr_qed_3_clk,
    output          i_hqm_qed_pipe_sr_qed_3_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_3_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_3_wdata,
    output          i_hqm_qed_pipe_sr_qed_3_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_4_addr,
    output          i_hqm_qed_pipe_sr_qed_4_clk,
    output          i_hqm_qed_pipe_sr_qed_4_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_4_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_4_wdata,
    output          i_hqm_qed_pipe_sr_qed_4_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_5_addr,
    output          i_hqm_qed_pipe_sr_qed_5_clk,
    output          i_hqm_qed_pipe_sr_qed_5_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_5_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_5_wdata,
    output          i_hqm_qed_pipe_sr_qed_5_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_6_addr,
    output          i_hqm_qed_pipe_sr_qed_6_clk,
    output          i_hqm_qed_pipe_sr_qed_6_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_6_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_6_wdata,
    output          i_hqm_qed_pipe_sr_qed_6_we,
    output  [10:0]  i_hqm_qed_pipe_sr_qed_7_addr,
    output          i_hqm_qed_pipe_sr_qed_7_clk,
    output          i_hqm_qed_pipe_sr_qed_7_clk_rst_n,
    output          i_hqm_qed_pipe_sr_qed_7_re,
    output  [138:0] i_hqm_qed_pipe_sr_qed_7_wdata,
    output          i_hqm_qed_pipe_sr_qed_7_we,
    output  [2:0]   i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_re,
    output  [2:0]   i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wclk_rst_n,
    output  [59:0]  i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_we,
    output  [2:0]   i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_re,
    output  [2:0]   i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wclk_rst_n,
    output  [59:0]  i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_we,
    output  [2:0]   i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_re,
    output  [2:0]   i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wclk_rst_n,
    output  [18:0]  i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_cnt_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_cnt_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_wclk_rst_n,
    output  [15:0]  i_hqm_reorder_pipe_rf_reord_cnt_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_cnt_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_dirhp_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_dirhp_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_wclk_rst_n,
    output  [16:0]  i_hqm_reorder_pipe_rf_reord_dirhp_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_dirhp_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_dirtp_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_dirtp_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_wclk_rst_n,
    output  [16:0]  i_hqm_reorder_pipe_rf_reord_dirtp_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_dirtp_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_lbhp_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_lbhp_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_wclk_rst_n,
    output  [16:0]  i_hqm_reorder_pipe_rf_reord_lbhp_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_lbhp_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_lbtp_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_lbtp_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_wclk_rst_n,
    output  [16:0]  i_hqm_reorder_pipe_rf_reord_lbtp_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_lbtp_mem_we,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_st_mem_raddr,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_rclk,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_re,
    output  [10:0]  i_hqm_reorder_pipe_rf_reord_st_mem_waddr,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_wclk,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_wclk_rst_n,
    output  [24:0]  i_hqm_reorder_pipe_rf_reord_st_mem_wdata,
    output          i_hqm_reorder_pipe_rf_reord_st_mem_we,
    output  [1:0]   i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_re,
    output  [1:0]   i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wclk_rst_n,
    output  [203:0] i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_we,
    output  [3:0]   i_hqm_reorder_pipe_rf_sn0_order_shft_mem_raddr,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rclk,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_re,
    output  [3:0]   i_hqm_reorder_pipe_rf_sn0_order_shft_mem_waddr,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wclk,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wclk_rst_n,
    output  [11:0]  i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wdata,
    output          i_hqm_reorder_pipe_rf_sn0_order_shft_mem_we,
    output  [3:0]   i_hqm_reorder_pipe_rf_sn1_order_shft_mem_raddr,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rclk,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_re,
    output  [3:0]   i_hqm_reorder_pipe_rf_sn1_order_shft_mem_waddr,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wclk,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wclk_rst_n,
    output  [11:0]  i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wdata,
    output          i_hqm_reorder_pipe_rf_sn1_order_shft_mem_we,
    output  [1:0]   i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_re,
    output  [1:0]   i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wclk_rst_n,
    output  [20:0]  i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_we,
    output  [4:0]   i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_raddr,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rclk,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rclk_rst_n,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_re,
    output  [4:0]   i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_waddr,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wclk,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wclk_rst_n,
    output  [12:0]  i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wdata,
    output          i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_we,
    output  [1:0]   i_hqm_reorder_pipe_rop_cfg_req_down_1_0,
    output  [1:0]   i_hqm_reorder_pipe_rop_cfg_rsp_down_5_4,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd0_raddr,
    output          i_hqm_system_rf_alarm_vf_synd0_rclk,
    output          i_hqm_system_rf_alarm_vf_synd0_rclk_rst_n,
    output          i_hqm_system_rf_alarm_vf_synd0_re,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd0_waddr,
    output          i_hqm_system_rf_alarm_vf_synd0_wclk,
    output          i_hqm_system_rf_alarm_vf_synd0_wclk_rst_n,
    output  [29:0]  i_hqm_system_rf_alarm_vf_synd0_wdata,
    output          i_hqm_system_rf_alarm_vf_synd0_we,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd1_raddr,
    output          i_hqm_system_rf_alarm_vf_synd1_rclk,
    output          i_hqm_system_rf_alarm_vf_synd1_rclk_rst_n,
    output          i_hqm_system_rf_alarm_vf_synd1_re,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd1_waddr,
    output          i_hqm_system_rf_alarm_vf_synd1_wclk,
    output          i_hqm_system_rf_alarm_vf_synd1_wclk_rst_n,
    output  [31:0]  i_hqm_system_rf_alarm_vf_synd1_wdata,
    output          i_hqm_system_rf_alarm_vf_synd1_we,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd2_raddr,
    output          i_hqm_system_rf_alarm_vf_synd2_rclk,
    output          i_hqm_system_rf_alarm_vf_synd2_rclk_rst_n,
    output          i_hqm_system_rf_alarm_vf_synd2_re,
    output  [3:0]   i_hqm_system_rf_alarm_vf_synd2_waddr,
    output          i_hqm_system_rf_alarm_vf_synd2_wclk,
    output          i_hqm_system_rf_alarm_vf_synd2_wclk_rst_n,
    output  [31:0]  i_hqm_system_rf_alarm_vf_synd2_wdata,
    output          i_hqm_system_rf_alarm_vf_synd2_we,
    output  [5:0]   i_hqm_system_rf_dir_wb0_raddr,
    output          i_hqm_system_rf_dir_wb0_rclk,
    output          i_hqm_system_rf_dir_wb0_rclk_rst_n,
    output          i_hqm_system_rf_dir_wb0_re,
    output  [5:0]   i_hqm_system_rf_dir_wb0_waddr,
    output          i_hqm_system_rf_dir_wb0_wclk,
    output          i_hqm_system_rf_dir_wb0_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_dir_wb0_wdata,
    output          i_hqm_system_rf_dir_wb0_we,
    output  [5:0]   i_hqm_system_rf_dir_wb1_raddr,
    output          i_hqm_system_rf_dir_wb1_rclk,
    output          i_hqm_system_rf_dir_wb1_rclk_rst_n,
    output          i_hqm_system_rf_dir_wb1_re,
    output  [5:0]   i_hqm_system_rf_dir_wb1_waddr,
    output          i_hqm_system_rf_dir_wb1_wclk,
    output          i_hqm_system_rf_dir_wb1_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_dir_wb1_wdata,
    output          i_hqm_system_rf_dir_wb1_we,
    output  [5:0]   i_hqm_system_rf_dir_wb2_raddr,
    output          i_hqm_system_rf_dir_wb2_rclk,
    output          i_hqm_system_rf_dir_wb2_rclk_rst_n,
    output          i_hqm_system_rf_dir_wb2_re,
    output  [5:0]   i_hqm_system_rf_dir_wb2_waddr,
    output          i_hqm_system_rf_dir_wb2_wclk,
    output          i_hqm_system_rf_dir_wb2_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_dir_wb2_wdata,
    output          i_hqm_system_rf_dir_wb2_we,
    output  [7:0]   i_hqm_system_rf_hcw_enq_fifo_raddr,
    output          i_hqm_system_rf_hcw_enq_fifo_rclk,
    output          i_hqm_system_rf_hcw_enq_fifo_rclk_rst_n,
    output          i_hqm_system_rf_hcw_enq_fifo_re,
    output  [7:0]   i_hqm_system_rf_hcw_enq_fifo_waddr,
    output          i_hqm_system_rf_hcw_enq_fifo_wclk,
    output          i_hqm_system_rf_hcw_enq_fifo_wclk_rst_n,
    output  [166:0] i_hqm_system_rf_hcw_enq_fifo_wdata,
    output          i_hqm_system_rf_hcw_enq_fifo_we,
    output  [5:0]   i_hqm_system_rf_ldb_wb0_raddr,
    output          i_hqm_system_rf_ldb_wb0_rclk,
    output          i_hqm_system_rf_ldb_wb0_rclk_rst_n,
    output          i_hqm_system_rf_ldb_wb0_re,
    output  [5:0]   i_hqm_system_rf_ldb_wb0_waddr,
    output          i_hqm_system_rf_ldb_wb0_wclk,
    output          i_hqm_system_rf_ldb_wb0_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_ldb_wb0_wdata,
    output          i_hqm_system_rf_ldb_wb0_we,
    output  [5:0]   i_hqm_system_rf_ldb_wb1_raddr,
    output          i_hqm_system_rf_ldb_wb1_rclk,
    output          i_hqm_system_rf_ldb_wb1_rclk_rst_n,
    output          i_hqm_system_rf_ldb_wb1_re,
    output  [5:0]   i_hqm_system_rf_ldb_wb1_waddr,
    output          i_hqm_system_rf_ldb_wb1_wclk,
    output          i_hqm_system_rf_ldb_wb1_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_ldb_wb1_wdata,
    output          i_hqm_system_rf_ldb_wb1_we,
    output  [5:0]   i_hqm_system_rf_ldb_wb2_raddr,
    output          i_hqm_system_rf_ldb_wb2_rclk,
    output          i_hqm_system_rf_ldb_wb2_rclk_rst_n,
    output          i_hqm_system_rf_ldb_wb2_re,
    output  [5:0]   i_hqm_system_rf_ldb_wb2_waddr,
    output          i_hqm_system_rf_ldb_wb2_wclk,
    output          i_hqm_system_rf_ldb_wb2_wclk_rst_n,
    output  [143:0] i_hqm_system_rf_ldb_wb2_wdata,
    output          i_hqm_system_rf_ldb_wb2_we,
    output  [4:0]   i_hqm_system_rf_lut_dir_cq2vf_pf_ro_raddr,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rclk,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_re,
    output  [4:0]   i_hqm_system_rf_lut_dir_cq2vf_pf_ro_waddr,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wclk,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wclk_rst_n,
    output  [12:0]  i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wdata,
    output          i_hqm_system_rf_lut_dir_cq2vf_pf_ro_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_addr_l_raddr,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_rclk,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_addr_l_waddr,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_wclk,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_wclk_rst_n,
    output  [26:0]  i_hqm_system_rf_lut_dir_cq_addr_l_wdata,
    output          i_hqm_system_rf_lut_dir_cq_addr_l_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_addr_u_raddr,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_rclk,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_addr_u_waddr,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_wclk,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_dir_cq_addr_u_wdata,
    output          i_hqm_system_rf_lut_dir_cq_addr_u_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_addr_l_raddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_rclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_addr_l_waddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_wclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_wclk_rst_n,
    output  [30:0]  i_hqm_system_rf_lut_dir_cq_ai_addr_l_wdata,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_l_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_addr_u_raddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_rclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_addr_u_waddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_wclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_dir_cq_ai_addr_u_wdata,
    output          i_hqm_system_rf_lut_dir_cq_ai_addr_u_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_data_raddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_rclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_ai_data_waddr,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_wclk,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_dir_cq_ai_data_wdata,
    output          i_hqm_system_rf_lut_dir_cq_ai_data_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_isr_raddr,
    output          i_hqm_system_rf_lut_dir_cq_isr_rclk,
    output          i_hqm_system_rf_lut_dir_cq_isr_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_isr_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_isr_waddr,
    output          i_hqm_system_rf_lut_dir_cq_isr_wclk,
    output          i_hqm_system_rf_lut_dir_cq_isr_wclk_rst_n,
    output  [12:0]  i_hqm_system_rf_lut_dir_cq_isr_wdata,
    output          i_hqm_system_rf_lut_dir_cq_isr_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_pasid_raddr,
    output          i_hqm_system_rf_lut_dir_cq_pasid_rclk,
    output          i_hqm_system_rf_lut_dir_cq_pasid_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_cq_pasid_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_cq_pasid_waddr,
    output          i_hqm_system_rf_lut_dir_cq_pasid_wclk,
    output          i_hqm_system_rf_lut_dir_cq_pasid_wclk_rst_n,
    output  [23:0]  i_hqm_system_rf_lut_dir_cq_pasid_wdata,
    output          i_hqm_system_rf_lut_dir_cq_pasid_we,
    output  [4:0]   i_hqm_system_rf_lut_dir_pp2vas_raddr,
    output          i_hqm_system_rf_lut_dir_pp2vas_rclk,
    output          i_hqm_system_rf_lut_dir_pp2vas_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_pp2vas_re,
    output  [4:0]   i_hqm_system_rf_lut_dir_pp2vas_waddr,
    output          i_hqm_system_rf_lut_dir_pp2vas_wclk,
    output          i_hqm_system_rf_lut_dir_pp2vas_wclk_rst_n,
    output  [10:0]  i_hqm_system_rf_lut_dir_pp2vas_wdata,
    output          i_hqm_system_rf_lut_dir_pp2vas_we,
    output  [1:0]   i_hqm_system_rf_lut_dir_pp_v_raddr,
    output          i_hqm_system_rf_lut_dir_pp_v_rclk,
    output          i_hqm_system_rf_lut_dir_pp_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_pp_v_re,
    output  [1:0]   i_hqm_system_rf_lut_dir_pp_v_waddr,
    output          i_hqm_system_rf_lut_dir_pp_v_wclk,
    output          i_hqm_system_rf_lut_dir_pp_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_dir_pp_v_wdata,
    output          i_hqm_system_rf_lut_dir_pp_v_we,
    output  [5:0]   i_hqm_system_rf_lut_dir_vasqid_v_raddr,
    output          i_hqm_system_rf_lut_dir_vasqid_v_rclk,
    output          i_hqm_system_rf_lut_dir_vasqid_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_dir_vasqid_v_re,
    output  [5:0]   i_hqm_system_rf_lut_dir_vasqid_v_waddr,
    output          i_hqm_system_rf_lut_dir_vasqid_v_wclk,
    output          i_hqm_system_rf_lut_dir_vasqid_v_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_dir_vasqid_v_wdata,
    output          i_hqm_system_rf_lut_dir_vasqid_v_we,
    output  [4:0]   i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_raddr,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rclk,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_re,
    output  [4:0]   i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_waddr,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wclk,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wclk_rst_n,
    output  [12:0]  i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wdata,
    output          i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_addr_l_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_addr_l_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_wclk_rst_n,
    output  [26:0]  i_hqm_system_rf_lut_ldb_cq_addr_l_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_addr_l_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_addr_u_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_addr_u_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_ldb_cq_addr_u_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_addr_u_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_addr_l_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_addr_l_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wclk_rst_n,
    output  [30:0]  i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_l_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_addr_u_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_addr_u_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_ai_addr_u_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_data_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_ai_data_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_lut_ldb_cq_ai_data_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_ai_data_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_isr_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_isr_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_isr_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_isr_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_isr_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_isr_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_isr_wclk_rst_n,
    output  [12:0]  i_hqm_system_rf_lut_ldb_cq_isr_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_isr_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_pasid_raddr,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_rclk,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_cq_pasid_waddr,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_wclk,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_wclk_rst_n,
    output  [23:0]  i_hqm_system_rf_lut_ldb_cq_pasid_wdata,
    output          i_hqm_system_rf_lut_ldb_cq_pasid_we,
    output  [4:0]   i_hqm_system_rf_lut_ldb_pp2vas_raddr,
    output          i_hqm_system_rf_lut_ldb_pp2vas_rclk,
    output          i_hqm_system_rf_lut_ldb_pp2vas_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_pp2vas_re,
    output  [4:0]   i_hqm_system_rf_lut_ldb_pp2vas_waddr,
    output          i_hqm_system_rf_lut_ldb_pp2vas_wclk,
    output          i_hqm_system_rf_lut_ldb_pp2vas_wclk_rst_n,
    output  [10:0]  i_hqm_system_rf_lut_ldb_pp2vas_wdata,
    output          i_hqm_system_rf_lut_ldb_pp2vas_we,
    output  [2:0]   i_hqm_system_rf_lut_ldb_qid2vqid_raddr,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_rclk,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_re,
    output  [2:0]   i_hqm_system_rf_lut_ldb_qid2vqid_waddr,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_wclk,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_wclk_rst_n,
    output  [20:0]  i_hqm_system_rf_lut_ldb_qid2vqid_wdata,
    output          i_hqm_system_rf_lut_ldb_qid2vqid_we,
    output  [5:0]   i_hqm_system_rf_lut_ldb_vasqid_v_raddr,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_rclk,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_re,
    output  [5:0]   i_hqm_system_rf_lut_ldb_vasqid_v_waddr,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_wclk,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_ldb_vasqid_v_wdata,
    output          i_hqm_system_rf_lut_ldb_vasqid_v_we,
    output  [7:0]   i_hqm_system_rf_lut_vf_dir_vpp2pp_raddr,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_rclk,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_re,
    output  [7:0]   i_hqm_system_rf_lut_vf_dir_vpp2pp_waddr,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_wclk,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_wclk_rst_n,
    output  [30:0]  i_hqm_system_rf_lut_vf_dir_vpp2pp_wdata,
    output          i_hqm_system_rf_lut_vf_dir_vpp2pp_we,
    output  [5:0]   i_hqm_system_rf_lut_vf_dir_vpp_v_raddr,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_rclk,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_re,
    output  [5:0]   i_hqm_system_rf_lut_vf_dir_vpp_v_waddr,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_wclk,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_vf_dir_vpp_v_wdata,
    output          i_hqm_system_rf_lut_vf_dir_vpp_v_we,
    output  [7:0]   i_hqm_system_rf_lut_vf_dir_vqid2qid_raddr,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_rclk,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_re,
    output  [7:0]   i_hqm_system_rf_lut_vf_dir_vqid2qid_waddr,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_wclk,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_wclk_rst_n,
    output  [30:0]  i_hqm_system_rf_lut_vf_dir_vqid2qid_wdata,
    output          i_hqm_system_rf_lut_vf_dir_vqid2qid_we,
    output  [5:0]   i_hqm_system_rf_lut_vf_dir_vqid_v_raddr,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_rclk,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_re,
    output  [5:0]   i_hqm_system_rf_lut_vf_dir_vqid_v_waddr,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_wclk,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_vf_dir_vqid_v_wdata,
    output          i_hqm_system_rf_lut_vf_dir_vqid_v_we,
    output  [7:0]   i_hqm_system_rf_lut_vf_ldb_vpp2pp_raddr,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_rclk,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_re,
    output  [7:0]   i_hqm_system_rf_lut_vf_ldb_vpp2pp_waddr,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_wclk,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_wclk_rst_n,
    output  [24:0]  i_hqm_system_rf_lut_vf_ldb_vpp2pp_wdata,
    output          i_hqm_system_rf_lut_vf_ldb_vpp2pp_we,
    output  [5:0]   i_hqm_system_rf_lut_vf_ldb_vpp_v_raddr,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_rclk,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_re,
    output  [5:0]   i_hqm_system_rf_lut_vf_ldb_vpp_v_waddr,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_wclk,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_vf_ldb_vpp_v_wdata,
    output          i_hqm_system_rf_lut_vf_ldb_vpp_v_we,
    output  [6:0]   i_hqm_system_rf_lut_vf_ldb_vqid2qid_raddr,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_rclk,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_re,
    output  [6:0]   i_hqm_system_rf_lut_vf_ldb_vqid2qid_waddr,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_wclk,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_wclk_rst_n,
    output  [26:0]  i_hqm_system_rf_lut_vf_ldb_vqid2qid_wdata,
    output          i_hqm_system_rf_lut_vf_ldb_vqid2qid_we,
    output  [4:0]   i_hqm_system_rf_lut_vf_ldb_vqid_v_raddr,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_rclk,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_rclk_rst_n,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_re,
    output  [4:0]   i_hqm_system_rf_lut_vf_ldb_vqid_v_waddr,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_wclk,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_wclk_rst_n,
    output  [16:0]  i_hqm_system_rf_lut_vf_ldb_vqid_v_wdata,
    output          i_hqm_system_rf_lut_vf_ldb_vqid_v_we,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word0_raddr,
    output          i_hqm_system_rf_msix_tbl_word0_rclk,
    output          i_hqm_system_rf_msix_tbl_word0_rclk_rst_n,
    output          i_hqm_system_rf_msix_tbl_word0_re,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word0_waddr,
    output          i_hqm_system_rf_msix_tbl_word0_wclk,
    output          i_hqm_system_rf_msix_tbl_word0_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_msix_tbl_word0_wdata,
    output          i_hqm_system_rf_msix_tbl_word0_we,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word1_raddr,
    output          i_hqm_system_rf_msix_tbl_word1_rclk,
    output          i_hqm_system_rf_msix_tbl_word1_rclk_rst_n,
    output          i_hqm_system_rf_msix_tbl_word1_re,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word1_waddr,
    output          i_hqm_system_rf_msix_tbl_word1_wclk,
    output          i_hqm_system_rf_msix_tbl_word1_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_msix_tbl_word1_wdata,
    output          i_hqm_system_rf_msix_tbl_word1_we,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word2_raddr,
    output          i_hqm_system_rf_msix_tbl_word2_rclk,
    output          i_hqm_system_rf_msix_tbl_word2_rclk_rst_n,
    output          i_hqm_system_rf_msix_tbl_word2_re,
    output  [5:0]   i_hqm_system_rf_msix_tbl_word2_waddr,
    output          i_hqm_system_rf_msix_tbl_word2_wclk,
    output          i_hqm_system_rf_msix_tbl_word2_wclk_rst_n,
    output  [32:0]  i_hqm_system_rf_msix_tbl_word2_wdata,
    output          i_hqm_system_rf_msix_tbl_word2_we,
    output  [6:0]   i_hqm_system_rf_sch_out_fifo_raddr,
    output          i_hqm_system_rf_sch_out_fifo_rclk,
    output          i_hqm_system_rf_sch_out_fifo_rclk_rst_n,
    output          i_hqm_system_rf_sch_out_fifo_re,
    output  [6:0]   i_hqm_system_rf_sch_out_fifo_waddr,
    output          i_hqm_system_rf_sch_out_fifo_wclk,
    output          i_hqm_system_rf_sch_out_fifo_wclk_rst_n,
    output  [269:0] i_hqm_system_rf_sch_out_fifo_wdata,
    output          i_hqm_system_rf_sch_out_fifo_we,
    output  [10:0]  i_hqm_system_sr_rob_mem_addr,
    output          i_hqm_system_sr_rob_mem_clk,
    output          i_hqm_system_sr_rob_mem_clk_rst_n,
    output          i_hqm_system_sr_rob_mem_re,
    output  [155:0] i_hqm_system_sr_rob_mem_wdata,
    output          i_hqm_system_sr_rob_mem_we,
    output  [1:0]   i_hqm_system_system_cfg_req_down_1_0,
    output  [1:0]   i_hqm_system_system_cfg_rsp_down_5_4,
    output          lsp_reset_done,
    output          lsp_unit_idle,
    output          lsp_unit_pipeidle,
    output          nalb_reset_done,
    output          nalb_unit_idle,
    output          nalb_unit_pipeidle,
    output          qed_reset_done,
    output          qed_unit_idle,
    output          qed_unit_pipeidle,
    output          rop_reset_done,
    output          rop_unit_pipeidle,
    output          sif_alarm_ready,
    output          system_idle,
    output          system_reset_done,
    output          visa_str_chp_lsp_cmp_data,
    output          wd_clkreq,
    output  [638:0] write_buffer_mstr,
    output          write_buffer_mstr_v
);

   wire [24:0]  ap_alarm_down_data;
   wire [44:0]  ap_aqed_data;
   wire [92:0]  ap_cfg_req_down;
   wire [38:0]  ap_cfg_rsp_down;
   wire [24:0]  aqed_alarm_down_data;
   wire [23:0]  aqed_ap_enq_data;
   wire [178:0] aqed_chp_sch_data;
   wire         aqed_clk_enable;
   wire         aqed_clk_idle;
   wire         aqed_lsp_dec_fid_cnt_v;
   wire [8:0]   aqed_lsp_deq_data;
   wire         aqed_lsp_deq_v;
   wire [6:0]   aqed_lsp_fid_cnt_upd_qid;
   wire         aqed_lsp_fid_cnt_upd_v;
   wire         aqed_lsp_fid_cnt_upd_val;
   wire [34:0]  aqed_lsp_sch_data;
   wire         aqed_lsp_stop_atqatm;
   wire [92:0]  chp_cfg_req_down;
   wire [38:0]  chp_cfg_rsp_down;
   wire [72:0]  chp_lsp_cmp_data;
   wire [63:0]  chp_lsp_ldb_cq_off;
   wire [28:0]  chp_lsp_token_data;
   wire [200:0] chp_rop_hcw_data;
   wire [7:0]   dp_lsp_enq_dir_data;
   wire [22:0]  dp_lsp_enq_rorply_data;
   wire [155:0] hcw_enq_w_req;
   wire [158:0] hcw_sched_w_req;
   wire [24:0]  hqm_alarm_data;
   wire         hqm_clk_rptr_rst_sync_b;
   wire         hqm_clk_rptr_rst_sync_bx;
   wire         hqm_clk_rptr_rst_sync_bxx;
   wire         hqm_clk_ungate_rptr;
   wire         hqm_clk_ungate_rptrx;
   wire         hqm_clk_ungate_rptrxx;
   wire         hqm_flr_prep_b;
   wire         hqm_flr_prep_rptr;
   wire         hqm_flr_prep_rptrx;
   wire         hqm_flr_prep_rptrxx;
   wire         hqm_gated_clk_chp;
   wire         hqm_gated_clk_dir;
   wire [0:0]   hqm_gated_clk_enable_and_chp;
   wire [0:0]   hqm_gated_clk_enable_and_dir;
   wire [0:0]   hqm_gated_clk_enable_and_lsp;
   wire [0:0]   hqm_gated_clk_enable_and_nalb;
   wire [0:0]   hqm_gated_clk_enable_and_qed;
   wire [0:0]   hqm_gated_clk_enable_and_sys;
   wire         hqm_gated_clk_enable_rptr_chp;
   wire         hqm_gated_clk_enable_rptr_dir;
   wire         hqm_gated_clk_enable_rptr_lsp;
   wire         hqm_gated_clk_enable_rptr_nalb;
   wire         hqm_gated_clk_enable_rptr_qed;
   wire         hqm_gated_clk_enable_rptr_sys;
   wire         hqm_gated_clk_lsp;
   wire         hqm_gated_clk_nalb;
   wire         hqm_gated_clk_qed;
   wire         hqm_gated_clk_sys;
   wire [0:0]   hqm_gated_local_clk_en_chp;
   wire [0:0]   hqm_gated_local_clk_en_dir;
   wire [0:0]   hqm_gated_local_clk_en_lsp;
   wire [0:0]   hqm_gated_local_clk_en_nalb;
   wire [0:0]   hqm_gated_local_clk_en_qed;
   wire [0:0]   hqm_gated_local_clk_en_sys;
   wire         hqm_gated_rst_b_active_aqed;
   wire         hqm_gated_rst_b_active_atm;
   wire         hqm_gated_rst_b_active_chp;
   wire         hqm_gated_rst_b_active_dir;
   wire         hqm_gated_rst_b_active_lsp;
   wire         hqm_gated_rst_b_active_nalb;
   wire         hqm_gated_rst_b_active_qed;
   wire         hqm_gated_rst_b_active_rop;
   wire         hqm_gated_rst_b_active_sys;
   wire [0:0]   hqm_gated_rst_b_aqed;
   wire [0:0]   hqm_gated_rst_b_atm;
   wire [0:0]   hqm_gated_rst_b_chp;
   wire [0:0]   hqm_gated_rst_b_dir;
   wire         hqm_gated_rst_b_done_aqed;
   wire         hqm_gated_rst_b_done_atm;
   wire         hqm_gated_rst_b_done_chp;
   wire         hqm_gated_rst_b_done_dir;
   wire         hqm_gated_rst_b_done_lsp;
   wire         hqm_gated_rst_b_done_nalb;
   wire         hqm_gated_rst_b_done_qed;
   wire         hqm_gated_rst_b_done_rop;
   wire         hqm_gated_rst_b_done_sys;
   wire [0:0]   hqm_gated_rst_b_lsp;
   wire [0:0]   hqm_gated_rst_b_nalb;
   wire         hqm_gated_rst_b_pgcb_sync_chp;
   wire [0:0]   hqm_gated_rst_b_qed;
   wire [0:0]   hqm_gated_rst_b_rop;
   wire         hqm_gated_rst_b_start_aqed;
   wire         hqm_gated_rst_b_start_atm;
   wire         hqm_gated_rst_b_start_chp;
   wire         hqm_gated_rst_b_start_dir;
   wire         hqm_gated_rst_b_start_lsp;
   wire         hqm_gated_rst_b_start_nalb;
   wire         hqm_gated_rst_b_start_qed;
   wire         hqm_gated_rst_b_start_rop;
   wire         hqm_gated_rst_b_start_sys;
   wire [0:0]   hqm_gated_rst_b_sys;
   wire         hqm_inp_gated_clk;
   wire         hqm_inp_gated_clk_enable_rptr;
   wire         hqm_inp_gated_clk_enable_rptrx;
   wire         hqm_inp_gated_clk_enable_rptrxx;
   wire         hqm_inp_gated_clkx;
   wire         hqm_inp_gated_clkxx;
   wire [0:0]   hqm_inp_gated_rst_b_aqed;
   wire [0:0]   hqm_inp_gated_rst_b_atm;
   wire [0:0]   hqm_inp_gated_rst_b_chp;
   wire [0:0]   hqm_inp_gated_rst_b_dir;
   wire [0:0]   hqm_inp_gated_rst_b_lsp;
   wire [0:0]   hqm_inp_gated_rst_b_nalb;
   wire [0:0]   hqm_inp_gated_rst_b_qed;
   wire [0:0]   hqm_inp_gated_rst_b_rop;
   wire [0:0]   hqm_inp_gated_rst_b_sys;
   wire [0:0]   hqm_pgcb_rst_b_chp;
   wire         hqm_pgcb_rst_b_start_chp;
   wire         hqm_proc_clk_en_qed_local;
   wire         hqm_rst_prep_aqed;
   wire         hqm_rst_prep_atm;
   wire         hqm_rst_prep_chp;
   wire         hqm_rst_prep_dir;
   wire         hqm_rst_prep_lsp;
   wire         hqm_rst_prep_nalb;
   wire         hqm_rst_prep_qed;
   wire         hqm_rst_prep_rop;
   wire         hqm_rst_prep_sys;
   wire         i_hqm_aqed_pipe_ap_aqed_ready;
   wire         i_hqm_aqed_pipe_aqed_alarm_down_v;
   wire         i_hqm_aqed_pipe_aqed_ap_enq_v;
   wire         i_hqm_aqed_pipe_aqed_chp_sch_v;
   wire         i_hqm_aqed_pipe_aqed_lsp_sch_v;
   wire         i_hqm_aqed_pipe_aqed_unit_idle;
   wire         i_hqm_aqed_pipe_qed_aqed_enq_ready;
   wire         i_hqm_credit_hist_pipe_aqed_chp_sch_ready;
   wire         i_hqm_credit_hist_pipe_chp_alarm_down_v;
   wire         i_hqm_credit_hist_pipe_chp_alarm_up_ready;
   wire         i_hqm_credit_hist_pipe_chp_cfg_req_down_read;
   wire         i_hqm_credit_hist_pipe_chp_cfg_req_down_write;
   wire         i_hqm_credit_hist_pipe_chp_cfg_rsp_down_ack;
   wire         i_hqm_credit_hist_pipe_chp_lsp_cmp_v;
   wire         i_hqm_credit_hist_pipe_chp_lsp_token_v;
   wire         i_hqm_credit_hist_pipe_chp_rop_hcw_v;
   wire         i_hqm_credit_hist_pipe_cwdi_interrupt_w_req_valid;
   wire         i_hqm_credit_hist_pipe_hcw_enq_w_req_ready;
   wire         i_hqm_credit_hist_pipe_hcw_sched_w_req_valid;
   wire         i_hqm_credit_hist_pipe_hqm_proc_clk_en_chp;
   wire         i_hqm_credit_hist_pipe_interrupt_w_req_valid;
   wire         i_hqm_credit_hist_pipe_qed_chp_sch_ready;
   wire         i_hqm_list_sel_pipe_ap_alarm_down_v;
   wire         i_hqm_list_sel_pipe_ap_alarm_up_ready;
   wire         i_hqm_list_sel_pipe_ap_aqed_v;
   wire         i_hqm_list_sel_pipe_ap_cfg_req_down_read;
   wire         i_hqm_list_sel_pipe_ap_cfg_req_down_write;
   wire         i_hqm_list_sel_pipe_ap_cfg_rsp_down_ack;
   wire         i_hqm_list_sel_pipe_aqed_ap_enq_ready;
   wire         i_hqm_list_sel_pipe_aqed_lsp_sch_ready;
   wire         i_hqm_list_sel_pipe_chp_lsp_cmp_ready;
   wire         i_hqm_list_sel_pipe_chp_lsp_token_ready;
   wire         i_hqm_list_sel_pipe_dp_lsp_enq_dir_ready;
   wire         i_hqm_list_sel_pipe_dp_lsp_enq_rorply_ready;
   wire         i_hqm_list_sel_pipe_hqm_proc_clk_en_lsp;
   wire         i_hqm_list_sel_pipe_lsp_alarm_down_v;
   wire         i_hqm_list_sel_pipe_lsp_alarm_up_ready;
   wire         i_hqm_list_sel_pipe_lsp_cfg_req_down_read;
   wire         i_hqm_list_sel_pipe_lsp_cfg_req_down_write;
   wire         i_hqm_list_sel_pipe_lsp_cfg_rsp_down_ack;
   wire         i_hqm_list_sel_pipe_lsp_dp_sch_dir_v;
   wire         i_hqm_list_sel_pipe_lsp_dp_sch_rorply_v;
   wire         i_hqm_list_sel_pipe_lsp_nalb_sch_atq_v;
   wire         i_hqm_list_sel_pipe_lsp_nalb_sch_rorply_v;
   wire         i_hqm_list_sel_pipe_lsp_nalb_sch_unoord_v;
   wire         i_hqm_list_sel_pipe_nalb_lsp_enq_lb_ready;
   wire         i_hqm_list_sel_pipe_nalb_lsp_enq_rorply_ready;
   wire         i_hqm_list_sel_pipe_rop_lsp_reordercmp_ready;
   wire         i_hqm_qed_pipe_dp_lsp_enq_dir_v;
   wire         i_hqm_qed_pipe_dp_lsp_enq_rorply_v;
   wire         i_hqm_qed_pipe_hqm_proc_clk_en_dir;
   wire         i_hqm_qed_pipe_hqm_proc_clk_en_nalb;
   wire         i_hqm_qed_pipe_lsp_dp_sch_dir_ready;
   wire         i_hqm_qed_pipe_lsp_dp_sch_rorply_ready;
   wire         i_hqm_qed_pipe_lsp_nalb_sch_atq_ready;
   wire         i_hqm_qed_pipe_lsp_nalb_sch_rorply_ready;
   wire         i_hqm_qed_pipe_lsp_nalb_sch_unoord_ready;
   wire         i_hqm_qed_pipe_nalb_lsp_enq_lb_v;
   wire         i_hqm_qed_pipe_nalb_lsp_enq_rorply_v;
   wire         i_hqm_qed_pipe_qed_alarm_down_v;
   wire         i_hqm_qed_pipe_qed_alarm_up_ready;
   wire         i_hqm_qed_pipe_qed_aqed_enq_v;
   wire         i_hqm_qed_pipe_qed_cfg_req_down_read;
   wire         i_hqm_qed_pipe_qed_cfg_req_down_write;
   wire         i_hqm_qed_pipe_qed_cfg_rsp_down_ack;
   wire         i_hqm_qed_pipe_qed_chp_sch_v;
   wire         i_hqm_qed_pipe_rop_dp_enq_ready;
   wire         i_hqm_qed_pipe_rop_dqed_enq_ready;
   wire         i_hqm_qed_pipe_rop_nalb_enq_ready;
   wire         i_hqm_qed_pipe_rop_qed_enq_ready;
   wire         i_hqm_reorder_pipe_chp_rop_hcw_ready;
   wire         i_hqm_reorder_pipe_rop_alarm_down_v;
   wire         i_hqm_reorder_pipe_rop_alarm_up_ready;
   wire         i_hqm_reorder_pipe_rop_cfg_req_down_read;
   wire         i_hqm_reorder_pipe_rop_cfg_req_down_write;
   wire         i_hqm_reorder_pipe_rop_cfg_rsp_down_ack;
   wire         i_hqm_reorder_pipe_rop_dp_enq_v;
   wire         i_hqm_reorder_pipe_rop_lsp_reordercmp_v;
   wire         i_hqm_reorder_pipe_rop_nalb_enq_v;
   wire         i_hqm_reorder_pipe_rop_qed_dqed_enq_v;
   wire         i_hqm_reorder_pipe_rop_qed_force_clockon;
   wire         i_hqm_reorder_pipe_rop_unit_idle;
   wire         i_hqm_system_cwdi_interrupt_w_req_ready;
   wire         i_hqm_system_hcw_enq_w_req_valid;
   wire         i_hqm_system_hcw_sched_w_req_ready;
   wire         i_hqm_system_hqm_alarm_ready;
   wire         i_hqm_system_hqm_proc_clk_en_sys;
   wire         i_hqm_system_interrupt_w_req_ready;
   wire         i_hqm_system_system_cfg_req_down_read;
   wire         i_hqm_system_system_cfg_req_down_write;
   wire         i_hqm_system_system_cfg_rsp_down_ack;
   wire [8:0]   interrupt_w_req;
   wire [24:0]  lsp_alarm_down_data;
   wire [36:0]  lsp_aqed_cmp_data;
   wire         lsp_aqed_cmp_ready;
   wire         lsp_aqed_cmp_v;
   wire [92:0]  lsp_cfg_req_down;
   wire [38:0]  lsp_cfg_rsp_down;
   wire [26:0]  lsp_dp_sch_dir_data;
   wire [7:0]   lsp_dp_sch_rorply_data;
   wire [7:0]   lsp_nalb_sch_atq_data;
   wire [7:0]   lsp_nalb_sch_rorply_data;
   wire [26:0]  lsp_nalb_sch_unoord_data;
   wire [9:0]   nalb_lsp_enq_lb_data;
   wire [26:0]  nalb_lsp_enq_rorply_data;
   wire         pgcb_clkx;
   wire         prim_clk_enable_rptr;
   wire         prim_clk_ungate_rptr_sys;
   wire         prim_gated_clk;
   wire [24:0]  qed_alarm_down_data;
   wire [138:0] qed_aqed_enq_data;
   wire [92:0]  qed_cfg_req_down;
   wire [38:0]  qed_cfg_rsp_down;
   wire [176:0] qed_chp_sch_data;
   wire [8:0]   qed_lsp_deq_data;
   wire         qed_lsp_deq_v;
   wire         qed_unit_idle_local;
   wire [0:0]   qed_unit_idle_qual;
   wire [24:0]  rop_alarm_down_data;
   wire [92:0]  rop_cfg_req_down;
   wire [38:0]  rop_cfg_rsp_down;
   wire         rop_clk_enable;
   wire         rop_clk_idle;
   wire [99:0]  rop_dp_enq_data;
   wire [16:0]  rop_lsp_reordercmp_data;
   wire [99:0]  rop_nalb_enq_data;
   wire [156:0] rop_qed_dqed_enq_data;
   wire         side_rst_sync_prim_n;
   wire [1:0]   spare_lsp_qed;
   wire [1:0]   spare_lsp_sys;
   wire [1:0]   spare_qed_lsp;
   wire [1:0]   spare_qed_sys;
   wire [1:0]   spare_sys_lsp;
   wire [1:0]   spare_sys_qed;
   wire [92:0]  system_cfg_req_down;
   wire [38:0]  system_cfg_rsp_down;

   hqm_aqed_pipe i_hqm_aqed_pipe
      (.hqm_gated_clk                            (hqm_gated_clk_lsp),
       .hqm_inp_gated_clk,
       .hqm_ungated_clk                          (hqm_clk_trunk),
       .hqm_rst_prep_aqed,
       .hqm_gated_rst_b_aqed,
       .hqm_inp_gated_rst_b_aqed,
       .hqm_gated_rst_b_start_aqed,
       .hqm_gated_rst_b_active_aqed,
       .hqm_gated_rst_b_done_aqed,
       .aqed_clk_idle,
       .aqed_clk_enable,
       .hqm_fullrate_clk                         (hqm_clk_trunk),
       .hqm_clk_rptr_rst_sync_b,
       .hqm_gatedclk_enable_and                  (hqm_gated_clk_enable_and_lsp),
       .hqm_clk_ungate                           (hqm_clk_ungate_rptr),
       .aqed_unit_idle                           (i_hqm_aqed_pipe_aqed_unit_idle),
       .aqed_unit_pipeidle,
       .aqed_reset_done,
       .aqed_cfg_req_up_read                     (i_hqm_list_sel_pipe_ap_cfg_req_down_read),
       .aqed_cfg_req_up_write                    (i_hqm_list_sel_pipe_ap_cfg_req_down_write),
       .aqed_cfg_req_up                          (ap_cfg_req_down),
       .aqed_cfg_rsp_up_ack                      (i_hqm_list_sel_pipe_ap_cfg_rsp_down_ack),
       .aqed_cfg_rsp_up                          (ap_cfg_rsp_down),
       .aqed_cfg_req_down_read,
       .aqed_cfg_req_down_write,
       .aqed_cfg_req_down,
       .aqed_cfg_rsp_down_ack,
       .aqed_cfg_rsp_down,
       // Tie to constant value: zero
       .aqed_alarm_up_v                          (1'b0),
       .aqed_alarm_up_ready                      (),
       // Tie to constant value: zero
       .aqed_alarm_up_data                       (25'b0),
       .aqed_alarm_down_v                        (i_hqm_aqed_pipe_aqed_alarm_down_v),
       .aqed_alarm_down_ready                    (i_hqm_list_sel_pipe_ap_alarm_up_ready),
       .aqed_alarm_down_data,
       .lsp_aqed_cmp_v,
       .lsp_aqed_cmp_ready,
       .lsp_aqed_cmp_data,
       .aqed_lsp_dec_fid_cnt_v,
       .aqed_lsp_fid_cnt_upd_v,
       .aqed_lsp_fid_cnt_upd_val,
       .aqed_lsp_fid_cnt_upd_qid,
       .aqed_lsp_stop_atqatm,
       .aqed_lsp_deq_v,
       .aqed_lsp_deq_data,
       .ap_aqed_v                                (i_hqm_list_sel_pipe_ap_aqed_v),
       .ap_aqed_ready                            (i_hqm_aqed_pipe_ap_aqed_ready),
       .ap_aqed_data,
       .qed_aqed_enq_v                           (i_hqm_qed_pipe_qed_aqed_enq_v),
       .qed_aqed_enq_ready                       (i_hqm_aqed_pipe_qed_aqed_enq_ready),
       .qed_aqed_enq_data,
       .aqed_ap_enq_v                            (i_hqm_aqed_pipe_aqed_ap_enq_v),
       .aqed_ap_enq_ready                        (i_hqm_list_sel_pipe_aqed_ap_enq_ready),
       .aqed_ap_enq_data,
       .aqed_chp_sch_v                           (i_hqm_aqed_pipe_aqed_chp_sch_v),
       .aqed_chp_sch_ready                       (i_hqm_credit_hist_pipe_aqed_chp_sch_ready),
       .aqed_chp_sch_data,
       .aqed_lsp_sch_v                           (i_hqm_aqed_pipe_aqed_lsp_sch_v),
       .aqed_lsp_sch_ready                       (i_hqm_list_sel_pipe_aqed_lsp_sch_ready),
       .aqed_lsp_sch_data,
       .bcam_AW_bcam_2048x26_wclk                (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_wclk),
       .bcam_AW_bcam_2048x26_rclk                (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_rclk),
       .bcam_AW_bcam_2048x26_cclk                (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cclk),
       .bcam_AW_bcam_2048x26_dfx_clk             (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_dfx_clk),
       .bcam_AW_bcam_2048x26_we                  (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_we),
       .bcam_AW_bcam_2048x26_waddr               (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_waddr),
       .bcam_AW_bcam_2048x26_wdata               (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_wdata),
       .bcam_AW_bcam_2048x26_ce                  (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_ce),
       .bcam_AW_bcam_2048x26_cdata               (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cdata),
       .bcam_AW_bcam_2048x26_cmatch              (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_cmatch),
       .bcam_AW_bcam_2048x26_re                  (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_re),
       .bcam_AW_bcam_2048x26_raddr               (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_raddr),
       .bcam_AW_bcam_2048x26_rdata               (i_hqm_aqed_pipe_bcam_AW_bcam_2048x26_rdata),
       .rf_aqed_fid_cnt_re                       (i_hqm_aqed_pipe_rf_aqed_fid_cnt_re),
       .rf_aqed_fid_cnt_rclk                     (i_hqm_aqed_pipe_rf_aqed_fid_cnt_rclk),
       .rf_aqed_fid_cnt_rclk_rst_n               (i_hqm_aqed_pipe_rf_aqed_fid_cnt_rclk_rst_n),
       .rf_aqed_fid_cnt_raddr                    (i_hqm_aqed_pipe_rf_aqed_fid_cnt_raddr),
       .rf_aqed_fid_cnt_waddr                    (i_hqm_aqed_pipe_rf_aqed_fid_cnt_waddr),
       .rf_aqed_fid_cnt_we                       (i_hqm_aqed_pipe_rf_aqed_fid_cnt_we),
       .rf_aqed_fid_cnt_wclk                     (i_hqm_aqed_pipe_rf_aqed_fid_cnt_wclk),
       .rf_aqed_fid_cnt_wclk_rst_n               (i_hqm_aqed_pipe_rf_aqed_fid_cnt_wclk_rst_n),
       .rf_aqed_fid_cnt_wdata                    (i_hqm_aqed_pipe_rf_aqed_fid_cnt_wdata),
       .rf_aqed_fid_cnt_rdata                    (i_hqm_aqed_pipe_rf_aqed_fid_cnt_rdata),
       .rf_aqed_fifo_ap_aqed_re                  (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_re),
       .rf_aqed_fifo_ap_aqed_rclk                (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rclk),
       .rf_aqed_fifo_ap_aqed_rclk_rst_n          (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rclk_rst_n),
       .rf_aqed_fifo_ap_aqed_raddr               (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_raddr),
       .rf_aqed_fifo_ap_aqed_waddr               (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_waddr),
       .rf_aqed_fifo_ap_aqed_we                  (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_we),
       .rf_aqed_fifo_ap_aqed_wclk                (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wclk),
       .rf_aqed_fifo_ap_aqed_wclk_rst_n          (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wclk_rst_n),
       .rf_aqed_fifo_ap_aqed_wdata               (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_wdata),
       .rf_aqed_fifo_ap_aqed_rdata               (i_hqm_aqed_pipe_rf_aqed_fifo_ap_aqed_rdata),
       .rf_aqed_fifo_aqed_ap_enq_re              (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_re),
       .rf_aqed_fifo_aqed_ap_enq_rclk            (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rclk),
       .rf_aqed_fifo_aqed_ap_enq_rclk_rst_n      (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rclk_rst_n),
       .rf_aqed_fifo_aqed_ap_enq_raddr           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_raddr),
       .rf_aqed_fifo_aqed_ap_enq_waddr           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_waddr),
       .rf_aqed_fifo_aqed_ap_enq_we              (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_we),
       .rf_aqed_fifo_aqed_ap_enq_wclk            (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wclk),
       .rf_aqed_fifo_aqed_ap_enq_wclk_rst_n      (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wclk_rst_n),
       .rf_aqed_fifo_aqed_ap_enq_wdata           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_wdata),
       .rf_aqed_fifo_aqed_ap_enq_rdata           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_ap_enq_rdata),
       .rf_aqed_fifo_aqed_chp_sch_re             (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_re),
       .rf_aqed_fifo_aqed_chp_sch_rclk           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rclk),
       .rf_aqed_fifo_aqed_chp_sch_rclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rclk_rst_n),
       .rf_aqed_fifo_aqed_chp_sch_raddr          (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_raddr),
       .rf_aqed_fifo_aqed_chp_sch_waddr          (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_waddr),
       .rf_aqed_fifo_aqed_chp_sch_we             (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_we),
       .rf_aqed_fifo_aqed_chp_sch_wclk           (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wclk),
       .rf_aqed_fifo_aqed_chp_sch_wclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wclk_rst_n),
       .rf_aqed_fifo_aqed_chp_sch_wdata          (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_wdata),
       .rf_aqed_fifo_aqed_chp_sch_rdata          (i_hqm_aqed_pipe_rf_aqed_fifo_aqed_chp_sch_rdata),
       .rf_aqed_fifo_freelist_return_re          (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_re),
       .rf_aqed_fifo_freelist_return_rclk        (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rclk),
       .rf_aqed_fifo_freelist_return_rclk_rst_n  (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rclk_rst_n),
       .rf_aqed_fifo_freelist_return_raddr       (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_raddr),
       .rf_aqed_fifo_freelist_return_waddr       (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_waddr),
       .rf_aqed_fifo_freelist_return_we          (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_we),
       .rf_aqed_fifo_freelist_return_wclk        (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wclk),
       .rf_aqed_fifo_freelist_return_wclk_rst_n  (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wclk_rst_n),
       .rf_aqed_fifo_freelist_return_wdata       (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_wdata),
       .rf_aqed_fifo_freelist_return_rdata       (i_hqm_aqed_pipe_rf_aqed_fifo_freelist_return_rdata),
       .rf_aqed_fifo_lsp_aqed_cmp_re             (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_re),
       .rf_aqed_fifo_lsp_aqed_cmp_rclk           (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rclk),
       .rf_aqed_fifo_lsp_aqed_cmp_rclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rclk_rst_n),
       .rf_aqed_fifo_lsp_aqed_cmp_raddr          (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_raddr),
       .rf_aqed_fifo_lsp_aqed_cmp_waddr          (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_waddr),
       .rf_aqed_fifo_lsp_aqed_cmp_we             (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_we),
       .rf_aqed_fifo_lsp_aqed_cmp_wclk           (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wclk),
       .rf_aqed_fifo_lsp_aqed_cmp_wclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wclk_rst_n),
       .rf_aqed_fifo_lsp_aqed_cmp_wdata          (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_wdata),
       .rf_aqed_fifo_lsp_aqed_cmp_rdata          (i_hqm_aqed_pipe_rf_aqed_fifo_lsp_aqed_cmp_rdata),
       .rf_aqed_fifo_qed_aqed_enq_re             (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_re),
       .rf_aqed_fifo_qed_aqed_enq_rclk           (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rclk),
       .rf_aqed_fifo_qed_aqed_enq_rclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rclk_rst_n),
       .rf_aqed_fifo_qed_aqed_enq_raddr          (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_raddr),
       .rf_aqed_fifo_qed_aqed_enq_waddr          (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_waddr),
       .rf_aqed_fifo_qed_aqed_enq_we             (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_we),
       .rf_aqed_fifo_qed_aqed_enq_wclk           (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wclk),
       .rf_aqed_fifo_qed_aqed_enq_wclk_rst_n     (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wclk_rst_n),
       .rf_aqed_fifo_qed_aqed_enq_wdata          (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_wdata),
       .rf_aqed_fifo_qed_aqed_enq_rdata          (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_rdata),
       .rf_aqed_fifo_qed_aqed_enq_fid_re         (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_re),
       .rf_aqed_fifo_qed_aqed_enq_fid_rclk       (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rclk),
       .rf_aqed_fifo_qed_aqed_enq_fid_rclk_rst_n (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rclk_rst_n),
       .rf_aqed_fifo_qed_aqed_enq_fid_raddr      (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_raddr),
       .rf_aqed_fifo_qed_aqed_enq_fid_waddr      (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_waddr),
       .rf_aqed_fifo_qed_aqed_enq_fid_we         (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_we),
       .rf_aqed_fifo_qed_aqed_enq_fid_wclk       (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wclk),
       .rf_aqed_fifo_qed_aqed_enq_fid_wclk_rst_n (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wclk_rst_n),
       .rf_aqed_fifo_qed_aqed_enq_fid_wdata      (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_wdata),
       .rf_aqed_fifo_qed_aqed_enq_fid_rdata      (i_hqm_aqed_pipe_rf_aqed_fifo_qed_aqed_enq_fid_rdata),
       .rf_aqed_ll_cnt_pri0_re                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_re),
       .rf_aqed_ll_cnt_pri0_rclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rclk),
       .rf_aqed_ll_cnt_pri0_rclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rclk_rst_n),
       .rf_aqed_ll_cnt_pri0_raddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_raddr),
       .rf_aqed_ll_cnt_pri0_waddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_waddr),
       .rf_aqed_ll_cnt_pri0_we                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_we),
       .rf_aqed_ll_cnt_pri0_wclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wclk),
       .rf_aqed_ll_cnt_pri0_wclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wclk_rst_n),
       .rf_aqed_ll_cnt_pri0_wdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_wdata),
       .rf_aqed_ll_cnt_pri0_rdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri0_rdata),
       .rf_aqed_ll_cnt_pri1_re                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_re),
       .rf_aqed_ll_cnt_pri1_rclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rclk),
       .rf_aqed_ll_cnt_pri1_rclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rclk_rst_n),
       .rf_aqed_ll_cnt_pri1_raddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_raddr),
       .rf_aqed_ll_cnt_pri1_waddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_waddr),
       .rf_aqed_ll_cnt_pri1_we                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_we),
       .rf_aqed_ll_cnt_pri1_wclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wclk),
       .rf_aqed_ll_cnt_pri1_wclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wclk_rst_n),
       .rf_aqed_ll_cnt_pri1_wdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_wdata),
       .rf_aqed_ll_cnt_pri1_rdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri1_rdata),
       .rf_aqed_ll_cnt_pri2_re                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_re),
       .rf_aqed_ll_cnt_pri2_rclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rclk),
       .rf_aqed_ll_cnt_pri2_rclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rclk_rst_n),
       .rf_aqed_ll_cnt_pri2_raddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_raddr),
       .rf_aqed_ll_cnt_pri2_waddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_waddr),
       .rf_aqed_ll_cnt_pri2_we                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_we),
       .rf_aqed_ll_cnt_pri2_wclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wclk),
       .rf_aqed_ll_cnt_pri2_wclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wclk_rst_n),
       .rf_aqed_ll_cnt_pri2_wdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_wdata),
       .rf_aqed_ll_cnt_pri2_rdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri2_rdata),
       .rf_aqed_ll_cnt_pri3_re                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_re),
       .rf_aqed_ll_cnt_pri3_rclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rclk),
       .rf_aqed_ll_cnt_pri3_rclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rclk_rst_n),
       .rf_aqed_ll_cnt_pri3_raddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_raddr),
       .rf_aqed_ll_cnt_pri3_waddr                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_waddr),
       .rf_aqed_ll_cnt_pri3_we                   (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_we),
       .rf_aqed_ll_cnt_pri3_wclk                 (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wclk),
       .rf_aqed_ll_cnt_pri3_wclk_rst_n           (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wclk_rst_n),
       .rf_aqed_ll_cnt_pri3_wdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_wdata),
       .rf_aqed_ll_cnt_pri3_rdata                (i_hqm_aqed_pipe_rf_aqed_ll_cnt_pri3_rdata),
       .rf_aqed_ll_qe_hp_pri0_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_re),
       .rf_aqed_ll_qe_hp_pri0_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rclk),
       .rf_aqed_ll_qe_hp_pri0_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rclk_rst_n),
       .rf_aqed_ll_qe_hp_pri0_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_raddr),
       .rf_aqed_ll_qe_hp_pri0_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_waddr),
       .rf_aqed_ll_qe_hp_pri0_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_we),
       .rf_aqed_ll_qe_hp_pri0_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wclk),
       .rf_aqed_ll_qe_hp_pri0_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wclk_rst_n),
       .rf_aqed_ll_qe_hp_pri0_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_wdata),
       .rf_aqed_ll_qe_hp_pri0_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri0_rdata),
       .rf_aqed_ll_qe_hp_pri1_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_re),
       .rf_aqed_ll_qe_hp_pri1_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rclk),
       .rf_aqed_ll_qe_hp_pri1_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rclk_rst_n),
       .rf_aqed_ll_qe_hp_pri1_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_raddr),
       .rf_aqed_ll_qe_hp_pri1_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_waddr),
       .rf_aqed_ll_qe_hp_pri1_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_we),
       .rf_aqed_ll_qe_hp_pri1_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wclk),
       .rf_aqed_ll_qe_hp_pri1_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wclk_rst_n),
       .rf_aqed_ll_qe_hp_pri1_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_wdata),
       .rf_aqed_ll_qe_hp_pri1_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri1_rdata),
       .rf_aqed_ll_qe_hp_pri2_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_re),
       .rf_aqed_ll_qe_hp_pri2_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rclk),
       .rf_aqed_ll_qe_hp_pri2_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rclk_rst_n),
       .rf_aqed_ll_qe_hp_pri2_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_raddr),
       .rf_aqed_ll_qe_hp_pri2_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_waddr),
       .rf_aqed_ll_qe_hp_pri2_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_we),
       .rf_aqed_ll_qe_hp_pri2_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wclk),
       .rf_aqed_ll_qe_hp_pri2_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wclk_rst_n),
       .rf_aqed_ll_qe_hp_pri2_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_wdata),
       .rf_aqed_ll_qe_hp_pri2_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri2_rdata),
       .rf_aqed_ll_qe_hp_pri3_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_re),
       .rf_aqed_ll_qe_hp_pri3_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rclk),
       .rf_aqed_ll_qe_hp_pri3_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rclk_rst_n),
       .rf_aqed_ll_qe_hp_pri3_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_raddr),
       .rf_aqed_ll_qe_hp_pri3_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_waddr),
       .rf_aqed_ll_qe_hp_pri3_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_we),
       .rf_aqed_ll_qe_hp_pri3_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wclk),
       .rf_aqed_ll_qe_hp_pri3_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wclk_rst_n),
       .rf_aqed_ll_qe_hp_pri3_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_wdata),
       .rf_aqed_ll_qe_hp_pri3_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_hp_pri3_rdata),
       .rf_aqed_ll_qe_tp_pri0_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_re),
       .rf_aqed_ll_qe_tp_pri0_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rclk),
       .rf_aqed_ll_qe_tp_pri0_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rclk_rst_n),
       .rf_aqed_ll_qe_tp_pri0_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_raddr),
       .rf_aqed_ll_qe_tp_pri0_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_waddr),
       .rf_aqed_ll_qe_tp_pri0_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_we),
       .rf_aqed_ll_qe_tp_pri0_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wclk),
       .rf_aqed_ll_qe_tp_pri0_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wclk_rst_n),
       .rf_aqed_ll_qe_tp_pri0_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_wdata),
       .rf_aqed_ll_qe_tp_pri0_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri0_rdata),
       .rf_aqed_ll_qe_tp_pri1_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_re),
       .rf_aqed_ll_qe_tp_pri1_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rclk),
       .rf_aqed_ll_qe_tp_pri1_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rclk_rst_n),
       .rf_aqed_ll_qe_tp_pri1_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_raddr),
       .rf_aqed_ll_qe_tp_pri1_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_waddr),
       .rf_aqed_ll_qe_tp_pri1_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_we),
       .rf_aqed_ll_qe_tp_pri1_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wclk),
       .rf_aqed_ll_qe_tp_pri1_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wclk_rst_n),
       .rf_aqed_ll_qe_tp_pri1_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_wdata),
       .rf_aqed_ll_qe_tp_pri1_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri1_rdata),
       .rf_aqed_ll_qe_tp_pri2_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_re),
       .rf_aqed_ll_qe_tp_pri2_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rclk),
       .rf_aqed_ll_qe_tp_pri2_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rclk_rst_n),
       .rf_aqed_ll_qe_tp_pri2_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_raddr),
       .rf_aqed_ll_qe_tp_pri2_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_waddr),
       .rf_aqed_ll_qe_tp_pri2_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_we),
       .rf_aqed_ll_qe_tp_pri2_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wclk),
       .rf_aqed_ll_qe_tp_pri2_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wclk_rst_n),
       .rf_aqed_ll_qe_tp_pri2_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_wdata),
       .rf_aqed_ll_qe_tp_pri2_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri2_rdata),
       .rf_aqed_ll_qe_tp_pri3_re                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_re),
       .rf_aqed_ll_qe_tp_pri3_rclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rclk),
       .rf_aqed_ll_qe_tp_pri3_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rclk_rst_n),
       .rf_aqed_ll_qe_tp_pri3_raddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_raddr),
       .rf_aqed_ll_qe_tp_pri3_waddr              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_waddr),
       .rf_aqed_ll_qe_tp_pri3_we                 (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_we),
       .rf_aqed_ll_qe_tp_pri3_wclk               (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wclk),
       .rf_aqed_ll_qe_tp_pri3_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wclk_rst_n),
       .rf_aqed_ll_qe_tp_pri3_wdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_wdata),
       .rf_aqed_ll_qe_tp_pri3_rdata              (i_hqm_aqed_pipe_rf_aqed_ll_qe_tp_pri3_rdata),
       .rf_aqed_qid_cnt_re                       (i_hqm_aqed_pipe_rf_aqed_qid_cnt_re),
       .rf_aqed_qid_cnt_rclk                     (i_hqm_aqed_pipe_rf_aqed_qid_cnt_rclk),
       .rf_aqed_qid_cnt_rclk_rst_n               (i_hqm_aqed_pipe_rf_aqed_qid_cnt_rclk_rst_n),
       .rf_aqed_qid_cnt_raddr                    (i_hqm_aqed_pipe_rf_aqed_qid_cnt_raddr),
       .rf_aqed_qid_cnt_waddr                    (i_hqm_aqed_pipe_rf_aqed_qid_cnt_waddr),
       .rf_aqed_qid_cnt_we                       (i_hqm_aqed_pipe_rf_aqed_qid_cnt_we),
       .rf_aqed_qid_cnt_wclk                     (i_hqm_aqed_pipe_rf_aqed_qid_cnt_wclk),
       .rf_aqed_qid_cnt_wclk_rst_n               (i_hqm_aqed_pipe_rf_aqed_qid_cnt_wclk_rst_n),
       .rf_aqed_qid_cnt_wdata                    (i_hqm_aqed_pipe_rf_aqed_qid_cnt_wdata),
       .rf_aqed_qid_cnt_rdata                    (i_hqm_aqed_pipe_rf_aqed_qid_cnt_rdata),
       .rf_aqed_qid_fid_limit_re                 (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_re),
       .rf_aqed_qid_fid_limit_rclk               (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rclk),
       .rf_aqed_qid_fid_limit_rclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rclk_rst_n),
       .rf_aqed_qid_fid_limit_raddr              (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_raddr),
       .rf_aqed_qid_fid_limit_waddr              (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_waddr),
       .rf_aqed_qid_fid_limit_we                 (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_we),
       .rf_aqed_qid_fid_limit_wclk               (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wclk),
       .rf_aqed_qid_fid_limit_wclk_rst_n         (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wclk_rst_n),
       .rf_aqed_qid_fid_limit_wdata              (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_wdata),
       .rf_aqed_qid_fid_limit_rdata              (i_hqm_aqed_pipe_rf_aqed_qid_fid_limit_rdata),
       .rf_rx_sync_qed_aqed_enq_re               (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_re),
       .rf_rx_sync_qed_aqed_enq_rclk             (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rclk),
       .rf_rx_sync_qed_aqed_enq_rclk_rst_n       (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rclk_rst_n),
       .rf_rx_sync_qed_aqed_enq_raddr            (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_raddr),
       .rf_rx_sync_qed_aqed_enq_waddr            (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_waddr),
       .rf_rx_sync_qed_aqed_enq_we               (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_we),
       .rf_rx_sync_qed_aqed_enq_wclk             (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wclk),
       .rf_rx_sync_qed_aqed_enq_wclk_rst_n       (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wclk_rst_n),
       .rf_rx_sync_qed_aqed_enq_wdata            (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_wdata),
       .rf_rx_sync_qed_aqed_enq_rdata            (i_hqm_aqed_pipe_rf_rx_sync_qed_aqed_enq_rdata),
       .sr_aqed_re                               (i_hqm_aqed_pipe_sr_aqed_re),
       .sr_aqed_clk                              (i_hqm_aqed_pipe_sr_aqed_clk),
       .sr_aqed_clk_rst_n                        (i_hqm_aqed_pipe_sr_aqed_clk_rst_n),
       .sr_aqed_addr                             (i_hqm_aqed_pipe_sr_aqed_addr),
       .sr_aqed_we                               (i_hqm_aqed_pipe_sr_aqed_we),
       .sr_aqed_wdata                            (i_hqm_aqed_pipe_sr_aqed_wdata),
       .sr_aqed_rdata                            (i_hqm_aqed_pipe_sr_aqed_rdata),
       .sr_aqed_freelist_re                      (i_hqm_aqed_pipe_sr_aqed_freelist_re),
       .sr_aqed_freelist_clk                     (i_hqm_aqed_pipe_sr_aqed_freelist_clk),
       .sr_aqed_freelist_clk_rst_n               (i_hqm_aqed_pipe_sr_aqed_freelist_clk_rst_n),
       .sr_aqed_freelist_addr                    (i_hqm_aqed_pipe_sr_aqed_freelist_addr),
       .sr_aqed_freelist_we                      (i_hqm_aqed_pipe_sr_aqed_freelist_we),
       .sr_aqed_freelist_wdata                   (i_hqm_aqed_pipe_sr_aqed_freelist_wdata),
       .sr_aqed_freelist_rdata                   (i_hqm_aqed_pipe_sr_aqed_freelist_rdata),
       .sr_aqed_ll_qe_hpnxt_re                   (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_re),
       .sr_aqed_ll_qe_hpnxt_clk                  (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_clk),
       .sr_aqed_ll_qe_hpnxt_clk_rst_n            (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_clk_rst_n),
       .sr_aqed_ll_qe_hpnxt_addr                 (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_addr),
       .sr_aqed_ll_qe_hpnxt_we                   (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_we),
       .sr_aqed_ll_qe_hpnxt_wdata                (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_wdata),
       .sr_aqed_ll_qe_hpnxt_rdata                (i_hqm_aqed_pipe_sr_aqed_ll_qe_hpnxt_rdata));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_aqed_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk,
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_aqed),
       .hqm_gated_clk          (hqm_gated_clk_lsp),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_aqed),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_aqed),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_aqed),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_aqed),
       .hqm_flr_prep           (hqm_flr_prep_rptr),
       .rst_prep               (hqm_rst_prep_aqed));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_atm_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk,
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_atm),
       .hqm_gated_clk          (hqm_gated_clk_lsp),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_atm),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_atm),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_atm),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_atm),
       .hqm_flr_prep           (hqm_flr_prep_rptr),
       .rst_prep               (hqm_rst_prep_atm));

   hqm_AW_clkgate i_hqm_chp_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_chp),
       .cfg_clkungate   (hqm_clk_ungate_rptrxx),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_chp));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_chp_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_chp),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_chp));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_chp_hqm_gated_clk_enable_or2
      (.clki0 (i_hqm_credit_hist_pipe_hqm_proc_clk_en_chp),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_chp));

   hqm_AW_flop i_hqm_chp_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bxx),
       .data   (hqm_gated_clk_enable_and_chp),
       .data_q (hqm_gated_clk_enable_rptr_chp));

   hqm_AW_reset_sync_scan i_hqm_chp_hqm_gated_rst_pgcb_sync_n
      (.clk            (pgcb_clk),
       .rst_n          (hqm_gated_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (hqm_gated_rst_b_pgcb_sync_chp));

   hqm_AW_clkgate i_hqm_chp_pgcb_clk
      (.clk             (pgcb_clk),
       .enable          (hqm_gated_rst_b_pgcb_sync_chp),
       // Tie to constant value: zero
       .cfg_clkungate   (1'b0),
       .fscan_clkungate,
       .gated_clk       (pgcb_clkx));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(0)) i_hqm_chp_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       .hqm_pgcb_clk           (pgcb_clkx),
       .hqm_pgcb_rst_n         (hqm_pgcb_rst_b_chp),
       .hqm_pgcb_rst_n_start   (hqm_pgcb_rst_b_start_chp),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkxx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_chp),
       .hqm_gated_clk          (hqm_gated_clk_chp),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_chp),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_chp),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_chp),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_chp),
       .hqm_flr_prep           (hqm_flr_prep_rptrxx),
       .rst_prep               (hqm_rst_prep_chp));

   hqm_credit_hist_pipe i_hqm_credit_hist_pipe
      (.hqm_gated_clk                                  (hqm_gated_clk_chp),
       .hqm_inp_gated_clk                              (hqm_inp_gated_clkxx),
       .hqm_proc_clk_en_chp                            (i_hqm_credit_hist_pipe_hqm_proc_clk_en_chp),
       .hqm_rst_prep_chp,
       .hqm_gated_rst_b_chp,
       .hqm_inp_gated_rst_b_chp,
       .hqm_pgcb_clk                                   (pgcb_clkx),
       .hqm_pgcb_rst_b_chp,
       .hqm_pgcb_rst_b_start_chp,
       .hqm_gated_rst_b_start_chp,
       .hqm_gated_rst_b_active_chp,
       .hqm_gated_rst_b_done_chp,
       .rop_unit_idle                                  (i_hqm_reorder_pipe_rop_unit_idle),
       .rop_clk_idle,
       .rop_clk_enable,
       .master_chp_timestamp,
       .hqm_proc_reset_done                            (hqm_proc_reset_done_sync_hqm),
       .chp_unit_idle,
       .chp_unit_pipeidle,
       .chp_reset_done,
       .chp_cfg_req_up_read                            (i_hqm_system_system_cfg_req_down_read),
       .chp_cfg_req_up_write                           (i_hqm_system_system_cfg_req_down_write),
       .chp_cfg_req_up                                 (system_cfg_req_down),
       .chp_cfg_rsp_up_ack                             (i_hqm_system_system_cfg_rsp_down_ack),
       .chp_cfg_rsp_up                                 (system_cfg_rsp_down),
       .chp_cfg_req_down_read                          (i_hqm_credit_hist_pipe_chp_cfg_req_down_read),
       .chp_cfg_req_down_write                         (i_hqm_credit_hist_pipe_chp_cfg_req_down_write),
       .chp_cfg_req_down,
       .chp_cfg_rsp_down_ack                           (i_hqm_credit_hist_pipe_chp_cfg_rsp_down_ack),
       .chp_cfg_rsp_down,
       .chp_alarm_up_v                                 (i_hqm_reorder_pipe_rop_alarm_down_v),
       .chp_alarm_up_ready                             (i_hqm_credit_hist_pipe_chp_alarm_up_ready),
       .chp_alarm_up_data                              (rop_alarm_down_data),
       .chp_alarm_down_v                               (i_hqm_credit_hist_pipe_chp_alarm_down_v),
       .chp_alarm_down_ready                           (i_hqm_system_hqm_alarm_ready),
       .chp_alarm_down_data                            (hqm_alarm_data),
       .hcw_enq_w_req,
       .hcw_enq_w_req_valid                            (i_hqm_system_hcw_enq_w_req_valid),
       .hcw_enq_w_req_ready                            (i_hqm_credit_hist_pipe_hcw_enq_w_req_ready),
       .hcw_sched_w_req,
       .hcw_sched_w_req_valid                          (i_hqm_credit_hist_pipe_hcw_sched_w_req_valid),
       .hcw_sched_w_req_ready                          (i_hqm_system_hcw_sched_w_req_ready),
       .interrupt_w_req,
       .interrupt_w_req_valid                          (i_hqm_credit_hist_pipe_interrupt_w_req_valid),
       .interrupt_w_req_ready                          (i_hqm_system_interrupt_w_req_ready),
       .cwdi_interrupt_w_req_valid                     (i_hqm_credit_hist_pipe_cwdi_interrupt_w_req_valid),
       .cwdi_interrupt_w_req_ready                     (i_hqm_system_cwdi_interrupt_w_req_ready),
       .chp_rop_hcw_v                                  (i_hqm_credit_hist_pipe_chp_rop_hcw_v),
       .chp_rop_hcw_ready                              (i_hqm_reorder_pipe_chp_rop_hcw_ready),
       .chp_rop_hcw_data,
       .chp_lsp_ldb_cq_off,
       .chp_lsp_cmp_v                                  (i_hqm_credit_hist_pipe_chp_lsp_cmp_v),
       .chp_lsp_cmp_ready                              (i_hqm_list_sel_pipe_chp_lsp_cmp_ready),
       .chp_lsp_cmp_data,
       .chp_lsp_token_v                                (i_hqm_credit_hist_pipe_chp_lsp_token_v),
       .chp_lsp_token_ready                            (i_hqm_list_sel_pipe_chp_lsp_token_ready),
       .chp_lsp_token_data,
       .qed_chp_sch_v                                  (i_hqm_qed_pipe_qed_chp_sch_v),
       .qed_chp_sch_ready                              (i_hqm_credit_hist_pipe_qed_chp_sch_ready),
       .qed_chp_sch_data,
       .aqed_chp_sch_v                                 (i_hqm_aqed_pipe_aqed_chp_sch_v),
       .aqed_chp_sch_ready                             (i_hqm_credit_hist_pipe_aqed_chp_sch_ready),
       .aqed_chp_sch_data,
       .visa_str_chp_lsp_cmp_data,
       .wd_clkreq,
       .rf_aqed_chp_sch_rx_sync_mem_re                 (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_re),
       .rf_aqed_chp_sch_rx_sync_mem_rclk               (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rclk),
       .rf_aqed_chp_sch_rx_sync_mem_rclk_rst_n         (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rclk_rst_n),
       .rf_aqed_chp_sch_rx_sync_mem_raddr              (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_raddr),
       .rf_aqed_chp_sch_rx_sync_mem_waddr              (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_waddr),
       .rf_aqed_chp_sch_rx_sync_mem_we                 (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_we),
       .rf_aqed_chp_sch_rx_sync_mem_wclk               (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wclk),
       .rf_aqed_chp_sch_rx_sync_mem_wclk_rst_n         (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wclk_rst_n),
       .rf_aqed_chp_sch_rx_sync_mem_wdata              (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_wdata),
       .rf_aqed_chp_sch_rx_sync_mem_rdata              (i_hqm_credit_hist_pipe_rf_aqed_chp_sch_rx_sync_mem_rdata),
       .rf_chp_chp_rop_hcw_fifo_mem_re                 (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_re),
       .rf_chp_chp_rop_hcw_fifo_mem_rclk               (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rclk),
       .rf_chp_chp_rop_hcw_fifo_mem_rclk_rst_n         (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rclk_rst_n),
       .rf_chp_chp_rop_hcw_fifo_mem_raddr              (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_raddr),
       .rf_chp_chp_rop_hcw_fifo_mem_waddr              (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_waddr),
       .rf_chp_chp_rop_hcw_fifo_mem_we                 (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_we),
       .rf_chp_chp_rop_hcw_fifo_mem_wclk               (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wclk),
       .rf_chp_chp_rop_hcw_fifo_mem_wclk_rst_n         (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wclk_rst_n),
       .rf_chp_chp_rop_hcw_fifo_mem_wdata              (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_wdata),
       .rf_chp_chp_rop_hcw_fifo_mem_rdata              (i_hqm_credit_hist_pipe_rf_chp_chp_rop_hcw_fifo_mem_rdata),
       .rf_chp_lsp_ap_cmp_fifo_mem_re                  (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_re),
       .rf_chp_lsp_ap_cmp_fifo_mem_rclk                (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rclk),
       .rf_chp_lsp_ap_cmp_fifo_mem_rclk_rst_n          (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rclk_rst_n),
       .rf_chp_lsp_ap_cmp_fifo_mem_raddr               (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_raddr),
       .rf_chp_lsp_ap_cmp_fifo_mem_waddr               (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_waddr),
       .rf_chp_lsp_ap_cmp_fifo_mem_we                  (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_we),
       .rf_chp_lsp_ap_cmp_fifo_mem_wclk                (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wclk),
       .rf_chp_lsp_ap_cmp_fifo_mem_wclk_rst_n          (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wclk_rst_n),
       .rf_chp_lsp_ap_cmp_fifo_mem_wdata               (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_wdata),
       .rf_chp_lsp_ap_cmp_fifo_mem_rdata               (i_hqm_credit_hist_pipe_rf_chp_lsp_ap_cmp_fifo_mem_rdata),
       .rf_chp_lsp_tok_fifo_mem_re                     (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_re),
       .rf_chp_lsp_tok_fifo_mem_rclk                   (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rclk),
       .rf_chp_lsp_tok_fifo_mem_rclk_rst_n             (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rclk_rst_n),
       .rf_chp_lsp_tok_fifo_mem_raddr                  (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_raddr),
       .rf_chp_lsp_tok_fifo_mem_waddr                  (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_waddr),
       .rf_chp_lsp_tok_fifo_mem_we                     (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_we),
       .rf_chp_lsp_tok_fifo_mem_wclk                   (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wclk),
       .rf_chp_lsp_tok_fifo_mem_wclk_rst_n             (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wclk_rst_n),
       .rf_chp_lsp_tok_fifo_mem_wdata                  (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_wdata),
       .rf_chp_lsp_tok_fifo_mem_rdata                  (i_hqm_credit_hist_pipe_rf_chp_lsp_tok_fifo_mem_rdata),
       .rf_chp_sys_tx_fifo_mem_re                      (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_re),
       .rf_chp_sys_tx_fifo_mem_rclk                    (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rclk),
       .rf_chp_sys_tx_fifo_mem_rclk_rst_n              (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rclk_rst_n),
       .rf_chp_sys_tx_fifo_mem_raddr                   (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_raddr),
       .rf_chp_sys_tx_fifo_mem_waddr                   (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_waddr),
       .rf_chp_sys_tx_fifo_mem_we                      (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_we),
       .rf_chp_sys_tx_fifo_mem_wclk                    (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wclk),
       .rf_chp_sys_tx_fifo_mem_wclk_rst_n              (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wclk_rst_n),
       .rf_chp_sys_tx_fifo_mem_wdata                   (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_wdata),
       .rf_chp_sys_tx_fifo_mem_rdata                   (i_hqm_credit_hist_pipe_rf_chp_sys_tx_fifo_mem_rdata),
       .rf_cmp_id_chk_enbl_mem_re                      (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_re),
       .rf_cmp_id_chk_enbl_mem_rclk                    (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rclk),
       .rf_cmp_id_chk_enbl_mem_rclk_rst_n              (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rclk_rst_n),
       .rf_cmp_id_chk_enbl_mem_raddr                   (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_raddr),
       .rf_cmp_id_chk_enbl_mem_waddr                   (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_waddr),
       .rf_cmp_id_chk_enbl_mem_we                      (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_we),
       .rf_cmp_id_chk_enbl_mem_wclk                    (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wclk),
       .rf_cmp_id_chk_enbl_mem_wclk_rst_n              (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wclk_rst_n),
       .rf_cmp_id_chk_enbl_mem_wdata                   (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_wdata),
       .rf_cmp_id_chk_enbl_mem_rdata                   (i_hqm_credit_hist_pipe_rf_cmp_id_chk_enbl_mem_rdata),
       .rf_count_rmw_pipe_dir_mem_re                   (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_re),
       .rf_count_rmw_pipe_dir_mem_rclk                 (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rclk),
       .rf_count_rmw_pipe_dir_mem_rclk_rst_n           (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rclk_rst_n),
       .rf_count_rmw_pipe_dir_mem_raddr                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_raddr),
       .rf_count_rmw_pipe_dir_mem_waddr                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_waddr),
       .rf_count_rmw_pipe_dir_mem_we                   (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_we),
       .rf_count_rmw_pipe_dir_mem_wclk                 (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wclk),
       .rf_count_rmw_pipe_dir_mem_wclk_rst_n           (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wclk_rst_n),
       .rf_count_rmw_pipe_dir_mem_wdata                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_wdata),
       .rf_count_rmw_pipe_dir_mem_rdata                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_dir_mem_rdata),
       .rf_count_rmw_pipe_ldb_mem_re                   (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_re),
       .rf_count_rmw_pipe_ldb_mem_rclk                 (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rclk),
       .rf_count_rmw_pipe_ldb_mem_rclk_rst_n           (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rclk_rst_n),
       .rf_count_rmw_pipe_ldb_mem_raddr                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_raddr),
       .rf_count_rmw_pipe_ldb_mem_waddr                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_waddr),
       .rf_count_rmw_pipe_ldb_mem_we                   (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_we),
       .rf_count_rmw_pipe_ldb_mem_wclk                 (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wclk),
       .rf_count_rmw_pipe_ldb_mem_wclk_rst_n           (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wclk_rst_n),
       .rf_count_rmw_pipe_ldb_mem_wdata                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_wdata),
       .rf_count_rmw_pipe_ldb_mem_rdata                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_ldb_mem_rdata),
       .rf_count_rmw_pipe_wd_dir_mem_re                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_re),
       .rf_count_rmw_pipe_wd_dir_mem_rclk              (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rclk),
       .rf_count_rmw_pipe_wd_dir_mem_rclk_rst_n        (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rclk_rst_n),
       .rf_count_rmw_pipe_wd_dir_mem_raddr             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_raddr),
       .rf_count_rmw_pipe_wd_dir_mem_waddr             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_waddr),
       .rf_count_rmw_pipe_wd_dir_mem_we                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_we),
       .rf_count_rmw_pipe_wd_dir_mem_wclk              (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wclk),
       .rf_count_rmw_pipe_wd_dir_mem_wclk_rst_n        (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wclk_rst_n),
       .rf_count_rmw_pipe_wd_dir_mem_wdata             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_wdata),
       .rf_count_rmw_pipe_wd_dir_mem_rdata             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_dir_mem_rdata),
       .rf_count_rmw_pipe_wd_ldb_mem_re                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_re),
       .rf_count_rmw_pipe_wd_ldb_mem_rclk              (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rclk),
       .rf_count_rmw_pipe_wd_ldb_mem_rclk_rst_n        (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rclk_rst_n),
       .rf_count_rmw_pipe_wd_ldb_mem_raddr             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_raddr),
       .rf_count_rmw_pipe_wd_ldb_mem_waddr             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_waddr),
       .rf_count_rmw_pipe_wd_ldb_mem_we                (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_we),
       .rf_count_rmw_pipe_wd_ldb_mem_wclk              (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wclk),
       .rf_count_rmw_pipe_wd_ldb_mem_wclk_rst_n        (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wclk_rst_n),
       .rf_count_rmw_pipe_wd_ldb_mem_wdata             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_wdata),
       .rf_count_rmw_pipe_wd_ldb_mem_rdata             (i_hqm_credit_hist_pipe_rf_count_rmw_pipe_wd_ldb_mem_rdata),
       .rf_dir_cq_depth_re                             (i_hqm_credit_hist_pipe_rf_dir_cq_depth_re),
       .rf_dir_cq_depth_rclk                           (i_hqm_credit_hist_pipe_rf_dir_cq_depth_rclk),
       .rf_dir_cq_depth_rclk_rst_n                     (i_hqm_credit_hist_pipe_rf_dir_cq_depth_rclk_rst_n),
       .rf_dir_cq_depth_raddr                          (i_hqm_credit_hist_pipe_rf_dir_cq_depth_raddr),
       .rf_dir_cq_depth_waddr                          (i_hqm_credit_hist_pipe_rf_dir_cq_depth_waddr),
       .rf_dir_cq_depth_we                             (i_hqm_credit_hist_pipe_rf_dir_cq_depth_we),
       .rf_dir_cq_depth_wclk                           (i_hqm_credit_hist_pipe_rf_dir_cq_depth_wclk),
       .rf_dir_cq_depth_wclk_rst_n                     (i_hqm_credit_hist_pipe_rf_dir_cq_depth_wclk_rst_n),
       .rf_dir_cq_depth_wdata                          (i_hqm_credit_hist_pipe_rf_dir_cq_depth_wdata),
       .rf_dir_cq_depth_rdata                          (i_hqm_credit_hist_pipe_rf_dir_cq_depth_rdata),
       .rf_dir_cq_intr_thresh_re                       (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_re),
       .rf_dir_cq_intr_thresh_rclk                     (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rclk),
       .rf_dir_cq_intr_thresh_rclk_rst_n               (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rclk_rst_n),
       .rf_dir_cq_intr_thresh_raddr                    (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_raddr),
       .rf_dir_cq_intr_thresh_waddr                    (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_waddr),
       .rf_dir_cq_intr_thresh_we                       (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_we),
       .rf_dir_cq_intr_thresh_wclk                     (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wclk),
       .rf_dir_cq_intr_thresh_wclk_rst_n               (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wclk_rst_n),
       .rf_dir_cq_intr_thresh_wdata                    (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_wdata),
       .rf_dir_cq_intr_thresh_rdata                    (i_hqm_credit_hist_pipe_rf_dir_cq_intr_thresh_rdata),
       .rf_dir_cq_token_depth_select_re                (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_re),
       .rf_dir_cq_token_depth_select_rclk              (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rclk),
       .rf_dir_cq_token_depth_select_rclk_rst_n        (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rclk_rst_n),
       .rf_dir_cq_token_depth_select_raddr             (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_raddr),
       .rf_dir_cq_token_depth_select_waddr             (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_waddr),
       .rf_dir_cq_token_depth_select_we                (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_we),
       .rf_dir_cq_token_depth_select_wclk              (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wclk),
       .rf_dir_cq_token_depth_select_wclk_rst_n        (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wclk_rst_n),
       .rf_dir_cq_token_depth_select_wdata             (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_wdata),
       .rf_dir_cq_token_depth_select_rdata             (i_hqm_credit_hist_pipe_rf_dir_cq_token_depth_select_rdata),
       .rf_dir_cq_wptr_re                              (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_re),
       .rf_dir_cq_wptr_rclk                            (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rclk),
       .rf_dir_cq_wptr_rclk_rst_n                      (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rclk_rst_n),
       .rf_dir_cq_wptr_raddr                           (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_raddr),
       .rf_dir_cq_wptr_waddr                           (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_waddr),
       .rf_dir_cq_wptr_we                              (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_we),
       .rf_dir_cq_wptr_wclk                            (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wclk),
       .rf_dir_cq_wptr_wclk_rst_n                      (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wclk_rst_n),
       .rf_dir_cq_wptr_wdata                           (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_wdata),
       .rf_dir_cq_wptr_rdata                           (i_hqm_credit_hist_pipe_rf_dir_cq_wptr_rdata),
       .rf_hcw_enq_w_rx_sync_mem_re                    (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_re),
       .rf_hcw_enq_w_rx_sync_mem_rclk                  (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rclk),
       .rf_hcw_enq_w_rx_sync_mem_rclk_rst_n            (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rclk_rst_n),
       .rf_hcw_enq_w_rx_sync_mem_raddr                 (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_raddr),
       .rf_hcw_enq_w_rx_sync_mem_waddr                 (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_waddr),
       .rf_hcw_enq_w_rx_sync_mem_we                    (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_we),
       .rf_hcw_enq_w_rx_sync_mem_wclk                  (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wclk),
       .rf_hcw_enq_w_rx_sync_mem_wclk_rst_n            (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wclk_rst_n),
       .rf_hcw_enq_w_rx_sync_mem_wdata                 (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_wdata),
       .rf_hcw_enq_w_rx_sync_mem_rdata                 (i_hqm_credit_hist_pipe_rf_hcw_enq_w_rx_sync_mem_rdata),
       .rf_hist_list_a_minmax_re                       (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_re),
       .rf_hist_list_a_minmax_rclk                     (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rclk),
       .rf_hist_list_a_minmax_rclk_rst_n               (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rclk_rst_n),
       .rf_hist_list_a_minmax_raddr                    (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_raddr),
       .rf_hist_list_a_minmax_waddr                    (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_waddr),
       .rf_hist_list_a_minmax_we                       (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_we),
       .rf_hist_list_a_minmax_wclk                     (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wclk),
       .rf_hist_list_a_minmax_wclk_rst_n               (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wclk_rst_n),
       .rf_hist_list_a_minmax_wdata                    (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_wdata),
       .rf_hist_list_a_minmax_rdata                    (i_hqm_credit_hist_pipe_rf_hist_list_a_minmax_rdata),
       .rf_hist_list_a_ptr_re                          (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_re),
       .rf_hist_list_a_ptr_rclk                        (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rclk),
       .rf_hist_list_a_ptr_rclk_rst_n                  (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rclk_rst_n),
       .rf_hist_list_a_ptr_raddr                       (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_raddr),
       .rf_hist_list_a_ptr_waddr                       (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_waddr),
       .rf_hist_list_a_ptr_we                          (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_we),
       .rf_hist_list_a_ptr_wclk                        (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wclk),
       .rf_hist_list_a_ptr_wclk_rst_n                  (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wclk_rst_n),
       .rf_hist_list_a_ptr_wdata                       (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_wdata),
       .rf_hist_list_a_ptr_rdata                       (i_hqm_credit_hist_pipe_rf_hist_list_a_ptr_rdata),
       .rf_hist_list_minmax_re                         (i_hqm_credit_hist_pipe_rf_hist_list_minmax_re),
       .rf_hist_list_minmax_rclk                       (i_hqm_credit_hist_pipe_rf_hist_list_minmax_rclk),
       .rf_hist_list_minmax_rclk_rst_n                 (i_hqm_credit_hist_pipe_rf_hist_list_minmax_rclk_rst_n),
       .rf_hist_list_minmax_raddr                      (i_hqm_credit_hist_pipe_rf_hist_list_minmax_raddr),
       .rf_hist_list_minmax_waddr                      (i_hqm_credit_hist_pipe_rf_hist_list_minmax_waddr),
       .rf_hist_list_minmax_we                         (i_hqm_credit_hist_pipe_rf_hist_list_minmax_we),
       .rf_hist_list_minmax_wclk                       (i_hqm_credit_hist_pipe_rf_hist_list_minmax_wclk),
       .rf_hist_list_minmax_wclk_rst_n                 (i_hqm_credit_hist_pipe_rf_hist_list_minmax_wclk_rst_n),
       .rf_hist_list_minmax_wdata                      (i_hqm_credit_hist_pipe_rf_hist_list_minmax_wdata),
       .rf_hist_list_minmax_rdata                      (i_hqm_credit_hist_pipe_rf_hist_list_minmax_rdata),
       .rf_hist_list_ptr_re                            (i_hqm_credit_hist_pipe_rf_hist_list_ptr_re),
       .rf_hist_list_ptr_rclk                          (i_hqm_credit_hist_pipe_rf_hist_list_ptr_rclk),
       .rf_hist_list_ptr_rclk_rst_n                    (i_hqm_credit_hist_pipe_rf_hist_list_ptr_rclk_rst_n),
       .rf_hist_list_ptr_raddr                         (i_hqm_credit_hist_pipe_rf_hist_list_ptr_raddr),
       .rf_hist_list_ptr_waddr                         (i_hqm_credit_hist_pipe_rf_hist_list_ptr_waddr),
       .rf_hist_list_ptr_we                            (i_hqm_credit_hist_pipe_rf_hist_list_ptr_we),
       .rf_hist_list_ptr_wclk                          (i_hqm_credit_hist_pipe_rf_hist_list_ptr_wclk),
       .rf_hist_list_ptr_wclk_rst_n                    (i_hqm_credit_hist_pipe_rf_hist_list_ptr_wclk_rst_n),
       .rf_hist_list_ptr_wdata                         (i_hqm_credit_hist_pipe_rf_hist_list_ptr_wdata),
       .rf_hist_list_ptr_rdata                         (i_hqm_credit_hist_pipe_rf_hist_list_ptr_rdata),
       .rf_ldb_cq_depth_re                             (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_re),
       .rf_ldb_cq_depth_rclk                           (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rclk),
       .rf_ldb_cq_depth_rclk_rst_n                     (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rclk_rst_n),
       .rf_ldb_cq_depth_raddr                          (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_raddr),
       .rf_ldb_cq_depth_waddr                          (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_waddr),
       .rf_ldb_cq_depth_we                             (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_we),
       .rf_ldb_cq_depth_wclk                           (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wclk),
       .rf_ldb_cq_depth_wclk_rst_n                     (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wclk_rst_n),
       .rf_ldb_cq_depth_wdata                          (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_wdata),
       .rf_ldb_cq_depth_rdata                          (i_hqm_credit_hist_pipe_rf_ldb_cq_depth_rdata),
       .rf_ldb_cq_intr_thresh_re                       (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_re),
       .rf_ldb_cq_intr_thresh_rclk                     (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rclk),
       .rf_ldb_cq_intr_thresh_rclk_rst_n               (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rclk_rst_n),
       .rf_ldb_cq_intr_thresh_raddr                    (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_raddr),
       .rf_ldb_cq_intr_thresh_waddr                    (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_waddr),
       .rf_ldb_cq_intr_thresh_we                       (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_we),
       .rf_ldb_cq_intr_thresh_wclk                     (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wclk),
       .rf_ldb_cq_intr_thresh_wclk_rst_n               (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wclk_rst_n),
       .rf_ldb_cq_intr_thresh_wdata                    (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_wdata),
       .rf_ldb_cq_intr_thresh_rdata                    (i_hqm_credit_hist_pipe_rf_ldb_cq_intr_thresh_rdata),
       .rf_ldb_cq_on_off_threshold_re                  (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_re),
       .rf_ldb_cq_on_off_threshold_rclk                (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rclk),
       .rf_ldb_cq_on_off_threshold_rclk_rst_n          (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rclk_rst_n),
       .rf_ldb_cq_on_off_threshold_raddr               (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_raddr),
       .rf_ldb_cq_on_off_threshold_waddr               (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_waddr),
       .rf_ldb_cq_on_off_threshold_we                  (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_we),
       .rf_ldb_cq_on_off_threshold_wclk                (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wclk),
       .rf_ldb_cq_on_off_threshold_wclk_rst_n          (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wclk_rst_n),
       .rf_ldb_cq_on_off_threshold_wdata               (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_wdata),
       .rf_ldb_cq_on_off_threshold_rdata               (i_hqm_credit_hist_pipe_rf_ldb_cq_on_off_threshold_rdata),
       .rf_ldb_cq_token_depth_select_re                (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_re),
       .rf_ldb_cq_token_depth_select_rclk              (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rclk),
       .rf_ldb_cq_token_depth_select_rclk_rst_n        (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rclk_rst_n),
       .rf_ldb_cq_token_depth_select_raddr             (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_raddr),
       .rf_ldb_cq_token_depth_select_waddr             (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_waddr),
       .rf_ldb_cq_token_depth_select_we                (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_we),
       .rf_ldb_cq_token_depth_select_wclk              (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wclk),
       .rf_ldb_cq_token_depth_select_wclk_rst_n        (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wclk_rst_n),
       .rf_ldb_cq_token_depth_select_wdata             (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_wdata),
       .rf_ldb_cq_token_depth_select_rdata             (i_hqm_credit_hist_pipe_rf_ldb_cq_token_depth_select_rdata),
       .rf_ldb_cq_wptr_re                              (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_re),
       .rf_ldb_cq_wptr_rclk                            (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rclk),
       .rf_ldb_cq_wptr_rclk_rst_n                      (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rclk_rst_n),
       .rf_ldb_cq_wptr_raddr                           (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_raddr),
       .rf_ldb_cq_wptr_waddr                           (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_waddr),
       .rf_ldb_cq_wptr_we                              (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_we),
       .rf_ldb_cq_wptr_wclk                            (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wclk),
       .rf_ldb_cq_wptr_wclk_rst_n                      (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wclk_rst_n),
       .rf_ldb_cq_wptr_wdata                           (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_wdata),
       .rf_ldb_cq_wptr_rdata                           (i_hqm_credit_hist_pipe_rf_ldb_cq_wptr_rdata),
       .rf_ord_qid_sn_re                               (i_hqm_credit_hist_pipe_rf_ord_qid_sn_re),
       .rf_ord_qid_sn_rclk                             (i_hqm_credit_hist_pipe_rf_ord_qid_sn_rclk),
       .rf_ord_qid_sn_rclk_rst_n                       (i_hqm_credit_hist_pipe_rf_ord_qid_sn_rclk_rst_n),
       .rf_ord_qid_sn_raddr                            (i_hqm_credit_hist_pipe_rf_ord_qid_sn_raddr),
       .rf_ord_qid_sn_waddr                            (i_hqm_credit_hist_pipe_rf_ord_qid_sn_waddr),
       .rf_ord_qid_sn_we                               (i_hqm_credit_hist_pipe_rf_ord_qid_sn_we),
       .rf_ord_qid_sn_wclk                             (i_hqm_credit_hist_pipe_rf_ord_qid_sn_wclk),
       .rf_ord_qid_sn_wclk_rst_n                       (i_hqm_credit_hist_pipe_rf_ord_qid_sn_wclk_rst_n),
       .rf_ord_qid_sn_wdata                            (i_hqm_credit_hist_pipe_rf_ord_qid_sn_wdata),
       .rf_ord_qid_sn_rdata                            (i_hqm_credit_hist_pipe_rf_ord_qid_sn_rdata),
       .rf_ord_qid_sn_map_re                           (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_re),
       .rf_ord_qid_sn_map_rclk                         (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rclk),
       .rf_ord_qid_sn_map_rclk_rst_n                   (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rclk_rst_n),
       .rf_ord_qid_sn_map_raddr                        (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_raddr),
       .rf_ord_qid_sn_map_waddr                        (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_waddr),
       .rf_ord_qid_sn_map_we                           (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_we),
       .rf_ord_qid_sn_map_wclk                         (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wclk),
       .rf_ord_qid_sn_map_wclk_rst_n                   (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wclk_rst_n),
       .rf_ord_qid_sn_map_wdata                        (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_wdata),
       .rf_ord_qid_sn_map_rdata                        (i_hqm_credit_hist_pipe_rf_ord_qid_sn_map_rdata),
       .rf_outbound_hcw_fifo_mem_re                    (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_re),
       .rf_outbound_hcw_fifo_mem_rclk                  (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rclk),
       .rf_outbound_hcw_fifo_mem_rclk_rst_n            (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rclk_rst_n),
       .rf_outbound_hcw_fifo_mem_raddr                 (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_raddr),
       .rf_outbound_hcw_fifo_mem_waddr                 (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_waddr),
       .rf_outbound_hcw_fifo_mem_we                    (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_we),
       .rf_outbound_hcw_fifo_mem_wclk                  (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wclk),
       .rf_outbound_hcw_fifo_mem_wclk_rst_n            (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wclk_rst_n),
       .rf_outbound_hcw_fifo_mem_wdata                 (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_wdata),
       .rf_outbound_hcw_fifo_mem_rdata                 (i_hqm_credit_hist_pipe_rf_outbound_hcw_fifo_mem_rdata),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_re         (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_re),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk       (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk_rst_n (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rclk_rst_n),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_raddr      (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_raddr),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_waddr      (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_waddr),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_we         (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_we),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk       (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk_rst_n (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wclk_rst_n),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_wdata      (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_wdata),
       .rf_qed_chp_sch_flid_ret_rx_sync_mem_rdata      (i_hqm_credit_hist_pipe_rf_qed_chp_sch_flid_ret_rx_sync_mem_rdata),
       .rf_qed_chp_sch_rx_sync_mem_re                  (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_re),
       .rf_qed_chp_sch_rx_sync_mem_rclk                (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rclk),
       .rf_qed_chp_sch_rx_sync_mem_rclk_rst_n          (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rclk_rst_n),
       .rf_qed_chp_sch_rx_sync_mem_raddr               (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_raddr),
       .rf_qed_chp_sch_rx_sync_mem_waddr               (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_waddr),
       .rf_qed_chp_sch_rx_sync_mem_we                  (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_we),
       .rf_qed_chp_sch_rx_sync_mem_wclk                (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wclk),
       .rf_qed_chp_sch_rx_sync_mem_wclk_rst_n          (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wclk_rst_n),
       .rf_qed_chp_sch_rx_sync_mem_wdata               (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_wdata),
       .rf_qed_chp_sch_rx_sync_mem_rdata               (i_hqm_credit_hist_pipe_rf_qed_chp_sch_rx_sync_mem_rdata),
       .rf_qed_to_cq_fifo_mem_re                       (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_re),
       .rf_qed_to_cq_fifo_mem_rclk                     (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rclk),
       .rf_qed_to_cq_fifo_mem_rclk_rst_n               (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rclk_rst_n),
       .rf_qed_to_cq_fifo_mem_raddr                    (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_raddr),
       .rf_qed_to_cq_fifo_mem_waddr                    (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_waddr),
       .rf_qed_to_cq_fifo_mem_we                       (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_we),
       .rf_qed_to_cq_fifo_mem_wclk                     (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wclk),
       .rf_qed_to_cq_fifo_mem_wclk_rst_n               (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wclk_rst_n),
       .rf_qed_to_cq_fifo_mem_wdata                    (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_wdata),
       .rf_qed_to_cq_fifo_mem_rdata                    (i_hqm_credit_hist_pipe_rf_qed_to_cq_fifo_mem_rdata),
       .rf_threshold_r_pipe_dir_mem_re                 (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_re),
       .rf_threshold_r_pipe_dir_mem_rclk               (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rclk),
       .rf_threshold_r_pipe_dir_mem_rclk_rst_n         (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rclk_rst_n),
       .rf_threshold_r_pipe_dir_mem_raddr              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_raddr),
       .rf_threshold_r_pipe_dir_mem_waddr              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_waddr),
       .rf_threshold_r_pipe_dir_mem_we                 (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_we),
       .rf_threshold_r_pipe_dir_mem_wclk               (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wclk),
       .rf_threshold_r_pipe_dir_mem_wclk_rst_n         (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wclk_rst_n),
       .rf_threshold_r_pipe_dir_mem_wdata              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_wdata),
       .rf_threshold_r_pipe_dir_mem_rdata              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_dir_mem_rdata),
       .rf_threshold_r_pipe_ldb_mem_re                 (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_re),
       .rf_threshold_r_pipe_ldb_mem_rclk               (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rclk),
       .rf_threshold_r_pipe_ldb_mem_rclk_rst_n         (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rclk_rst_n),
       .rf_threshold_r_pipe_ldb_mem_raddr              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_raddr),
       .rf_threshold_r_pipe_ldb_mem_waddr              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_waddr),
       .rf_threshold_r_pipe_ldb_mem_we                 (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_we),
       .rf_threshold_r_pipe_ldb_mem_wclk               (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wclk),
       .rf_threshold_r_pipe_ldb_mem_wclk_rst_n         (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wclk_rst_n),
       .rf_threshold_r_pipe_ldb_mem_wdata              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_wdata),
       .rf_threshold_r_pipe_ldb_mem_rdata              (i_hqm_credit_hist_pipe_rf_threshold_r_pipe_ldb_mem_rdata),
       .sr_freelist_0_re                               (i_hqm_credit_hist_pipe_sr_freelist_0_re),
       .sr_freelist_0_clk                              (i_hqm_credit_hist_pipe_sr_freelist_0_clk),
       .sr_freelist_0_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_0_clk_rst_n),
       .sr_freelist_0_addr                             (i_hqm_credit_hist_pipe_sr_freelist_0_addr),
       .sr_freelist_0_we                               (i_hqm_credit_hist_pipe_sr_freelist_0_we),
       .sr_freelist_0_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_0_wdata),
       .sr_freelist_0_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_0_rdata),
       .sr_freelist_1_re                               (i_hqm_credit_hist_pipe_sr_freelist_1_re),
       .sr_freelist_1_clk                              (i_hqm_credit_hist_pipe_sr_freelist_1_clk),
       .sr_freelist_1_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_1_clk_rst_n),
       .sr_freelist_1_addr                             (i_hqm_credit_hist_pipe_sr_freelist_1_addr),
       .sr_freelist_1_we                               (i_hqm_credit_hist_pipe_sr_freelist_1_we),
       .sr_freelist_1_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_1_wdata),
       .sr_freelist_1_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_1_rdata),
       .sr_freelist_2_re                               (i_hqm_credit_hist_pipe_sr_freelist_2_re),
       .sr_freelist_2_clk                              (i_hqm_credit_hist_pipe_sr_freelist_2_clk),
       .sr_freelist_2_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_2_clk_rst_n),
       .sr_freelist_2_addr                             (i_hqm_credit_hist_pipe_sr_freelist_2_addr),
       .sr_freelist_2_we                               (i_hqm_credit_hist_pipe_sr_freelist_2_we),
       .sr_freelist_2_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_2_wdata),
       .sr_freelist_2_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_2_rdata),
       .sr_freelist_3_re                               (i_hqm_credit_hist_pipe_sr_freelist_3_re),
       .sr_freelist_3_clk                              (i_hqm_credit_hist_pipe_sr_freelist_3_clk),
       .sr_freelist_3_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_3_clk_rst_n),
       .sr_freelist_3_addr                             (i_hqm_credit_hist_pipe_sr_freelist_3_addr),
       .sr_freelist_3_we                               (i_hqm_credit_hist_pipe_sr_freelist_3_we),
       .sr_freelist_3_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_3_wdata),
       .sr_freelist_3_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_3_rdata),
       .sr_freelist_4_re                               (i_hqm_credit_hist_pipe_sr_freelist_4_re),
       .sr_freelist_4_clk                              (i_hqm_credit_hist_pipe_sr_freelist_4_clk),
       .sr_freelist_4_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_4_clk_rst_n),
       .sr_freelist_4_addr                             (i_hqm_credit_hist_pipe_sr_freelist_4_addr),
       .sr_freelist_4_we                               (i_hqm_credit_hist_pipe_sr_freelist_4_we),
       .sr_freelist_4_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_4_wdata),
       .sr_freelist_4_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_4_rdata),
       .sr_freelist_5_re                               (i_hqm_credit_hist_pipe_sr_freelist_5_re),
       .sr_freelist_5_clk                              (i_hqm_credit_hist_pipe_sr_freelist_5_clk),
       .sr_freelist_5_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_5_clk_rst_n),
       .sr_freelist_5_addr                             (i_hqm_credit_hist_pipe_sr_freelist_5_addr),
       .sr_freelist_5_we                               (i_hqm_credit_hist_pipe_sr_freelist_5_we),
       .sr_freelist_5_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_5_wdata),
       .sr_freelist_5_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_5_rdata),
       .sr_freelist_6_re                               (i_hqm_credit_hist_pipe_sr_freelist_6_re),
       .sr_freelist_6_clk                              (i_hqm_credit_hist_pipe_sr_freelist_6_clk),
       .sr_freelist_6_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_6_clk_rst_n),
       .sr_freelist_6_addr                             (i_hqm_credit_hist_pipe_sr_freelist_6_addr),
       .sr_freelist_6_we                               (i_hqm_credit_hist_pipe_sr_freelist_6_we),
       .sr_freelist_6_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_6_wdata),
       .sr_freelist_6_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_6_rdata),
       .sr_freelist_7_re                               (i_hqm_credit_hist_pipe_sr_freelist_7_re),
       .sr_freelist_7_clk                              (i_hqm_credit_hist_pipe_sr_freelist_7_clk),
       .sr_freelist_7_clk_rst_n                        (i_hqm_credit_hist_pipe_sr_freelist_7_clk_rst_n),
       .sr_freelist_7_addr                             (i_hqm_credit_hist_pipe_sr_freelist_7_addr),
       .sr_freelist_7_we                               (i_hqm_credit_hist_pipe_sr_freelist_7_we),
       .sr_freelist_7_wdata                            (i_hqm_credit_hist_pipe_sr_freelist_7_wdata),
       .sr_freelist_7_rdata                            (i_hqm_credit_hist_pipe_sr_freelist_7_rdata),
       .sr_hist_list_re                                (i_hqm_credit_hist_pipe_sr_hist_list_re),
       .sr_hist_list_clk                               (i_hqm_credit_hist_pipe_sr_hist_list_clk),
       .sr_hist_list_clk_rst_n                         (i_hqm_credit_hist_pipe_sr_hist_list_clk_rst_n),
       .sr_hist_list_addr                              (i_hqm_credit_hist_pipe_sr_hist_list_addr),
       .sr_hist_list_we                                (i_hqm_credit_hist_pipe_sr_hist_list_we),
       .sr_hist_list_wdata                             (i_hqm_credit_hist_pipe_sr_hist_list_wdata),
       .sr_hist_list_rdata                             (i_hqm_credit_hist_pipe_sr_hist_list_rdata),
       .sr_hist_list_a_re                              (i_hqm_credit_hist_pipe_sr_hist_list_a_re),
       .sr_hist_list_a_clk                             (i_hqm_credit_hist_pipe_sr_hist_list_a_clk),
       .sr_hist_list_a_clk_rst_n                       (i_hqm_credit_hist_pipe_sr_hist_list_a_clk_rst_n),
       .sr_hist_list_a_addr                            (i_hqm_credit_hist_pipe_sr_hist_list_a_addr),
       .sr_hist_list_a_we                              (i_hqm_credit_hist_pipe_sr_hist_list_a_we),
       .sr_hist_list_a_wdata                           (i_hqm_credit_hist_pipe_sr_hist_list_a_wdata),
       .sr_hist_list_a_rdata                           (i_hqm_credit_hist_pipe_sr_hist_list_a_rdata));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_dir_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_dir),
       .hqm_gated_clk          (hqm_gated_clk_dir),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_dir),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_dir),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_dir),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_dir),
       .hqm_flr_prep           (hqm_flr_prep_rptrx),
       .rst_prep               (hqm_rst_prep_dir));

   hqm_AW_clkgate i_hqm_dp_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_dir),
       .cfg_clkungate   (hqm_clk_ungate_rptrx),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_dir));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_dp_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_dir),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_dir));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_dp_hqm_gated_clk_enable_or2
      (.clki0 (i_hqm_qed_pipe_hqm_proc_clk_en_dir),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_dir));

   hqm_AW_flop i_hqm_dp_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_gated_clk_enable_and_dir),
       .data_q (hqm_gated_clk_enable_rptr_dir));

   hqm_list_sel_pipe i_hqm_list_sel_pipe
      (.hqm_gated_clk                                      (hqm_gated_clk_lsp),
       .hqm_inp_gated_clk,
       .hqm_proc_clk_en_lsp                                (i_hqm_list_sel_pipe_hqm_proc_clk_en_lsp),
       .hqm_rst_prep_lsp,
       .hqm_gated_rst_b_lsp,
       .hqm_inp_gated_rst_b_lsp,
       .hqm_rst_prep_atm,
       .hqm_gated_rst_b_atm,
       .hqm_inp_gated_rst_b_atm,
       .hqm_gated_rst_b_start_lsp,
       .hqm_gated_rst_b_active_lsp,
       .hqm_gated_rst_b_done_lsp,
       .hqm_gated_rst_b_start_atm,
       .hqm_gated_rst_b_active_atm,
       .hqm_gated_rst_b_done_atm,
       .aqed_clk_idle,
       .aqed_unit_idle                                     (i_hqm_aqed_pipe_aqed_unit_idle),
       .aqed_clk_enable,
       .lsp_unit_idle,
       .lsp_unit_pipeidle,
       .lsp_reset_done,
       .ap_unit_idle,
       .ap_unit_pipeidle,
       .ap_reset_done,
       .lsp_cfg_req_up_read                                (i_hqm_qed_pipe_qed_cfg_req_down_read),
       .lsp_cfg_req_up_write                               (i_hqm_qed_pipe_qed_cfg_req_down_write),
       .lsp_cfg_req_up                                     (qed_cfg_req_down),
       .lsp_cfg_rsp_up_ack                                 (i_hqm_qed_pipe_qed_cfg_rsp_down_ack),
       .lsp_cfg_rsp_up                                     (qed_cfg_rsp_down),
       .lsp_cfg_req_down_read                              (i_hqm_list_sel_pipe_lsp_cfg_req_down_read),
       .lsp_cfg_req_down_write                             (i_hqm_list_sel_pipe_lsp_cfg_req_down_write),
       .lsp_cfg_req_down,
       .lsp_cfg_rsp_down_ack                               (i_hqm_list_sel_pipe_lsp_cfg_rsp_down_ack),
       .lsp_cfg_rsp_down,
       .ap_cfg_req_up_read                                 (i_hqm_list_sel_pipe_lsp_cfg_req_down_read),
       .ap_cfg_req_up_write                                (i_hqm_list_sel_pipe_lsp_cfg_req_down_write),
       .ap_cfg_req_up                                      (lsp_cfg_req_down),
       .ap_cfg_rsp_up_ack                                  (i_hqm_list_sel_pipe_lsp_cfg_rsp_down_ack),
       .ap_cfg_rsp_up                                      (lsp_cfg_rsp_down),
       .ap_cfg_req_down_read                               (i_hqm_list_sel_pipe_ap_cfg_req_down_read),
       .ap_cfg_req_down_write                              (i_hqm_list_sel_pipe_ap_cfg_req_down_write),
       .ap_cfg_req_down,
       .ap_cfg_rsp_down_ack                                (i_hqm_list_sel_pipe_ap_cfg_rsp_down_ack),
       .ap_cfg_rsp_down,
       .lsp_alarm_up_v                                     (i_hqm_list_sel_pipe_ap_alarm_down_v),
       .lsp_alarm_up_ready                                 (i_hqm_list_sel_pipe_lsp_alarm_up_ready),
       .lsp_alarm_up_data                                  (ap_alarm_down_data),
       .lsp_alarm_down_v                                   (i_hqm_list_sel_pipe_lsp_alarm_down_v),
       .lsp_alarm_down_ready                               (i_hqm_qed_pipe_qed_alarm_up_ready),
       .lsp_alarm_down_data,
       .ap_alarm_up_v                                      (i_hqm_aqed_pipe_aqed_alarm_down_v),
       .ap_alarm_up_ready                                  (i_hqm_list_sel_pipe_ap_alarm_up_ready),
       .ap_alarm_up_data                                   (aqed_alarm_down_data),
       .ap_alarm_down_v                                    (i_hqm_list_sel_pipe_ap_alarm_down_v),
       .ap_alarm_down_ready                                (i_hqm_list_sel_pipe_lsp_alarm_up_ready),
       .ap_alarm_down_data,
       .lsp_aqed_cmp_v,
       .lsp_aqed_cmp_ready,
       .lsp_aqed_cmp_data,
       .aqed_lsp_dec_fid_cnt_v,
       .chp_lsp_ldb_cq_off,
       .chp_lsp_cmp_v                                      (i_hqm_credit_hist_pipe_chp_lsp_cmp_v),
       .chp_lsp_cmp_ready                                  (i_hqm_list_sel_pipe_chp_lsp_cmp_ready),
       .chp_lsp_cmp_data,
       .qed_lsp_deq_v,
       .qed_lsp_deq_data,
       .aqed_lsp_deq_v,
       .aqed_lsp_deq_data,
       .chp_lsp_token_v                                    (i_hqm_credit_hist_pipe_chp_lsp_token_v),
       .chp_lsp_token_ready                                (i_hqm_list_sel_pipe_chp_lsp_token_ready),
       .chp_lsp_token_data,
       .lsp_nalb_sch_unoord_v                              (i_hqm_list_sel_pipe_lsp_nalb_sch_unoord_v),
       .lsp_nalb_sch_unoord_ready                          (i_hqm_qed_pipe_lsp_nalb_sch_unoord_ready),
       .lsp_nalb_sch_unoord_data,
       .lsp_dp_sch_dir_v                                   (i_hqm_list_sel_pipe_lsp_dp_sch_dir_v),
       .lsp_dp_sch_dir_ready                               (i_hqm_qed_pipe_lsp_dp_sch_dir_ready),
       .lsp_dp_sch_dir_data,
       .lsp_nalb_sch_rorply_v                              (i_hqm_list_sel_pipe_lsp_nalb_sch_rorply_v),
       .lsp_nalb_sch_rorply_ready                          (i_hqm_qed_pipe_lsp_nalb_sch_rorply_ready),
       .lsp_nalb_sch_rorply_data,
       .lsp_dp_sch_rorply_v                                (i_hqm_list_sel_pipe_lsp_dp_sch_rorply_v),
       .lsp_dp_sch_rorply_ready                            (i_hqm_qed_pipe_lsp_dp_sch_rorply_ready),
       .lsp_dp_sch_rorply_data,
       .lsp_nalb_sch_atq_v                                 (i_hqm_list_sel_pipe_lsp_nalb_sch_atq_v),
       .lsp_nalb_sch_atq_ready                             (i_hqm_qed_pipe_lsp_nalb_sch_atq_ready),
       .lsp_nalb_sch_atq_data,
       .nalb_lsp_enq_lb_v                                  (i_hqm_qed_pipe_nalb_lsp_enq_lb_v),
       .nalb_lsp_enq_lb_ready                              (i_hqm_list_sel_pipe_nalb_lsp_enq_lb_ready),
       .nalb_lsp_enq_lb_data,
       .nalb_lsp_enq_rorply_v                              (i_hqm_qed_pipe_nalb_lsp_enq_rorply_v),
       .nalb_lsp_enq_rorply_ready                          (i_hqm_list_sel_pipe_nalb_lsp_enq_rorply_ready),
       .nalb_lsp_enq_rorply_data,
       .dp_lsp_enq_dir_v                                   (i_hqm_qed_pipe_dp_lsp_enq_dir_v),
       .dp_lsp_enq_dir_ready                               (i_hqm_list_sel_pipe_dp_lsp_enq_dir_ready),
       .dp_lsp_enq_dir_data,
       .dp_lsp_enq_rorply_v                                (i_hqm_qed_pipe_dp_lsp_enq_rorply_v),
       .dp_lsp_enq_rorply_ready                            (i_hqm_list_sel_pipe_dp_lsp_enq_rorply_ready),
       .dp_lsp_enq_rorply_data,
       .rop_lsp_reordercmp_v                               (i_hqm_reorder_pipe_rop_lsp_reordercmp_v),
       .rop_lsp_reordercmp_ready                           (i_hqm_list_sel_pipe_rop_lsp_reordercmp_ready),
       .rop_lsp_reordercmp_data,
       .aqed_lsp_sch_v                                     (i_hqm_aqed_pipe_aqed_lsp_sch_v),
       .aqed_lsp_sch_ready                                 (i_hqm_list_sel_pipe_aqed_lsp_sch_ready),
       .aqed_lsp_sch_data,
       .ap_aqed_v                                          (i_hqm_list_sel_pipe_ap_aqed_v),
       .ap_aqed_ready                                      (i_hqm_aqed_pipe_ap_aqed_ready),
       .ap_aqed_data,
       .aqed_ap_enq_v                                      (i_hqm_aqed_pipe_aqed_ap_enq_v),
       .aqed_ap_enq_ready                                  (i_hqm_list_sel_pipe_aqed_ap_enq_ready),
       .aqed_ap_enq_data,
       .aqed_lsp_fid_cnt_upd_v,
       .aqed_lsp_fid_cnt_upd_val,
       .aqed_lsp_fid_cnt_upd_qid,
       .aqed_lsp_stop_atqatm,
       .spare_qed_lsp,
       .spare_sys_lsp,
       .spare_lsp_qed,
       .spare_lsp_sys,
       .rf_aqed_lsp_deq_fifo_mem_re                        (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_re),
       .rf_aqed_lsp_deq_fifo_mem_rclk                      (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rclk),
       .rf_aqed_lsp_deq_fifo_mem_rclk_rst_n                (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rclk_rst_n),
       .rf_aqed_lsp_deq_fifo_mem_raddr                     (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_raddr),
       .rf_aqed_lsp_deq_fifo_mem_waddr                     (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_waddr),
       .rf_aqed_lsp_deq_fifo_mem_we                        (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_we),
       .rf_aqed_lsp_deq_fifo_mem_wclk                      (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wclk),
       .rf_aqed_lsp_deq_fifo_mem_wclk_rst_n                (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wclk_rst_n),
       .rf_aqed_lsp_deq_fifo_mem_wdata                     (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_wdata),
       .rf_aqed_lsp_deq_fifo_mem_rdata                     (i_hqm_list_sel_pipe_rf_aqed_lsp_deq_fifo_mem_rdata),
       .rf_atm_cmp_fifo_mem_re                             (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_re),
       .rf_atm_cmp_fifo_mem_rclk                           (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rclk),
       .rf_atm_cmp_fifo_mem_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rclk_rst_n),
       .rf_atm_cmp_fifo_mem_raddr                          (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_raddr),
       .rf_atm_cmp_fifo_mem_waddr                          (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_waddr),
       .rf_atm_cmp_fifo_mem_we                             (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_we),
       .rf_atm_cmp_fifo_mem_wclk                           (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wclk),
       .rf_atm_cmp_fifo_mem_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wclk_rst_n),
       .rf_atm_cmp_fifo_mem_wdata                          (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_wdata),
       .rf_atm_cmp_fifo_mem_rdata                          (i_hqm_list_sel_pipe_rf_atm_cmp_fifo_mem_rdata),
       .rf_cfg_atm_qid_dpth_thrsh_mem_re                   (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_re),
       .rf_cfg_atm_qid_dpth_thrsh_mem_rclk                 (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rclk),
       .rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rclk_rst_n),
       .rf_cfg_atm_qid_dpth_thrsh_mem_raddr                (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_raddr),
       .rf_cfg_atm_qid_dpth_thrsh_mem_waddr                (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_waddr),
       .rf_cfg_atm_qid_dpth_thrsh_mem_we                   (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_we),
       .rf_cfg_atm_qid_dpth_thrsh_mem_wclk                 (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wclk),
       .rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wclk_rst_n),
       .rf_cfg_atm_qid_dpth_thrsh_mem_wdata                (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_wdata),
       .rf_cfg_atm_qid_dpth_thrsh_mem_rdata                (i_hqm_list_sel_pipe_rf_cfg_atm_qid_dpth_thrsh_mem_rdata),
       .rf_cfg_cq2priov_mem_re                             (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_re),
       .rf_cfg_cq2priov_mem_rclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rclk),
       .rf_cfg_cq2priov_mem_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rclk_rst_n),
       .rf_cfg_cq2priov_mem_raddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_raddr),
       .rf_cfg_cq2priov_mem_waddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_waddr),
       .rf_cfg_cq2priov_mem_we                             (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_we),
       .rf_cfg_cq2priov_mem_wclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wclk),
       .rf_cfg_cq2priov_mem_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wclk_rst_n),
       .rf_cfg_cq2priov_mem_wdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_wdata),
       .rf_cfg_cq2priov_mem_rdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2priov_mem_rdata),
       .rf_cfg_cq2priov_odd_mem_re                         (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_re),
       .rf_cfg_cq2priov_odd_mem_rclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rclk),
       .rf_cfg_cq2priov_odd_mem_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rclk_rst_n),
       .rf_cfg_cq2priov_odd_mem_raddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_raddr),
       .rf_cfg_cq2priov_odd_mem_waddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_waddr),
       .rf_cfg_cq2priov_odd_mem_we                         (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_we),
       .rf_cfg_cq2priov_odd_mem_wclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wclk),
       .rf_cfg_cq2priov_odd_mem_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wclk_rst_n),
       .rf_cfg_cq2priov_odd_mem_wdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_wdata),
       .rf_cfg_cq2priov_odd_mem_rdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2priov_odd_mem_rdata),
       .rf_cfg_cq2qid_0_mem_re                             (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_re),
       .rf_cfg_cq2qid_0_mem_rclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rclk),
       .rf_cfg_cq2qid_0_mem_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rclk_rst_n),
       .rf_cfg_cq2qid_0_mem_raddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_raddr),
       .rf_cfg_cq2qid_0_mem_waddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_waddr),
       .rf_cfg_cq2qid_0_mem_we                             (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_we),
       .rf_cfg_cq2qid_0_mem_wclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wclk),
       .rf_cfg_cq2qid_0_mem_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wclk_rst_n),
       .rf_cfg_cq2qid_0_mem_wdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_wdata),
       .rf_cfg_cq2qid_0_mem_rdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_mem_rdata),
       .rf_cfg_cq2qid_0_odd_mem_re                         (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_re),
       .rf_cfg_cq2qid_0_odd_mem_rclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rclk),
       .rf_cfg_cq2qid_0_odd_mem_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rclk_rst_n),
       .rf_cfg_cq2qid_0_odd_mem_raddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_raddr),
       .rf_cfg_cq2qid_0_odd_mem_waddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_waddr),
       .rf_cfg_cq2qid_0_odd_mem_we                         (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_we),
       .rf_cfg_cq2qid_0_odd_mem_wclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wclk),
       .rf_cfg_cq2qid_0_odd_mem_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wclk_rst_n),
       .rf_cfg_cq2qid_0_odd_mem_wdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_wdata),
       .rf_cfg_cq2qid_0_odd_mem_rdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_0_odd_mem_rdata),
       .rf_cfg_cq2qid_1_mem_re                             (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_re),
       .rf_cfg_cq2qid_1_mem_rclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rclk),
       .rf_cfg_cq2qid_1_mem_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rclk_rst_n),
       .rf_cfg_cq2qid_1_mem_raddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_raddr),
       .rf_cfg_cq2qid_1_mem_waddr                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_waddr),
       .rf_cfg_cq2qid_1_mem_we                             (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_we),
       .rf_cfg_cq2qid_1_mem_wclk                           (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wclk),
       .rf_cfg_cq2qid_1_mem_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wclk_rst_n),
       .rf_cfg_cq2qid_1_mem_wdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_wdata),
       .rf_cfg_cq2qid_1_mem_rdata                          (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_mem_rdata),
       .rf_cfg_cq2qid_1_odd_mem_re                         (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_re),
       .rf_cfg_cq2qid_1_odd_mem_rclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rclk),
       .rf_cfg_cq2qid_1_odd_mem_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rclk_rst_n),
       .rf_cfg_cq2qid_1_odd_mem_raddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_raddr),
       .rf_cfg_cq2qid_1_odd_mem_waddr                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_waddr),
       .rf_cfg_cq2qid_1_odd_mem_we                         (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_we),
       .rf_cfg_cq2qid_1_odd_mem_wclk                       (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wclk),
       .rf_cfg_cq2qid_1_odd_mem_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wclk_rst_n),
       .rf_cfg_cq2qid_1_odd_mem_wdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_wdata),
       .rf_cfg_cq2qid_1_odd_mem_rdata                      (i_hqm_list_sel_pipe_rf_cfg_cq2qid_1_odd_mem_rdata),
       .rf_cfg_cq_ldb_inflight_limit_mem_re                (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_re),
       .rf_cfg_cq_ldb_inflight_limit_mem_rclk              (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rclk),
       .rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n        (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rclk_rst_n),
       .rf_cfg_cq_ldb_inflight_limit_mem_raddr             (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_raddr),
       .rf_cfg_cq_ldb_inflight_limit_mem_waddr             (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_waddr),
       .rf_cfg_cq_ldb_inflight_limit_mem_we                (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_we),
       .rf_cfg_cq_ldb_inflight_limit_mem_wclk              (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wclk),
       .rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n        (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wclk_rst_n),
       .rf_cfg_cq_ldb_inflight_limit_mem_wdata             (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_wdata),
       .rf_cfg_cq_ldb_inflight_limit_mem_rdata             (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_limit_mem_rdata),
       .rf_cfg_cq_ldb_inflight_threshold_mem_re            (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_re),
       .rf_cfg_cq_ldb_inflight_threshold_mem_rclk          (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rclk),
       .rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rclk_rst_n),
       .rf_cfg_cq_ldb_inflight_threshold_mem_raddr         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_raddr),
       .rf_cfg_cq_ldb_inflight_threshold_mem_waddr         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_waddr),
       .rf_cfg_cq_ldb_inflight_threshold_mem_we            (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_we),
       .rf_cfg_cq_ldb_inflight_threshold_mem_wclk          (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wclk),
       .rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wclk_rst_n),
       .rf_cfg_cq_ldb_inflight_threshold_mem_wdata         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_wdata),
       .rf_cfg_cq_ldb_inflight_threshold_mem_rdata         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_inflight_threshold_mem_rdata),
       .rf_cfg_cq_ldb_token_depth_select_mem_re            (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_re),
       .rf_cfg_cq_ldb_token_depth_select_mem_rclk          (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rclk),
       .rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rclk_rst_n),
       .rf_cfg_cq_ldb_token_depth_select_mem_raddr         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_raddr),
       .rf_cfg_cq_ldb_token_depth_select_mem_waddr         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_waddr),
       .rf_cfg_cq_ldb_token_depth_select_mem_we            (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_we),
       .rf_cfg_cq_ldb_token_depth_select_mem_wclk          (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wclk),
       .rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wclk_rst_n),
       .rf_cfg_cq_ldb_token_depth_select_mem_wdata         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_wdata),
       .rf_cfg_cq_ldb_token_depth_select_mem_rdata         (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_token_depth_select_mem_rdata),
       .rf_cfg_cq_ldb_wu_limit_mem_re                      (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_re),
       .rf_cfg_cq_ldb_wu_limit_mem_rclk                    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rclk),
       .rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n              (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rclk_rst_n),
       .rf_cfg_cq_ldb_wu_limit_mem_raddr                   (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_raddr),
       .rf_cfg_cq_ldb_wu_limit_mem_waddr                   (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_waddr),
       .rf_cfg_cq_ldb_wu_limit_mem_we                      (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_we),
       .rf_cfg_cq_ldb_wu_limit_mem_wclk                    (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wclk),
       .rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n              (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wclk_rst_n),
       .rf_cfg_cq_ldb_wu_limit_mem_wdata                   (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_wdata),
       .rf_cfg_cq_ldb_wu_limit_mem_rdata                   (i_hqm_list_sel_pipe_rf_cfg_cq_ldb_wu_limit_mem_rdata),
       .rf_cfg_dir_qid_dpth_thrsh_mem_re                   (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_re),
       .rf_cfg_dir_qid_dpth_thrsh_mem_rclk                 (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rclk),
       .rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rclk_rst_n),
       .rf_cfg_dir_qid_dpth_thrsh_mem_raddr                (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_raddr),
       .rf_cfg_dir_qid_dpth_thrsh_mem_waddr                (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_waddr),
       .rf_cfg_dir_qid_dpth_thrsh_mem_we                   (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_we),
       .rf_cfg_dir_qid_dpth_thrsh_mem_wclk                 (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wclk),
       .rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wclk_rst_n),
       .rf_cfg_dir_qid_dpth_thrsh_mem_wdata                (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_wdata),
       .rf_cfg_dir_qid_dpth_thrsh_mem_rdata                (i_hqm_list_sel_pipe_rf_cfg_dir_qid_dpth_thrsh_mem_rdata),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_re                  (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_re),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_rclk                (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rclk),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n          (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rclk_rst_n),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_raddr               (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_raddr),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_waddr               (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_waddr),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_we                  (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_we),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_wclk                (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wclk),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n          (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wclk_rst_n),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_wdata               (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_wdata),
       .rf_cfg_nalb_qid_dpth_thrsh_mem_rdata               (i_hqm_list_sel_pipe_rf_cfg_nalb_qid_dpth_thrsh_mem_rdata),
       .rf_cfg_qid_aqed_active_limit_mem_re                (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_re),
       .rf_cfg_qid_aqed_active_limit_mem_rclk              (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rclk),
       .rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n        (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rclk_rst_n),
       .rf_cfg_qid_aqed_active_limit_mem_raddr             (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_raddr),
       .rf_cfg_qid_aqed_active_limit_mem_waddr             (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_waddr),
       .rf_cfg_qid_aqed_active_limit_mem_we                (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_we),
       .rf_cfg_qid_aqed_active_limit_mem_wclk              (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wclk),
       .rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n        (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wclk_rst_n),
       .rf_cfg_qid_aqed_active_limit_mem_wdata             (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_wdata),
       .rf_cfg_qid_aqed_active_limit_mem_rdata             (i_hqm_list_sel_pipe_rf_cfg_qid_aqed_active_limit_mem_rdata),
       .rf_cfg_qid_ldb_inflight_limit_mem_re               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_re),
       .rf_cfg_qid_ldb_inflight_limit_mem_rclk             (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rclk),
       .rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n       (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rclk_rst_n),
       .rf_cfg_qid_ldb_inflight_limit_mem_raddr            (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_raddr),
       .rf_cfg_qid_ldb_inflight_limit_mem_waddr            (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_waddr),
       .rf_cfg_qid_ldb_inflight_limit_mem_we               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_we),
       .rf_cfg_qid_ldb_inflight_limit_mem_wclk             (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wclk),
       .rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n       (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wclk_rst_n),
       .rf_cfg_qid_ldb_inflight_limit_mem_wdata            (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_wdata),
       .rf_cfg_qid_ldb_inflight_limit_mem_rdata            (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_inflight_limit_mem_rdata),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_re                  (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_re),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_rclk                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rclk),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n          (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rclk_rst_n),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_raddr               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_raddr),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_waddr               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_waddr),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_we                  (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_we),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_wclk                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wclk),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n          (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wclk_rst_n),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_wdata               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_wdata),
       .rf_cfg_qid_ldb_qid2cqidix2_mem_rdata               (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix2_mem_rdata),
       .rf_cfg_qid_ldb_qid2cqidix_mem_re                   (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_re),
       .rf_cfg_qid_ldb_qid2cqidix_mem_rclk                 (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rclk),
       .rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rclk_rst_n),
       .rf_cfg_qid_ldb_qid2cqidix_mem_raddr                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_raddr),
       .rf_cfg_qid_ldb_qid2cqidix_mem_waddr                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_waddr),
       .rf_cfg_qid_ldb_qid2cqidix_mem_we                   (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_we),
       .rf_cfg_qid_ldb_qid2cqidix_mem_wclk                 (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wclk),
       .rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n           (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wclk_rst_n),
       .rf_cfg_qid_ldb_qid2cqidix_mem_wdata                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_wdata),
       .rf_cfg_qid_ldb_qid2cqidix_mem_rdata                (i_hqm_list_sel_pipe_rf_cfg_qid_ldb_qid2cqidix_mem_rdata),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_re                 (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_re),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk               (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n         (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rclk_rst_n),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr              (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_raddr),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr              (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_waddr),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_we                 (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_we),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk               (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n         (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wclk_rst_n),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata              (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_wdata),
       .rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata              (i_hqm_list_sel_pipe_rf_chp_lsp_cmp_rx_sync_fifo_mem_rdata),
       .rf_chp_lsp_token_rx_sync_fifo_mem_re               (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_re),
       .rf_chp_lsp_token_rx_sync_fifo_mem_rclk             (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rclk),
       .rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n       (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rclk_rst_n),
       .rf_chp_lsp_token_rx_sync_fifo_mem_raddr            (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_raddr),
       .rf_chp_lsp_token_rx_sync_fifo_mem_waddr            (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_waddr),
       .rf_chp_lsp_token_rx_sync_fifo_mem_we               (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_we),
       .rf_chp_lsp_token_rx_sync_fifo_mem_wclk             (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wclk),
       .rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n       (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wclk_rst_n),
       .rf_chp_lsp_token_rx_sync_fifo_mem_wdata            (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_wdata),
       .rf_chp_lsp_token_rx_sync_fifo_mem_rdata            (i_hqm_list_sel_pipe_rf_chp_lsp_token_rx_sync_fifo_mem_rdata),
       .rf_cq_atm_pri_arbindex_mem_re                      (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_re),
       .rf_cq_atm_pri_arbindex_mem_rclk                    (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rclk),
       .rf_cq_atm_pri_arbindex_mem_rclk_rst_n              (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rclk_rst_n),
       .rf_cq_atm_pri_arbindex_mem_raddr                   (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_raddr),
       .rf_cq_atm_pri_arbindex_mem_waddr                   (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_waddr),
       .rf_cq_atm_pri_arbindex_mem_we                      (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_we),
       .rf_cq_atm_pri_arbindex_mem_wclk                    (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wclk),
       .rf_cq_atm_pri_arbindex_mem_wclk_rst_n              (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wclk_rst_n),
       .rf_cq_atm_pri_arbindex_mem_wdata                   (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_wdata),
       .rf_cq_atm_pri_arbindex_mem_rdata                   (i_hqm_list_sel_pipe_rf_cq_atm_pri_arbindex_mem_rdata),
       .rf_cq_dir_tot_sch_cnt_mem_re                       (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_re),
       .rf_cq_dir_tot_sch_cnt_mem_rclk                     (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rclk),
       .rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rclk_rst_n),
       .rf_cq_dir_tot_sch_cnt_mem_raddr                    (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_raddr),
       .rf_cq_dir_tot_sch_cnt_mem_waddr                    (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_waddr),
       .rf_cq_dir_tot_sch_cnt_mem_we                       (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_we),
       .rf_cq_dir_tot_sch_cnt_mem_wclk                     (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wclk),
       .rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wclk_rst_n),
       .rf_cq_dir_tot_sch_cnt_mem_wdata                    (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_wdata),
       .rf_cq_dir_tot_sch_cnt_mem_rdata                    (i_hqm_list_sel_pipe_rf_cq_dir_tot_sch_cnt_mem_rdata),
       .rf_cq_ldb_inflight_count_mem_re                    (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_re),
       .rf_cq_ldb_inflight_count_mem_rclk                  (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rclk),
       .rf_cq_ldb_inflight_count_mem_rclk_rst_n            (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rclk_rst_n),
       .rf_cq_ldb_inflight_count_mem_raddr                 (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_raddr),
       .rf_cq_ldb_inflight_count_mem_waddr                 (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_waddr),
       .rf_cq_ldb_inflight_count_mem_we                    (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_we),
       .rf_cq_ldb_inflight_count_mem_wclk                  (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wclk),
       .rf_cq_ldb_inflight_count_mem_wclk_rst_n            (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wclk_rst_n),
       .rf_cq_ldb_inflight_count_mem_wdata                 (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_wdata),
       .rf_cq_ldb_inflight_count_mem_rdata                 (i_hqm_list_sel_pipe_rf_cq_ldb_inflight_count_mem_rdata),
       .rf_cq_ldb_token_count_mem_re                       (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_re),
       .rf_cq_ldb_token_count_mem_rclk                     (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rclk),
       .rf_cq_ldb_token_count_mem_rclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rclk_rst_n),
       .rf_cq_ldb_token_count_mem_raddr                    (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_raddr),
       .rf_cq_ldb_token_count_mem_waddr                    (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_waddr),
       .rf_cq_ldb_token_count_mem_we                       (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_we),
       .rf_cq_ldb_token_count_mem_wclk                     (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wclk),
       .rf_cq_ldb_token_count_mem_wclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wclk_rst_n),
       .rf_cq_ldb_token_count_mem_wdata                    (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_wdata),
       .rf_cq_ldb_token_count_mem_rdata                    (i_hqm_list_sel_pipe_rf_cq_ldb_token_count_mem_rdata),
       .rf_cq_ldb_tot_sch_cnt_mem_re                       (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_re),
       .rf_cq_ldb_tot_sch_cnt_mem_rclk                     (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rclk),
       .rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rclk_rst_n),
       .rf_cq_ldb_tot_sch_cnt_mem_raddr                    (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_raddr),
       .rf_cq_ldb_tot_sch_cnt_mem_waddr                    (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_waddr),
       .rf_cq_ldb_tot_sch_cnt_mem_we                       (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_we),
       .rf_cq_ldb_tot_sch_cnt_mem_wclk                     (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wclk),
       .rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n               (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wclk_rst_n),
       .rf_cq_ldb_tot_sch_cnt_mem_wdata                    (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_wdata),
       .rf_cq_ldb_tot_sch_cnt_mem_rdata                    (i_hqm_list_sel_pipe_rf_cq_ldb_tot_sch_cnt_mem_rdata),
       .rf_cq_ldb_wu_count_mem_re                          (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_re),
       .rf_cq_ldb_wu_count_mem_rclk                        (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rclk),
       .rf_cq_ldb_wu_count_mem_rclk_rst_n                  (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rclk_rst_n),
       .rf_cq_ldb_wu_count_mem_raddr                       (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_raddr),
       .rf_cq_ldb_wu_count_mem_waddr                       (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_waddr),
       .rf_cq_ldb_wu_count_mem_we                          (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_we),
       .rf_cq_ldb_wu_count_mem_wclk                        (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wclk),
       .rf_cq_ldb_wu_count_mem_wclk_rst_n                  (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wclk_rst_n),
       .rf_cq_ldb_wu_count_mem_wdata                       (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_wdata),
       .rf_cq_ldb_wu_count_mem_rdata                       (i_hqm_list_sel_pipe_rf_cq_ldb_wu_count_mem_rdata),
       .rf_cq_nalb_pri_arbindex_mem_re                     (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_re),
       .rf_cq_nalb_pri_arbindex_mem_rclk                   (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rclk),
       .rf_cq_nalb_pri_arbindex_mem_rclk_rst_n             (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rclk_rst_n),
       .rf_cq_nalb_pri_arbindex_mem_raddr                  (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_raddr),
       .rf_cq_nalb_pri_arbindex_mem_waddr                  (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_waddr),
       .rf_cq_nalb_pri_arbindex_mem_we                     (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_we),
       .rf_cq_nalb_pri_arbindex_mem_wclk                   (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wclk),
       .rf_cq_nalb_pri_arbindex_mem_wclk_rst_n             (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wclk_rst_n),
       .rf_cq_nalb_pri_arbindex_mem_wdata                  (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_wdata),
       .rf_cq_nalb_pri_arbindex_mem_rdata                  (i_hqm_list_sel_pipe_rf_cq_nalb_pri_arbindex_mem_rdata),
       .rf_dir_enq_cnt_mem_re                              (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_re),
       .rf_dir_enq_cnt_mem_rclk                            (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rclk),
       .rf_dir_enq_cnt_mem_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rclk_rst_n),
       .rf_dir_enq_cnt_mem_raddr                           (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_raddr),
       .rf_dir_enq_cnt_mem_waddr                           (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_waddr),
       .rf_dir_enq_cnt_mem_we                              (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_we),
       .rf_dir_enq_cnt_mem_wclk                            (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wclk),
       .rf_dir_enq_cnt_mem_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wclk_rst_n),
       .rf_dir_enq_cnt_mem_wdata                           (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_wdata),
       .rf_dir_enq_cnt_mem_rdata                           (i_hqm_list_sel_pipe_rf_dir_enq_cnt_mem_rdata),
       .rf_dir_tok_cnt_mem_re                              (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_re),
       .rf_dir_tok_cnt_mem_rclk                            (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rclk),
       .rf_dir_tok_cnt_mem_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rclk_rst_n),
       .rf_dir_tok_cnt_mem_raddr                           (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_raddr),
       .rf_dir_tok_cnt_mem_waddr                           (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_waddr),
       .rf_dir_tok_cnt_mem_we                              (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_we),
       .rf_dir_tok_cnt_mem_wclk                            (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wclk),
       .rf_dir_tok_cnt_mem_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wclk_rst_n),
       .rf_dir_tok_cnt_mem_wdata                           (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_wdata),
       .rf_dir_tok_cnt_mem_rdata                           (i_hqm_list_sel_pipe_rf_dir_tok_cnt_mem_rdata),
       .rf_dir_tok_lim_mem_re                              (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_re),
       .rf_dir_tok_lim_mem_rclk                            (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rclk),
       .rf_dir_tok_lim_mem_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rclk_rst_n),
       .rf_dir_tok_lim_mem_raddr                           (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_raddr),
       .rf_dir_tok_lim_mem_waddr                           (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_waddr),
       .rf_dir_tok_lim_mem_we                              (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_we),
       .rf_dir_tok_lim_mem_wclk                            (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wclk),
       .rf_dir_tok_lim_mem_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wclk_rst_n),
       .rf_dir_tok_lim_mem_wdata                           (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_wdata),
       .rf_dir_tok_lim_mem_rdata                           (i_hqm_list_sel_pipe_rf_dir_tok_lim_mem_rdata),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re              (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_re),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk            (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n      (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rclk_rst_n),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_raddr),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_waddr),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we              (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_we),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk            (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n      (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wclk_rst_n),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_wdata),
       .rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_dir_rx_sync_fifo_mem_rdata),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_re),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk         (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n   (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr        (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_raddr),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr        (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_waddr),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we           (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_we),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk         (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n   (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata        (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_wdata),
       .rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata        (i_hqm_list_sel_pipe_rf_dp_lsp_enq_rorply_rx_sync_fifo_mem_rdata),
       .rf_enq_nalb_fifo_mem_re                            (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_re),
       .rf_enq_nalb_fifo_mem_rclk                          (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rclk),
       .rf_enq_nalb_fifo_mem_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rclk_rst_n),
       .rf_enq_nalb_fifo_mem_raddr                         (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_raddr),
       .rf_enq_nalb_fifo_mem_waddr                         (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_waddr),
       .rf_enq_nalb_fifo_mem_we                            (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_we),
       .rf_enq_nalb_fifo_mem_wclk                          (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wclk),
       .rf_enq_nalb_fifo_mem_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wclk_rst_n),
       .rf_enq_nalb_fifo_mem_wdata                         (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_wdata),
       .rf_enq_nalb_fifo_mem_rdata                         (i_hqm_list_sel_pipe_rf_enq_nalb_fifo_mem_rdata),
       .rf_ldb_token_rtn_fifo_mem_re                       (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_re),
       .rf_ldb_token_rtn_fifo_mem_rclk                     (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rclk),
       .rf_ldb_token_rtn_fifo_mem_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rclk_rst_n),
       .rf_ldb_token_rtn_fifo_mem_raddr                    (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_raddr),
       .rf_ldb_token_rtn_fifo_mem_waddr                    (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_waddr),
       .rf_ldb_token_rtn_fifo_mem_we                       (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_we),
       .rf_ldb_token_rtn_fifo_mem_wclk                     (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wclk),
       .rf_ldb_token_rtn_fifo_mem_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wclk_rst_n),
       .rf_ldb_token_rtn_fifo_mem_wdata                    (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_wdata),
       .rf_ldb_token_rtn_fifo_mem_rdata                    (i_hqm_list_sel_pipe_rf_ldb_token_rtn_fifo_mem_rdata),
       .rf_nalb_cmp_fifo_mem_re                            (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_re),
       .rf_nalb_cmp_fifo_mem_rclk                          (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rclk),
       .rf_nalb_cmp_fifo_mem_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rclk_rst_n),
       .rf_nalb_cmp_fifo_mem_raddr                         (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_raddr),
       .rf_nalb_cmp_fifo_mem_waddr                         (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_waddr),
       .rf_nalb_cmp_fifo_mem_we                            (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_we),
       .rf_nalb_cmp_fifo_mem_wclk                          (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wclk),
       .rf_nalb_cmp_fifo_mem_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wclk_rst_n),
       .rf_nalb_cmp_fifo_mem_wdata                         (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_wdata),
       .rf_nalb_cmp_fifo_mem_rdata                         (i_hqm_list_sel_pipe_rf_nalb_cmp_fifo_mem_rdata),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re             (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_re),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk           (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n     (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rclk_rst_n),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr          (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_raddr),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr          (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_waddr),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we             (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_we),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk           (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n     (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wclk_rst_n),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata          (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_wdata),
       .rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata          (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_lb_rx_sync_fifo_mem_rdata),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re         (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_re),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk       (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rclk_rst_n),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr      (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_raddr),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr      (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_waddr),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we         (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_we),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk       (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wclk_rst_n),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata      (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_wdata),
       .rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata      (i_hqm_list_sel_pipe_rf_nalb_lsp_enq_rorply_rx_sync_fifo_mem_rdata),
       .rf_nalb_sel_nalb_fifo_mem_re                       (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_re),
       .rf_nalb_sel_nalb_fifo_mem_rclk                     (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rclk),
       .rf_nalb_sel_nalb_fifo_mem_rclk_rst_n               (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rclk_rst_n),
       .rf_nalb_sel_nalb_fifo_mem_raddr                    (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_raddr),
       .rf_nalb_sel_nalb_fifo_mem_waddr                    (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_waddr),
       .rf_nalb_sel_nalb_fifo_mem_we                       (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_we),
       .rf_nalb_sel_nalb_fifo_mem_wclk                     (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wclk),
       .rf_nalb_sel_nalb_fifo_mem_wclk_rst_n               (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wclk_rst_n),
       .rf_nalb_sel_nalb_fifo_mem_wdata                    (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_wdata),
       .rf_nalb_sel_nalb_fifo_mem_rdata                    (i_hqm_list_sel_pipe_rf_nalb_sel_nalb_fifo_mem_rdata),
       .rf_qed_lsp_deq_fifo_mem_re                         (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_re),
       .rf_qed_lsp_deq_fifo_mem_rclk                       (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rclk),
       .rf_qed_lsp_deq_fifo_mem_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rclk_rst_n),
       .rf_qed_lsp_deq_fifo_mem_raddr                      (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_raddr),
       .rf_qed_lsp_deq_fifo_mem_waddr                      (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_waddr),
       .rf_qed_lsp_deq_fifo_mem_we                         (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_we),
       .rf_qed_lsp_deq_fifo_mem_wclk                       (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wclk),
       .rf_qed_lsp_deq_fifo_mem_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wclk_rst_n),
       .rf_qed_lsp_deq_fifo_mem_wdata                      (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_wdata),
       .rf_qed_lsp_deq_fifo_mem_rdata                      (i_hqm_list_sel_pipe_rf_qed_lsp_deq_fifo_mem_rdata),
       .rf_qid_aqed_active_count_mem_re                    (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_re),
       .rf_qid_aqed_active_count_mem_rclk                  (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rclk),
       .rf_qid_aqed_active_count_mem_rclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rclk_rst_n),
       .rf_qid_aqed_active_count_mem_raddr                 (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_raddr),
       .rf_qid_aqed_active_count_mem_waddr                 (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_waddr),
       .rf_qid_aqed_active_count_mem_we                    (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_we),
       .rf_qid_aqed_active_count_mem_wclk                  (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wclk),
       .rf_qid_aqed_active_count_mem_wclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wclk_rst_n),
       .rf_qid_aqed_active_count_mem_wdata                 (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_wdata),
       .rf_qid_aqed_active_count_mem_rdata                 (i_hqm_list_sel_pipe_rf_qid_aqed_active_count_mem_rdata),
       .rf_qid_atm_active_mem_re                           (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_re),
       .rf_qid_atm_active_mem_rclk                         (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rclk),
       .rf_qid_atm_active_mem_rclk_rst_n                   (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rclk_rst_n),
       .rf_qid_atm_active_mem_raddr                        (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_raddr),
       .rf_qid_atm_active_mem_waddr                        (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_waddr),
       .rf_qid_atm_active_mem_we                           (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_we),
       .rf_qid_atm_active_mem_wclk                         (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wclk),
       .rf_qid_atm_active_mem_wclk_rst_n                   (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wclk_rst_n),
       .rf_qid_atm_active_mem_wdata                        (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_wdata),
       .rf_qid_atm_active_mem_rdata                        (i_hqm_list_sel_pipe_rf_qid_atm_active_mem_rdata),
       .rf_qid_atm_tot_enq_cnt_mem_re                      (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_re),
       .rf_qid_atm_tot_enq_cnt_mem_rclk                    (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rclk),
       .rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rclk_rst_n),
       .rf_qid_atm_tot_enq_cnt_mem_raddr                   (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_raddr),
       .rf_qid_atm_tot_enq_cnt_mem_waddr                   (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_waddr),
       .rf_qid_atm_tot_enq_cnt_mem_we                      (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_we),
       .rf_qid_atm_tot_enq_cnt_mem_wclk                    (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wclk),
       .rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wclk_rst_n),
       .rf_qid_atm_tot_enq_cnt_mem_wdata                   (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_wdata),
       .rf_qid_atm_tot_enq_cnt_mem_rdata                   (i_hqm_list_sel_pipe_rf_qid_atm_tot_enq_cnt_mem_rdata),
       .rf_qid_atq_enqueue_count_mem_re                    (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_re),
       .rf_qid_atq_enqueue_count_mem_rclk                  (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rclk),
       .rf_qid_atq_enqueue_count_mem_rclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rclk_rst_n),
       .rf_qid_atq_enqueue_count_mem_raddr                 (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_raddr),
       .rf_qid_atq_enqueue_count_mem_waddr                 (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_waddr),
       .rf_qid_atq_enqueue_count_mem_we                    (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_we),
       .rf_qid_atq_enqueue_count_mem_wclk                  (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wclk),
       .rf_qid_atq_enqueue_count_mem_wclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wclk_rst_n),
       .rf_qid_atq_enqueue_count_mem_wdata                 (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_wdata),
       .rf_qid_atq_enqueue_count_mem_rdata                 (i_hqm_list_sel_pipe_rf_qid_atq_enqueue_count_mem_rdata),
       .rf_qid_dir_max_depth_mem_re                        (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_re),
       .rf_qid_dir_max_depth_mem_rclk                      (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rclk),
       .rf_qid_dir_max_depth_mem_rclk_rst_n                (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rclk_rst_n),
       .rf_qid_dir_max_depth_mem_raddr                     (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_raddr),
       .rf_qid_dir_max_depth_mem_waddr                     (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_waddr),
       .rf_qid_dir_max_depth_mem_we                        (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_we),
       .rf_qid_dir_max_depth_mem_wclk                      (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wclk),
       .rf_qid_dir_max_depth_mem_wclk_rst_n                (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wclk_rst_n),
       .rf_qid_dir_max_depth_mem_wdata                     (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_wdata),
       .rf_qid_dir_max_depth_mem_rdata                     (i_hqm_list_sel_pipe_rf_qid_dir_max_depth_mem_rdata),
       .rf_qid_dir_replay_count_mem_re                     (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_re),
       .rf_qid_dir_replay_count_mem_rclk                   (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rclk),
       .rf_qid_dir_replay_count_mem_rclk_rst_n             (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rclk_rst_n),
       .rf_qid_dir_replay_count_mem_raddr                  (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_raddr),
       .rf_qid_dir_replay_count_mem_waddr                  (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_waddr),
       .rf_qid_dir_replay_count_mem_we                     (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_we),
       .rf_qid_dir_replay_count_mem_wclk                   (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wclk),
       .rf_qid_dir_replay_count_mem_wclk_rst_n             (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wclk_rst_n),
       .rf_qid_dir_replay_count_mem_wdata                  (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_wdata),
       .rf_qid_dir_replay_count_mem_rdata                  (i_hqm_list_sel_pipe_rf_qid_dir_replay_count_mem_rdata),
       .rf_qid_dir_tot_enq_cnt_mem_re                      (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_re),
       .rf_qid_dir_tot_enq_cnt_mem_rclk                    (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rclk),
       .rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rclk_rst_n),
       .rf_qid_dir_tot_enq_cnt_mem_raddr                   (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_raddr),
       .rf_qid_dir_tot_enq_cnt_mem_waddr                   (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_waddr),
       .rf_qid_dir_tot_enq_cnt_mem_we                      (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_we),
       .rf_qid_dir_tot_enq_cnt_mem_wclk                    (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wclk),
       .rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wclk_rst_n),
       .rf_qid_dir_tot_enq_cnt_mem_wdata                   (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_wdata),
       .rf_qid_dir_tot_enq_cnt_mem_rdata                   (i_hqm_list_sel_pipe_rf_qid_dir_tot_enq_cnt_mem_rdata),
       .rf_qid_ldb_enqueue_count_mem_re                    (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_re),
       .rf_qid_ldb_enqueue_count_mem_rclk                  (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rclk),
       .rf_qid_ldb_enqueue_count_mem_rclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rclk_rst_n),
       .rf_qid_ldb_enqueue_count_mem_raddr                 (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_raddr),
       .rf_qid_ldb_enqueue_count_mem_waddr                 (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_waddr),
       .rf_qid_ldb_enqueue_count_mem_we                    (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_we),
       .rf_qid_ldb_enqueue_count_mem_wclk                  (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wclk),
       .rf_qid_ldb_enqueue_count_mem_wclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wclk_rst_n),
       .rf_qid_ldb_enqueue_count_mem_wdata                 (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_wdata),
       .rf_qid_ldb_enqueue_count_mem_rdata                 (i_hqm_list_sel_pipe_rf_qid_ldb_enqueue_count_mem_rdata),
       .rf_qid_ldb_inflight_count_mem_re                   (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_re),
       .rf_qid_ldb_inflight_count_mem_rclk                 (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rclk),
       .rf_qid_ldb_inflight_count_mem_rclk_rst_n           (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rclk_rst_n),
       .rf_qid_ldb_inflight_count_mem_raddr                (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_raddr),
       .rf_qid_ldb_inflight_count_mem_waddr                (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_waddr),
       .rf_qid_ldb_inflight_count_mem_we                   (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_we),
       .rf_qid_ldb_inflight_count_mem_wclk                 (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wclk),
       .rf_qid_ldb_inflight_count_mem_wclk_rst_n           (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wclk_rst_n),
       .rf_qid_ldb_inflight_count_mem_wdata                (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_wdata),
       .rf_qid_ldb_inflight_count_mem_rdata                (i_hqm_list_sel_pipe_rf_qid_ldb_inflight_count_mem_rdata),
       .rf_qid_ldb_replay_count_mem_re                     (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_re),
       .rf_qid_ldb_replay_count_mem_rclk                   (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rclk),
       .rf_qid_ldb_replay_count_mem_rclk_rst_n             (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rclk_rst_n),
       .rf_qid_ldb_replay_count_mem_raddr                  (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_raddr),
       .rf_qid_ldb_replay_count_mem_waddr                  (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_waddr),
       .rf_qid_ldb_replay_count_mem_we                     (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_we),
       .rf_qid_ldb_replay_count_mem_wclk                   (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wclk),
       .rf_qid_ldb_replay_count_mem_wclk_rst_n             (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wclk_rst_n),
       .rf_qid_ldb_replay_count_mem_wdata                  (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_wdata),
       .rf_qid_ldb_replay_count_mem_rdata                  (i_hqm_list_sel_pipe_rf_qid_ldb_replay_count_mem_rdata),
       .rf_qid_naldb_max_depth_mem_re                      (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_re),
       .rf_qid_naldb_max_depth_mem_rclk                    (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rclk),
       .rf_qid_naldb_max_depth_mem_rclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rclk_rst_n),
       .rf_qid_naldb_max_depth_mem_raddr                   (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_raddr),
       .rf_qid_naldb_max_depth_mem_waddr                   (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_waddr),
       .rf_qid_naldb_max_depth_mem_we                      (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_we),
       .rf_qid_naldb_max_depth_mem_wclk                    (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wclk),
       .rf_qid_naldb_max_depth_mem_wclk_rst_n              (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wclk_rst_n),
       .rf_qid_naldb_max_depth_mem_wdata                   (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_wdata),
       .rf_qid_naldb_max_depth_mem_rdata                   (i_hqm_list_sel_pipe_rf_qid_naldb_max_depth_mem_rdata),
       .rf_qid_naldb_tot_enq_cnt_mem_re                    (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_re),
       .rf_qid_naldb_tot_enq_cnt_mem_rclk                  (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rclk),
       .rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rclk_rst_n),
       .rf_qid_naldb_tot_enq_cnt_mem_raddr                 (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_raddr),
       .rf_qid_naldb_tot_enq_cnt_mem_waddr                 (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_waddr),
       .rf_qid_naldb_tot_enq_cnt_mem_we                    (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_we),
       .rf_qid_naldb_tot_enq_cnt_mem_wclk                  (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wclk),
       .rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n            (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wclk_rst_n),
       .rf_qid_naldb_tot_enq_cnt_mem_wdata                 (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_wdata),
       .rf_qid_naldb_tot_enq_cnt_mem_rdata                 (i_hqm_list_sel_pipe_rf_qid_naldb_tot_enq_cnt_mem_rdata),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re          (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_re),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk        (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n  (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rclk_rst_n),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr       (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_raddr),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr       (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_waddr),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we          (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_we),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk        (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n  (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wclk_rst_n),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata       (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_wdata),
       .rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata       (i_hqm_list_sel_pipe_rf_rop_lsp_reordercmp_rx_sync_fifo_mem_rdata),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_re              (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_re),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_rclk            (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rclk),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n      (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rclk_rst_n),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_raddr           (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_raddr),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_waddr           (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_waddr),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_we              (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_we),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_wclk            (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wclk),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n      (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wclk_rst_n),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_wdata           (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_wdata),
       .rf_send_atm_to_cq_rx_sync_fifo_mem_rdata           (i_hqm_list_sel_pipe_rf_send_atm_to_cq_rx_sync_fifo_mem_rdata),
       .rf_uno_atm_cmp_fifo_mem_re                         (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_re),
       .rf_uno_atm_cmp_fifo_mem_rclk                       (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rclk),
       .rf_uno_atm_cmp_fifo_mem_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rclk_rst_n),
       .rf_uno_atm_cmp_fifo_mem_raddr                      (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_raddr),
       .rf_uno_atm_cmp_fifo_mem_waddr                      (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_waddr),
       .rf_uno_atm_cmp_fifo_mem_we                         (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_we),
       .rf_uno_atm_cmp_fifo_mem_wclk                       (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wclk),
       .rf_uno_atm_cmp_fifo_mem_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wclk_rst_n),
       .rf_uno_atm_cmp_fifo_mem_wdata                      (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_wdata),
       .rf_uno_atm_cmp_fifo_mem_rdata                      (i_hqm_list_sel_pipe_rf_uno_atm_cmp_fifo_mem_rdata),
       .rf_aqed_qid2cqidix_re                              (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_re),
       .rf_aqed_qid2cqidix_rclk                            (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rclk),
       .rf_aqed_qid2cqidix_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rclk_rst_n),
       .rf_aqed_qid2cqidix_raddr                           (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_raddr),
       .rf_aqed_qid2cqidix_waddr                           (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_waddr),
       .rf_aqed_qid2cqidix_we                              (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_we),
       .rf_aqed_qid2cqidix_wclk                            (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wclk),
       .rf_aqed_qid2cqidix_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wclk_rst_n),
       .rf_aqed_qid2cqidix_wdata                           (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_wdata),
       .rf_aqed_qid2cqidix_rdata                           (i_hqm_list_sel_pipe_rf_aqed_qid2cqidix_rdata),
       .rf_atm_fifo_ap_aqed_re                             (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_re),
       .rf_atm_fifo_ap_aqed_rclk                           (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rclk),
       .rf_atm_fifo_ap_aqed_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rclk_rst_n),
       .rf_atm_fifo_ap_aqed_raddr                          (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_raddr),
       .rf_atm_fifo_ap_aqed_waddr                          (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_waddr),
       .rf_atm_fifo_ap_aqed_we                             (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_we),
       .rf_atm_fifo_ap_aqed_wclk                           (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wclk),
       .rf_atm_fifo_ap_aqed_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wclk_rst_n),
       .rf_atm_fifo_ap_aqed_wdata                          (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_wdata),
       .rf_atm_fifo_ap_aqed_rdata                          (i_hqm_list_sel_pipe_rf_atm_fifo_ap_aqed_rdata),
       .rf_atm_fifo_aqed_ap_enq_re                         (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_re),
       .rf_atm_fifo_aqed_ap_enq_rclk                       (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rclk),
       .rf_atm_fifo_aqed_ap_enq_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rclk_rst_n),
       .rf_atm_fifo_aqed_ap_enq_raddr                      (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_raddr),
       .rf_atm_fifo_aqed_ap_enq_waddr                      (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_waddr),
       .rf_atm_fifo_aqed_ap_enq_we                         (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_we),
       .rf_atm_fifo_aqed_ap_enq_wclk                       (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wclk),
       .rf_atm_fifo_aqed_ap_enq_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wclk_rst_n),
       .rf_atm_fifo_aqed_ap_enq_wdata                      (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_wdata),
       .rf_atm_fifo_aqed_ap_enq_rdata                      (i_hqm_list_sel_pipe_rf_atm_fifo_aqed_ap_enq_rdata),
       .rf_fid2cqqidix_re                                  (i_hqm_list_sel_pipe_rf_fid2cqqidix_re),
       .rf_fid2cqqidix_rclk                                (i_hqm_list_sel_pipe_rf_fid2cqqidix_rclk),
       .rf_fid2cqqidix_rclk_rst_n                          (i_hqm_list_sel_pipe_rf_fid2cqqidix_rclk_rst_n),
       .rf_fid2cqqidix_raddr                               (i_hqm_list_sel_pipe_rf_fid2cqqidix_raddr),
       .rf_fid2cqqidix_waddr                               (i_hqm_list_sel_pipe_rf_fid2cqqidix_waddr),
       .rf_fid2cqqidix_we                                  (i_hqm_list_sel_pipe_rf_fid2cqqidix_we),
       .rf_fid2cqqidix_wclk                                (i_hqm_list_sel_pipe_rf_fid2cqqidix_wclk),
       .rf_fid2cqqidix_wclk_rst_n                          (i_hqm_list_sel_pipe_rf_fid2cqqidix_wclk_rst_n),
       .rf_fid2cqqidix_wdata                               (i_hqm_list_sel_pipe_rf_fid2cqqidix_wdata),
       .rf_fid2cqqidix_rdata                               (i_hqm_list_sel_pipe_rf_fid2cqqidix_rdata),
       .rf_ll_enq_cnt_r_bin0_dup0_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_re),
       .rf_ll_enq_cnt_r_bin0_dup0_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rclk),
       .rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup0_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_raddr),
       .rf_ll_enq_cnt_r_bin0_dup0_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_waddr),
       .rf_ll_enq_cnt_r_bin0_dup0_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_we),
       .rf_ll_enq_cnt_r_bin0_dup0_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wclk),
       .rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup0_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_wdata),
       .rf_ll_enq_cnt_r_bin0_dup0_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup0_rdata),
       .rf_ll_enq_cnt_r_bin0_dup1_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_re),
       .rf_ll_enq_cnt_r_bin0_dup1_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rclk),
       .rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup1_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_raddr),
       .rf_ll_enq_cnt_r_bin0_dup1_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_waddr),
       .rf_ll_enq_cnt_r_bin0_dup1_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_we),
       .rf_ll_enq_cnt_r_bin0_dup1_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wclk),
       .rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup1_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_wdata),
       .rf_ll_enq_cnt_r_bin0_dup1_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup1_rdata),
       .rf_ll_enq_cnt_r_bin0_dup2_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_re),
       .rf_ll_enq_cnt_r_bin0_dup2_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rclk),
       .rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup2_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_raddr),
       .rf_ll_enq_cnt_r_bin0_dup2_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_waddr),
       .rf_ll_enq_cnt_r_bin0_dup2_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_we),
       .rf_ll_enq_cnt_r_bin0_dup2_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wclk),
       .rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup2_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_wdata),
       .rf_ll_enq_cnt_r_bin0_dup2_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup2_rdata),
       .rf_ll_enq_cnt_r_bin0_dup3_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_re),
       .rf_ll_enq_cnt_r_bin0_dup3_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rclk),
       .rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup3_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_raddr),
       .rf_ll_enq_cnt_r_bin0_dup3_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_waddr),
       .rf_ll_enq_cnt_r_bin0_dup3_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_we),
       .rf_ll_enq_cnt_r_bin0_dup3_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wclk),
       .rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin0_dup3_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_wdata),
       .rf_ll_enq_cnt_r_bin0_dup3_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin0_dup3_rdata),
       .rf_ll_enq_cnt_r_bin1_dup0_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_re),
       .rf_ll_enq_cnt_r_bin1_dup0_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rclk),
       .rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup0_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_raddr),
       .rf_ll_enq_cnt_r_bin1_dup0_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_waddr),
       .rf_ll_enq_cnt_r_bin1_dup0_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_we),
       .rf_ll_enq_cnt_r_bin1_dup0_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wclk),
       .rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup0_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_wdata),
       .rf_ll_enq_cnt_r_bin1_dup0_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup0_rdata),
       .rf_ll_enq_cnt_r_bin1_dup1_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_re),
       .rf_ll_enq_cnt_r_bin1_dup1_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rclk),
       .rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup1_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_raddr),
       .rf_ll_enq_cnt_r_bin1_dup1_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_waddr),
       .rf_ll_enq_cnt_r_bin1_dup1_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_we),
       .rf_ll_enq_cnt_r_bin1_dup1_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wclk),
       .rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup1_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_wdata),
       .rf_ll_enq_cnt_r_bin1_dup1_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup1_rdata),
       .rf_ll_enq_cnt_r_bin1_dup2_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_re),
       .rf_ll_enq_cnt_r_bin1_dup2_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rclk),
       .rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup2_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_raddr),
       .rf_ll_enq_cnt_r_bin1_dup2_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_waddr),
       .rf_ll_enq_cnt_r_bin1_dup2_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_we),
       .rf_ll_enq_cnt_r_bin1_dup2_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wclk),
       .rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup2_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_wdata),
       .rf_ll_enq_cnt_r_bin1_dup2_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup2_rdata),
       .rf_ll_enq_cnt_r_bin1_dup3_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_re),
       .rf_ll_enq_cnt_r_bin1_dup3_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rclk),
       .rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup3_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_raddr),
       .rf_ll_enq_cnt_r_bin1_dup3_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_waddr),
       .rf_ll_enq_cnt_r_bin1_dup3_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_we),
       .rf_ll_enq_cnt_r_bin1_dup3_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wclk),
       .rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin1_dup3_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_wdata),
       .rf_ll_enq_cnt_r_bin1_dup3_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin1_dup3_rdata),
       .rf_ll_enq_cnt_r_bin2_dup0_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_re),
       .rf_ll_enq_cnt_r_bin2_dup0_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rclk),
       .rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup0_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_raddr),
       .rf_ll_enq_cnt_r_bin2_dup0_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_waddr),
       .rf_ll_enq_cnt_r_bin2_dup0_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_we),
       .rf_ll_enq_cnt_r_bin2_dup0_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wclk),
       .rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup0_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_wdata),
       .rf_ll_enq_cnt_r_bin2_dup0_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup0_rdata),
       .rf_ll_enq_cnt_r_bin2_dup1_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_re),
       .rf_ll_enq_cnt_r_bin2_dup1_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rclk),
       .rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup1_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_raddr),
       .rf_ll_enq_cnt_r_bin2_dup1_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_waddr),
       .rf_ll_enq_cnt_r_bin2_dup1_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_we),
       .rf_ll_enq_cnt_r_bin2_dup1_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wclk),
       .rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup1_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_wdata),
       .rf_ll_enq_cnt_r_bin2_dup1_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup1_rdata),
       .rf_ll_enq_cnt_r_bin2_dup2_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_re),
       .rf_ll_enq_cnt_r_bin2_dup2_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rclk),
       .rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup2_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_raddr),
       .rf_ll_enq_cnt_r_bin2_dup2_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_waddr),
       .rf_ll_enq_cnt_r_bin2_dup2_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_we),
       .rf_ll_enq_cnt_r_bin2_dup2_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wclk),
       .rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup2_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_wdata),
       .rf_ll_enq_cnt_r_bin2_dup2_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup2_rdata),
       .rf_ll_enq_cnt_r_bin2_dup3_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_re),
       .rf_ll_enq_cnt_r_bin2_dup3_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rclk),
       .rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup3_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_raddr),
       .rf_ll_enq_cnt_r_bin2_dup3_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_waddr),
       .rf_ll_enq_cnt_r_bin2_dup3_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_we),
       .rf_ll_enq_cnt_r_bin2_dup3_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wclk),
       .rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin2_dup3_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_wdata),
       .rf_ll_enq_cnt_r_bin2_dup3_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin2_dup3_rdata),
       .rf_ll_enq_cnt_r_bin3_dup0_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_re),
       .rf_ll_enq_cnt_r_bin3_dup0_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rclk),
       .rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup0_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_raddr),
       .rf_ll_enq_cnt_r_bin3_dup0_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_waddr),
       .rf_ll_enq_cnt_r_bin3_dup0_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_we),
       .rf_ll_enq_cnt_r_bin3_dup0_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wclk),
       .rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup0_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_wdata),
       .rf_ll_enq_cnt_r_bin3_dup0_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup0_rdata),
       .rf_ll_enq_cnt_r_bin3_dup1_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_re),
       .rf_ll_enq_cnt_r_bin3_dup1_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rclk),
       .rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup1_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_raddr),
       .rf_ll_enq_cnt_r_bin3_dup1_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_waddr),
       .rf_ll_enq_cnt_r_bin3_dup1_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_we),
       .rf_ll_enq_cnt_r_bin3_dup1_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wclk),
       .rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup1_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_wdata),
       .rf_ll_enq_cnt_r_bin3_dup1_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup1_rdata),
       .rf_ll_enq_cnt_r_bin3_dup2_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_re),
       .rf_ll_enq_cnt_r_bin3_dup2_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rclk),
       .rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup2_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_raddr),
       .rf_ll_enq_cnt_r_bin3_dup2_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_waddr),
       .rf_ll_enq_cnt_r_bin3_dup2_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_we),
       .rf_ll_enq_cnt_r_bin3_dup2_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wclk),
       .rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup2_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_wdata),
       .rf_ll_enq_cnt_r_bin3_dup2_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup2_rdata),
       .rf_ll_enq_cnt_r_bin3_dup3_re                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_re),
       .rf_ll_enq_cnt_r_bin3_dup3_rclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rclk),
       .rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup3_raddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_raddr),
       .rf_ll_enq_cnt_r_bin3_dup3_waddr                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_waddr),
       .rf_ll_enq_cnt_r_bin3_dup3_we                       (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_we),
       .rf_ll_enq_cnt_r_bin3_dup3_wclk                     (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wclk),
       .rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n               (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wclk_rst_n),
       .rf_ll_enq_cnt_r_bin3_dup3_wdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_wdata),
       .rf_ll_enq_cnt_r_bin3_dup3_rdata                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_r_bin3_dup3_rdata),
       .rf_ll_enq_cnt_s_bin0_re                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_re),
       .rf_ll_enq_cnt_s_bin0_rclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rclk),
       .rf_ll_enq_cnt_s_bin0_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rclk_rst_n),
       .rf_ll_enq_cnt_s_bin0_raddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_raddr),
       .rf_ll_enq_cnt_s_bin0_waddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_waddr),
       .rf_ll_enq_cnt_s_bin0_we                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_we),
       .rf_ll_enq_cnt_s_bin0_wclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wclk),
       .rf_ll_enq_cnt_s_bin0_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wclk_rst_n),
       .rf_ll_enq_cnt_s_bin0_wdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_wdata),
       .rf_ll_enq_cnt_s_bin0_rdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin0_rdata),
       .rf_ll_enq_cnt_s_bin1_re                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_re),
       .rf_ll_enq_cnt_s_bin1_rclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rclk),
       .rf_ll_enq_cnt_s_bin1_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rclk_rst_n),
       .rf_ll_enq_cnt_s_bin1_raddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_raddr),
       .rf_ll_enq_cnt_s_bin1_waddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_waddr),
       .rf_ll_enq_cnt_s_bin1_we                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_we),
       .rf_ll_enq_cnt_s_bin1_wclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wclk),
       .rf_ll_enq_cnt_s_bin1_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wclk_rst_n),
       .rf_ll_enq_cnt_s_bin1_wdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_wdata),
       .rf_ll_enq_cnt_s_bin1_rdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin1_rdata),
       .rf_ll_enq_cnt_s_bin2_re                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_re),
       .rf_ll_enq_cnt_s_bin2_rclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rclk),
       .rf_ll_enq_cnt_s_bin2_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rclk_rst_n),
       .rf_ll_enq_cnt_s_bin2_raddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_raddr),
       .rf_ll_enq_cnt_s_bin2_waddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_waddr),
       .rf_ll_enq_cnt_s_bin2_we                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_we),
       .rf_ll_enq_cnt_s_bin2_wclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wclk),
       .rf_ll_enq_cnt_s_bin2_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wclk_rst_n),
       .rf_ll_enq_cnt_s_bin2_wdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_wdata),
       .rf_ll_enq_cnt_s_bin2_rdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin2_rdata),
       .rf_ll_enq_cnt_s_bin3_re                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_re),
       .rf_ll_enq_cnt_s_bin3_rclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rclk),
       .rf_ll_enq_cnt_s_bin3_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rclk_rst_n),
       .rf_ll_enq_cnt_s_bin3_raddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_raddr),
       .rf_ll_enq_cnt_s_bin3_waddr                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_waddr),
       .rf_ll_enq_cnt_s_bin3_we                            (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_we),
       .rf_ll_enq_cnt_s_bin3_wclk                          (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wclk),
       .rf_ll_enq_cnt_s_bin3_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wclk_rst_n),
       .rf_ll_enq_cnt_s_bin3_wdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_wdata),
       .rf_ll_enq_cnt_s_bin3_rdata                         (i_hqm_list_sel_pipe_rf_ll_enq_cnt_s_bin3_rdata),
       .rf_ll_rdylst_hp_bin0_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_re),
       .rf_ll_rdylst_hp_bin0_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rclk),
       .rf_ll_rdylst_hp_bin0_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rclk_rst_n),
       .rf_ll_rdylst_hp_bin0_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_raddr),
       .rf_ll_rdylst_hp_bin0_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_waddr),
       .rf_ll_rdylst_hp_bin0_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_we),
       .rf_ll_rdylst_hp_bin0_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wclk),
       .rf_ll_rdylst_hp_bin0_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wclk_rst_n),
       .rf_ll_rdylst_hp_bin0_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_wdata),
       .rf_ll_rdylst_hp_bin0_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin0_rdata),
       .rf_ll_rdylst_hp_bin1_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_re),
       .rf_ll_rdylst_hp_bin1_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rclk),
       .rf_ll_rdylst_hp_bin1_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rclk_rst_n),
       .rf_ll_rdylst_hp_bin1_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_raddr),
       .rf_ll_rdylst_hp_bin1_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_waddr),
       .rf_ll_rdylst_hp_bin1_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_we),
       .rf_ll_rdylst_hp_bin1_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wclk),
       .rf_ll_rdylst_hp_bin1_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wclk_rst_n),
       .rf_ll_rdylst_hp_bin1_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_wdata),
       .rf_ll_rdylst_hp_bin1_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin1_rdata),
       .rf_ll_rdylst_hp_bin2_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_re),
       .rf_ll_rdylst_hp_bin2_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rclk),
       .rf_ll_rdylst_hp_bin2_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rclk_rst_n),
       .rf_ll_rdylst_hp_bin2_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_raddr),
       .rf_ll_rdylst_hp_bin2_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_waddr),
       .rf_ll_rdylst_hp_bin2_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_we),
       .rf_ll_rdylst_hp_bin2_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wclk),
       .rf_ll_rdylst_hp_bin2_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wclk_rst_n),
       .rf_ll_rdylst_hp_bin2_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_wdata),
       .rf_ll_rdylst_hp_bin2_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin2_rdata),
       .rf_ll_rdylst_hp_bin3_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_re),
       .rf_ll_rdylst_hp_bin3_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rclk),
       .rf_ll_rdylst_hp_bin3_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rclk_rst_n),
       .rf_ll_rdylst_hp_bin3_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_raddr),
       .rf_ll_rdylst_hp_bin3_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_waddr),
       .rf_ll_rdylst_hp_bin3_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_we),
       .rf_ll_rdylst_hp_bin3_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wclk),
       .rf_ll_rdylst_hp_bin3_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wclk_rst_n),
       .rf_ll_rdylst_hp_bin3_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_wdata),
       .rf_ll_rdylst_hp_bin3_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hp_bin3_rdata),
       .rf_ll_rdylst_hpnxt_bin0_re                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_re),
       .rf_ll_rdylst_hpnxt_bin0_rclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rclk),
       .rf_ll_rdylst_hpnxt_bin0_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin0_raddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_raddr),
       .rf_ll_rdylst_hpnxt_bin0_waddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_waddr),
       .rf_ll_rdylst_hpnxt_bin0_we                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_we),
       .rf_ll_rdylst_hpnxt_bin0_wclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wclk),
       .rf_ll_rdylst_hpnxt_bin0_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin0_wdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_wdata),
       .rf_ll_rdylst_hpnxt_bin0_rdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin0_rdata),
       .rf_ll_rdylst_hpnxt_bin1_re                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_re),
       .rf_ll_rdylst_hpnxt_bin1_rclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rclk),
       .rf_ll_rdylst_hpnxt_bin1_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin1_raddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_raddr),
       .rf_ll_rdylst_hpnxt_bin1_waddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_waddr),
       .rf_ll_rdylst_hpnxt_bin1_we                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_we),
       .rf_ll_rdylst_hpnxt_bin1_wclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wclk),
       .rf_ll_rdylst_hpnxt_bin1_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin1_wdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_wdata),
       .rf_ll_rdylst_hpnxt_bin1_rdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin1_rdata),
       .rf_ll_rdylst_hpnxt_bin2_re                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_re),
       .rf_ll_rdylst_hpnxt_bin2_rclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rclk),
       .rf_ll_rdylst_hpnxt_bin2_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin2_raddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_raddr),
       .rf_ll_rdylst_hpnxt_bin2_waddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_waddr),
       .rf_ll_rdylst_hpnxt_bin2_we                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_we),
       .rf_ll_rdylst_hpnxt_bin2_wclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wclk),
       .rf_ll_rdylst_hpnxt_bin2_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin2_wdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_wdata),
       .rf_ll_rdylst_hpnxt_bin2_rdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin2_rdata),
       .rf_ll_rdylst_hpnxt_bin3_re                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_re),
       .rf_ll_rdylst_hpnxt_bin3_rclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rclk),
       .rf_ll_rdylst_hpnxt_bin3_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin3_raddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_raddr),
       .rf_ll_rdylst_hpnxt_bin3_waddr                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_waddr),
       .rf_ll_rdylst_hpnxt_bin3_we                         (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_we),
       .rf_ll_rdylst_hpnxt_bin3_wclk                       (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wclk),
       .rf_ll_rdylst_hpnxt_bin3_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wclk_rst_n),
       .rf_ll_rdylst_hpnxt_bin3_wdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_wdata),
       .rf_ll_rdylst_hpnxt_bin3_rdata                      (i_hqm_list_sel_pipe_rf_ll_rdylst_hpnxt_bin3_rdata),
       .rf_ll_rdylst_tp_bin0_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_re),
       .rf_ll_rdylst_tp_bin0_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rclk),
       .rf_ll_rdylst_tp_bin0_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rclk_rst_n),
       .rf_ll_rdylst_tp_bin0_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_raddr),
       .rf_ll_rdylst_tp_bin0_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_waddr),
       .rf_ll_rdylst_tp_bin0_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_we),
       .rf_ll_rdylst_tp_bin0_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wclk),
       .rf_ll_rdylst_tp_bin0_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wclk_rst_n),
       .rf_ll_rdylst_tp_bin0_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_wdata),
       .rf_ll_rdylst_tp_bin0_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin0_rdata),
       .rf_ll_rdylst_tp_bin1_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_re),
       .rf_ll_rdylst_tp_bin1_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rclk),
       .rf_ll_rdylst_tp_bin1_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rclk_rst_n),
       .rf_ll_rdylst_tp_bin1_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_raddr),
       .rf_ll_rdylst_tp_bin1_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_waddr),
       .rf_ll_rdylst_tp_bin1_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_we),
       .rf_ll_rdylst_tp_bin1_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wclk),
       .rf_ll_rdylst_tp_bin1_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wclk_rst_n),
       .rf_ll_rdylst_tp_bin1_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_wdata),
       .rf_ll_rdylst_tp_bin1_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin1_rdata),
       .rf_ll_rdylst_tp_bin2_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_re),
       .rf_ll_rdylst_tp_bin2_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rclk),
       .rf_ll_rdylst_tp_bin2_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rclk_rst_n),
       .rf_ll_rdylst_tp_bin2_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_raddr),
       .rf_ll_rdylst_tp_bin2_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_waddr),
       .rf_ll_rdylst_tp_bin2_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_we),
       .rf_ll_rdylst_tp_bin2_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wclk),
       .rf_ll_rdylst_tp_bin2_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wclk_rst_n),
       .rf_ll_rdylst_tp_bin2_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_wdata),
       .rf_ll_rdylst_tp_bin2_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin2_rdata),
       .rf_ll_rdylst_tp_bin3_re                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_re),
       .rf_ll_rdylst_tp_bin3_rclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rclk),
       .rf_ll_rdylst_tp_bin3_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rclk_rst_n),
       .rf_ll_rdylst_tp_bin3_raddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_raddr),
       .rf_ll_rdylst_tp_bin3_waddr                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_waddr),
       .rf_ll_rdylst_tp_bin3_we                            (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_we),
       .rf_ll_rdylst_tp_bin3_wclk                          (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wclk),
       .rf_ll_rdylst_tp_bin3_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wclk_rst_n),
       .rf_ll_rdylst_tp_bin3_wdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_wdata),
       .rf_ll_rdylst_tp_bin3_rdata                         (i_hqm_list_sel_pipe_rf_ll_rdylst_tp_bin3_rdata),
       .rf_ll_rlst_cnt_re                                  (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_re),
       .rf_ll_rlst_cnt_rclk                                (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rclk),
       .rf_ll_rlst_cnt_rclk_rst_n                          (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rclk_rst_n),
       .rf_ll_rlst_cnt_raddr                               (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_raddr),
       .rf_ll_rlst_cnt_waddr                               (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_waddr),
       .rf_ll_rlst_cnt_we                                  (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_we),
       .rf_ll_rlst_cnt_wclk                                (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wclk),
       .rf_ll_rlst_cnt_wclk_rst_n                          (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wclk_rst_n),
       .rf_ll_rlst_cnt_wdata                               (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_wdata),
       .rf_ll_rlst_cnt_rdata                               (i_hqm_list_sel_pipe_rf_ll_rlst_cnt_rdata),
       .rf_ll_sch_cnt_dup0_re                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_re),
       .rf_ll_sch_cnt_dup0_rclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rclk),
       .rf_ll_sch_cnt_dup0_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rclk_rst_n),
       .rf_ll_sch_cnt_dup0_raddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_raddr),
       .rf_ll_sch_cnt_dup0_waddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_waddr),
       .rf_ll_sch_cnt_dup0_we                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_we),
       .rf_ll_sch_cnt_dup0_wclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wclk),
       .rf_ll_sch_cnt_dup0_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wclk_rst_n),
       .rf_ll_sch_cnt_dup0_wdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_wdata),
       .rf_ll_sch_cnt_dup0_rdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup0_rdata),
       .rf_ll_sch_cnt_dup1_re                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_re),
       .rf_ll_sch_cnt_dup1_rclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rclk),
       .rf_ll_sch_cnt_dup1_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rclk_rst_n),
       .rf_ll_sch_cnt_dup1_raddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_raddr),
       .rf_ll_sch_cnt_dup1_waddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_waddr),
       .rf_ll_sch_cnt_dup1_we                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_we),
       .rf_ll_sch_cnt_dup1_wclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wclk),
       .rf_ll_sch_cnt_dup1_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wclk_rst_n),
       .rf_ll_sch_cnt_dup1_wdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_wdata),
       .rf_ll_sch_cnt_dup1_rdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup1_rdata),
       .rf_ll_sch_cnt_dup2_re                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_re),
       .rf_ll_sch_cnt_dup2_rclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rclk),
       .rf_ll_sch_cnt_dup2_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rclk_rst_n),
       .rf_ll_sch_cnt_dup2_raddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_raddr),
       .rf_ll_sch_cnt_dup2_waddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_waddr),
       .rf_ll_sch_cnt_dup2_we                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_we),
       .rf_ll_sch_cnt_dup2_wclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wclk),
       .rf_ll_sch_cnt_dup2_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wclk_rst_n),
       .rf_ll_sch_cnt_dup2_wdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_wdata),
       .rf_ll_sch_cnt_dup2_rdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup2_rdata),
       .rf_ll_sch_cnt_dup3_re                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_re),
       .rf_ll_sch_cnt_dup3_rclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rclk),
       .rf_ll_sch_cnt_dup3_rclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rclk_rst_n),
       .rf_ll_sch_cnt_dup3_raddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_raddr),
       .rf_ll_sch_cnt_dup3_waddr                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_waddr),
       .rf_ll_sch_cnt_dup3_we                              (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_we),
       .rf_ll_sch_cnt_dup3_wclk                            (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wclk),
       .rf_ll_sch_cnt_dup3_wclk_rst_n                      (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wclk_rst_n),
       .rf_ll_sch_cnt_dup3_wdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_wdata),
       .rf_ll_sch_cnt_dup3_rdata                           (i_hqm_list_sel_pipe_rf_ll_sch_cnt_dup3_rdata),
       .rf_ll_schlst_hp_bin0_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_re),
       .rf_ll_schlst_hp_bin0_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rclk),
       .rf_ll_schlst_hp_bin0_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rclk_rst_n),
       .rf_ll_schlst_hp_bin0_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_raddr),
       .rf_ll_schlst_hp_bin0_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_waddr),
       .rf_ll_schlst_hp_bin0_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_we),
       .rf_ll_schlst_hp_bin0_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wclk),
       .rf_ll_schlst_hp_bin0_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wclk_rst_n),
       .rf_ll_schlst_hp_bin0_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_wdata),
       .rf_ll_schlst_hp_bin0_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin0_rdata),
       .rf_ll_schlst_hp_bin1_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_re),
       .rf_ll_schlst_hp_bin1_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rclk),
       .rf_ll_schlst_hp_bin1_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rclk_rst_n),
       .rf_ll_schlst_hp_bin1_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_raddr),
       .rf_ll_schlst_hp_bin1_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_waddr),
       .rf_ll_schlst_hp_bin1_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_we),
       .rf_ll_schlst_hp_bin1_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wclk),
       .rf_ll_schlst_hp_bin1_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wclk_rst_n),
       .rf_ll_schlst_hp_bin1_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_wdata),
       .rf_ll_schlst_hp_bin1_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin1_rdata),
       .rf_ll_schlst_hp_bin2_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_re),
       .rf_ll_schlst_hp_bin2_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rclk),
       .rf_ll_schlst_hp_bin2_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rclk_rst_n),
       .rf_ll_schlst_hp_bin2_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_raddr),
       .rf_ll_schlst_hp_bin2_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_waddr),
       .rf_ll_schlst_hp_bin2_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_we),
       .rf_ll_schlst_hp_bin2_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wclk),
       .rf_ll_schlst_hp_bin2_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wclk_rst_n),
       .rf_ll_schlst_hp_bin2_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_wdata),
       .rf_ll_schlst_hp_bin2_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin2_rdata),
       .rf_ll_schlst_hp_bin3_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_re),
       .rf_ll_schlst_hp_bin3_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rclk),
       .rf_ll_schlst_hp_bin3_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rclk_rst_n),
       .rf_ll_schlst_hp_bin3_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_raddr),
       .rf_ll_schlst_hp_bin3_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_waddr),
       .rf_ll_schlst_hp_bin3_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_we),
       .rf_ll_schlst_hp_bin3_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wclk),
       .rf_ll_schlst_hp_bin3_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wclk_rst_n),
       .rf_ll_schlst_hp_bin3_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_wdata),
       .rf_ll_schlst_hp_bin3_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_hp_bin3_rdata),
       .rf_ll_schlst_hpnxt_bin0_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_re),
       .rf_ll_schlst_hpnxt_bin0_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rclk),
       .rf_ll_schlst_hpnxt_bin0_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rclk_rst_n),
       .rf_ll_schlst_hpnxt_bin0_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_raddr),
       .rf_ll_schlst_hpnxt_bin0_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_waddr),
       .rf_ll_schlst_hpnxt_bin0_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_we),
       .rf_ll_schlst_hpnxt_bin0_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wclk),
       .rf_ll_schlst_hpnxt_bin0_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wclk_rst_n),
       .rf_ll_schlst_hpnxt_bin0_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_wdata),
       .rf_ll_schlst_hpnxt_bin0_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin0_rdata),
       .rf_ll_schlst_hpnxt_bin1_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_re),
       .rf_ll_schlst_hpnxt_bin1_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rclk),
       .rf_ll_schlst_hpnxt_bin1_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rclk_rst_n),
       .rf_ll_schlst_hpnxt_bin1_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_raddr),
       .rf_ll_schlst_hpnxt_bin1_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_waddr),
       .rf_ll_schlst_hpnxt_bin1_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_we),
       .rf_ll_schlst_hpnxt_bin1_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wclk),
       .rf_ll_schlst_hpnxt_bin1_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wclk_rst_n),
       .rf_ll_schlst_hpnxt_bin1_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_wdata),
       .rf_ll_schlst_hpnxt_bin1_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin1_rdata),
       .rf_ll_schlst_hpnxt_bin2_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_re),
       .rf_ll_schlst_hpnxt_bin2_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rclk),
       .rf_ll_schlst_hpnxt_bin2_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rclk_rst_n),
       .rf_ll_schlst_hpnxt_bin2_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_raddr),
       .rf_ll_schlst_hpnxt_bin2_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_waddr),
       .rf_ll_schlst_hpnxt_bin2_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_we),
       .rf_ll_schlst_hpnxt_bin2_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wclk),
       .rf_ll_schlst_hpnxt_bin2_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wclk_rst_n),
       .rf_ll_schlst_hpnxt_bin2_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_wdata),
       .rf_ll_schlst_hpnxt_bin2_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin2_rdata),
       .rf_ll_schlst_hpnxt_bin3_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_re),
       .rf_ll_schlst_hpnxt_bin3_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rclk),
       .rf_ll_schlst_hpnxt_bin3_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rclk_rst_n),
       .rf_ll_schlst_hpnxt_bin3_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_raddr),
       .rf_ll_schlst_hpnxt_bin3_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_waddr),
       .rf_ll_schlst_hpnxt_bin3_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_we),
       .rf_ll_schlst_hpnxt_bin3_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wclk),
       .rf_ll_schlst_hpnxt_bin3_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wclk_rst_n),
       .rf_ll_schlst_hpnxt_bin3_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_wdata),
       .rf_ll_schlst_hpnxt_bin3_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_hpnxt_bin3_rdata),
       .rf_ll_schlst_tp_bin0_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_re),
       .rf_ll_schlst_tp_bin0_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rclk),
       .rf_ll_schlst_tp_bin0_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rclk_rst_n),
       .rf_ll_schlst_tp_bin0_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_raddr),
       .rf_ll_schlst_tp_bin0_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_waddr),
       .rf_ll_schlst_tp_bin0_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_we),
       .rf_ll_schlst_tp_bin0_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wclk),
       .rf_ll_schlst_tp_bin0_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wclk_rst_n),
       .rf_ll_schlst_tp_bin0_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_wdata),
       .rf_ll_schlst_tp_bin0_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin0_rdata),
       .rf_ll_schlst_tp_bin1_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_re),
       .rf_ll_schlst_tp_bin1_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rclk),
       .rf_ll_schlst_tp_bin1_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rclk_rst_n),
       .rf_ll_schlst_tp_bin1_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_raddr),
       .rf_ll_schlst_tp_bin1_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_waddr),
       .rf_ll_schlst_tp_bin1_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_we),
       .rf_ll_schlst_tp_bin1_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wclk),
       .rf_ll_schlst_tp_bin1_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wclk_rst_n),
       .rf_ll_schlst_tp_bin1_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_wdata),
       .rf_ll_schlst_tp_bin1_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin1_rdata),
       .rf_ll_schlst_tp_bin2_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_re),
       .rf_ll_schlst_tp_bin2_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rclk),
       .rf_ll_schlst_tp_bin2_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rclk_rst_n),
       .rf_ll_schlst_tp_bin2_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_raddr),
       .rf_ll_schlst_tp_bin2_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_waddr),
       .rf_ll_schlst_tp_bin2_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_we),
       .rf_ll_schlst_tp_bin2_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wclk),
       .rf_ll_schlst_tp_bin2_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wclk_rst_n),
       .rf_ll_schlst_tp_bin2_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_wdata),
       .rf_ll_schlst_tp_bin2_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin2_rdata),
       .rf_ll_schlst_tp_bin3_re                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_re),
       .rf_ll_schlst_tp_bin3_rclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rclk),
       .rf_ll_schlst_tp_bin3_rclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rclk_rst_n),
       .rf_ll_schlst_tp_bin3_raddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_raddr),
       .rf_ll_schlst_tp_bin3_waddr                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_waddr),
       .rf_ll_schlst_tp_bin3_we                            (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_we),
       .rf_ll_schlst_tp_bin3_wclk                          (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wclk),
       .rf_ll_schlst_tp_bin3_wclk_rst_n                    (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wclk_rst_n),
       .rf_ll_schlst_tp_bin3_wdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_wdata),
       .rf_ll_schlst_tp_bin3_rdata                         (i_hqm_list_sel_pipe_rf_ll_schlst_tp_bin3_rdata),
       .rf_ll_schlst_tpprv_bin0_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_re),
       .rf_ll_schlst_tpprv_bin0_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rclk),
       .rf_ll_schlst_tpprv_bin0_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rclk_rst_n),
       .rf_ll_schlst_tpprv_bin0_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_raddr),
       .rf_ll_schlst_tpprv_bin0_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_waddr),
       .rf_ll_schlst_tpprv_bin0_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_we),
       .rf_ll_schlst_tpprv_bin0_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wclk),
       .rf_ll_schlst_tpprv_bin0_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wclk_rst_n),
       .rf_ll_schlst_tpprv_bin0_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_wdata),
       .rf_ll_schlst_tpprv_bin0_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin0_rdata),
       .rf_ll_schlst_tpprv_bin1_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_re),
       .rf_ll_schlst_tpprv_bin1_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rclk),
       .rf_ll_schlst_tpprv_bin1_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rclk_rst_n),
       .rf_ll_schlst_tpprv_bin1_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_raddr),
       .rf_ll_schlst_tpprv_bin1_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_waddr),
       .rf_ll_schlst_tpprv_bin1_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_we),
       .rf_ll_schlst_tpprv_bin1_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wclk),
       .rf_ll_schlst_tpprv_bin1_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wclk_rst_n),
       .rf_ll_schlst_tpprv_bin1_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_wdata),
       .rf_ll_schlst_tpprv_bin1_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin1_rdata),
       .rf_ll_schlst_tpprv_bin2_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_re),
       .rf_ll_schlst_tpprv_bin2_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rclk),
       .rf_ll_schlst_tpprv_bin2_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rclk_rst_n),
       .rf_ll_schlst_tpprv_bin2_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_raddr),
       .rf_ll_schlst_tpprv_bin2_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_waddr),
       .rf_ll_schlst_tpprv_bin2_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_we),
       .rf_ll_schlst_tpprv_bin2_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wclk),
       .rf_ll_schlst_tpprv_bin2_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wclk_rst_n),
       .rf_ll_schlst_tpprv_bin2_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_wdata),
       .rf_ll_schlst_tpprv_bin2_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin2_rdata),
       .rf_ll_schlst_tpprv_bin3_re                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_re),
       .rf_ll_schlst_tpprv_bin3_rclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rclk),
       .rf_ll_schlst_tpprv_bin3_rclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rclk_rst_n),
       .rf_ll_schlst_tpprv_bin3_raddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_raddr),
       .rf_ll_schlst_tpprv_bin3_waddr                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_waddr),
       .rf_ll_schlst_tpprv_bin3_we                         (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_we),
       .rf_ll_schlst_tpprv_bin3_wclk                       (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wclk),
       .rf_ll_schlst_tpprv_bin3_wclk_rst_n                 (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wclk_rst_n),
       .rf_ll_schlst_tpprv_bin3_wdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_wdata),
       .rf_ll_schlst_tpprv_bin3_rdata                      (i_hqm_list_sel_pipe_rf_ll_schlst_tpprv_bin3_rdata),
       .rf_ll_slst_cnt_re                                  (i_hqm_list_sel_pipe_rf_ll_slst_cnt_re),
       .rf_ll_slst_cnt_rclk                                (i_hqm_list_sel_pipe_rf_ll_slst_cnt_rclk),
       .rf_ll_slst_cnt_rclk_rst_n                          (i_hqm_list_sel_pipe_rf_ll_slst_cnt_rclk_rst_n),
       .rf_ll_slst_cnt_raddr                               (i_hqm_list_sel_pipe_rf_ll_slst_cnt_raddr),
       .rf_ll_slst_cnt_waddr                               (i_hqm_list_sel_pipe_rf_ll_slst_cnt_waddr),
       .rf_ll_slst_cnt_we                                  (i_hqm_list_sel_pipe_rf_ll_slst_cnt_we),
       .rf_ll_slst_cnt_wclk                                (i_hqm_list_sel_pipe_rf_ll_slst_cnt_wclk),
       .rf_ll_slst_cnt_wclk_rst_n                          (i_hqm_list_sel_pipe_rf_ll_slst_cnt_wclk_rst_n),
       .rf_ll_slst_cnt_wdata                               (i_hqm_list_sel_pipe_rf_ll_slst_cnt_wdata),
       .rf_ll_slst_cnt_rdata                               (i_hqm_list_sel_pipe_rf_ll_slst_cnt_rdata),
       .rf_qid_rdylst_clamp_re                             (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_re),
       .rf_qid_rdylst_clamp_rclk                           (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rclk),
       .rf_qid_rdylst_clamp_rclk_rst_n                     (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rclk_rst_n),
       .rf_qid_rdylst_clamp_raddr                          (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_raddr),
       .rf_qid_rdylst_clamp_waddr                          (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_waddr),
       .rf_qid_rdylst_clamp_we                             (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_we),
       .rf_qid_rdylst_clamp_wclk                           (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wclk),
       .rf_qid_rdylst_clamp_wclk_rst_n                     (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wclk_rst_n),
       .rf_qid_rdylst_clamp_wdata                          (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_wdata),
       .rf_qid_rdylst_clamp_rdata                          (i_hqm_list_sel_pipe_rf_qid_rdylst_clamp_rdata));

   hqm_AW_flop i_hqm_lsp_clk_ungate_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_clk_ungate),
       .data_q (hqm_clk_ungate_rptr));

   hqm_AW_clkgate i_hqm_lsp_clkgate
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_inp_gated_clk_enable_rptr),
       .cfg_clkungate   (hqm_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (hqm_inp_gated_clk));

   hqm_AW_clkgate i_hqm_lsp_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_lsp),
       .cfg_clkungate   (hqm_clk_ungate_rptr),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_lsp));

   hqm_AW_flop_set i_hqm_lsp_flr_prep_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_flr_prep),
       .data_q (hqm_flr_prep_rptr));

   hqm_AW_reset_sync_scan i_hqm_lsp_hqm_clk_rptr_rst_sync_n
      (.clk            (hqm_clk_trunk),
       .rst_n          (hqm_clk_rptr_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (hqm_clk_rptr_rst_sync_b));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_lsp_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_lsp),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_lsp));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_lsp_hqm_gated_clk_enable_or2
      (.clki0 (i_hqm_list_sel_pipe_hqm_proc_clk_en_lsp),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_lsp));

   hqm_AW_flop i_hqm_lsp_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_gated_clk_enable_and_lsp),
       .data_q (hqm_gated_clk_enable_rptr_lsp));

   hqm_AW_flop i_hqm_lsp_hqm_inp_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_b),
       .data   (hqm_clk_enable),
       .data_q (hqm_inp_gated_clk_enable_rptr));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_lsp_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk,
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_lsp),
       .hqm_gated_clk          (hqm_gated_clk_lsp),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_lsp),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_lsp),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_lsp),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_lsp),
       .hqm_flr_prep           (hqm_flr_prep_rptr),
       .rst_prep               (hqm_rst_prep_lsp));

   hqm_AW_clkgate i_hqm_nalb_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_nalb),
       .cfg_clkungate   (hqm_clk_ungate_rptrx),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_nalb));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_nalb_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_nalb),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_nalb));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_nalb_hqm_gated_clk_enable_or2
      (.clki0 (i_hqm_qed_pipe_hqm_proc_clk_en_nalb),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_nalb));

   hqm_AW_flop i_hqm_nalb_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_gated_clk_enable_and_nalb),
       .data_q (hqm_gated_clk_enable_rptr_nalb));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_nalb_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_nalb),
       .hqm_gated_clk          (hqm_gated_clk_nalb),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_nalb),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_nalb),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_nalb),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_nalb),
       .hqm_flr_prep           (hqm_flr_prep_rptrx),
       .rst_prep               (hqm_rst_prep_nalb));

   hqm_AW_flop i_hqm_qed_clk_en_proc_ft_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_proc_clk_en_qed_local),
       .data_q (hqm_proc_clk_en_qed));

   hqm_AW_flop i_hqm_qed_clk_ungate_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_clk_ungate),
       .data_q (hqm_clk_ungate_rptrx));

   hqm_AW_clkgate i_hqm_qed_clkgate
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_inp_gated_clk_enable_rptrx),
       .cfg_clkungate   (hqm_clk_ungate_rptrx),
       .fscan_clkungate,
       .gated_clk       (hqm_inp_gated_clkx));

   hqm_AW_clkgate i_hqm_qed_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_qed),
       .cfg_clkungate   (hqm_clk_ungate_rptrx),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_qed));

   hqm_AW_inv i_hqm_qed_flr_prep_inv
      (.a (hqm_flr_prep_rptrx),
       .o (hqm_flr_prep_b));

   hqm_AW_flop_set i_hqm_qed_flr_prep_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_flr_prep),
       .data_q (hqm_flr_prep_rptrx));

   hqm_AW_reset_sync_scan i_hqm_qed_hqm_clk_rptr_rst_sync_n
      (.clk            (hqm_clk_trunk),
       .rst_n          (hqm_clk_rptr_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (hqm_clk_rptr_rst_sync_bx));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_qed_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_qed),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_qed));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_qed_hqm_gated_clk_enable_or2
      (.clki0 (hqm_proc_clk_en_qed_local),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_qed));

   hqm_AW_flop i_hqm_qed_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_gated_clk_enable_and_qed),
       .data_q (hqm_gated_clk_enable_rptr_qed));

   hqm_AW_flop i_hqm_qed_hqm_inp_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (hqm_clk_enable),
       .data_q (hqm_inp_gated_clk_enable_rptrx));

   hqm_qed_pipe i_hqm_qed_pipe
      (.hqm_gated_clk_qed,
       .hqm_proc_clk_en_qed                       (hqm_proc_clk_en_qed_local),
       .hqm_rst_prep_qed,
       .hqm_gated_rst_b_qed,
       .hqm_inp_gated_rst_b_qed,
       .hqm_gated_clk_nalb,
       .hqm_proc_clk_en_nalb                      (i_hqm_qed_pipe_hqm_proc_clk_en_nalb),
       .hqm_rst_prep_nalb,
       .hqm_gated_rst_b_nalb,
       .hqm_inp_gated_rst_b_nalb,
       .hqm_gated_clk_dir,
       .hqm_proc_clk_en_dir                       (i_hqm_qed_pipe_hqm_proc_clk_en_dir),
       .hqm_rst_prep_dir,
       .hqm_gated_rst_b_dir,
       .hqm_inp_gated_rst_b_dir,
       .hqm_inp_gated_clk                         (hqm_inp_gated_clkx),
       .hqm_gated_rst_b_start_qed,
       .hqm_gated_rst_b_active_qed,
       .hqm_gated_rst_b_done_qed,
       .hqm_gated_rst_b_start_nalb,
       .hqm_gated_rst_b_active_nalb,
       .hqm_gated_rst_b_done_nalb,
       .hqm_gated_rst_b_start_dir,
       .hqm_gated_rst_b_active_dir,
       .hqm_gated_rst_b_done_dir,
       .rop_qed_force_clockon                     (i_hqm_reorder_pipe_rop_qed_force_clockon),
       .qed_lsp_deq_v,
       .qed_lsp_deq_data,
       .qed_unit_idle                             (qed_unit_idle_local),
       .qed_unit_pipeidle,
       .qed_reset_done,
       .nalb_unit_idle,
       .nalb_unit_pipeidle,
       .nalb_reset_done,
       .dp_unit_idle,
       .dp_unit_pipeidle,
       .dp_reset_done,
       .qed_cfg_req_up_read                       (i_hqm_reorder_pipe_rop_cfg_req_down_read),
       .qed_cfg_req_up_write                      (i_hqm_reorder_pipe_rop_cfg_req_down_write),
       .qed_cfg_req_up                            (rop_cfg_req_down),
       .qed_cfg_rsp_up_ack                        (i_hqm_reorder_pipe_rop_cfg_rsp_down_ack),
       .qed_cfg_rsp_up                            (rop_cfg_rsp_down),
       .qed_cfg_req_down_read                     (i_hqm_qed_pipe_qed_cfg_req_down_read),
       .qed_cfg_req_down_write                    (i_hqm_qed_pipe_qed_cfg_req_down_write),
       .qed_cfg_req_down,
       .qed_cfg_rsp_down_ack                      (i_hqm_qed_pipe_qed_cfg_rsp_down_ack),
       .qed_cfg_rsp_down,
       .qed_alarm_up_v                            (i_hqm_list_sel_pipe_lsp_alarm_down_v),
       .qed_alarm_up_ready                        (i_hqm_qed_pipe_qed_alarm_up_ready),
       .qed_alarm_up_data                         (lsp_alarm_down_data),
       .qed_alarm_down_v                          (i_hqm_qed_pipe_qed_alarm_down_v),
       .qed_alarm_down_ready                      (i_hqm_reorder_pipe_rop_alarm_up_ready),
       .qed_alarm_down_data,
       .rop_qed_dqed_enq_v                        (i_hqm_reorder_pipe_rop_qed_dqed_enq_v),
       .rop_qed_enq_ready                         (i_hqm_qed_pipe_rop_qed_enq_ready),
       .rop_dqed_enq_ready                        (i_hqm_qed_pipe_rop_dqed_enq_ready),
       .rop_qed_dqed_enq_data,
       .qed_chp_sch_v                             (i_hqm_qed_pipe_qed_chp_sch_v),
       .qed_chp_sch_ready                         (i_hqm_credit_hist_pipe_qed_chp_sch_ready),
       .qed_chp_sch_data,
       .qed_aqed_enq_v                            (i_hqm_qed_pipe_qed_aqed_enq_v),
       .qed_aqed_enq_ready                        (i_hqm_aqed_pipe_qed_aqed_enq_ready),
       .qed_aqed_enq_data,
       .rop_dp_enq_v                              (i_hqm_reorder_pipe_rop_dp_enq_v),
       .rop_dp_enq_ready                          (i_hqm_qed_pipe_rop_dp_enq_ready),
       .rop_dp_enq_data,
       .lsp_dp_sch_dir_v                          (i_hqm_list_sel_pipe_lsp_dp_sch_dir_v),
       .lsp_dp_sch_dir_ready                      (i_hqm_qed_pipe_lsp_dp_sch_dir_ready),
       .lsp_dp_sch_dir_data,
       .lsp_dp_sch_rorply_v                       (i_hqm_list_sel_pipe_lsp_dp_sch_rorply_v),
       .lsp_dp_sch_rorply_ready                   (i_hqm_qed_pipe_lsp_dp_sch_rorply_ready),
       .lsp_dp_sch_rorply_data,
       .dp_lsp_enq_dir_v                          (i_hqm_qed_pipe_dp_lsp_enq_dir_v),
       .dp_lsp_enq_dir_ready                      (i_hqm_list_sel_pipe_dp_lsp_enq_dir_ready),
       .dp_lsp_enq_dir_data,
       .dp_lsp_enq_rorply_v                       (i_hqm_qed_pipe_dp_lsp_enq_rorply_v),
       .dp_lsp_enq_rorply_ready                   (i_hqm_list_sel_pipe_dp_lsp_enq_rorply_ready),
       .dp_lsp_enq_rorply_data,
       .rop_nalb_enq_v                            (i_hqm_reorder_pipe_rop_nalb_enq_v),
       .rop_nalb_enq_ready                        (i_hqm_qed_pipe_rop_nalb_enq_ready),
       .rop_nalb_enq_data,
       .lsp_nalb_sch_unoord_v                     (i_hqm_list_sel_pipe_lsp_nalb_sch_unoord_v),
       .lsp_nalb_sch_unoord_ready                 (i_hqm_qed_pipe_lsp_nalb_sch_unoord_ready),
       .lsp_nalb_sch_unoord_data,
       .lsp_nalb_sch_rorply_v                     (i_hqm_list_sel_pipe_lsp_nalb_sch_rorply_v),
       .lsp_nalb_sch_rorply_ready                 (i_hqm_qed_pipe_lsp_nalb_sch_rorply_ready),
       .lsp_nalb_sch_rorply_data,
       .lsp_nalb_sch_atq_v                        (i_hqm_list_sel_pipe_lsp_nalb_sch_atq_v),
       .lsp_nalb_sch_atq_ready                    (i_hqm_qed_pipe_lsp_nalb_sch_atq_ready),
       .lsp_nalb_sch_atq_data,
       .nalb_lsp_enq_lb_v                         (i_hqm_qed_pipe_nalb_lsp_enq_lb_v),
       .nalb_lsp_enq_lb_ready                     (i_hqm_list_sel_pipe_nalb_lsp_enq_lb_ready),
       .nalb_lsp_enq_lb_data,
       .nalb_lsp_enq_rorply_v                     (i_hqm_qed_pipe_nalb_lsp_enq_rorply_v),
       .nalb_lsp_enq_rorply_ready                 (i_hqm_list_sel_pipe_nalb_lsp_enq_rorply_ready),
       .nalb_lsp_enq_rorply_data,
       .spare_lsp_qed,
       .spare_sys_qed,
       .spare_qed_lsp,
       .spare_qed_sys,
       .rf_qed_chp_sch_data_re                    (i_hqm_qed_pipe_rf_qed_chp_sch_data_re),
       .rf_qed_chp_sch_data_rclk                  (i_hqm_qed_pipe_rf_qed_chp_sch_data_rclk),
       .rf_qed_chp_sch_data_rclk_rst_n            (i_hqm_qed_pipe_rf_qed_chp_sch_data_rclk_rst_n),
       .rf_qed_chp_sch_data_raddr                 (i_hqm_qed_pipe_rf_qed_chp_sch_data_raddr),
       .rf_qed_chp_sch_data_waddr                 (i_hqm_qed_pipe_rf_qed_chp_sch_data_waddr),
       .rf_qed_chp_sch_data_we                    (i_hqm_qed_pipe_rf_qed_chp_sch_data_we),
       .rf_qed_chp_sch_data_wclk                  (i_hqm_qed_pipe_rf_qed_chp_sch_data_wclk),
       .rf_qed_chp_sch_data_wclk_rst_n            (i_hqm_qed_pipe_rf_qed_chp_sch_data_wclk_rst_n),
       .rf_qed_chp_sch_data_wdata                 (i_hqm_qed_pipe_rf_qed_chp_sch_data_wdata),
       .rf_qed_chp_sch_data_rdata                 (i_hqm_qed_pipe_rf_qed_chp_sch_data_rdata),
       .rf_rx_sync_dp_dqed_data_re                (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_re),
       .rf_rx_sync_dp_dqed_data_rclk              (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rclk),
       .rf_rx_sync_dp_dqed_data_rclk_rst_n        (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rclk_rst_n),
       .rf_rx_sync_dp_dqed_data_raddr             (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_raddr),
       .rf_rx_sync_dp_dqed_data_waddr             (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_waddr),
       .rf_rx_sync_dp_dqed_data_we                (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_we),
       .rf_rx_sync_dp_dqed_data_wclk              (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wclk),
       .rf_rx_sync_dp_dqed_data_wclk_rst_n        (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wclk_rst_n),
       .rf_rx_sync_dp_dqed_data_wdata             (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_wdata),
       .rf_rx_sync_dp_dqed_data_rdata             (i_hqm_qed_pipe_rf_rx_sync_dp_dqed_data_rdata),
       .rf_rx_sync_nalb_qed_data_re               (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_re),
       .rf_rx_sync_nalb_qed_data_rclk             (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rclk),
       .rf_rx_sync_nalb_qed_data_rclk_rst_n       (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rclk_rst_n),
       .rf_rx_sync_nalb_qed_data_raddr            (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_raddr),
       .rf_rx_sync_nalb_qed_data_waddr            (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_waddr),
       .rf_rx_sync_nalb_qed_data_we               (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_we),
       .rf_rx_sync_nalb_qed_data_wclk             (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wclk),
       .rf_rx_sync_nalb_qed_data_wclk_rst_n       (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wclk_rst_n),
       .rf_rx_sync_nalb_qed_data_wdata            (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_wdata),
       .rf_rx_sync_nalb_qed_data_rdata            (i_hqm_qed_pipe_rf_rx_sync_nalb_qed_data_rdata),
       .rf_rx_sync_rop_qed_dqed_enq_re            (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_re),
       .rf_rx_sync_rop_qed_dqed_enq_rclk          (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rclk),
       .rf_rx_sync_rop_qed_dqed_enq_rclk_rst_n    (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rclk_rst_n),
       .rf_rx_sync_rop_qed_dqed_enq_raddr         (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_raddr),
       .rf_rx_sync_rop_qed_dqed_enq_waddr         (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_waddr),
       .rf_rx_sync_rop_qed_dqed_enq_we            (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_we),
       .rf_rx_sync_rop_qed_dqed_enq_wclk          (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wclk),
       .rf_rx_sync_rop_qed_dqed_enq_wclk_rst_n    (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wclk_rst_n),
       .rf_rx_sync_rop_qed_dqed_enq_wdata         (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_wdata),
       .rf_rx_sync_rop_qed_dqed_enq_rdata         (i_hqm_qed_pipe_rf_rx_sync_rop_qed_dqed_enq_rdata),
       .sr_qed_0_re                               (i_hqm_qed_pipe_sr_qed_0_re),
       .sr_qed_0_clk                              (i_hqm_qed_pipe_sr_qed_0_clk),
       .sr_qed_0_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_0_clk_rst_n),
       .sr_qed_0_addr                             (i_hqm_qed_pipe_sr_qed_0_addr),
       .sr_qed_0_we                               (i_hqm_qed_pipe_sr_qed_0_we),
       .sr_qed_0_wdata                            (i_hqm_qed_pipe_sr_qed_0_wdata),
       .sr_qed_0_rdata                            (i_hqm_qed_pipe_sr_qed_0_rdata),
       .sr_qed_1_re                               (i_hqm_qed_pipe_sr_qed_1_re),
       .sr_qed_1_clk                              (i_hqm_qed_pipe_sr_qed_1_clk),
       .sr_qed_1_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_1_clk_rst_n),
       .sr_qed_1_addr                             (i_hqm_qed_pipe_sr_qed_1_addr),
       .sr_qed_1_we                               (i_hqm_qed_pipe_sr_qed_1_we),
       .sr_qed_1_wdata                            (i_hqm_qed_pipe_sr_qed_1_wdata),
       .sr_qed_1_rdata                            (i_hqm_qed_pipe_sr_qed_1_rdata),
       .sr_qed_2_re                               (i_hqm_qed_pipe_sr_qed_2_re),
       .sr_qed_2_clk                              (i_hqm_qed_pipe_sr_qed_2_clk),
       .sr_qed_2_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_2_clk_rst_n),
       .sr_qed_2_addr                             (i_hqm_qed_pipe_sr_qed_2_addr),
       .sr_qed_2_we                               (i_hqm_qed_pipe_sr_qed_2_we),
       .sr_qed_2_wdata                            (i_hqm_qed_pipe_sr_qed_2_wdata),
       .sr_qed_2_rdata                            (i_hqm_qed_pipe_sr_qed_2_rdata),
       .sr_qed_3_re                               (i_hqm_qed_pipe_sr_qed_3_re),
       .sr_qed_3_clk                              (i_hqm_qed_pipe_sr_qed_3_clk),
       .sr_qed_3_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_3_clk_rst_n),
       .sr_qed_3_addr                             (i_hqm_qed_pipe_sr_qed_3_addr),
       .sr_qed_3_we                               (i_hqm_qed_pipe_sr_qed_3_we),
       .sr_qed_3_wdata                            (i_hqm_qed_pipe_sr_qed_3_wdata),
       .sr_qed_3_rdata                            (i_hqm_qed_pipe_sr_qed_3_rdata),
       .sr_qed_4_re                               (i_hqm_qed_pipe_sr_qed_4_re),
       .sr_qed_4_clk                              (i_hqm_qed_pipe_sr_qed_4_clk),
       .sr_qed_4_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_4_clk_rst_n),
       .sr_qed_4_addr                             (i_hqm_qed_pipe_sr_qed_4_addr),
       .sr_qed_4_we                               (i_hqm_qed_pipe_sr_qed_4_we),
       .sr_qed_4_wdata                            (i_hqm_qed_pipe_sr_qed_4_wdata),
       .sr_qed_4_rdata                            (i_hqm_qed_pipe_sr_qed_4_rdata),
       .sr_qed_5_re                               (i_hqm_qed_pipe_sr_qed_5_re),
       .sr_qed_5_clk                              (i_hqm_qed_pipe_sr_qed_5_clk),
       .sr_qed_5_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_5_clk_rst_n),
       .sr_qed_5_addr                             (i_hqm_qed_pipe_sr_qed_5_addr),
       .sr_qed_5_we                               (i_hqm_qed_pipe_sr_qed_5_we),
       .sr_qed_5_wdata                            (i_hqm_qed_pipe_sr_qed_5_wdata),
       .sr_qed_5_rdata                            (i_hqm_qed_pipe_sr_qed_5_rdata),
       .sr_qed_6_re                               (i_hqm_qed_pipe_sr_qed_6_re),
       .sr_qed_6_clk                              (i_hqm_qed_pipe_sr_qed_6_clk),
       .sr_qed_6_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_6_clk_rst_n),
       .sr_qed_6_addr                             (i_hqm_qed_pipe_sr_qed_6_addr),
       .sr_qed_6_we                               (i_hqm_qed_pipe_sr_qed_6_we),
       .sr_qed_6_wdata                            (i_hqm_qed_pipe_sr_qed_6_wdata),
       .sr_qed_6_rdata                            (i_hqm_qed_pipe_sr_qed_6_rdata),
       .sr_qed_7_re                               (i_hqm_qed_pipe_sr_qed_7_re),
       .sr_qed_7_clk                              (i_hqm_qed_pipe_sr_qed_7_clk),
       .sr_qed_7_clk_rst_n                        (i_hqm_qed_pipe_sr_qed_7_clk_rst_n),
       .sr_qed_7_addr                             (i_hqm_qed_pipe_sr_qed_7_addr),
       .sr_qed_7_we                               (i_hqm_qed_pipe_sr_qed_7_we),
       .sr_qed_7_wdata                            (i_hqm_qed_pipe_sr_qed_7_wdata),
       .sr_qed_7_rdata                            (i_hqm_qed_pipe_sr_qed_7_rdata),
       .rf_atq_cnt_re                             (i_hqm_qed_pipe_rf_atq_cnt_re),
       .rf_atq_cnt_rclk                           (i_hqm_qed_pipe_rf_atq_cnt_rclk),
       .rf_atq_cnt_rclk_rst_n                     (i_hqm_qed_pipe_rf_atq_cnt_rclk_rst_n),
       .rf_atq_cnt_raddr                          (i_hqm_qed_pipe_rf_atq_cnt_raddr),
       .rf_atq_cnt_waddr                          (i_hqm_qed_pipe_rf_atq_cnt_waddr),
       .rf_atq_cnt_we                             (i_hqm_qed_pipe_rf_atq_cnt_we),
       .rf_atq_cnt_wclk                           (i_hqm_qed_pipe_rf_atq_cnt_wclk),
       .rf_atq_cnt_wclk_rst_n                     (i_hqm_qed_pipe_rf_atq_cnt_wclk_rst_n),
       .rf_atq_cnt_wdata                          (i_hqm_qed_pipe_rf_atq_cnt_wdata),
       .rf_atq_cnt_rdata                          (i_hqm_qed_pipe_rf_atq_cnt_rdata),
       .rf_atq_hp_re                              (i_hqm_qed_pipe_rf_atq_hp_re),
       .rf_atq_hp_rclk                            (i_hqm_qed_pipe_rf_atq_hp_rclk),
       .rf_atq_hp_rclk_rst_n                      (i_hqm_qed_pipe_rf_atq_hp_rclk_rst_n),
       .rf_atq_hp_raddr                           (i_hqm_qed_pipe_rf_atq_hp_raddr),
       .rf_atq_hp_waddr                           (i_hqm_qed_pipe_rf_atq_hp_waddr),
       .rf_atq_hp_we                              (i_hqm_qed_pipe_rf_atq_hp_we),
       .rf_atq_hp_wclk                            (i_hqm_qed_pipe_rf_atq_hp_wclk),
       .rf_atq_hp_wclk_rst_n                      (i_hqm_qed_pipe_rf_atq_hp_wclk_rst_n),
       .rf_atq_hp_wdata                           (i_hqm_qed_pipe_rf_atq_hp_wdata),
       .rf_atq_hp_rdata                           (i_hqm_qed_pipe_rf_atq_hp_rdata),
       .rf_atq_tp_re                              (i_hqm_qed_pipe_rf_atq_tp_re),
       .rf_atq_tp_rclk                            (i_hqm_qed_pipe_rf_atq_tp_rclk),
       .rf_atq_tp_rclk_rst_n                      (i_hqm_qed_pipe_rf_atq_tp_rclk_rst_n),
       .rf_atq_tp_raddr                           (i_hqm_qed_pipe_rf_atq_tp_raddr),
       .rf_atq_tp_waddr                           (i_hqm_qed_pipe_rf_atq_tp_waddr),
       .rf_atq_tp_we                              (i_hqm_qed_pipe_rf_atq_tp_we),
       .rf_atq_tp_wclk                            (i_hqm_qed_pipe_rf_atq_tp_wclk),
       .rf_atq_tp_wclk_rst_n                      (i_hqm_qed_pipe_rf_atq_tp_wclk_rst_n),
       .rf_atq_tp_wdata                           (i_hqm_qed_pipe_rf_atq_tp_wdata),
       .rf_atq_tp_rdata                           (i_hqm_qed_pipe_rf_atq_tp_rdata),
       .rf_lsp_nalb_sch_atq_re                    (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_re),
       .rf_lsp_nalb_sch_atq_rclk                  (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rclk),
       .rf_lsp_nalb_sch_atq_rclk_rst_n            (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rclk_rst_n),
       .rf_lsp_nalb_sch_atq_raddr                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_raddr),
       .rf_lsp_nalb_sch_atq_waddr                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_waddr),
       .rf_lsp_nalb_sch_atq_we                    (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_we),
       .rf_lsp_nalb_sch_atq_wclk                  (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wclk),
       .rf_lsp_nalb_sch_atq_wclk_rst_n            (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wclk_rst_n),
       .rf_lsp_nalb_sch_atq_wdata                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_wdata),
       .rf_lsp_nalb_sch_atq_rdata                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_atq_rdata),
       .rf_lsp_nalb_sch_rorply_re                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_re),
       .rf_lsp_nalb_sch_rorply_rclk               (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rclk),
       .rf_lsp_nalb_sch_rorply_rclk_rst_n         (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rclk_rst_n),
       .rf_lsp_nalb_sch_rorply_raddr              (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_raddr),
       .rf_lsp_nalb_sch_rorply_waddr              (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_waddr),
       .rf_lsp_nalb_sch_rorply_we                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_we),
       .rf_lsp_nalb_sch_rorply_wclk               (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wclk),
       .rf_lsp_nalb_sch_rorply_wclk_rst_n         (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wclk_rst_n),
       .rf_lsp_nalb_sch_rorply_wdata              (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_wdata),
       .rf_lsp_nalb_sch_rorply_rdata              (i_hqm_qed_pipe_rf_lsp_nalb_sch_rorply_rdata),
       .rf_lsp_nalb_sch_unoord_re                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_re),
       .rf_lsp_nalb_sch_unoord_rclk               (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rclk),
       .rf_lsp_nalb_sch_unoord_rclk_rst_n         (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rclk_rst_n),
       .rf_lsp_nalb_sch_unoord_raddr              (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_raddr),
       .rf_lsp_nalb_sch_unoord_waddr              (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_waddr),
       .rf_lsp_nalb_sch_unoord_we                 (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_we),
       .rf_lsp_nalb_sch_unoord_wclk               (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wclk),
       .rf_lsp_nalb_sch_unoord_wclk_rst_n         (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wclk_rst_n),
       .rf_lsp_nalb_sch_unoord_wdata              (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_wdata),
       .rf_lsp_nalb_sch_unoord_rdata              (i_hqm_qed_pipe_rf_lsp_nalb_sch_unoord_rdata),
       .rf_nalb_cnt_re                            (i_hqm_qed_pipe_rf_nalb_cnt_re),
       .rf_nalb_cnt_rclk                          (i_hqm_qed_pipe_rf_nalb_cnt_rclk),
       .rf_nalb_cnt_rclk_rst_n                    (i_hqm_qed_pipe_rf_nalb_cnt_rclk_rst_n),
       .rf_nalb_cnt_raddr                         (i_hqm_qed_pipe_rf_nalb_cnt_raddr),
       .rf_nalb_cnt_waddr                         (i_hqm_qed_pipe_rf_nalb_cnt_waddr),
       .rf_nalb_cnt_we                            (i_hqm_qed_pipe_rf_nalb_cnt_we),
       .rf_nalb_cnt_wclk                          (i_hqm_qed_pipe_rf_nalb_cnt_wclk),
       .rf_nalb_cnt_wclk_rst_n                    (i_hqm_qed_pipe_rf_nalb_cnt_wclk_rst_n),
       .rf_nalb_cnt_wdata                         (i_hqm_qed_pipe_rf_nalb_cnt_wdata),
       .rf_nalb_cnt_rdata                         (i_hqm_qed_pipe_rf_nalb_cnt_rdata),
       .rf_nalb_hp_re                             (i_hqm_qed_pipe_rf_nalb_hp_re),
       .rf_nalb_hp_rclk                           (i_hqm_qed_pipe_rf_nalb_hp_rclk),
       .rf_nalb_hp_rclk_rst_n                     (i_hqm_qed_pipe_rf_nalb_hp_rclk_rst_n),
       .rf_nalb_hp_raddr                          (i_hqm_qed_pipe_rf_nalb_hp_raddr),
       .rf_nalb_hp_waddr                          (i_hqm_qed_pipe_rf_nalb_hp_waddr),
       .rf_nalb_hp_we                             (i_hqm_qed_pipe_rf_nalb_hp_we),
       .rf_nalb_hp_wclk                           (i_hqm_qed_pipe_rf_nalb_hp_wclk),
       .rf_nalb_hp_wclk_rst_n                     (i_hqm_qed_pipe_rf_nalb_hp_wclk_rst_n),
       .rf_nalb_hp_wdata                          (i_hqm_qed_pipe_rf_nalb_hp_wdata),
       .rf_nalb_hp_rdata                          (i_hqm_qed_pipe_rf_nalb_hp_rdata),
       .rf_nalb_lsp_enq_rorply_re                 (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_re),
       .rf_nalb_lsp_enq_rorply_rclk               (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rclk),
       .rf_nalb_lsp_enq_rorply_rclk_rst_n         (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rclk_rst_n),
       .rf_nalb_lsp_enq_rorply_raddr              (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_raddr),
       .rf_nalb_lsp_enq_rorply_waddr              (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_waddr),
       .rf_nalb_lsp_enq_rorply_we                 (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_we),
       .rf_nalb_lsp_enq_rorply_wclk               (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wclk),
       .rf_nalb_lsp_enq_rorply_wclk_rst_n         (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wclk_rst_n),
       .rf_nalb_lsp_enq_rorply_wdata              (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_wdata),
       .rf_nalb_lsp_enq_rorply_rdata              (i_hqm_qed_pipe_rf_nalb_lsp_enq_rorply_rdata),
       .rf_nalb_lsp_enq_unoord_re                 (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_re),
       .rf_nalb_lsp_enq_unoord_rclk               (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rclk),
       .rf_nalb_lsp_enq_unoord_rclk_rst_n         (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rclk_rst_n),
       .rf_nalb_lsp_enq_unoord_raddr              (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_raddr),
       .rf_nalb_lsp_enq_unoord_waddr              (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_waddr),
       .rf_nalb_lsp_enq_unoord_we                 (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_we),
       .rf_nalb_lsp_enq_unoord_wclk               (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wclk),
       .rf_nalb_lsp_enq_unoord_wclk_rst_n         (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wclk_rst_n),
       .rf_nalb_lsp_enq_unoord_wdata              (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_wdata),
       .rf_nalb_lsp_enq_unoord_rdata              (i_hqm_qed_pipe_rf_nalb_lsp_enq_unoord_rdata),
       .rf_nalb_qed_re                            (i_hqm_qed_pipe_rf_nalb_qed_re),
       .rf_nalb_qed_rclk                          (i_hqm_qed_pipe_rf_nalb_qed_rclk),
       .rf_nalb_qed_rclk_rst_n                    (i_hqm_qed_pipe_rf_nalb_qed_rclk_rst_n),
       .rf_nalb_qed_raddr                         (i_hqm_qed_pipe_rf_nalb_qed_raddr),
       .rf_nalb_qed_waddr                         (i_hqm_qed_pipe_rf_nalb_qed_waddr),
       .rf_nalb_qed_we                            (i_hqm_qed_pipe_rf_nalb_qed_we),
       .rf_nalb_qed_wclk                          (i_hqm_qed_pipe_rf_nalb_qed_wclk),
       .rf_nalb_qed_wclk_rst_n                    (i_hqm_qed_pipe_rf_nalb_qed_wclk_rst_n),
       .rf_nalb_qed_wdata                         (i_hqm_qed_pipe_rf_nalb_qed_wdata),
       .rf_nalb_qed_rdata                         (i_hqm_qed_pipe_rf_nalb_qed_rdata),
       .rf_nalb_replay_cnt_re                     (i_hqm_qed_pipe_rf_nalb_replay_cnt_re),
       .rf_nalb_replay_cnt_rclk                   (i_hqm_qed_pipe_rf_nalb_replay_cnt_rclk),
       .rf_nalb_replay_cnt_rclk_rst_n             (i_hqm_qed_pipe_rf_nalb_replay_cnt_rclk_rst_n),
       .rf_nalb_replay_cnt_raddr                  (i_hqm_qed_pipe_rf_nalb_replay_cnt_raddr),
       .rf_nalb_replay_cnt_waddr                  (i_hqm_qed_pipe_rf_nalb_replay_cnt_waddr),
       .rf_nalb_replay_cnt_we                     (i_hqm_qed_pipe_rf_nalb_replay_cnt_we),
       .rf_nalb_replay_cnt_wclk                   (i_hqm_qed_pipe_rf_nalb_replay_cnt_wclk),
       .rf_nalb_replay_cnt_wclk_rst_n             (i_hqm_qed_pipe_rf_nalb_replay_cnt_wclk_rst_n),
       .rf_nalb_replay_cnt_wdata                  (i_hqm_qed_pipe_rf_nalb_replay_cnt_wdata),
       .rf_nalb_replay_cnt_rdata                  (i_hqm_qed_pipe_rf_nalb_replay_cnt_rdata),
       .rf_nalb_replay_hp_re                      (i_hqm_qed_pipe_rf_nalb_replay_hp_re),
       .rf_nalb_replay_hp_rclk                    (i_hqm_qed_pipe_rf_nalb_replay_hp_rclk),
       .rf_nalb_replay_hp_rclk_rst_n              (i_hqm_qed_pipe_rf_nalb_replay_hp_rclk_rst_n),
       .rf_nalb_replay_hp_raddr                   (i_hqm_qed_pipe_rf_nalb_replay_hp_raddr),
       .rf_nalb_replay_hp_waddr                   (i_hqm_qed_pipe_rf_nalb_replay_hp_waddr),
       .rf_nalb_replay_hp_we                      (i_hqm_qed_pipe_rf_nalb_replay_hp_we),
       .rf_nalb_replay_hp_wclk                    (i_hqm_qed_pipe_rf_nalb_replay_hp_wclk),
       .rf_nalb_replay_hp_wclk_rst_n              (i_hqm_qed_pipe_rf_nalb_replay_hp_wclk_rst_n),
       .rf_nalb_replay_hp_wdata                   (i_hqm_qed_pipe_rf_nalb_replay_hp_wdata),
       .rf_nalb_replay_hp_rdata                   (i_hqm_qed_pipe_rf_nalb_replay_hp_rdata),
       .rf_nalb_replay_tp_re                      (i_hqm_qed_pipe_rf_nalb_replay_tp_re),
       .rf_nalb_replay_tp_rclk                    (i_hqm_qed_pipe_rf_nalb_replay_tp_rclk),
       .rf_nalb_replay_tp_rclk_rst_n              (i_hqm_qed_pipe_rf_nalb_replay_tp_rclk_rst_n),
       .rf_nalb_replay_tp_raddr                   (i_hqm_qed_pipe_rf_nalb_replay_tp_raddr),
       .rf_nalb_replay_tp_waddr                   (i_hqm_qed_pipe_rf_nalb_replay_tp_waddr),
       .rf_nalb_replay_tp_we                      (i_hqm_qed_pipe_rf_nalb_replay_tp_we),
       .rf_nalb_replay_tp_wclk                    (i_hqm_qed_pipe_rf_nalb_replay_tp_wclk),
       .rf_nalb_replay_tp_wclk_rst_n              (i_hqm_qed_pipe_rf_nalb_replay_tp_wclk_rst_n),
       .rf_nalb_replay_tp_wdata                   (i_hqm_qed_pipe_rf_nalb_replay_tp_wdata),
       .rf_nalb_replay_tp_rdata                   (i_hqm_qed_pipe_rf_nalb_replay_tp_rdata),
       .rf_nalb_rofrag_cnt_re                     (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_re),
       .rf_nalb_rofrag_cnt_rclk                   (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rclk),
       .rf_nalb_rofrag_cnt_rclk_rst_n             (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rclk_rst_n),
       .rf_nalb_rofrag_cnt_raddr                  (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_raddr),
       .rf_nalb_rofrag_cnt_waddr                  (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_waddr),
       .rf_nalb_rofrag_cnt_we                     (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_we),
       .rf_nalb_rofrag_cnt_wclk                   (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wclk),
       .rf_nalb_rofrag_cnt_wclk_rst_n             (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wclk_rst_n),
       .rf_nalb_rofrag_cnt_wdata                  (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_wdata),
       .rf_nalb_rofrag_cnt_rdata                  (i_hqm_qed_pipe_rf_nalb_rofrag_cnt_rdata),
       .rf_nalb_rofrag_hp_re                      (i_hqm_qed_pipe_rf_nalb_rofrag_hp_re),
       .rf_nalb_rofrag_hp_rclk                    (i_hqm_qed_pipe_rf_nalb_rofrag_hp_rclk),
       .rf_nalb_rofrag_hp_rclk_rst_n              (i_hqm_qed_pipe_rf_nalb_rofrag_hp_rclk_rst_n),
       .rf_nalb_rofrag_hp_raddr                   (i_hqm_qed_pipe_rf_nalb_rofrag_hp_raddr),
       .rf_nalb_rofrag_hp_waddr                   (i_hqm_qed_pipe_rf_nalb_rofrag_hp_waddr),
       .rf_nalb_rofrag_hp_we                      (i_hqm_qed_pipe_rf_nalb_rofrag_hp_we),
       .rf_nalb_rofrag_hp_wclk                    (i_hqm_qed_pipe_rf_nalb_rofrag_hp_wclk),
       .rf_nalb_rofrag_hp_wclk_rst_n              (i_hqm_qed_pipe_rf_nalb_rofrag_hp_wclk_rst_n),
       .rf_nalb_rofrag_hp_wdata                   (i_hqm_qed_pipe_rf_nalb_rofrag_hp_wdata),
       .rf_nalb_rofrag_hp_rdata                   (i_hqm_qed_pipe_rf_nalb_rofrag_hp_rdata),
       .rf_nalb_rofrag_tp_re                      (i_hqm_qed_pipe_rf_nalb_rofrag_tp_re),
       .rf_nalb_rofrag_tp_rclk                    (i_hqm_qed_pipe_rf_nalb_rofrag_tp_rclk),
       .rf_nalb_rofrag_tp_rclk_rst_n              (i_hqm_qed_pipe_rf_nalb_rofrag_tp_rclk_rst_n),
       .rf_nalb_rofrag_tp_raddr                   (i_hqm_qed_pipe_rf_nalb_rofrag_tp_raddr),
       .rf_nalb_rofrag_tp_waddr                   (i_hqm_qed_pipe_rf_nalb_rofrag_tp_waddr),
       .rf_nalb_rofrag_tp_we                      (i_hqm_qed_pipe_rf_nalb_rofrag_tp_we),
       .rf_nalb_rofrag_tp_wclk                    (i_hqm_qed_pipe_rf_nalb_rofrag_tp_wclk),
       .rf_nalb_rofrag_tp_wclk_rst_n              (i_hqm_qed_pipe_rf_nalb_rofrag_tp_wclk_rst_n),
       .rf_nalb_rofrag_tp_wdata                   (i_hqm_qed_pipe_rf_nalb_rofrag_tp_wdata),
       .rf_nalb_rofrag_tp_rdata                   (i_hqm_qed_pipe_rf_nalb_rofrag_tp_rdata),
       .rf_nalb_tp_re                             (i_hqm_qed_pipe_rf_nalb_tp_re),
       .rf_nalb_tp_rclk                           (i_hqm_qed_pipe_rf_nalb_tp_rclk),
       .rf_nalb_tp_rclk_rst_n                     (i_hqm_qed_pipe_rf_nalb_tp_rclk_rst_n),
       .rf_nalb_tp_raddr                          (i_hqm_qed_pipe_rf_nalb_tp_raddr),
       .rf_nalb_tp_waddr                          (i_hqm_qed_pipe_rf_nalb_tp_waddr),
       .rf_nalb_tp_we                             (i_hqm_qed_pipe_rf_nalb_tp_we),
       .rf_nalb_tp_wclk                           (i_hqm_qed_pipe_rf_nalb_tp_wclk),
       .rf_nalb_tp_wclk_rst_n                     (i_hqm_qed_pipe_rf_nalb_tp_wclk_rst_n),
       .rf_nalb_tp_wdata                          (i_hqm_qed_pipe_rf_nalb_tp_wdata),
       .rf_nalb_tp_rdata                          (i_hqm_qed_pipe_rf_nalb_tp_rdata),
       .rf_rop_nalb_enq_ro_re                     (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_re),
       .rf_rop_nalb_enq_ro_rclk                   (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rclk),
       .rf_rop_nalb_enq_ro_rclk_rst_n             (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rclk_rst_n),
       .rf_rop_nalb_enq_ro_raddr                  (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_raddr),
       .rf_rop_nalb_enq_ro_waddr                  (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_waddr),
       .rf_rop_nalb_enq_ro_we                     (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_we),
       .rf_rop_nalb_enq_ro_wclk                   (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wclk),
       .rf_rop_nalb_enq_ro_wclk_rst_n             (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wclk_rst_n),
       .rf_rop_nalb_enq_ro_wdata                  (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_wdata),
       .rf_rop_nalb_enq_ro_rdata                  (i_hqm_qed_pipe_rf_rop_nalb_enq_ro_rdata),
       .rf_rop_nalb_enq_unoord_re                 (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_re),
       .rf_rop_nalb_enq_unoord_rclk               (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rclk),
       .rf_rop_nalb_enq_unoord_rclk_rst_n         (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rclk_rst_n),
       .rf_rop_nalb_enq_unoord_raddr              (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_raddr),
       .rf_rop_nalb_enq_unoord_waddr              (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_waddr),
       .rf_rop_nalb_enq_unoord_we                 (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_we),
       .rf_rop_nalb_enq_unoord_wclk               (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wclk),
       .rf_rop_nalb_enq_unoord_wclk_rst_n         (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wclk_rst_n),
       .rf_rop_nalb_enq_unoord_wdata              (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_wdata),
       .rf_rop_nalb_enq_unoord_rdata              (i_hqm_qed_pipe_rf_rop_nalb_enq_unoord_rdata),
       .rf_rx_sync_lsp_nalb_sch_atq_re            (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_re),
       .rf_rx_sync_lsp_nalb_sch_atq_rclk          (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rclk),
       .rf_rx_sync_lsp_nalb_sch_atq_rclk_rst_n    (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_atq_raddr         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_raddr),
       .rf_rx_sync_lsp_nalb_sch_atq_waddr         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_waddr),
       .rf_rx_sync_lsp_nalb_sch_atq_we            (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_we),
       .rf_rx_sync_lsp_nalb_sch_atq_wclk          (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wclk),
       .rf_rx_sync_lsp_nalb_sch_atq_wclk_rst_n    (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_atq_wdata         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_wdata),
       .rf_rx_sync_lsp_nalb_sch_atq_rdata         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_atq_rdata),
       .rf_rx_sync_lsp_nalb_sch_rorply_re         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_re),
       .rf_rx_sync_lsp_nalb_sch_rorply_rclk       (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rclk),
       .rf_rx_sync_lsp_nalb_sch_rorply_rclk_rst_n (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_rorply_raddr      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_raddr),
       .rf_rx_sync_lsp_nalb_sch_rorply_waddr      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_waddr),
       .rf_rx_sync_lsp_nalb_sch_rorply_we         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_we),
       .rf_rx_sync_lsp_nalb_sch_rorply_wclk       (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wclk),
       .rf_rx_sync_lsp_nalb_sch_rorply_wclk_rst_n (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_rorply_wdata      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_wdata),
       .rf_rx_sync_lsp_nalb_sch_rorply_rdata      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_rorply_rdata),
       .rf_rx_sync_lsp_nalb_sch_unoord_re         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_re),
       .rf_rx_sync_lsp_nalb_sch_unoord_rclk       (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rclk),
       .rf_rx_sync_lsp_nalb_sch_unoord_rclk_rst_n (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_unoord_raddr      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_raddr),
       .rf_rx_sync_lsp_nalb_sch_unoord_waddr      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_waddr),
       .rf_rx_sync_lsp_nalb_sch_unoord_we         (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_we),
       .rf_rx_sync_lsp_nalb_sch_unoord_wclk       (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wclk),
       .rf_rx_sync_lsp_nalb_sch_unoord_wclk_rst_n (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wclk_rst_n),
       .rf_rx_sync_lsp_nalb_sch_unoord_wdata      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_wdata),
       .rf_rx_sync_lsp_nalb_sch_unoord_rdata      (i_hqm_qed_pipe_rf_rx_sync_lsp_nalb_sch_unoord_rdata),
       .rf_rx_sync_rop_nalb_enq_re                (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_re),
       .rf_rx_sync_rop_nalb_enq_rclk              (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rclk),
       .rf_rx_sync_rop_nalb_enq_rclk_rst_n        (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rclk_rst_n),
       .rf_rx_sync_rop_nalb_enq_raddr             (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_raddr),
       .rf_rx_sync_rop_nalb_enq_waddr             (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_waddr),
       .rf_rx_sync_rop_nalb_enq_we                (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_we),
       .rf_rx_sync_rop_nalb_enq_wclk              (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wclk),
       .rf_rx_sync_rop_nalb_enq_wclk_rst_n        (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wclk_rst_n),
       .rf_rx_sync_rop_nalb_enq_wdata             (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_wdata),
       .rf_rx_sync_rop_nalb_enq_rdata             (i_hqm_qed_pipe_rf_rx_sync_rop_nalb_enq_rdata),
       .sr_nalb_nxthp_re                          (i_hqm_qed_pipe_sr_nalb_nxthp_re),
       .sr_nalb_nxthp_clk                         (i_hqm_qed_pipe_sr_nalb_nxthp_clk),
       .sr_nalb_nxthp_clk_rst_n                   (i_hqm_qed_pipe_sr_nalb_nxthp_clk_rst_n),
       .sr_nalb_nxthp_addr                        (i_hqm_qed_pipe_sr_nalb_nxthp_addr),
       .sr_nalb_nxthp_we                          (i_hqm_qed_pipe_sr_nalb_nxthp_we),
       .sr_nalb_nxthp_wdata                       (i_hqm_qed_pipe_sr_nalb_nxthp_wdata),
       .sr_nalb_nxthp_rdata                       (i_hqm_qed_pipe_sr_nalb_nxthp_rdata),
       .rf_dir_cnt_re                             (i_hqm_qed_pipe_rf_dir_cnt_re),
       .rf_dir_cnt_rclk                           (i_hqm_qed_pipe_rf_dir_cnt_rclk),
       .rf_dir_cnt_rclk_rst_n                     (i_hqm_qed_pipe_rf_dir_cnt_rclk_rst_n),
       .rf_dir_cnt_raddr                          (i_hqm_qed_pipe_rf_dir_cnt_raddr),
       .rf_dir_cnt_waddr                          (i_hqm_qed_pipe_rf_dir_cnt_waddr),
       .rf_dir_cnt_we                             (i_hqm_qed_pipe_rf_dir_cnt_we),
       .rf_dir_cnt_wclk                           (i_hqm_qed_pipe_rf_dir_cnt_wclk),
       .rf_dir_cnt_wclk_rst_n                     (i_hqm_qed_pipe_rf_dir_cnt_wclk_rst_n),
       .rf_dir_cnt_wdata                          (i_hqm_qed_pipe_rf_dir_cnt_wdata),
       .rf_dir_cnt_rdata                          (i_hqm_qed_pipe_rf_dir_cnt_rdata),
       .rf_dir_hp_re                              (i_hqm_qed_pipe_rf_dir_hp_re),
       .rf_dir_hp_rclk                            (i_hqm_qed_pipe_rf_dir_hp_rclk),
       .rf_dir_hp_rclk_rst_n                      (i_hqm_qed_pipe_rf_dir_hp_rclk_rst_n),
       .rf_dir_hp_raddr                           (i_hqm_qed_pipe_rf_dir_hp_raddr),
       .rf_dir_hp_waddr                           (i_hqm_qed_pipe_rf_dir_hp_waddr),
       .rf_dir_hp_we                              (i_hqm_qed_pipe_rf_dir_hp_we),
       .rf_dir_hp_wclk                            (i_hqm_qed_pipe_rf_dir_hp_wclk),
       .rf_dir_hp_wclk_rst_n                      (i_hqm_qed_pipe_rf_dir_hp_wclk_rst_n),
       .rf_dir_hp_wdata                           (i_hqm_qed_pipe_rf_dir_hp_wdata),
       .rf_dir_hp_rdata                           (i_hqm_qed_pipe_rf_dir_hp_rdata),
       .rf_dir_replay_cnt_re                      (i_hqm_qed_pipe_rf_dir_replay_cnt_re),
       .rf_dir_replay_cnt_rclk                    (i_hqm_qed_pipe_rf_dir_replay_cnt_rclk),
       .rf_dir_replay_cnt_rclk_rst_n              (i_hqm_qed_pipe_rf_dir_replay_cnt_rclk_rst_n),
       .rf_dir_replay_cnt_raddr                   (i_hqm_qed_pipe_rf_dir_replay_cnt_raddr),
       .rf_dir_replay_cnt_waddr                   (i_hqm_qed_pipe_rf_dir_replay_cnt_waddr),
       .rf_dir_replay_cnt_we                      (i_hqm_qed_pipe_rf_dir_replay_cnt_we),
       .rf_dir_replay_cnt_wclk                    (i_hqm_qed_pipe_rf_dir_replay_cnt_wclk),
       .rf_dir_replay_cnt_wclk_rst_n              (i_hqm_qed_pipe_rf_dir_replay_cnt_wclk_rst_n),
       .rf_dir_replay_cnt_wdata                   (i_hqm_qed_pipe_rf_dir_replay_cnt_wdata),
       .rf_dir_replay_cnt_rdata                   (i_hqm_qed_pipe_rf_dir_replay_cnt_rdata),
       .rf_dir_replay_hp_re                       (i_hqm_qed_pipe_rf_dir_replay_hp_re),
       .rf_dir_replay_hp_rclk                     (i_hqm_qed_pipe_rf_dir_replay_hp_rclk),
       .rf_dir_replay_hp_rclk_rst_n               (i_hqm_qed_pipe_rf_dir_replay_hp_rclk_rst_n),
       .rf_dir_replay_hp_raddr                    (i_hqm_qed_pipe_rf_dir_replay_hp_raddr),
       .rf_dir_replay_hp_waddr                    (i_hqm_qed_pipe_rf_dir_replay_hp_waddr),
       .rf_dir_replay_hp_we                       (i_hqm_qed_pipe_rf_dir_replay_hp_we),
       .rf_dir_replay_hp_wclk                     (i_hqm_qed_pipe_rf_dir_replay_hp_wclk),
       .rf_dir_replay_hp_wclk_rst_n               (i_hqm_qed_pipe_rf_dir_replay_hp_wclk_rst_n),
       .rf_dir_replay_hp_wdata                    (i_hqm_qed_pipe_rf_dir_replay_hp_wdata),
       .rf_dir_replay_hp_rdata                    (i_hqm_qed_pipe_rf_dir_replay_hp_rdata),
       .rf_dir_replay_tp_re                       (i_hqm_qed_pipe_rf_dir_replay_tp_re),
       .rf_dir_replay_tp_rclk                     (i_hqm_qed_pipe_rf_dir_replay_tp_rclk),
       .rf_dir_replay_tp_rclk_rst_n               (i_hqm_qed_pipe_rf_dir_replay_tp_rclk_rst_n),
       .rf_dir_replay_tp_raddr                    (i_hqm_qed_pipe_rf_dir_replay_tp_raddr),
       .rf_dir_replay_tp_waddr                    (i_hqm_qed_pipe_rf_dir_replay_tp_waddr),
       .rf_dir_replay_tp_we                       (i_hqm_qed_pipe_rf_dir_replay_tp_we),
       .rf_dir_replay_tp_wclk                     (i_hqm_qed_pipe_rf_dir_replay_tp_wclk),
       .rf_dir_replay_tp_wclk_rst_n               (i_hqm_qed_pipe_rf_dir_replay_tp_wclk_rst_n),
       .rf_dir_replay_tp_wdata                    (i_hqm_qed_pipe_rf_dir_replay_tp_wdata),
       .rf_dir_replay_tp_rdata                    (i_hqm_qed_pipe_rf_dir_replay_tp_rdata),
       .rf_dir_rofrag_cnt_re                      (i_hqm_qed_pipe_rf_dir_rofrag_cnt_re),
       .rf_dir_rofrag_cnt_rclk                    (i_hqm_qed_pipe_rf_dir_rofrag_cnt_rclk),
       .rf_dir_rofrag_cnt_rclk_rst_n              (i_hqm_qed_pipe_rf_dir_rofrag_cnt_rclk_rst_n),
       .rf_dir_rofrag_cnt_raddr                   (i_hqm_qed_pipe_rf_dir_rofrag_cnt_raddr),
       .rf_dir_rofrag_cnt_waddr                   (i_hqm_qed_pipe_rf_dir_rofrag_cnt_waddr),
       .rf_dir_rofrag_cnt_we                      (i_hqm_qed_pipe_rf_dir_rofrag_cnt_we),
       .rf_dir_rofrag_cnt_wclk                    (i_hqm_qed_pipe_rf_dir_rofrag_cnt_wclk),
       .rf_dir_rofrag_cnt_wclk_rst_n              (i_hqm_qed_pipe_rf_dir_rofrag_cnt_wclk_rst_n),
       .rf_dir_rofrag_cnt_wdata                   (i_hqm_qed_pipe_rf_dir_rofrag_cnt_wdata),
       .rf_dir_rofrag_cnt_rdata                   (i_hqm_qed_pipe_rf_dir_rofrag_cnt_rdata),
       .rf_dir_rofrag_hp_re                       (i_hqm_qed_pipe_rf_dir_rofrag_hp_re),
       .rf_dir_rofrag_hp_rclk                     (i_hqm_qed_pipe_rf_dir_rofrag_hp_rclk),
       .rf_dir_rofrag_hp_rclk_rst_n               (i_hqm_qed_pipe_rf_dir_rofrag_hp_rclk_rst_n),
       .rf_dir_rofrag_hp_raddr                    (i_hqm_qed_pipe_rf_dir_rofrag_hp_raddr),
       .rf_dir_rofrag_hp_waddr                    (i_hqm_qed_pipe_rf_dir_rofrag_hp_waddr),
       .rf_dir_rofrag_hp_we                       (i_hqm_qed_pipe_rf_dir_rofrag_hp_we),
       .rf_dir_rofrag_hp_wclk                     (i_hqm_qed_pipe_rf_dir_rofrag_hp_wclk),
       .rf_dir_rofrag_hp_wclk_rst_n               (i_hqm_qed_pipe_rf_dir_rofrag_hp_wclk_rst_n),
       .rf_dir_rofrag_hp_wdata                    (i_hqm_qed_pipe_rf_dir_rofrag_hp_wdata),
       .rf_dir_rofrag_hp_rdata                    (i_hqm_qed_pipe_rf_dir_rofrag_hp_rdata),
       .rf_dir_rofrag_tp_re                       (i_hqm_qed_pipe_rf_dir_rofrag_tp_re),
       .rf_dir_rofrag_tp_rclk                     (i_hqm_qed_pipe_rf_dir_rofrag_tp_rclk),
       .rf_dir_rofrag_tp_rclk_rst_n               (i_hqm_qed_pipe_rf_dir_rofrag_tp_rclk_rst_n),
       .rf_dir_rofrag_tp_raddr                    (i_hqm_qed_pipe_rf_dir_rofrag_tp_raddr),
       .rf_dir_rofrag_tp_waddr                    (i_hqm_qed_pipe_rf_dir_rofrag_tp_waddr),
       .rf_dir_rofrag_tp_we                       (i_hqm_qed_pipe_rf_dir_rofrag_tp_we),
       .rf_dir_rofrag_tp_wclk                     (i_hqm_qed_pipe_rf_dir_rofrag_tp_wclk),
       .rf_dir_rofrag_tp_wclk_rst_n               (i_hqm_qed_pipe_rf_dir_rofrag_tp_wclk_rst_n),
       .rf_dir_rofrag_tp_wdata                    (i_hqm_qed_pipe_rf_dir_rofrag_tp_wdata),
       .rf_dir_rofrag_tp_rdata                    (i_hqm_qed_pipe_rf_dir_rofrag_tp_rdata),
       .rf_dir_tp_re                              (i_hqm_qed_pipe_rf_dir_tp_re),
       .rf_dir_tp_rclk                            (i_hqm_qed_pipe_rf_dir_tp_rclk),
       .rf_dir_tp_rclk_rst_n                      (i_hqm_qed_pipe_rf_dir_tp_rclk_rst_n),
       .rf_dir_tp_raddr                           (i_hqm_qed_pipe_rf_dir_tp_raddr),
       .rf_dir_tp_waddr                           (i_hqm_qed_pipe_rf_dir_tp_waddr),
       .rf_dir_tp_we                              (i_hqm_qed_pipe_rf_dir_tp_we),
       .rf_dir_tp_wclk                            (i_hqm_qed_pipe_rf_dir_tp_wclk),
       .rf_dir_tp_wclk_rst_n                      (i_hqm_qed_pipe_rf_dir_tp_wclk_rst_n),
       .rf_dir_tp_wdata                           (i_hqm_qed_pipe_rf_dir_tp_wdata),
       .rf_dir_tp_rdata                           (i_hqm_qed_pipe_rf_dir_tp_rdata),
       .rf_dp_dqed_re                             (i_hqm_qed_pipe_rf_dp_dqed_re),
       .rf_dp_dqed_rclk                           (i_hqm_qed_pipe_rf_dp_dqed_rclk),
       .rf_dp_dqed_rclk_rst_n                     (i_hqm_qed_pipe_rf_dp_dqed_rclk_rst_n),
       .rf_dp_dqed_raddr                          (i_hqm_qed_pipe_rf_dp_dqed_raddr),
       .rf_dp_dqed_waddr                          (i_hqm_qed_pipe_rf_dp_dqed_waddr),
       .rf_dp_dqed_we                             (i_hqm_qed_pipe_rf_dp_dqed_we),
       .rf_dp_dqed_wclk                           (i_hqm_qed_pipe_rf_dp_dqed_wclk),
       .rf_dp_dqed_wclk_rst_n                     (i_hqm_qed_pipe_rf_dp_dqed_wclk_rst_n),
       .rf_dp_dqed_wdata                          (i_hqm_qed_pipe_rf_dp_dqed_wdata),
       .rf_dp_dqed_rdata                          (i_hqm_qed_pipe_rf_dp_dqed_rdata),
       .rf_dp_lsp_enq_dir_re                      (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_re),
       .rf_dp_lsp_enq_dir_rclk                    (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rclk),
       .rf_dp_lsp_enq_dir_rclk_rst_n              (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rclk_rst_n),
       .rf_dp_lsp_enq_dir_raddr                   (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_raddr),
       .rf_dp_lsp_enq_dir_waddr                   (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_waddr),
       .rf_dp_lsp_enq_dir_we                      (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_we),
       .rf_dp_lsp_enq_dir_wclk                    (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wclk),
       .rf_dp_lsp_enq_dir_wclk_rst_n              (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wclk_rst_n),
       .rf_dp_lsp_enq_dir_wdata                   (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_wdata),
       .rf_dp_lsp_enq_dir_rdata                   (i_hqm_qed_pipe_rf_dp_lsp_enq_dir_rdata),
       .rf_dp_lsp_enq_rorply_re                   (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_re),
       .rf_dp_lsp_enq_rorply_rclk                 (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rclk),
       .rf_dp_lsp_enq_rorply_rclk_rst_n           (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rclk_rst_n),
       .rf_dp_lsp_enq_rorply_raddr                (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_raddr),
       .rf_dp_lsp_enq_rorply_waddr                (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_waddr),
       .rf_dp_lsp_enq_rorply_we                   (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_we),
       .rf_dp_lsp_enq_rorply_wclk                 (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wclk),
       .rf_dp_lsp_enq_rorply_wclk_rst_n           (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wclk_rst_n),
       .rf_dp_lsp_enq_rorply_wdata                (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_wdata),
       .rf_dp_lsp_enq_rorply_rdata                (i_hqm_qed_pipe_rf_dp_lsp_enq_rorply_rdata),
       .rf_lsp_dp_sch_dir_re                      (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_re),
       .rf_lsp_dp_sch_dir_rclk                    (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rclk),
       .rf_lsp_dp_sch_dir_rclk_rst_n              (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rclk_rst_n),
       .rf_lsp_dp_sch_dir_raddr                   (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_raddr),
       .rf_lsp_dp_sch_dir_waddr                   (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_waddr),
       .rf_lsp_dp_sch_dir_we                      (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_we),
       .rf_lsp_dp_sch_dir_wclk                    (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wclk),
       .rf_lsp_dp_sch_dir_wclk_rst_n              (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wclk_rst_n),
       .rf_lsp_dp_sch_dir_wdata                   (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_wdata),
       .rf_lsp_dp_sch_dir_rdata                   (i_hqm_qed_pipe_rf_lsp_dp_sch_dir_rdata),
       .rf_lsp_dp_sch_rorply_re                   (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_re),
       .rf_lsp_dp_sch_rorply_rclk                 (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rclk),
       .rf_lsp_dp_sch_rorply_rclk_rst_n           (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rclk_rst_n),
       .rf_lsp_dp_sch_rorply_raddr                (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_raddr),
       .rf_lsp_dp_sch_rorply_waddr                (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_waddr),
       .rf_lsp_dp_sch_rorply_we                   (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_we),
       .rf_lsp_dp_sch_rorply_wclk                 (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wclk),
       .rf_lsp_dp_sch_rorply_wclk_rst_n           (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wclk_rst_n),
       .rf_lsp_dp_sch_rorply_wdata                (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_wdata),
       .rf_lsp_dp_sch_rorply_rdata                (i_hqm_qed_pipe_rf_lsp_dp_sch_rorply_rdata),
       .rf_rop_dp_enq_dir_re                      (i_hqm_qed_pipe_rf_rop_dp_enq_dir_re),
       .rf_rop_dp_enq_dir_rclk                    (i_hqm_qed_pipe_rf_rop_dp_enq_dir_rclk),
       .rf_rop_dp_enq_dir_rclk_rst_n              (i_hqm_qed_pipe_rf_rop_dp_enq_dir_rclk_rst_n),
       .rf_rop_dp_enq_dir_raddr                   (i_hqm_qed_pipe_rf_rop_dp_enq_dir_raddr),
       .rf_rop_dp_enq_dir_waddr                   (i_hqm_qed_pipe_rf_rop_dp_enq_dir_waddr),
       .rf_rop_dp_enq_dir_we                      (i_hqm_qed_pipe_rf_rop_dp_enq_dir_we),
       .rf_rop_dp_enq_dir_wclk                    (i_hqm_qed_pipe_rf_rop_dp_enq_dir_wclk),
       .rf_rop_dp_enq_dir_wclk_rst_n              (i_hqm_qed_pipe_rf_rop_dp_enq_dir_wclk_rst_n),
       .rf_rop_dp_enq_dir_wdata                   (i_hqm_qed_pipe_rf_rop_dp_enq_dir_wdata),
       .rf_rop_dp_enq_dir_rdata                   (i_hqm_qed_pipe_rf_rop_dp_enq_dir_rdata),
       .rf_rop_dp_enq_ro_re                       (i_hqm_qed_pipe_rf_rop_dp_enq_ro_re),
       .rf_rop_dp_enq_ro_rclk                     (i_hqm_qed_pipe_rf_rop_dp_enq_ro_rclk),
       .rf_rop_dp_enq_ro_rclk_rst_n               (i_hqm_qed_pipe_rf_rop_dp_enq_ro_rclk_rst_n),
       .rf_rop_dp_enq_ro_raddr                    (i_hqm_qed_pipe_rf_rop_dp_enq_ro_raddr),
       .rf_rop_dp_enq_ro_waddr                    (i_hqm_qed_pipe_rf_rop_dp_enq_ro_waddr),
       .rf_rop_dp_enq_ro_we                       (i_hqm_qed_pipe_rf_rop_dp_enq_ro_we),
       .rf_rop_dp_enq_ro_wclk                     (i_hqm_qed_pipe_rf_rop_dp_enq_ro_wclk),
       .rf_rop_dp_enq_ro_wclk_rst_n               (i_hqm_qed_pipe_rf_rop_dp_enq_ro_wclk_rst_n),
       .rf_rop_dp_enq_ro_wdata                    (i_hqm_qed_pipe_rf_rop_dp_enq_ro_wdata),
       .rf_rop_dp_enq_ro_rdata                    (i_hqm_qed_pipe_rf_rop_dp_enq_ro_rdata),
       .rf_rx_sync_lsp_dp_sch_dir_re              (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_re),
       .rf_rx_sync_lsp_dp_sch_dir_rclk            (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rclk),
       .rf_rx_sync_lsp_dp_sch_dir_rclk_rst_n      (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rclk_rst_n),
       .rf_rx_sync_lsp_dp_sch_dir_raddr           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_raddr),
       .rf_rx_sync_lsp_dp_sch_dir_waddr           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_waddr),
       .rf_rx_sync_lsp_dp_sch_dir_we              (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_we),
       .rf_rx_sync_lsp_dp_sch_dir_wclk            (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wclk),
       .rf_rx_sync_lsp_dp_sch_dir_wclk_rst_n      (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wclk_rst_n),
       .rf_rx_sync_lsp_dp_sch_dir_wdata           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_wdata),
       .rf_rx_sync_lsp_dp_sch_dir_rdata           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_dir_rdata),
       .rf_rx_sync_lsp_dp_sch_rorply_re           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_re),
       .rf_rx_sync_lsp_dp_sch_rorply_rclk         (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rclk),
       .rf_rx_sync_lsp_dp_sch_rorply_rclk_rst_n   (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rclk_rst_n),
       .rf_rx_sync_lsp_dp_sch_rorply_raddr        (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_raddr),
       .rf_rx_sync_lsp_dp_sch_rorply_waddr        (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_waddr),
       .rf_rx_sync_lsp_dp_sch_rorply_we           (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_we),
       .rf_rx_sync_lsp_dp_sch_rorply_wclk         (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wclk),
       .rf_rx_sync_lsp_dp_sch_rorply_wclk_rst_n   (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wclk_rst_n),
       .rf_rx_sync_lsp_dp_sch_rorply_wdata        (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_wdata),
       .rf_rx_sync_lsp_dp_sch_rorply_rdata        (i_hqm_qed_pipe_rf_rx_sync_lsp_dp_sch_rorply_rdata),
       .rf_rx_sync_rop_dp_enq_re                  (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_re),
       .rf_rx_sync_rop_dp_enq_rclk                (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rclk),
       .rf_rx_sync_rop_dp_enq_rclk_rst_n          (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rclk_rst_n),
       .rf_rx_sync_rop_dp_enq_raddr               (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_raddr),
       .rf_rx_sync_rop_dp_enq_waddr               (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_waddr),
       .rf_rx_sync_rop_dp_enq_we                  (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_we),
       .rf_rx_sync_rop_dp_enq_wclk                (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wclk),
       .rf_rx_sync_rop_dp_enq_wclk_rst_n          (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wclk_rst_n),
       .rf_rx_sync_rop_dp_enq_wdata               (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_wdata),
       .rf_rx_sync_rop_dp_enq_rdata               (i_hqm_qed_pipe_rf_rx_sync_rop_dp_enq_rdata),
       .sr_dir_nxthp_re                           (i_hqm_qed_pipe_sr_dir_nxthp_re),
       .sr_dir_nxthp_clk                          (i_hqm_qed_pipe_sr_dir_nxthp_clk),
       .sr_dir_nxthp_clk_rst_n                    (i_hqm_qed_pipe_sr_dir_nxthp_clk_rst_n),
       .sr_dir_nxthp_addr                         (i_hqm_qed_pipe_sr_dir_nxthp_addr),
       .sr_dir_nxthp_we                           (i_hqm_qed_pipe_sr_dir_nxthp_we),
       .sr_dir_nxthp_wdata                        (i_hqm_qed_pipe_sr_dir_nxthp_wdata),
       .sr_dir_nxthp_rdata                        (i_hqm_qed_pipe_sr_dir_nxthp_rdata));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_qed_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_qed),
       .hqm_gated_clk          (hqm_gated_clk_qed),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_qed),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_qed),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_qed),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_qed),
       .hqm_flr_prep           (hqm_flr_prep_rptrx),
       .rst_prep               (hqm_rst_prep_qed));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_qed_unit_idle_and2
      (.clki0 (qed_unit_idle_local),
       .clki1 (hqm_flr_prep_b),
       .clko  (qed_unit_idle_qual));

   hqm_AW_flop i_hqm_qed_unit_idle_ft_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bx),
       .data   (qed_unit_idle_qual),
       .data_q (qed_unit_idle));

   hqm_reorder_pipe i_hqm_reorder_pipe
      (.hqm_gated_clk                          (hqm_gated_clk_chp),
       .hqm_inp_gated_clk                      (hqm_inp_gated_clkxx),
       .hqm_rst_prep_rop,
       .hqm_gated_rst_b_rop,
       .hqm_inp_gated_rst_b_rop,
       .hqm_gated_rst_b_start_rop,
       .hqm_gated_rst_b_active_rop,
       .hqm_gated_rst_b_done_rop,
       .rop_clk_idle,
       .rop_clk_enable,
       .rop_unit_idle                          (i_hqm_reorder_pipe_rop_unit_idle),
       .rop_unit_pipeidle,
       .rop_reset_done,
       .rop_cfg_req_up_read                    (i_hqm_credit_hist_pipe_chp_cfg_req_down_read),
       .rop_cfg_req_up_write                   (i_hqm_credit_hist_pipe_chp_cfg_req_down_write),
       .rop_cfg_req_up                         (chp_cfg_req_down),
       .rop_cfg_rsp_up_ack                     (i_hqm_credit_hist_pipe_chp_cfg_rsp_down_ack),
       .rop_cfg_rsp_up                         (chp_cfg_rsp_down),
       .rop_cfg_req_down_read                  (i_hqm_reorder_pipe_rop_cfg_req_down_read),
       .rop_cfg_req_down_write                 (i_hqm_reorder_pipe_rop_cfg_req_down_write),
       .rop_cfg_req_down,
       .rop_cfg_rsp_down_ack                   (i_hqm_reorder_pipe_rop_cfg_rsp_down_ack),
       .rop_cfg_rsp_down,
       .rop_alarm_up_v                         (i_hqm_qed_pipe_qed_alarm_down_v),
       .rop_alarm_up_ready                     (i_hqm_reorder_pipe_rop_alarm_up_ready),
       .rop_alarm_up_data                      (qed_alarm_down_data),
       .rop_alarm_down_v                       (i_hqm_reorder_pipe_rop_alarm_down_v),
       .rop_alarm_down_ready                   (i_hqm_credit_hist_pipe_chp_alarm_up_ready),
       .rop_alarm_down_data,
       .chp_rop_hcw_v                          (i_hqm_credit_hist_pipe_chp_rop_hcw_v),
       .chp_rop_hcw_ready                      (i_hqm_reorder_pipe_chp_rop_hcw_ready),
       .chp_rop_hcw_data,
       .rop_dp_enq_v                           (i_hqm_reorder_pipe_rop_dp_enq_v),
       .rop_dp_enq_ready                       (i_hqm_qed_pipe_rop_dp_enq_ready),
       .rop_dp_enq_data,
       .rop_nalb_enq_v                         (i_hqm_reorder_pipe_rop_nalb_enq_v),
       .rop_nalb_enq_ready                     (i_hqm_qed_pipe_rop_nalb_enq_ready),
       .rop_nalb_enq_data,
       .rop_qed_dqed_enq_v                     (i_hqm_reorder_pipe_rop_qed_dqed_enq_v),
       .rop_qed_enq_ready                      (i_hqm_qed_pipe_rop_qed_enq_ready),
       .rop_dqed_enq_ready                     (i_hqm_qed_pipe_rop_dqed_enq_ready),
       .rop_qed_dqed_enq_data,
       .rop_qed_force_clockon                  (i_hqm_reorder_pipe_rop_qed_force_clockon),
       .rop_lsp_reordercmp_v                   (i_hqm_reorder_pipe_rop_lsp_reordercmp_v),
       .rop_lsp_reordercmp_ready               (i_hqm_list_sel_pipe_rop_lsp_reordercmp_ready),
       .rop_lsp_reordercmp_data,
       .rf_dir_rply_req_fifo_mem_re            (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_re),
       .rf_dir_rply_req_fifo_mem_rclk          (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rclk),
       .rf_dir_rply_req_fifo_mem_rclk_rst_n    (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rclk_rst_n),
       .rf_dir_rply_req_fifo_mem_raddr         (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_raddr),
       .rf_dir_rply_req_fifo_mem_waddr         (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_waddr),
       .rf_dir_rply_req_fifo_mem_we            (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_we),
       .rf_dir_rply_req_fifo_mem_wclk          (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wclk),
       .rf_dir_rply_req_fifo_mem_wclk_rst_n    (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wclk_rst_n),
       .rf_dir_rply_req_fifo_mem_wdata         (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_wdata),
       .rf_dir_rply_req_fifo_mem_rdata         (i_hqm_reorder_pipe_rf_dir_rply_req_fifo_mem_rdata),
       .rf_ldb_rply_req_fifo_mem_re            (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_re),
       .rf_ldb_rply_req_fifo_mem_rclk          (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rclk),
       .rf_ldb_rply_req_fifo_mem_rclk_rst_n    (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rclk_rst_n),
       .rf_ldb_rply_req_fifo_mem_raddr         (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_raddr),
       .rf_ldb_rply_req_fifo_mem_waddr         (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_waddr),
       .rf_ldb_rply_req_fifo_mem_we            (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_we),
       .rf_ldb_rply_req_fifo_mem_wclk          (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wclk),
       .rf_ldb_rply_req_fifo_mem_wclk_rst_n    (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wclk_rst_n),
       .rf_ldb_rply_req_fifo_mem_wdata         (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_wdata),
       .rf_ldb_rply_req_fifo_mem_rdata         (i_hqm_reorder_pipe_rf_ldb_rply_req_fifo_mem_rdata),
       .rf_lsp_reordercmp_fifo_mem_re          (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_re),
       .rf_lsp_reordercmp_fifo_mem_rclk        (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rclk),
       .rf_lsp_reordercmp_fifo_mem_rclk_rst_n  (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rclk_rst_n),
       .rf_lsp_reordercmp_fifo_mem_raddr       (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_raddr),
       .rf_lsp_reordercmp_fifo_mem_waddr       (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_waddr),
       .rf_lsp_reordercmp_fifo_mem_we          (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_we),
       .rf_lsp_reordercmp_fifo_mem_wclk        (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wclk),
       .rf_lsp_reordercmp_fifo_mem_wclk_rst_n  (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wclk_rst_n),
       .rf_lsp_reordercmp_fifo_mem_wdata       (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_wdata),
       .rf_lsp_reordercmp_fifo_mem_rdata       (i_hqm_reorder_pipe_rf_lsp_reordercmp_fifo_mem_rdata),
       .rf_reord_cnt_mem_re                    (i_hqm_reorder_pipe_rf_reord_cnt_mem_re),
       .rf_reord_cnt_mem_rclk                  (i_hqm_reorder_pipe_rf_reord_cnt_mem_rclk),
       .rf_reord_cnt_mem_rclk_rst_n            (i_hqm_reorder_pipe_rf_reord_cnt_mem_rclk_rst_n),
       .rf_reord_cnt_mem_raddr                 (i_hqm_reorder_pipe_rf_reord_cnt_mem_raddr),
       .rf_reord_cnt_mem_waddr                 (i_hqm_reorder_pipe_rf_reord_cnt_mem_waddr),
       .rf_reord_cnt_mem_we                    (i_hqm_reorder_pipe_rf_reord_cnt_mem_we),
       .rf_reord_cnt_mem_wclk                  (i_hqm_reorder_pipe_rf_reord_cnt_mem_wclk),
       .rf_reord_cnt_mem_wclk_rst_n            (i_hqm_reorder_pipe_rf_reord_cnt_mem_wclk_rst_n),
       .rf_reord_cnt_mem_wdata                 (i_hqm_reorder_pipe_rf_reord_cnt_mem_wdata),
       .rf_reord_cnt_mem_rdata                 (i_hqm_reorder_pipe_rf_reord_cnt_mem_rdata),
       .rf_reord_dirhp_mem_re                  (i_hqm_reorder_pipe_rf_reord_dirhp_mem_re),
       .rf_reord_dirhp_mem_rclk                (i_hqm_reorder_pipe_rf_reord_dirhp_mem_rclk),
       .rf_reord_dirhp_mem_rclk_rst_n          (i_hqm_reorder_pipe_rf_reord_dirhp_mem_rclk_rst_n),
       .rf_reord_dirhp_mem_raddr               (i_hqm_reorder_pipe_rf_reord_dirhp_mem_raddr),
       .rf_reord_dirhp_mem_waddr               (i_hqm_reorder_pipe_rf_reord_dirhp_mem_waddr),
       .rf_reord_dirhp_mem_we                  (i_hqm_reorder_pipe_rf_reord_dirhp_mem_we),
       .rf_reord_dirhp_mem_wclk                (i_hqm_reorder_pipe_rf_reord_dirhp_mem_wclk),
       .rf_reord_dirhp_mem_wclk_rst_n          (i_hqm_reorder_pipe_rf_reord_dirhp_mem_wclk_rst_n),
       .rf_reord_dirhp_mem_wdata               (i_hqm_reorder_pipe_rf_reord_dirhp_mem_wdata),
       .rf_reord_dirhp_mem_rdata               (i_hqm_reorder_pipe_rf_reord_dirhp_mem_rdata),
       .rf_reord_dirtp_mem_re                  (i_hqm_reorder_pipe_rf_reord_dirtp_mem_re),
       .rf_reord_dirtp_mem_rclk                (i_hqm_reorder_pipe_rf_reord_dirtp_mem_rclk),
       .rf_reord_dirtp_mem_rclk_rst_n          (i_hqm_reorder_pipe_rf_reord_dirtp_mem_rclk_rst_n),
       .rf_reord_dirtp_mem_raddr               (i_hqm_reorder_pipe_rf_reord_dirtp_mem_raddr),
       .rf_reord_dirtp_mem_waddr               (i_hqm_reorder_pipe_rf_reord_dirtp_mem_waddr),
       .rf_reord_dirtp_mem_we                  (i_hqm_reorder_pipe_rf_reord_dirtp_mem_we),
       .rf_reord_dirtp_mem_wclk                (i_hqm_reorder_pipe_rf_reord_dirtp_mem_wclk),
       .rf_reord_dirtp_mem_wclk_rst_n          (i_hqm_reorder_pipe_rf_reord_dirtp_mem_wclk_rst_n),
       .rf_reord_dirtp_mem_wdata               (i_hqm_reorder_pipe_rf_reord_dirtp_mem_wdata),
       .rf_reord_dirtp_mem_rdata               (i_hqm_reorder_pipe_rf_reord_dirtp_mem_rdata),
       .rf_reord_lbhp_mem_re                   (i_hqm_reorder_pipe_rf_reord_lbhp_mem_re),
       .rf_reord_lbhp_mem_rclk                 (i_hqm_reorder_pipe_rf_reord_lbhp_mem_rclk),
       .rf_reord_lbhp_mem_rclk_rst_n           (i_hqm_reorder_pipe_rf_reord_lbhp_mem_rclk_rst_n),
       .rf_reord_lbhp_mem_raddr                (i_hqm_reorder_pipe_rf_reord_lbhp_mem_raddr),
       .rf_reord_lbhp_mem_waddr                (i_hqm_reorder_pipe_rf_reord_lbhp_mem_waddr),
       .rf_reord_lbhp_mem_we                   (i_hqm_reorder_pipe_rf_reord_lbhp_mem_we),
       .rf_reord_lbhp_mem_wclk                 (i_hqm_reorder_pipe_rf_reord_lbhp_mem_wclk),
       .rf_reord_lbhp_mem_wclk_rst_n           (i_hqm_reorder_pipe_rf_reord_lbhp_mem_wclk_rst_n),
       .rf_reord_lbhp_mem_wdata                (i_hqm_reorder_pipe_rf_reord_lbhp_mem_wdata),
       .rf_reord_lbhp_mem_rdata                (i_hqm_reorder_pipe_rf_reord_lbhp_mem_rdata),
       .rf_reord_lbtp_mem_re                   (i_hqm_reorder_pipe_rf_reord_lbtp_mem_re),
       .rf_reord_lbtp_mem_rclk                 (i_hqm_reorder_pipe_rf_reord_lbtp_mem_rclk),
       .rf_reord_lbtp_mem_rclk_rst_n           (i_hqm_reorder_pipe_rf_reord_lbtp_mem_rclk_rst_n),
       .rf_reord_lbtp_mem_raddr                (i_hqm_reorder_pipe_rf_reord_lbtp_mem_raddr),
       .rf_reord_lbtp_mem_waddr                (i_hqm_reorder_pipe_rf_reord_lbtp_mem_waddr),
       .rf_reord_lbtp_mem_we                   (i_hqm_reorder_pipe_rf_reord_lbtp_mem_we),
       .rf_reord_lbtp_mem_wclk                 (i_hqm_reorder_pipe_rf_reord_lbtp_mem_wclk),
       .rf_reord_lbtp_mem_wclk_rst_n           (i_hqm_reorder_pipe_rf_reord_lbtp_mem_wclk_rst_n),
       .rf_reord_lbtp_mem_wdata                (i_hqm_reorder_pipe_rf_reord_lbtp_mem_wdata),
       .rf_reord_lbtp_mem_rdata                (i_hqm_reorder_pipe_rf_reord_lbtp_mem_rdata),
       .rf_reord_st_mem_re                     (i_hqm_reorder_pipe_rf_reord_st_mem_re),
       .rf_reord_st_mem_rclk                   (i_hqm_reorder_pipe_rf_reord_st_mem_rclk),
       .rf_reord_st_mem_rclk_rst_n             (i_hqm_reorder_pipe_rf_reord_st_mem_rclk_rst_n),
       .rf_reord_st_mem_raddr                  (i_hqm_reorder_pipe_rf_reord_st_mem_raddr),
       .rf_reord_st_mem_waddr                  (i_hqm_reorder_pipe_rf_reord_st_mem_waddr),
       .rf_reord_st_mem_we                     (i_hqm_reorder_pipe_rf_reord_st_mem_we),
       .rf_reord_st_mem_wclk                   (i_hqm_reorder_pipe_rf_reord_st_mem_wclk),
       .rf_reord_st_mem_wclk_rst_n             (i_hqm_reorder_pipe_rf_reord_st_mem_wclk_rst_n),
       .rf_reord_st_mem_wdata                  (i_hqm_reorder_pipe_rf_reord_st_mem_wdata),
       .rf_reord_st_mem_rdata                  (i_hqm_reorder_pipe_rf_reord_st_mem_rdata),
       .rf_rop_chp_rop_hcw_fifo_mem_re         (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_re),
       .rf_rop_chp_rop_hcw_fifo_mem_rclk       (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rclk),
       .rf_rop_chp_rop_hcw_fifo_mem_rclk_rst_n (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rclk_rst_n),
       .rf_rop_chp_rop_hcw_fifo_mem_raddr      (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_raddr),
       .rf_rop_chp_rop_hcw_fifo_mem_waddr      (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_waddr),
       .rf_rop_chp_rop_hcw_fifo_mem_we         (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_we),
       .rf_rop_chp_rop_hcw_fifo_mem_wclk       (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wclk),
       .rf_rop_chp_rop_hcw_fifo_mem_wclk_rst_n (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wclk_rst_n),
       .rf_rop_chp_rop_hcw_fifo_mem_wdata      (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_wdata),
       .rf_rop_chp_rop_hcw_fifo_mem_rdata      (i_hqm_reorder_pipe_rf_rop_chp_rop_hcw_fifo_mem_rdata),
       .rf_sn0_order_shft_mem_re               (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_re),
       .rf_sn0_order_shft_mem_rclk             (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rclk),
       .rf_sn0_order_shft_mem_rclk_rst_n       (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rclk_rst_n),
       .rf_sn0_order_shft_mem_raddr            (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_raddr),
       .rf_sn0_order_shft_mem_waddr            (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_waddr),
       .rf_sn0_order_shft_mem_we               (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_we),
       .rf_sn0_order_shft_mem_wclk             (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wclk),
       .rf_sn0_order_shft_mem_wclk_rst_n       (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wclk_rst_n),
       .rf_sn0_order_shft_mem_wdata            (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_wdata),
       .rf_sn0_order_shft_mem_rdata            (i_hqm_reorder_pipe_rf_sn0_order_shft_mem_rdata),
       .rf_sn1_order_shft_mem_re               (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_re),
       .rf_sn1_order_shft_mem_rclk             (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rclk),
       .rf_sn1_order_shft_mem_rclk_rst_n       (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rclk_rst_n),
       .rf_sn1_order_shft_mem_raddr            (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_raddr),
       .rf_sn1_order_shft_mem_waddr            (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_waddr),
       .rf_sn1_order_shft_mem_we               (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_we),
       .rf_sn1_order_shft_mem_wclk             (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wclk),
       .rf_sn1_order_shft_mem_wclk_rst_n       (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wclk_rst_n),
       .rf_sn1_order_shft_mem_wdata            (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_wdata),
       .rf_sn1_order_shft_mem_rdata            (i_hqm_reorder_pipe_rf_sn1_order_shft_mem_rdata),
       .rf_sn_complete_fifo_mem_re             (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_re),
       .rf_sn_complete_fifo_mem_rclk           (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rclk),
       .rf_sn_complete_fifo_mem_rclk_rst_n     (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rclk_rst_n),
       .rf_sn_complete_fifo_mem_raddr          (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_raddr),
       .rf_sn_complete_fifo_mem_waddr          (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_waddr),
       .rf_sn_complete_fifo_mem_we             (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_we),
       .rf_sn_complete_fifo_mem_wclk           (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wclk),
       .rf_sn_complete_fifo_mem_wclk_rst_n     (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wclk_rst_n),
       .rf_sn_complete_fifo_mem_wdata          (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_wdata),
       .rf_sn_complete_fifo_mem_rdata          (i_hqm_reorder_pipe_rf_sn_complete_fifo_mem_rdata),
       .rf_sn_ordered_fifo_mem_re              (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_re),
       .rf_sn_ordered_fifo_mem_rclk            (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rclk),
       .rf_sn_ordered_fifo_mem_rclk_rst_n      (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rclk_rst_n),
       .rf_sn_ordered_fifo_mem_raddr           (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_raddr),
       .rf_sn_ordered_fifo_mem_waddr           (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_waddr),
       .rf_sn_ordered_fifo_mem_we              (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_we),
       .rf_sn_ordered_fifo_mem_wclk            (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wclk),
       .rf_sn_ordered_fifo_mem_wclk_rst_n      (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wclk_rst_n),
       .rf_sn_ordered_fifo_mem_wdata           (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_wdata),
       .rf_sn_ordered_fifo_mem_rdata           (i_hqm_reorder_pipe_rf_sn_ordered_fifo_mem_rdata));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_rop_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkxx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_rop),
       .hqm_gated_clk          (hqm_gated_clk_chp),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_rop),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_rop),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_rop),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_rop),
       .hqm_flr_prep           (hqm_flr_prep_rptrxx),
       .rst_prep               (hqm_rst_prep_rop));

   hqm_system i_hqm_system
      (.prim_gated_clk,
       .hqm_inp_gated_clk                  (hqm_inp_gated_clkxx),
       .hqm_inp_gated_rst_b                (hqm_gated_rst_b),
       .hqm_inp_gated_rst_b_sys,
       .hqm_gated_clk                      (hqm_gated_clk_sys),
       .hqm_gated_rst_b_sys,
       .hqm_proc_clk_en_sys                (i_hqm_system_hqm_proc_clk_en_sys),
       .hqm_gated_rst_b_start_sys,
       .hqm_gated_rst_b_active_sys,
       .hqm_gated_rst_b_done_sys,
       .hcw_enq_in_ready,
       .hcw_enq_in_v,
       .hcw_enq_in_data,
       .write_buffer_mstr_ready,
       .write_buffer_mstr_v,
       .write_buffer_mstr,
       .sif_alarm_ready,
       .sif_alarm_v,
       .sif_alarm_data,
       .pci_cfg_sciov_en,
       .pci_cfg_pmsixctl_msie,
       .pci_cfg_pmsixctl_fm,
       .hqm_rst_prep_sys,
       .system_reset_done,
       .system_idle,
       .system_cfg_req_up_write            (mstr_cfg_req_down_write),
       .system_cfg_req_up_read             (mstr_cfg_req_down_read),
       .system_cfg_req_up                  (mstr_cfg_req_down),
       .system_cfg_req_down_write          (i_hqm_system_system_cfg_req_down_write),
       .system_cfg_req_down_read           (i_hqm_system_system_cfg_req_down_read),
       .system_cfg_req_down,
       .system_cfg_rsp_down_ack            (i_hqm_system_system_cfg_rsp_down_ack),
       .system_cfg_rsp_down,
       .hqm_alarm_ready                    (i_hqm_system_hqm_alarm_ready),
       .hqm_alarm_v                        (i_hqm_credit_hist_pipe_chp_alarm_down_v),
       .hqm_alarm_data,
       .hcw_enq_w_req_ready                (i_hqm_credit_hist_pipe_hcw_enq_w_req_ready),
       .hcw_enq_w_req_valid                (i_hqm_system_hcw_enq_w_req_valid),
       .hcw_enq_w_req,
       .hcw_sched_w_req_ready              (i_hqm_system_hcw_sched_w_req_ready),
       .hcw_sched_w_req_valid              (i_hqm_credit_hist_pipe_hcw_sched_w_req_valid),
       .hcw_sched_w_req,
       .interrupt_w_req_ready              (i_hqm_system_interrupt_w_req_ready),
       .interrupt_w_req_valid              (i_hqm_credit_hist_pipe_interrupt_w_req_valid),
       .interrupt_w_req,
       .cwdi_interrupt_w_req_ready         (i_hqm_system_cwdi_interrupt_w_req_ready),
       .cwdi_interrupt_w_req_valid         (i_hqm_credit_hist_pipe_cwdi_interrupt_w_req_valid),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .hqm_system_visa                    (hqm_system_visa_str),
       .spare_lsp_sys,
       .spare_qed_sys,
       .spare_sys_lsp,
       .spare_sys_qed,
       .rf_alarm_vf_synd0_re               (i_hqm_system_rf_alarm_vf_synd0_re),
       .rf_alarm_vf_synd0_rclk             (i_hqm_system_rf_alarm_vf_synd0_rclk),
       .rf_alarm_vf_synd0_rclk_rst_n       (i_hqm_system_rf_alarm_vf_synd0_rclk_rst_n),
       .rf_alarm_vf_synd0_raddr            (i_hqm_system_rf_alarm_vf_synd0_raddr),
       .rf_alarm_vf_synd0_waddr            (i_hqm_system_rf_alarm_vf_synd0_waddr),
       .rf_alarm_vf_synd0_we               (i_hqm_system_rf_alarm_vf_synd0_we),
       .rf_alarm_vf_synd0_wclk             (i_hqm_system_rf_alarm_vf_synd0_wclk),
       .rf_alarm_vf_synd0_wclk_rst_n       (i_hqm_system_rf_alarm_vf_synd0_wclk_rst_n),
       .rf_alarm_vf_synd0_wdata            (i_hqm_system_rf_alarm_vf_synd0_wdata),
       .rf_alarm_vf_synd0_rdata            (i_hqm_system_rf_alarm_vf_synd0_rdata),
       .rf_alarm_vf_synd1_re               (i_hqm_system_rf_alarm_vf_synd1_re),
       .rf_alarm_vf_synd1_rclk             (i_hqm_system_rf_alarm_vf_synd1_rclk),
       .rf_alarm_vf_synd1_rclk_rst_n       (i_hqm_system_rf_alarm_vf_synd1_rclk_rst_n),
       .rf_alarm_vf_synd1_raddr            (i_hqm_system_rf_alarm_vf_synd1_raddr),
       .rf_alarm_vf_synd1_waddr            (i_hqm_system_rf_alarm_vf_synd1_waddr),
       .rf_alarm_vf_synd1_we               (i_hqm_system_rf_alarm_vf_synd1_we),
       .rf_alarm_vf_synd1_wclk             (i_hqm_system_rf_alarm_vf_synd1_wclk),
       .rf_alarm_vf_synd1_wclk_rst_n       (i_hqm_system_rf_alarm_vf_synd1_wclk_rst_n),
       .rf_alarm_vf_synd1_wdata            (i_hqm_system_rf_alarm_vf_synd1_wdata),
       .rf_alarm_vf_synd1_rdata            (i_hqm_system_rf_alarm_vf_synd1_rdata),
       .rf_alarm_vf_synd2_re               (i_hqm_system_rf_alarm_vf_synd2_re),
       .rf_alarm_vf_synd2_rclk             (i_hqm_system_rf_alarm_vf_synd2_rclk),
       .rf_alarm_vf_synd2_rclk_rst_n       (i_hqm_system_rf_alarm_vf_synd2_rclk_rst_n),
       .rf_alarm_vf_synd2_raddr            (i_hqm_system_rf_alarm_vf_synd2_raddr),
       .rf_alarm_vf_synd2_waddr            (i_hqm_system_rf_alarm_vf_synd2_waddr),
       .rf_alarm_vf_synd2_we               (i_hqm_system_rf_alarm_vf_synd2_we),
       .rf_alarm_vf_synd2_wclk             (i_hqm_system_rf_alarm_vf_synd2_wclk),
       .rf_alarm_vf_synd2_wclk_rst_n       (i_hqm_system_rf_alarm_vf_synd2_wclk_rst_n),
       .rf_alarm_vf_synd2_wdata            (i_hqm_system_rf_alarm_vf_synd2_wdata),
       .rf_alarm_vf_synd2_rdata            (i_hqm_system_rf_alarm_vf_synd2_rdata),
       .rf_dir_wb0_re                      (i_hqm_system_rf_dir_wb0_re),
       .rf_dir_wb0_rclk                    (i_hqm_system_rf_dir_wb0_rclk),
       .rf_dir_wb0_rclk_rst_n              (i_hqm_system_rf_dir_wb0_rclk_rst_n),
       .rf_dir_wb0_raddr                   (i_hqm_system_rf_dir_wb0_raddr),
       .rf_dir_wb0_waddr                   (i_hqm_system_rf_dir_wb0_waddr),
       .rf_dir_wb0_we                      (i_hqm_system_rf_dir_wb0_we),
       .rf_dir_wb0_wclk                    (i_hqm_system_rf_dir_wb0_wclk),
       .rf_dir_wb0_wclk_rst_n              (i_hqm_system_rf_dir_wb0_wclk_rst_n),
       .rf_dir_wb0_wdata                   (i_hqm_system_rf_dir_wb0_wdata),
       .rf_dir_wb0_rdata                   (i_hqm_system_rf_dir_wb0_rdata),
       .rf_dir_wb1_re                      (i_hqm_system_rf_dir_wb1_re),
       .rf_dir_wb1_rclk                    (i_hqm_system_rf_dir_wb1_rclk),
       .rf_dir_wb1_rclk_rst_n              (i_hqm_system_rf_dir_wb1_rclk_rst_n),
       .rf_dir_wb1_raddr                   (i_hqm_system_rf_dir_wb1_raddr),
       .rf_dir_wb1_waddr                   (i_hqm_system_rf_dir_wb1_waddr),
       .rf_dir_wb1_we                      (i_hqm_system_rf_dir_wb1_we),
       .rf_dir_wb1_wclk                    (i_hqm_system_rf_dir_wb1_wclk),
       .rf_dir_wb1_wclk_rst_n              (i_hqm_system_rf_dir_wb1_wclk_rst_n),
       .rf_dir_wb1_wdata                   (i_hqm_system_rf_dir_wb1_wdata),
       .rf_dir_wb1_rdata                   (i_hqm_system_rf_dir_wb1_rdata),
       .rf_dir_wb2_re                      (i_hqm_system_rf_dir_wb2_re),
       .rf_dir_wb2_rclk                    (i_hqm_system_rf_dir_wb2_rclk),
       .rf_dir_wb2_rclk_rst_n              (i_hqm_system_rf_dir_wb2_rclk_rst_n),
       .rf_dir_wb2_raddr                   (i_hqm_system_rf_dir_wb2_raddr),
       .rf_dir_wb2_waddr                   (i_hqm_system_rf_dir_wb2_waddr),
       .rf_dir_wb2_we                      (i_hqm_system_rf_dir_wb2_we),
       .rf_dir_wb2_wclk                    (i_hqm_system_rf_dir_wb2_wclk),
       .rf_dir_wb2_wclk_rst_n              (i_hqm_system_rf_dir_wb2_wclk_rst_n),
       .rf_dir_wb2_wdata                   (i_hqm_system_rf_dir_wb2_wdata),
       .rf_dir_wb2_rdata                   (i_hqm_system_rf_dir_wb2_rdata),
       .rf_hcw_enq_fifo_re                 (i_hqm_system_rf_hcw_enq_fifo_re),
       .rf_hcw_enq_fifo_rclk               (i_hqm_system_rf_hcw_enq_fifo_rclk),
       .rf_hcw_enq_fifo_rclk_rst_n         (i_hqm_system_rf_hcw_enq_fifo_rclk_rst_n),
       .rf_hcw_enq_fifo_raddr              (i_hqm_system_rf_hcw_enq_fifo_raddr),
       .rf_hcw_enq_fifo_waddr              (i_hqm_system_rf_hcw_enq_fifo_waddr),
       .rf_hcw_enq_fifo_we                 (i_hqm_system_rf_hcw_enq_fifo_we),
       .rf_hcw_enq_fifo_wclk               (i_hqm_system_rf_hcw_enq_fifo_wclk),
       .rf_hcw_enq_fifo_wclk_rst_n         (i_hqm_system_rf_hcw_enq_fifo_wclk_rst_n),
       .rf_hcw_enq_fifo_wdata              (i_hqm_system_rf_hcw_enq_fifo_wdata),
       .rf_hcw_enq_fifo_rdata              (i_hqm_system_rf_hcw_enq_fifo_rdata),
       .rf_ldb_wb0_re                      (i_hqm_system_rf_ldb_wb0_re),
       .rf_ldb_wb0_rclk                    (i_hqm_system_rf_ldb_wb0_rclk),
       .rf_ldb_wb0_rclk_rst_n              (i_hqm_system_rf_ldb_wb0_rclk_rst_n),
       .rf_ldb_wb0_raddr                   (i_hqm_system_rf_ldb_wb0_raddr),
       .rf_ldb_wb0_waddr                   (i_hqm_system_rf_ldb_wb0_waddr),
       .rf_ldb_wb0_we                      (i_hqm_system_rf_ldb_wb0_we),
       .rf_ldb_wb0_wclk                    (i_hqm_system_rf_ldb_wb0_wclk),
       .rf_ldb_wb0_wclk_rst_n              (i_hqm_system_rf_ldb_wb0_wclk_rst_n),
       .rf_ldb_wb0_wdata                   (i_hqm_system_rf_ldb_wb0_wdata),
       .rf_ldb_wb0_rdata                   (i_hqm_system_rf_ldb_wb0_rdata),
       .rf_ldb_wb1_re                      (i_hqm_system_rf_ldb_wb1_re),
       .rf_ldb_wb1_rclk                    (i_hqm_system_rf_ldb_wb1_rclk),
       .rf_ldb_wb1_rclk_rst_n              (i_hqm_system_rf_ldb_wb1_rclk_rst_n),
       .rf_ldb_wb1_raddr                   (i_hqm_system_rf_ldb_wb1_raddr),
       .rf_ldb_wb1_waddr                   (i_hqm_system_rf_ldb_wb1_waddr),
       .rf_ldb_wb1_we                      (i_hqm_system_rf_ldb_wb1_we),
       .rf_ldb_wb1_wclk                    (i_hqm_system_rf_ldb_wb1_wclk),
       .rf_ldb_wb1_wclk_rst_n              (i_hqm_system_rf_ldb_wb1_wclk_rst_n),
       .rf_ldb_wb1_wdata                   (i_hqm_system_rf_ldb_wb1_wdata),
       .rf_ldb_wb1_rdata                   (i_hqm_system_rf_ldb_wb1_rdata),
       .rf_ldb_wb2_re                      (i_hqm_system_rf_ldb_wb2_re),
       .rf_ldb_wb2_rclk                    (i_hqm_system_rf_ldb_wb2_rclk),
       .rf_ldb_wb2_rclk_rst_n              (i_hqm_system_rf_ldb_wb2_rclk_rst_n),
       .rf_ldb_wb2_raddr                   (i_hqm_system_rf_ldb_wb2_raddr),
       .rf_ldb_wb2_waddr                   (i_hqm_system_rf_ldb_wb2_waddr),
       .rf_ldb_wb2_we                      (i_hqm_system_rf_ldb_wb2_we),
       .rf_ldb_wb2_wclk                    (i_hqm_system_rf_ldb_wb2_wclk),
       .rf_ldb_wb2_wclk_rst_n              (i_hqm_system_rf_ldb_wb2_wclk_rst_n),
       .rf_ldb_wb2_wdata                   (i_hqm_system_rf_ldb_wb2_wdata),
       .rf_ldb_wb2_rdata                   (i_hqm_system_rf_ldb_wb2_rdata),
       .rf_lut_dir_cq2vf_pf_ro_re          (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_re),
       .rf_lut_dir_cq2vf_pf_ro_rclk        (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rclk),
       .rf_lut_dir_cq2vf_pf_ro_rclk_rst_n  (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rclk_rst_n),
       .rf_lut_dir_cq2vf_pf_ro_raddr       (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_raddr),
       .rf_lut_dir_cq2vf_pf_ro_waddr       (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_waddr),
       .rf_lut_dir_cq2vf_pf_ro_we          (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_we),
       .rf_lut_dir_cq2vf_pf_ro_wclk        (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wclk),
       .rf_lut_dir_cq2vf_pf_ro_wclk_rst_n  (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wclk_rst_n),
       .rf_lut_dir_cq2vf_pf_ro_wdata       (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_wdata),
       .rf_lut_dir_cq2vf_pf_ro_rdata       (i_hqm_system_rf_lut_dir_cq2vf_pf_ro_rdata),
       .rf_lut_dir_cq_addr_l_re            (i_hqm_system_rf_lut_dir_cq_addr_l_re),
       .rf_lut_dir_cq_addr_l_rclk          (i_hqm_system_rf_lut_dir_cq_addr_l_rclk),
       .rf_lut_dir_cq_addr_l_rclk_rst_n    (i_hqm_system_rf_lut_dir_cq_addr_l_rclk_rst_n),
       .rf_lut_dir_cq_addr_l_raddr         (i_hqm_system_rf_lut_dir_cq_addr_l_raddr),
       .rf_lut_dir_cq_addr_l_waddr         (i_hqm_system_rf_lut_dir_cq_addr_l_waddr),
       .rf_lut_dir_cq_addr_l_we            (i_hqm_system_rf_lut_dir_cq_addr_l_we),
       .rf_lut_dir_cq_addr_l_wclk          (i_hqm_system_rf_lut_dir_cq_addr_l_wclk),
       .rf_lut_dir_cq_addr_l_wclk_rst_n    (i_hqm_system_rf_lut_dir_cq_addr_l_wclk_rst_n),
       .rf_lut_dir_cq_addr_l_wdata         (i_hqm_system_rf_lut_dir_cq_addr_l_wdata),
       .rf_lut_dir_cq_addr_l_rdata         (i_hqm_system_rf_lut_dir_cq_addr_l_rdata),
       .rf_lut_dir_cq_addr_u_re            (i_hqm_system_rf_lut_dir_cq_addr_u_re),
       .rf_lut_dir_cq_addr_u_rclk          (i_hqm_system_rf_lut_dir_cq_addr_u_rclk),
       .rf_lut_dir_cq_addr_u_rclk_rst_n    (i_hqm_system_rf_lut_dir_cq_addr_u_rclk_rst_n),
       .rf_lut_dir_cq_addr_u_raddr         (i_hqm_system_rf_lut_dir_cq_addr_u_raddr),
       .rf_lut_dir_cq_addr_u_waddr         (i_hqm_system_rf_lut_dir_cq_addr_u_waddr),
       .rf_lut_dir_cq_addr_u_we            (i_hqm_system_rf_lut_dir_cq_addr_u_we),
       .rf_lut_dir_cq_addr_u_wclk          (i_hqm_system_rf_lut_dir_cq_addr_u_wclk),
       .rf_lut_dir_cq_addr_u_wclk_rst_n    (i_hqm_system_rf_lut_dir_cq_addr_u_wclk_rst_n),
       .rf_lut_dir_cq_addr_u_wdata         (i_hqm_system_rf_lut_dir_cq_addr_u_wdata),
       .rf_lut_dir_cq_addr_u_rdata         (i_hqm_system_rf_lut_dir_cq_addr_u_rdata),
       .rf_lut_dir_cq_ai_addr_l_re         (i_hqm_system_rf_lut_dir_cq_ai_addr_l_re),
       .rf_lut_dir_cq_ai_addr_l_rclk       (i_hqm_system_rf_lut_dir_cq_ai_addr_l_rclk),
       .rf_lut_dir_cq_ai_addr_l_rclk_rst_n (i_hqm_system_rf_lut_dir_cq_ai_addr_l_rclk_rst_n),
       .rf_lut_dir_cq_ai_addr_l_raddr      (i_hqm_system_rf_lut_dir_cq_ai_addr_l_raddr),
       .rf_lut_dir_cq_ai_addr_l_waddr      (i_hqm_system_rf_lut_dir_cq_ai_addr_l_waddr),
       .rf_lut_dir_cq_ai_addr_l_we         (i_hqm_system_rf_lut_dir_cq_ai_addr_l_we),
       .rf_lut_dir_cq_ai_addr_l_wclk       (i_hqm_system_rf_lut_dir_cq_ai_addr_l_wclk),
       .rf_lut_dir_cq_ai_addr_l_wclk_rst_n (i_hqm_system_rf_lut_dir_cq_ai_addr_l_wclk_rst_n),
       .rf_lut_dir_cq_ai_addr_l_wdata      (i_hqm_system_rf_lut_dir_cq_ai_addr_l_wdata),
       .rf_lut_dir_cq_ai_addr_l_rdata      (i_hqm_system_rf_lut_dir_cq_ai_addr_l_rdata),
       .rf_lut_dir_cq_ai_addr_u_re         (i_hqm_system_rf_lut_dir_cq_ai_addr_u_re),
       .rf_lut_dir_cq_ai_addr_u_rclk       (i_hqm_system_rf_lut_dir_cq_ai_addr_u_rclk),
       .rf_lut_dir_cq_ai_addr_u_rclk_rst_n (i_hqm_system_rf_lut_dir_cq_ai_addr_u_rclk_rst_n),
       .rf_lut_dir_cq_ai_addr_u_raddr      (i_hqm_system_rf_lut_dir_cq_ai_addr_u_raddr),
       .rf_lut_dir_cq_ai_addr_u_waddr      (i_hqm_system_rf_lut_dir_cq_ai_addr_u_waddr),
       .rf_lut_dir_cq_ai_addr_u_we         (i_hqm_system_rf_lut_dir_cq_ai_addr_u_we),
       .rf_lut_dir_cq_ai_addr_u_wclk       (i_hqm_system_rf_lut_dir_cq_ai_addr_u_wclk),
       .rf_lut_dir_cq_ai_addr_u_wclk_rst_n (i_hqm_system_rf_lut_dir_cq_ai_addr_u_wclk_rst_n),
       .rf_lut_dir_cq_ai_addr_u_wdata      (i_hqm_system_rf_lut_dir_cq_ai_addr_u_wdata),
       .rf_lut_dir_cq_ai_addr_u_rdata      (i_hqm_system_rf_lut_dir_cq_ai_addr_u_rdata),
       .rf_lut_dir_cq_ai_data_re           (i_hqm_system_rf_lut_dir_cq_ai_data_re),
       .rf_lut_dir_cq_ai_data_rclk         (i_hqm_system_rf_lut_dir_cq_ai_data_rclk),
       .rf_lut_dir_cq_ai_data_rclk_rst_n   (i_hqm_system_rf_lut_dir_cq_ai_data_rclk_rst_n),
       .rf_lut_dir_cq_ai_data_raddr        (i_hqm_system_rf_lut_dir_cq_ai_data_raddr),
       .rf_lut_dir_cq_ai_data_waddr        (i_hqm_system_rf_lut_dir_cq_ai_data_waddr),
       .rf_lut_dir_cq_ai_data_we           (i_hqm_system_rf_lut_dir_cq_ai_data_we),
       .rf_lut_dir_cq_ai_data_wclk         (i_hqm_system_rf_lut_dir_cq_ai_data_wclk),
       .rf_lut_dir_cq_ai_data_wclk_rst_n   (i_hqm_system_rf_lut_dir_cq_ai_data_wclk_rst_n),
       .rf_lut_dir_cq_ai_data_wdata        (i_hqm_system_rf_lut_dir_cq_ai_data_wdata),
       .rf_lut_dir_cq_ai_data_rdata        (i_hqm_system_rf_lut_dir_cq_ai_data_rdata),
       .rf_lut_dir_cq_isr_re               (i_hqm_system_rf_lut_dir_cq_isr_re),
       .rf_lut_dir_cq_isr_rclk             (i_hqm_system_rf_lut_dir_cq_isr_rclk),
       .rf_lut_dir_cq_isr_rclk_rst_n       (i_hqm_system_rf_lut_dir_cq_isr_rclk_rst_n),
       .rf_lut_dir_cq_isr_raddr            (i_hqm_system_rf_lut_dir_cq_isr_raddr),
       .rf_lut_dir_cq_isr_waddr            (i_hqm_system_rf_lut_dir_cq_isr_waddr),
       .rf_lut_dir_cq_isr_we               (i_hqm_system_rf_lut_dir_cq_isr_we),
       .rf_lut_dir_cq_isr_wclk             (i_hqm_system_rf_lut_dir_cq_isr_wclk),
       .rf_lut_dir_cq_isr_wclk_rst_n       (i_hqm_system_rf_lut_dir_cq_isr_wclk_rst_n),
       .rf_lut_dir_cq_isr_wdata            (i_hqm_system_rf_lut_dir_cq_isr_wdata),
       .rf_lut_dir_cq_isr_rdata            (i_hqm_system_rf_lut_dir_cq_isr_rdata),
       .rf_lut_dir_cq_pasid_re             (i_hqm_system_rf_lut_dir_cq_pasid_re),
       .rf_lut_dir_cq_pasid_rclk           (i_hqm_system_rf_lut_dir_cq_pasid_rclk),
       .rf_lut_dir_cq_pasid_rclk_rst_n     (i_hqm_system_rf_lut_dir_cq_pasid_rclk_rst_n),
       .rf_lut_dir_cq_pasid_raddr          (i_hqm_system_rf_lut_dir_cq_pasid_raddr),
       .rf_lut_dir_cq_pasid_waddr          (i_hqm_system_rf_lut_dir_cq_pasid_waddr),
       .rf_lut_dir_cq_pasid_we             (i_hqm_system_rf_lut_dir_cq_pasid_we),
       .rf_lut_dir_cq_pasid_wclk           (i_hqm_system_rf_lut_dir_cq_pasid_wclk),
       .rf_lut_dir_cq_pasid_wclk_rst_n     (i_hqm_system_rf_lut_dir_cq_pasid_wclk_rst_n),
       .rf_lut_dir_cq_pasid_wdata          (i_hqm_system_rf_lut_dir_cq_pasid_wdata),
       .rf_lut_dir_cq_pasid_rdata          (i_hqm_system_rf_lut_dir_cq_pasid_rdata),
       .rf_lut_dir_pp2vas_re               (i_hqm_system_rf_lut_dir_pp2vas_re),
       .rf_lut_dir_pp2vas_rclk             (i_hqm_system_rf_lut_dir_pp2vas_rclk),
       .rf_lut_dir_pp2vas_rclk_rst_n       (i_hqm_system_rf_lut_dir_pp2vas_rclk_rst_n),
       .rf_lut_dir_pp2vas_raddr            (i_hqm_system_rf_lut_dir_pp2vas_raddr),
       .rf_lut_dir_pp2vas_waddr            (i_hqm_system_rf_lut_dir_pp2vas_waddr),
       .rf_lut_dir_pp2vas_we               (i_hqm_system_rf_lut_dir_pp2vas_we),
       .rf_lut_dir_pp2vas_wclk             (i_hqm_system_rf_lut_dir_pp2vas_wclk),
       .rf_lut_dir_pp2vas_wclk_rst_n       (i_hqm_system_rf_lut_dir_pp2vas_wclk_rst_n),
       .rf_lut_dir_pp2vas_wdata            (i_hqm_system_rf_lut_dir_pp2vas_wdata),
       .rf_lut_dir_pp2vas_rdata            (i_hqm_system_rf_lut_dir_pp2vas_rdata),
       .rf_lut_dir_pp_v_re                 (i_hqm_system_rf_lut_dir_pp_v_re),
       .rf_lut_dir_pp_v_rclk               (i_hqm_system_rf_lut_dir_pp_v_rclk),
       .rf_lut_dir_pp_v_rclk_rst_n         (i_hqm_system_rf_lut_dir_pp_v_rclk_rst_n),
       .rf_lut_dir_pp_v_raddr              (i_hqm_system_rf_lut_dir_pp_v_raddr),
       .rf_lut_dir_pp_v_waddr              (i_hqm_system_rf_lut_dir_pp_v_waddr),
       .rf_lut_dir_pp_v_we                 (i_hqm_system_rf_lut_dir_pp_v_we),
       .rf_lut_dir_pp_v_wclk               (i_hqm_system_rf_lut_dir_pp_v_wclk),
       .rf_lut_dir_pp_v_wclk_rst_n         (i_hqm_system_rf_lut_dir_pp_v_wclk_rst_n),
       .rf_lut_dir_pp_v_wdata              (i_hqm_system_rf_lut_dir_pp_v_wdata),
       .rf_lut_dir_pp_v_rdata              (i_hqm_system_rf_lut_dir_pp_v_rdata),
       .rf_lut_dir_vasqid_v_re             (i_hqm_system_rf_lut_dir_vasqid_v_re),
       .rf_lut_dir_vasqid_v_rclk           (i_hqm_system_rf_lut_dir_vasqid_v_rclk),
       .rf_lut_dir_vasqid_v_rclk_rst_n     (i_hqm_system_rf_lut_dir_vasqid_v_rclk_rst_n),
       .rf_lut_dir_vasqid_v_raddr          (i_hqm_system_rf_lut_dir_vasqid_v_raddr),
       .rf_lut_dir_vasqid_v_waddr          (i_hqm_system_rf_lut_dir_vasqid_v_waddr),
       .rf_lut_dir_vasqid_v_we             (i_hqm_system_rf_lut_dir_vasqid_v_we),
       .rf_lut_dir_vasqid_v_wclk           (i_hqm_system_rf_lut_dir_vasqid_v_wclk),
       .rf_lut_dir_vasqid_v_wclk_rst_n     (i_hqm_system_rf_lut_dir_vasqid_v_wclk_rst_n),
       .rf_lut_dir_vasqid_v_wdata          (i_hqm_system_rf_lut_dir_vasqid_v_wdata),
       .rf_lut_dir_vasqid_v_rdata          (i_hqm_system_rf_lut_dir_vasqid_v_rdata),
       .rf_lut_ldb_cq2vf_pf_ro_re          (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_re),
       .rf_lut_ldb_cq2vf_pf_ro_rclk        (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rclk),
       .rf_lut_ldb_cq2vf_pf_ro_rclk_rst_n  (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rclk_rst_n),
       .rf_lut_ldb_cq2vf_pf_ro_raddr       (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_raddr),
       .rf_lut_ldb_cq2vf_pf_ro_waddr       (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_waddr),
       .rf_lut_ldb_cq2vf_pf_ro_we          (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_we),
       .rf_lut_ldb_cq2vf_pf_ro_wclk        (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wclk),
       .rf_lut_ldb_cq2vf_pf_ro_wclk_rst_n  (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wclk_rst_n),
       .rf_lut_ldb_cq2vf_pf_ro_wdata       (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_wdata),
       .rf_lut_ldb_cq2vf_pf_ro_rdata       (i_hqm_system_rf_lut_ldb_cq2vf_pf_ro_rdata),
       .rf_lut_ldb_cq_addr_l_re            (i_hqm_system_rf_lut_ldb_cq_addr_l_re),
       .rf_lut_ldb_cq_addr_l_rclk          (i_hqm_system_rf_lut_ldb_cq_addr_l_rclk),
       .rf_lut_ldb_cq_addr_l_rclk_rst_n    (i_hqm_system_rf_lut_ldb_cq_addr_l_rclk_rst_n),
       .rf_lut_ldb_cq_addr_l_raddr         (i_hqm_system_rf_lut_ldb_cq_addr_l_raddr),
       .rf_lut_ldb_cq_addr_l_waddr         (i_hqm_system_rf_lut_ldb_cq_addr_l_waddr),
       .rf_lut_ldb_cq_addr_l_we            (i_hqm_system_rf_lut_ldb_cq_addr_l_we),
       .rf_lut_ldb_cq_addr_l_wclk          (i_hqm_system_rf_lut_ldb_cq_addr_l_wclk),
       .rf_lut_ldb_cq_addr_l_wclk_rst_n    (i_hqm_system_rf_lut_ldb_cq_addr_l_wclk_rst_n),
       .rf_lut_ldb_cq_addr_l_wdata         (i_hqm_system_rf_lut_ldb_cq_addr_l_wdata),
       .rf_lut_ldb_cq_addr_l_rdata         (i_hqm_system_rf_lut_ldb_cq_addr_l_rdata),
       .rf_lut_ldb_cq_addr_u_re            (i_hqm_system_rf_lut_ldb_cq_addr_u_re),
       .rf_lut_ldb_cq_addr_u_rclk          (i_hqm_system_rf_lut_ldb_cq_addr_u_rclk),
       .rf_lut_ldb_cq_addr_u_rclk_rst_n    (i_hqm_system_rf_lut_ldb_cq_addr_u_rclk_rst_n),
       .rf_lut_ldb_cq_addr_u_raddr         (i_hqm_system_rf_lut_ldb_cq_addr_u_raddr),
       .rf_lut_ldb_cq_addr_u_waddr         (i_hqm_system_rf_lut_ldb_cq_addr_u_waddr),
       .rf_lut_ldb_cq_addr_u_we            (i_hqm_system_rf_lut_ldb_cq_addr_u_we),
       .rf_lut_ldb_cq_addr_u_wclk          (i_hqm_system_rf_lut_ldb_cq_addr_u_wclk),
       .rf_lut_ldb_cq_addr_u_wclk_rst_n    (i_hqm_system_rf_lut_ldb_cq_addr_u_wclk_rst_n),
       .rf_lut_ldb_cq_addr_u_wdata         (i_hqm_system_rf_lut_ldb_cq_addr_u_wdata),
       .rf_lut_ldb_cq_addr_u_rdata         (i_hqm_system_rf_lut_ldb_cq_addr_u_rdata),
       .rf_lut_ldb_cq_ai_addr_l_re         (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_re),
       .rf_lut_ldb_cq_ai_addr_l_rclk       (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rclk),
       .rf_lut_ldb_cq_ai_addr_l_rclk_rst_n (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rclk_rst_n),
       .rf_lut_ldb_cq_ai_addr_l_raddr      (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_raddr),
       .rf_lut_ldb_cq_ai_addr_l_waddr      (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_waddr),
       .rf_lut_ldb_cq_ai_addr_l_we         (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_we),
       .rf_lut_ldb_cq_ai_addr_l_wclk       (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wclk),
       .rf_lut_ldb_cq_ai_addr_l_wclk_rst_n (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wclk_rst_n),
       .rf_lut_ldb_cq_ai_addr_l_wdata      (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_wdata),
       .rf_lut_ldb_cq_ai_addr_l_rdata      (i_hqm_system_rf_lut_ldb_cq_ai_addr_l_rdata),
       .rf_lut_ldb_cq_ai_addr_u_re         (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_re),
       .rf_lut_ldb_cq_ai_addr_u_rclk       (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rclk),
       .rf_lut_ldb_cq_ai_addr_u_rclk_rst_n (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rclk_rst_n),
       .rf_lut_ldb_cq_ai_addr_u_raddr      (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_raddr),
       .rf_lut_ldb_cq_ai_addr_u_waddr      (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_waddr),
       .rf_lut_ldb_cq_ai_addr_u_we         (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_we),
       .rf_lut_ldb_cq_ai_addr_u_wclk       (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wclk),
       .rf_lut_ldb_cq_ai_addr_u_wclk_rst_n (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wclk_rst_n),
       .rf_lut_ldb_cq_ai_addr_u_wdata      (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_wdata),
       .rf_lut_ldb_cq_ai_addr_u_rdata      (i_hqm_system_rf_lut_ldb_cq_ai_addr_u_rdata),
       .rf_lut_ldb_cq_ai_data_re           (i_hqm_system_rf_lut_ldb_cq_ai_data_re),
       .rf_lut_ldb_cq_ai_data_rclk         (i_hqm_system_rf_lut_ldb_cq_ai_data_rclk),
       .rf_lut_ldb_cq_ai_data_rclk_rst_n   (i_hqm_system_rf_lut_ldb_cq_ai_data_rclk_rst_n),
       .rf_lut_ldb_cq_ai_data_raddr        (i_hqm_system_rf_lut_ldb_cq_ai_data_raddr),
       .rf_lut_ldb_cq_ai_data_waddr        (i_hqm_system_rf_lut_ldb_cq_ai_data_waddr),
       .rf_lut_ldb_cq_ai_data_we           (i_hqm_system_rf_lut_ldb_cq_ai_data_we),
       .rf_lut_ldb_cq_ai_data_wclk         (i_hqm_system_rf_lut_ldb_cq_ai_data_wclk),
       .rf_lut_ldb_cq_ai_data_wclk_rst_n   (i_hqm_system_rf_lut_ldb_cq_ai_data_wclk_rst_n),
       .rf_lut_ldb_cq_ai_data_wdata        (i_hqm_system_rf_lut_ldb_cq_ai_data_wdata),
       .rf_lut_ldb_cq_ai_data_rdata        (i_hqm_system_rf_lut_ldb_cq_ai_data_rdata),
       .rf_lut_ldb_cq_isr_re               (i_hqm_system_rf_lut_ldb_cq_isr_re),
       .rf_lut_ldb_cq_isr_rclk             (i_hqm_system_rf_lut_ldb_cq_isr_rclk),
       .rf_lut_ldb_cq_isr_rclk_rst_n       (i_hqm_system_rf_lut_ldb_cq_isr_rclk_rst_n),
       .rf_lut_ldb_cq_isr_raddr            (i_hqm_system_rf_lut_ldb_cq_isr_raddr),
       .rf_lut_ldb_cq_isr_waddr            (i_hqm_system_rf_lut_ldb_cq_isr_waddr),
       .rf_lut_ldb_cq_isr_we               (i_hqm_system_rf_lut_ldb_cq_isr_we),
       .rf_lut_ldb_cq_isr_wclk             (i_hqm_system_rf_lut_ldb_cq_isr_wclk),
       .rf_lut_ldb_cq_isr_wclk_rst_n       (i_hqm_system_rf_lut_ldb_cq_isr_wclk_rst_n),
       .rf_lut_ldb_cq_isr_wdata            (i_hqm_system_rf_lut_ldb_cq_isr_wdata),
       .rf_lut_ldb_cq_isr_rdata            (i_hqm_system_rf_lut_ldb_cq_isr_rdata),
       .rf_lut_ldb_cq_pasid_re             (i_hqm_system_rf_lut_ldb_cq_pasid_re),
       .rf_lut_ldb_cq_pasid_rclk           (i_hqm_system_rf_lut_ldb_cq_pasid_rclk),
       .rf_lut_ldb_cq_pasid_rclk_rst_n     (i_hqm_system_rf_lut_ldb_cq_pasid_rclk_rst_n),
       .rf_lut_ldb_cq_pasid_raddr          (i_hqm_system_rf_lut_ldb_cq_pasid_raddr),
       .rf_lut_ldb_cq_pasid_waddr          (i_hqm_system_rf_lut_ldb_cq_pasid_waddr),
       .rf_lut_ldb_cq_pasid_we             (i_hqm_system_rf_lut_ldb_cq_pasid_we),
       .rf_lut_ldb_cq_pasid_wclk           (i_hqm_system_rf_lut_ldb_cq_pasid_wclk),
       .rf_lut_ldb_cq_pasid_wclk_rst_n     (i_hqm_system_rf_lut_ldb_cq_pasid_wclk_rst_n),
       .rf_lut_ldb_cq_pasid_wdata          (i_hqm_system_rf_lut_ldb_cq_pasid_wdata),
       .rf_lut_ldb_cq_pasid_rdata          (i_hqm_system_rf_lut_ldb_cq_pasid_rdata),
       .rf_lut_ldb_pp2vas_re               (i_hqm_system_rf_lut_ldb_pp2vas_re),
       .rf_lut_ldb_pp2vas_rclk             (i_hqm_system_rf_lut_ldb_pp2vas_rclk),
       .rf_lut_ldb_pp2vas_rclk_rst_n       (i_hqm_system_rf_lut_ldb_pp2vas_rclk_rst_n),
       .rf_lut_ldb_pp2vas_raddr            (i_hqm_system_rf_lut_ldb_pp2vas_raddr),
       .rf_lut_ldb_pp2vas_waddr            (i_hqm_system_rf_lut_ldb_pp2vas_waddr),
       .rf_lut_ldb_pp2vas_we               (i_hqm_system_rf_lut_ldb_pp2vas_we),
       .rf_lut_ldb_pp2vas_wclk             (i_hqm_system_rf_lut_ldb_pp2vas_wclk),
       .rf_lut_ldb_pp2vas_wclk_rst_n       (i_hqm_system_rf_lut_ldb_pp2vas_wclk_rst_n),
       .rf_lut_ldb_pp2vas_wdata            (i_hqm_system_rf_lut_ldb_pp2vas_wdata),
       .rf_lut_ldb_pp2vas_rdata            (i_hqm_system_rf_lut_ldb_pp2vas_rdata),
       .rf_lut_ldb_qid2vqid_re             (i_hqm_system_rf_lut_ldb_qid2vqid_re),
       .rf_lut_ldb_qid2vqid_rclk           (i_hqm_system_rf_lut_ldb_qid2vqid_rclk),
       .rf_lut_ldb_qid2vqid_rclk_rst_n     (i_hqm_system_rf_lut_ldb_qid2vqid_rclk_rst_n),
       .rf_lut_ldb_qid2vqid_raddr          (i_hqm_system_rf_lut_ldb_qid2vqid_raddr),
       .rf_lut_ldb_qid2vqid_waddr          (i_hqm_system_rf_lut_ldb_qid2vqid_waddr),
       .rf_lut_ldb_qid2vqid_we             (i_hqm_system_rf_lut_ldb_qid2vqid_we),
       .rf_lut_ldb_qid2vqid_wclk           (i_hqm_system_rf_lut_ldb_qid2vqid_wclk),
       .rf_lut_ldb_qid2vqid_wclk_rst_n     (i_hqm_system_rf_lut_ldb_qid2vqid_wclk_rst_n),
       .rf_lut_ldb_qid2vqid_wdata          (i_hqm_system_rf_lut_ldb_qid2vqid_wdata),
       .rf_lut_ldb_qid2vqid_rdata          (i_hqm_system_rf_lut_ldb_qid2vqid_rdata),
       .rf_lut_ldb_vasqid_v_re             (i_hqm_system_rf_lut_ldb_vasqid_v_re),
       .rf_lut_ldb_vasqid_v_rclk           (i_hqm_system_rf_lut_ldb_vasqid_v_rclk),
       .rf_lut_ldb_vasqid_v_rclk_rst_n     (i_hqm_system_rf_lut_ldb_vasqid_v_rclk_rst_n),
       .rf_lut_ldb_vasqid_v_raddr          (i_hqm_system_rf_lut_ldb_vasqid_v_raddr),
       .rf_lut_ldb_vasqid_v_waddr          (i_hqm_system_rf_lut_ldb_vasqid_v_waddr),
       .rf_lut_ldb_vasqid_v_we             (i_hqm_system_rf_lut_ldb_vasqid_v_we),
       .rf_lut_ldb_vasqid_v_wclk           (i_hqm_system_rf_lut_ldb_vasqid_v_wclk),
       .rf_lut_ldb_vasqid_v_wclk_rst_n     (i_hqm_system_rf_lut_ldb_vasqid_v_wclk_rst_n),
       .rf_lut_ldb_vasqid_v_wdata          (i_hqm_system_rf_lut_ldb_vasqid_v_wdata),
       .rf_lut_ldb_vasqid_v_rdata          (i_hqm_system_rf_lut_ldb_vasqid_v_rdata),
       .rf_lut_vf_dir_vpp2pp_re            (i_hqm_system_rf_lut_vf_dir_vpp2pp_re),
       .rf_lut_vf_dir_vpp2pp_rclk          (i_hqm_system_rf_lut_vf_dir_vpp2pp_rclk),
       .rf_lut_vf_dir_vpp2pp_rclk_rst_n    (i_hqm_system_rf_lut_vf_dir_vpp2pp_rclk_rst_n),
       .rf_lut_vf_dir_vpp2pp_raddr         (i_hqm_system_rf_lut_vf_dir_vpp2pp_raddr),
       .rf_lut_vf_dir_vpp2pp_waddr         (i_hqm_system_rf_lut_vf_dir_vpp2pp_waddr),
       .rf_lut_vf_dir_vpp2pp_we            (i_hqm_system_rf_lut_vf_dir_vpp2pp_we),
       .rf_lut_vf_dir_vpp2pp_wclk          (i_hqm_system_rf_lut_vf_dir_vpp2pp_wclk),
       .rf_lut_vf_dir_vpp2pp_wclk_rst_n    (i_hqm_system_rf_lut_vf_dir_vpp2pp_wclk_rst_n),
       .rf_lut_vf_dir_vpp2pp_wdata         (i_hqm_system_rf_lut_vf_dir_vpp2pp_wdata),
       .rf_lut_vf_dir_vpp2pp_rdata         (i_hqm_system_rf_lut_vf_dir_vpp2pp_rdata),
       .rf_lut_vf_dir_vpp_v_re             (i_hqm_system_rf_lut_vf_dir_vpp_v_re),
       .rf_lut_vf_dir_vpp_v_rclk           (i_hqm_system_rf_lut_vf_dir_vpp_v_rclk),
       .rf_lut_vf_dir_vpp_v_rclk_rst_n     (i_hqm_system_rf_lut_vf_dir_vpp_v_rclk_rst_n),
       .rf_lut_vf_dir_vpp_v_raddr          (i_hqm_system_rf_lut_vf_dir_vpp_v_raddr),
       .rf_lut_vf_dir_vpp_v_waddr          (i_hqm_system_rf_lut_vf_dir_vpp_v_waddr),
       .rf_lut_vf_dir_vpp_v_we             (i_hqm_system_rf_lut_vf_dir_vpp_v_we),
       .rf_lut_vf_dir_vpp_v_wclk           (i_hqm_system_rf_lut_vf_dir_vpp_v_wclk),
       .rf_lut_vf_dir_vpp_v_wclk_rst_n     (i_hqm_system_rf_lut_vf_dir_vpp_v_wclk_rst_n),
       .rf_lut_vf_dir_vpp_v_wdata          (i_hqm_system_rf_lut_vf_dir_vpp_v_wdata),
       .rf_lut_vf_dir_vpp_v_rdata          (i_hqm_system_rf_lut_vf_dir_vpp_v_rdata),
       .rf_lut_vf_dir_vqid2qid_re          (i_hqm_system_rf_lut_vf_dir_vqid2qid_re),
       .rf_lut_vf_dir_vqid2qid_rclk        (i_hqm_system_rf_lut_vf_dir_vqid2qid_rclk),
       .rf_lut_vf_dir_vqid2qid_rclk_rst_n  (i_hqm_system_rf_lut_vf_dir_vqid2qid_rclk_rst_n),
       .rf_lut_vf_dir_vqid2qid_raddr       (i_hqm_system_rf_lut_vf_dir_vqid2qid_raddr),
       .rf_lut_vf_dir_vqid2qid_waddr       (i_hqm_system_rf_lut_vf_dir_vqid2qid_waddr),
       .rf_lut_vf_dir_vqid2qid_we          (i_hqm_system_rf_lut_vf_dir_vqid2qid_we),
       .rf_lut_vf_dir_vqid2qid_wclk        (i_hqm_system_rf_lut_vf_dir_vqid2qid_wclk),
       .rf_lut_vf_dir_vqid2qid_wclk_rst_n  (i_hqm_system_rf_lut_vf_dir_vqid2qid_wclk_rst_n),
       .rf_lut_vf_dir_vqid2qid_wdata       (i_hqm_system_rf_lut_vf_dir_vqid2qid_wdata),
       .rf_lut_vf_dir_vqid2qid_rdata       (i_hqm_system_rf_lut_vf_dir_vqid2qid_rdata),
       .rf_lut_vf_dir_vqid_v_re            (i_hqm_system_rf_lut_vf_dir_vqid_v_re),
       .rf_lut_vf_dir_vqid_v_rclk          (i_hqm_system_rf_lut_vf_dir_vqid_v_rclk),
       .rf_lut_vf_dir_vqid_v_rclk_rst_n    (i_hqm_system_rf_lut_vf_dir_vqid_v_rclk_rst_n),
       .rf_lut_vf_dir_vqid_v_raddr         (i_hqm_system_rf_lut_vf_dir_vqid_v_raddr),
       .rf_lut_vf_dir_vqid_v_waddr         (i_hqm_system_rf_lut_vf_dir_vqid_v_waddr),
       .rf_lut_vf_dir_vqid_v_we            (i_hqm_system_rf_lut_vf_dir_vqid_v_we),
       .rf_lut_vf_dir_vqid_v_wclk          (i_hqm_system_rf_lut_vf_dir_vqid_v_wclk),
       .rf_lut_vf_dir_vqid_v_wclk_rst_n    (i_hqm_system_rf_lut_vf_dir_vqid_v_wclk_rst_n),
       .rf_lut_vf_dir_vqid_v_wdata         (i_hqm_system_rf_lut_vf_dir_vqid_v_wdata),
       .rf_lut_vf_dir_vqid_v_rdata         (i_hqm_system_rf_lut_vf_dir_vqid_v_rdata),
       .rf_lut_vf_ldb_vpp2pp_re            (i_hqm_system_rf_lut_vf_ldb_vpp2pp_re),
       .rf_lut_vf_ldb_vpp2pp_rclk          (i_hqm_system_rf_lut_vf_ldb_vpp2pp_rclk),
       .rf_lut_vf_ldb_vpp2pp_rclk_rst_n    (i_hqm_system_rf_lut_vf_ldb_vpp2pp_rclk_rst_n),
       .rf_lut_vf_ldb_vpp2pp_raddr         (i_hqm_system_rf_lut_vf_ldb_vpp2pp_raddr),
       .rf_lut_vf_ldb_vpp2pp_waddr         (i_hqm_system_rf_lut_vf_ldb_vpp2pp_waddr),
       .rf_lut_vf_ldb_vpp2pp_we            (i_hqm_system_rf_lut_vf_ldb_vpp2pp_we),
       .rf_lut_vf_ldb_vpp2pp_wclk          (i_hqm_system_rf_lut_vf_ldb_vpp2pp_wclk),
       .rf_lut_vf_ldb_vpp2pp_wclk_rst_n    (i_hqm_system_rf_lut_vf_ldb_vpp2pp_wclk_rst_n),
       .rf_lut_vf_ldb_vpp2pp_wdata         (i_hqm_system_rf_lut_vf_ldb_vpp2pp_wdata),
       .rf_lut_vf_ldb_vpp2pp_rdata         (i_hqm_system_rf_lut_vf_ldb_vpp2pp_rdata),
       .rf_lut_vf_ldb_vpp_v_re             (i_hqm_system_rf_lut_vf_ldb_vpp_v_re),
       .rf_lut_vf_ldb_vpp_v_rclk           (i_hqm_system_rf_lut_vf_ldb_vpp_v_rclk),
       .rf_lut_vf_ldb_vpp_v_rclk_rst_n     (i_hqm_system_rf_lut_vf_ldb_vpp_v_rclk_rst_n),
       .rf_lut_vf_ldb_vpp_v_raddr          (i_hqm_system_rf_lut_vf_ldb_vpp_v_raddr),
       .rf_lut_vf_ldb_vpp_v_waddr          (i_hqm_system_rf_lut_vf_ldb_vpp_v_waddr),
       .rf_lut_vf_ldb_vpp_v_we             (i_hqm_system_rf_lut_vf_ldb_vpp_v_we),
       .rf_lut_vf_ldb_vpp_v_wclk           (i_hqm_system_rf_lut_vf_ldb_vpp_v_wclk),
       .rf_lut_vf_ldb_vpp_v_wclk_rst_n     (i_hqm_system_rf_lut_vf_ldb_vpp_v_wclk_rst_n),
       .rf_lut_vf_ldb_vpp_v_wdata          (i_hqm_system_rf_lut_vf_ldb_vpp_v_wdata),
       .rf_lut_vf_ldb_vpp_v_rdata          (i_hqm_system_rf_lut_vf_ldb_vpp_v_rdata),
       .rf_lut_vf_ldb_vqid2qid_re          (i_hqm_system_rf_lut_vf_ldb_vqid2qid_re),
       .rf_lut_vf_ldb_vqid2qid_rclk        (i_hqm_system_rf_lut_vf_ldb_vqid2qid_rclk),
       .rf_lut_vf_ldb_vqid2qid_rclk_rst_n  (i_hqm_system_rf_lut_vf_ldb_vqid2qid_rclk_rst_n),
       .rf_lut_vf_ldb_vqid2qid_raddr       (i_hqm_system_rf_lut_vf_ldb_vqid2qid_raddr),
       .rf_lut_vf_ldb_vqid2qid_waddr       (i_hqm_system_rf_lut_vf_ldb_vqid2qid_waddr),
       .rf_lut_vf_ldb_vqid2qid_we          (i_hqm_system_rf_lut_vf_ldb_vqid2qid_we),
       .rf_lut_vf_ldb_vqid2qid_wclk        (i_hqm_system_rf_lut_vf_ldb_vqid2qid_wclk),
       .rf_lut_vf_ldb_vqid2qid_wclk_rst_n  (i_hqm_system_rf_lut_vf_ldb_vqid2qid_wclk_rst_n),
       .rf_lut_vf_ldb_vqid2qid_wdata       (i_hqm_system_rf_lut_vf_ldb_vqid2qid_wdata),
       .rf_lut_vf_ldb_vqid2qid_rdata       (i_hqm_system_rf_lut_vf_ldb_vqid2qid_rdata),
       .rf_lut_vf_ldb_vqid_v_re            (i_hqm_system_rf_lut_vf_ldb_vqid_v_re),
       .rf_lut_vf_ldb_vqid_v_rclk          (i_hqm_system_rf_lut_vf_ldb_vqid_v_rclk),
       .rf_lut_vf_ldb_vqid_v_rclk_rst_n    (i_hqm_system_rf_lut_vf_ldb_vqid_v_rclk_rst_n),
       .rf_lut_vf_ldb_vqid_v_raddr         (i_hqm_system_rf_lut_vf_ldb_vqid_v_raddr),
       .rf_lut_vf_ldb_vqid_v_waddr         (i_hqm_system_rf_lut_vf_ldb_vqid_v_waddr),
       .rf_lut_vf_ldb_vqid_v_we            (i_hqm_system_rf_lut_vf_ldb_vqid_v_we),
       .rf_lut_vf_ldb_vqid_v_wclk          (i_hqm_system_rf_lut_vf_ldb_vqid_v_wclk),
       .rf_lut_vf_ldb_vqid_v_wclk_rst_n    (i_hqm_system_rf_lut_vf_ldb_vqid_v_wclk_rst_n),
       .rf_lut_vf_ldb_vqid_v_wdata         (i_hqm_system_rf_lut_vf_ldb_vqid_v_wdata),
       .rf_lut_vf_ldb_vqid_v_rdata         (i_hqm_system_rf_lut_vf_ldb_vqid_v_rdata),
       .rf_msix_tbl_word0_re               (i_hqm_system_rf_msix_tbl_word0_re),
       .rf_msix_tbl_word0_rclk             (i_hqm_system_rf_msix_tbl_word0_rclk),
       .rf_msix_tbl_word0_rclk_rst_n       (i_hqm_system_rf_msix_tbl_word0_rclk_rst_n),
       .rf_msix_tbl_word0_raddr            (i_hqm_system_rf_msix_tbl_word0_raddr),
       .rf_msix_tbl_word0_waddr            (i_hqm_system_rf_msix_tbl_word0_waddr),
       .rf_msix_tbl_word0_we               (i_hqm_system_rf_msix_tbl_word0_we),
       .rf_msix_tbl_word0_wclk             (i_hqm_system_rf_msix_tbl_word0_wclk),
       .rf_msix_tbl_word0_wclk_rst_n       (i_hqm_system_rf_msix_tbl_word0_wclk_rst_n),
       .rf_msix_tbl_word0_wdata            (i_hqm_system_rf_msix_tbl_word0_wdata),
       .rf_msix_tbl_word0_rdata            (i_hqm_system_rf_msix_tbl_word0_rdata),
       .rf_msix_tbl_word1_re               (i_hqm_system_rf_msix_tbl_word1_re),
       .rf_msix_tbl_word1_rclk             (i_hqm_system_rf_msix_tbl_word1_rclk),
       .rf_msix_tbl_word1_rclk_rst_n       (i_hqm_system_rf_msix_tbl_word1_rclk_rst_n),
       .rf_msix_tbl_word1_raddr            (i_hqm_system_rf_msix_tbl_word1_raddr),
       .rf_msix_tbl_word1_waddr            (i_hqm_system_rf_msix_tbl_word1_waddr),
       .rf_msix_tbl_word1_we               (i_hqm_system_rf_msix_tbl_word1_we),
       .rf_msix_tbl_word1_wclk             (i_hqm_system_rf_msix_tbl_word1_wclk),
       .rf_msix_tbl_word1_wclk_rst_n       (i_hqm_system_rf_msix_tbl_word1_wclk_rst_n),
       .rf_msix_tbl_word1_wdata            (i_hqm_system_rf_msix_tbl_word1_wdata),
       .rf_msix_tbl_word1_rdata            (i_hqm_system_rf_msix_tbl_word1_rdata),
       .rf_msix_tbl_word2_re               (i_hqm_system_rf_msix_tbl_word2_re),
       .rf_msix_tbl_word2_rclk             (i_hqm_system_rf_msix_tbl_word2_rclk),
       .rf_msix_tbl_word2_rclk_rst_n       (i_hqm_system_rf_msix_tbl_word2_rclk_rst_n),
       .rf_msix_tbl_word2_raddr            (i_hqm_system_rf_msix_tbl_word2_raddr),
       .rf_msix_tbl_word2_waddr            (i_hqm_system_rf_msix_tbl_word2_waddr),
       .rf_msix_tbl_word2_we               (i_hqm_system_rf_msix_tbl_word2_we),
       .rf_msix_tbl_word2_wclk             (i_hqm_system_rf_msix_tbl_word2_wclk),
       .rf_msix_tbl_word2_wclk_rst_n       (i_hqm_system_rf_msix_tbl_word2_wclk_rst_n),
       .rf_msix_tbl_word2_wdata            (i_hqm_system_rf_msix_tbl_word2_wdata),
       .rf_msix_tbl_word2_rdata            (i_hqm_system_rf_msix_tbl_word2_rdata),
       .rf_sch_out_fifo_re                 (i_hqm_system_rf_sch_out_fifo_re),
       .rf_sch_out_fifo_rclk               (i_hqm_system_rf_sch_out_fifo_rclk),
       .rf_sch_out_fifo_rclk_rst_n         (i_hqm_system_rf_sch_out_fifo_rclk_rst_n),
       .rf_sch_out_fifo_raddr              (i_hqm_system_rf_sch_out_fifo_raddr),
       .rf_sch_out_fifo_waddr              (i_hqm_system_rf_sch_out_fifo_waddr),
       .rf_sch_out_fifo_we                 (i_hqm_system_rf_sch_out_fifo_we),
       .rf_sch_out_fifo_wclk               (i_hqm_system_rf_sch_out_fifo_wclk),
       .rf_sch_out_fifo_wclk_rst_n         (i_hqm_system_rf_sch_out_fifo_wclk_rst_n),
       .rf_sch_out_fifo_wdata              (i_hqm_system_rf_sch_out_fifo_wdata),
       .rf_sch_out_fifo_rdata              (i_hqm_system_rf_sch_out_fifo_rdata),
       .sr_rob_mem_re                      (i_hqm_system_sr_rob_mem_re),
       .sr_rob_mem_clk                     (i_hqm_system_sr_rob_mem_clk),
       .sr_rob_mem_clk_rst_n               (i_hqm_system_sr_rob_mem_clk_rst_n),
       .sr_rob_mem_addr                    (i_hqm_system_sr_rob_mem_addr),
       .sr_rob_mem_we                      (i_hqm_system_sr_rob_mem_we),
       .sr_rob_mem_wdata                   (i_hqm_system_sr_rob_mem_wdata),
       .sr_rob_mem_rdata                   (i_hqm_system_sr_rob_mem_rdata));

   hqm_AW_flop i_hqm_system_clk_ungate_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bxx),
       .data   (hqm_clk_ungate),
       .data_q (hqm_clk_ungate_rptrxx));

   hqm_AW_clkgate i_hqm_system_clkgate
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_inp_gated_clk_enable_rptrxx),
       .cfg_clkungate   (hqm_clk_ungate_rptrxx),
       .fscan_clkungate,
       .gated_clk       (hqm_inp_gated_clkxx));

   hqm_AW_clkgate i_hqm_system_clkproc
      (.clk             (hqm_clk_trunk),
       .enable          (hqm_gated_clk_enable_rptr_sys),
       .cfg_clkungate   (hqm_clk_ungate_rptrxx),
       .fscan_clkungate,
       .gated_clk       (hqm_gated_clk_sys));

   hqm_AW_flop_set i_hqm_system_flr_prep_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bxx),
       .data   (hqm_flr_prep),
       .data_q (hqm_flr_prep_rptrxx));

   hqm_AW_reset_sync_scan i_hqm_system_hqm_clk_rptr_rst_sync_n
      (.clk            (hqm_clk_trunk),
       .rst_n          (hqm_clk_rptr_rst_b),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (hqm_clk_rptr_rst_sync_bxx));

   hqm_AW_clkand2_comb
      #(.WIDTH(1)) i_hqm_system_hqm_gated_clk_enable_and2
      (.clki0 (hqm_gated_local_clk_en_sys),
       .clki1 (hqm_clk_enable),
       .clko  (hqm_gated_clk_enable_and_sys));

   hqm_AW_clkor2_comb
      #(.WIDTH(1)) i_hqm_system_hqm_gated_clk_enable_or2
      (.clki0 (i_hqm_system_hqm_proc_clk_en_sys),
       .clki1 (hqm_gated_local_override),
       .clko  (hqm_gated_local_clk_en_sys));

   hqm_AW_flop i_hqm_system_hqm_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bxx),
       .data   (hqm_gated_clk_enable_and_sys),
       .data_q (hqm_gated_clk_enable_rptr_sys));

   hqm_AW_flop i_hqm_system_hqm_inp_gated_clk_enable_rptr
      (.clk    (hqm_clk_trunk),
       .rst_n  (hqm_clk_rptr_rst_sync_bxx),
       .data   (hqm_clk_enable),
       .data_q (hqm_inp_gated_clk_enable_rptrxx));

   hqm_AW_flop i_hqm_system_prim_clk_enable_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (prim_clk_enable),
       .data_q (prim_clk_enable_rptr));

   hqm_AW_flop i_hqm_system_prim_clk_ungate_rptr
      (.clk    (prim_clk),
       .rst_n  (side_rst_sync_prim_n),
       .data   (prim_clk_ungate),
       .data_q (prim_clk_ungate_rptr_sys));

   hqm_AW_clkgate i_hqm_system_prim_clkgate
      (.clk             (prim_clk),
       .enable          (prim_clk_enable_rptr),
       .cfg_clkungate   (prim_clk_ungate_rptr_sys),
       .fscan_clkungate,
       .gated_clk       (prim_gated_clk));

   hqm_AW_reset_core
      #(.NUM_GATED(1),
        .NUM_INP_GATED(1),
        .NUM_PATCH_GATED(1),
        .NUM_PGSB(1),
        .NO_PGCB(1)) i_hqm_system_reset_core
      (.fscan_rstbypen,
       .fscan_byprst_b,
       // Tie to constant value: zero
       .hqm_pgcb_clk           (1'b0),
       .hqm_pgcb_rst_n         (),
       .hqm_pgcb_rst_n_start   (),
       .hqm_inp_gated_clk      (hqm_inp_gated_clkxx),
       .hqm_inp_gated_rst_b    (hqm_gated_rst_b),
       .hqm_inp_gated_rst_n    (hqm_inp_gated_rst_b_sys),
       .hqm_gated_clk          (hqm_gated_clk_sys),
       .hqm_gated_rst_b,
       .hqm_gated_rst_n        (hqm_gated_rst_b_sys),
       .hqm_gated_rst_n_start  (hqm_gated_rst_b_start_sys),
       .hqm_gated_rst_n_active (hqm_gated_rst_b_active_sys),
       .hqm_gated_rst_n_done   (hqm_gated_rst_b_done_sys),
       .hqm_flr_prep           (hqm_flr_prep_rptrxx),
       .rst_prep               (hqm_rst_prep_sys));

   hqm_AW_reset_sync_scan i_hqm_system_side_rst_sync_prim_n
      (.clk            (prim_clk),
       .rst_n          (i_hqm_system_side_rst_sync_prim_n_rst_n),
       .fscan_rstbypen,
       .fscan_byprst_b,
       .rst_n_sync     (side_rst_sync_prim_n));

   assign ap_alarm_down_v                                   = i_hqm_list_sel_pipe_ap_alarm_down_v;
   assign ap_alarm_up_ready                                 = i_hqm_list_sel_pipe_ap_alarm_up_ready;
   assign ap_aqed_ready                                     = i_hqm_aqed_pipe_ap_aqed_ready;
   assign ap_aqed_v                                         = i_hqm_list_sel_pipe_ap_aqed_v;
   assign ap_cfg_req_down_read                              = i_hqm_list_sel_pipe_ap_cfg_req_down_read;
   assign ap_cfg_req_down_write                             = i_hqm_list_sel_pipe_ap_cfg_req_down_write;
   assign ap_cfg_rsp_down_ack                               = i_hqm_list_sel_pipe_ap_cfg_rsp_down_ack;
   assign aqed_alarm_down_v                                 = i_hqm_aqed_pipe_aqed_alarm_down_v;
   assign aqed_ap_enq_ready                                 = i_hqm_list_sel_pipe_aqed_ap_enq_ready;
   assign aqed_ap_enq_v                                     = i_hqm_aqed_pipe_aqed_ap_enq_v;
   assign aqed_chp_sch_ready                                = i_hqm_credit_hist_pipe_aqed_chp_sch_ready;
   assign aqed_chp_sch_v                                    = i_hqm_aqed_pipe_aqed_chp_sch_v;
   assign aqed_lsp_sch_ready                                = i_hqm_list_sel_pipe_aqed_lsp_sch_ready;
   assign aqed_lsp_sch_v                                    = i_hqm_aqed_pipe_aqed_lsp_sch_v;
   assign aqed_unit_idle                                    = i_hqm_aqed_pipe_aqed_unit_idle;
   assign chp_alarm_up_ready                                = i_hqm_credit_hist_pipe_chp_alarm_up_ready;
   assign chp_cfg_req_down_read                             = i_hqm_credit_hist_pipe_chp_cfg_req_down_read;
   assign chp_cfg_req_down_write                            = i_hqm_credit_hist_pipe_chp_cfg_req_down_write;
   assign chp_cfg_rsp_down_ack                              = i_hqm_credit_hist_pipe_chp_cfg_rsp_down_ack;
   assign chp_lsp_cmp_ready                                 = i_hqm_list_sel_pipe_chp_lsp_cmp_ready;
   assign chp_lsp_cmp_v                                     = i_hqm_credit_hist_pipe_chp_lsp_cmp_v;
   assign chp_lsp_token_ready                               = i_hqm_list_sel_pipe_chp_lsp_token_ready;
   assign chp_lsp_token_v                                   = i_hqm_credit_hist_pipe_chp_lsp_token_v;
   assign chp_rop_hcw_ready                                 = i_hqm_reorder_pipe_chp_rop_hcw_ready;
   assign chp_rop_hcw_v                                     = i_hqm_credit_hist_pipe_chp_rop_hcw_v;
   assign cwdi_interrupt_w_req_ready                        = i_hqm_system_cwdi_interrupt_w_req_ready;
   assign cwdi_interrupt_w_req_valid                        = i_hqm_credit_hist_pipe_cwdi_interrupt_w_req_valid;
   assign dp_lsp_enq_dir_ready                              = i_hqm_list_sel_pipe_dp_lsp_enq_dir_ready;
   assign dp_lsp_enq_dir_v                                  = i_hqm_qed_pipe_dp_lsp_enq_dir_v;
   assign dp_lsp_enq_rorply_ready                           = i_hqm_list_sel_pipe_dp_lsp_enq_rorply_ready;
   assign dp_lsp_enq_rorply_v                               = i_hqm_qed_pipe_dp_lsp_enq_rorply_v;
   assign hcw_enq_w_req_ready                               = i_hqm_credit_hist_pipe_hcw_enq_w_req_ready;
   assign hcw_enq_w_req_valid                               = i_hqm_system_hcw_enq_w_req_valid;
   assign hcw_sched_w_req_ready                             = i_hqm_system_hcw_sched_w_req_ready;
   assign hcw_sched_w_req_valid                             = i_hqm_credit_hist_pipe_hcw_sched_w_req_valid;
   assign hqm_alarm_ready                                   = i_hqm_system_hqm_alarm_ready;
   assign hqm_alarm_v                                       = i_hqm_credit_hist_pipe_chp_alarm_down_v;
   assign hqm_proc_clk_en_chp                               = i_hqm_credit_hist_pipe_hqm_proc_clk_en_chp;
   assign hqm_proc_clk_en_dir                               = i_hqm_qed_pipe_hqm_proc_clk_en_dir;
   assign hqm_proc_clk_en_lsp                               = i_hqm_list_sel_pipe_hqm_proc_clk_en_lsp;
   assign hqm_proc_clk_en_nalb                              = i_hqm_qed_pipe_hqm_proc_clk_en_nalb;
   assign hqm_proc_clk_en_sys                               = i_hqm_system_hqm_proc_clk_en_sys;
   assign interrupt_w_req_ready                             = i_hqm_system_interrupt_w_req_ready;
   assign interrupt_w_req_valid                             = i_hqm_credit_hist_pipe_interrupt_w_req_valid;
   assign lsp_alarm_down_v                                  = i_hqm_list_sel_pipe_lsp_alarm_down_v;
   assign lsp_alarm_up_ready                                = i_hqm_list_sel_pipe_lsp_alarm_up_ready;
   assign lsp_cfg_req_down_read                             = i_hqm_list_sel_pipe_lsp_cfg_req_down_read;
   assign lsp_cfg_req_down_write                            = i_hqm_list_sel_pipe_lsp_cfg_req_down_write;
   assign lsp_cfg_rsp_down_ack                              = i_hqm_list_sel_pipe_lsp_cfg_rsp_down_ack;
   assign lsp_dp_sch_dir_ready                              = i_hqm_qed_pipe_lsp_dp_sch_dir_ready;
   assign lsp_dp_sch_dir_v                                  = i_hqm_list_sel_pipe_lsp_dp_sch_dir_v;
   assign lsp_dp_sch_rorply_ready                           = i_hqm_qed_pipe_lsp_dp_sch_rorply_ready;
   assign lsp_dp_sch_rorply_v                               = i_hqm_list_sel_pipe_lsp_dp_sch_rorply_v;
   assign lsp_nalb_sch_atq_ready                            = i_hqm_qed_pipe_lsp_nalb_sch_atq_ready;
   assign lsp_nalb_sch_atq_v                                = i_hqm_list_sel_pipe_lsp_nalb_sch_atq_v;
   assign lsp_nalb_sch_rorply_ready                         = i_hqm_qed_pipe_lsp_nalb_sch_rorply_ready;
   assign lsp_nalb_sch_rorply_v                             = i_hqm_list_sel_pipe_lsp_nalb_sch_rorply_v;
   assign lsp_nalb_sch_unoord_ready                         = i_hqm_qed_pipe_lsp_nalb_sch_unoord_ready;
   assign lsp_nalb_sch_unoord_v                             = i_hqm_list_sel_pipe_lsp_nalb_sch_unoord_v;
   assign nalb_lsp_enq_lb_ready                             = i_hqm_list_sel_pipe_nalb_lsp_enq_lb_ready;
   assign nalb_lsp_enq_lb_v                                 = i_hqm_qed_pipe_nalb_lsp_enq_lb_v;
   assign nalb_lsp_enq_rorply_ready                         = i_hqm_list_sel_pipe_nalb_lsp_enq_rorply_ready;
   assign nalb_lsp_enq_rorply_v                             = i_hqm_qed_pipe_nalb_lsp_enq_rorply_v;
   assign qed_alarm_down_v                                  = i_hqm_qed_pipe_qed_alarm_down_v;
   assign qed_alarm_up_ready                                = i_hqm_qed_pipe_qed_alarm_up_ready;
   assign qed_aqed_enq_ready                                = i_hqm_aqed_pipe_qed_aqed_enq_ready;
   assign qed_aqed_enq_v                                    = i_hqm_qed_pipe_qed_aqed_enq_v;
   assign qed_cfg_req_down_read                             = i_hqm_qed_pipe_qed_cfg_req_down_read;
   assign qed_cfg_req_down_write                            = i_hqm_qed_pipe_qed_cfg_req_down_write;
   assign qed_cfg_rsp_down_ack                              = i_hqm_qed_pipe_qed_cfg_rsp_down_ack;
   assign qed_chp_sch_ready                                 = i_hqm_credit_hist_pipe_qed_chp_sch_ready;
   assign qed_chp_sch_v                                     = i_hqm_qed_pipe_qed_chp_sch_v;
   assign rop_alarm_down_v                                  = i_hqm_reorder_pipe_rop_alarm_down_v;
   assign rop_alarm_up_ready                                = i_hqm_reorder_pipe_rop_alarm_up_ready;
   assign rop_cfg_req_down_read                             = i_hqm_reorder_pipe_rop_cfg_req_down_read;
   assign rop_cfg_req_down_write                            = i_hqm_reorder_pipe_rop_cfg_req_down_write;
   assign rop_cfg_rsp_down_ack                              = i_hqm_reorder_pipe_rop_cfg_rsp_down_ack;
   assign rop_dp_enq_ready                                  = i_hqm_qed_pipe_rop_dp_enq_ready;
   assign rop_dp_enq_v                                      = i_hqm_reorder_pipe_rop_dp_enq_v;
   assign rop_dqed_enq_ready                                = i_hqm_qed_pipe_rop_dqed_enq_ready;
   assign rop_lsp_reordercmp_ready                          = i_hqm_list_sel_pipe_rop_lsp_reordercmp_ready;
   assign rop_lsp_reordercmp_v                              = i_hqm_reorder_pipe_rop_lsp_reordercmp_v;
   assign rop_nalb_enq_ready                                = i_hqm_qed_pipe_rop_nalb_enq_ready;
   assign rop_nalb_enq_v                                    = i_hqm_reorder_pipe_rop_nalb_enq_v;
   assign rop_qed_dqed_enq_v                                = i_hqm_reorder_pipe_rop_qed_dqed_enq_v;
   assign rop_qed_enq_ready                                 = i_hqm_qed_pipe_rop_qed_enq_ready;
   assign rop_qed_force_clockon                             = i_hqm_reorder_pipe_rop_qed_force_clockon;
   assign rop_unit_idle                                     = i_hqm_reorder_pipe_rop_unit_idle;
   assign system_cfg_req_down_read                          = i_hqm_system_system_cfg_req_down_read;
   assign system_cfg_req_down_write                         = i_hqm_system_system_cfg_req_down_write;
   assign system_cfg_rsp_down_ack                           = i_hqm_system_system_cfg_rsp_down_ack;
   assign i_hqm_aqed_pipe_aqed_lsp_deq_v                    = aqed_lsp_deq_v;
   assign i_hqm_credit_hist_pipe_chp_cfg_req_down_1_0       = chp_cfg_req_down[1:0];
   assign i_hqm_credit_hist_pipe_chp_cfg_rsp_down_5_4       = chp_cfg_rsp_down[5:4];
   assign i_hqm_list_sel_pipe_ap_cfg_req_down_1_0           = ap_cfg_req_down[1:0];
   assign i_hqm_list_sel_pipe_ap_cfg_rsp_down_5_4           = ap_cfg_rsp_down[5:4];
   assign i_hqm_list_sel_pipe_lsp_cfg_req_down_1_0          = lsp_cfg_req_down[1:0];
   assign i_hqm_list_sel_pipe_lsp_cfg_rsp_down_5_4          = lsp_cfg_rsp_down[5:4];
   assign i_hqm_qed_pipe_qed_cfg_req_down_1_0               = qed_cfg_req_down[1:0];
   assign i_hqm_qed_pipe_qed_cfg_rsp_down_5_4               = qed_cfg_rsp_down[5:4];
   assign i_hqm_qed_pipe_qed_lsp_deq_v                      = qed_lsp_deq_v;
   assign i_hqm_reorder_pipe_rop_cfg_req_down_1_0           = rop_cfg_req_down[1:0];
   assign i_hqm_reorder_pipe_rop_cfg_rsp_down_5_4           = rop_cfg_rsp_down[5:4];
   assign i_hqm_system_system_cfg_req_down_1_0              = system_cfg_req_down[1:0];
   assign i_hqm_system_system_cfg_rsp_down_5_4              = system_cfg_rsp_down[5:4];


endmodule
