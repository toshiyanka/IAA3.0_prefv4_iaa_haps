module ctech_lib_msff (
   input logic clk,
   input logic d,
   output logic o
);
   d04fkn00ld0b5 ctech_lib_dcszo (.clk(clk), .d(d), .o(o));
endmodule
