//------------------------------------------------------------------------------------------------------------------------
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2023 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code ("Material") are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//
//------------------------------------------------------------------------------------------------------------------------
// Intel Proprietary        Intel Confidential        Intel Proprietary        Intel Confidential        Intel Proprietary
//------------------------------------------------------------------------------------------------------------------------
// Generated by                  : cudoming
// Generated on                  : April 19, 2023
//------------------------------------------------------------------------------------------------------------------------
// General Information:
// ------------------------------
// 1r1w0c standard array DFX wrapper for SDG server designs.
// Synthesizable RTL for array DFX wrapper.
// RTL is written in SystemVerilog.
//------------------------------------------------------------------------------------------------------------------------
// Detail Information:
// ------------------------------
// Addresses        : RD/WR addresses are encoded.
//                    Input addresses will be valid at the array in 1 phases after being driven.
//                    Address latency of 1 is corresponding to a B-latch.
// Enables          : RD/WR enables are used to condition the clock and wordlines.
//                  : Input enables will be valid at the array in 1 phases after being driven.
//                    Enable latency of 1 is corresponding to a B-latch.
// Write Data       : Write data will be valid at the array 2 phases after being driven.
//                    Write data latency of 2 is corresponding to a rising-edge flop. 
// Read Data        : Read data will be valid at the output of a SDL 1 phase after being read.
//                    Read data latency of 1 is corresponding to a B-latch.
// Address Offset   : 
//------------------------------------------------------------------------------------------------------------------------
//
//------------------------------------------------------------------------------------------------------------------------
// Other Information:
// ------------------------------
// SDG RFIP RTL Release Path:
// /p/hdk/rtl/ip_releases/shdk74/array_macro_module
//
//------------------------------------------------------------------------------------------------------------------------


`ifdef INTC_MEM_DISABLE_CTECH_SCAN_FEATURES
  `define INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
`endif // INTC_MEM_DISABLE_CTECH_SCAN_FEATURES

`ifndef ARF124B256E1R1W0CBBEHCAA4ACW_DFX_WRAPPER_SV
`define ARF124B256E1R1W0CBBEHCAA4ACW_DFX_WRAPPER_SV

///------------------------------------------------------------------------------------------------------------------------
/// Parent Module    : n\a
/// Child Module     : arf124b256e1r1w0cbbehcaa4acw
///------------------------------------------------------------------------------------------------------------------------


// LV_pragma translate_off
// LV_pragma translate_on

//------------------------------------------------------------------------------------------------------------------------
// module arf124b256e1r1w0cbbehcaa4acw_dfx_wrapper
//------------------------------------------------------------------------------------------------------------------------
module arf124b256e1r1w0cbbehcaa4acw_dfx_wrapper #
(

//------------------------------------------------------------------------------------------------------------------------
// parameters
//------------------------------------------------------------------------------------------------------------------------
  parameter MODULE                                = "arf124b256e1r1w0cbbehcaa4acw_dfx_wrapper",
  parameter BITS                                  = 124,
  parameter ENTRIES                               = 256,
  parameter AWIDTH                                = 8,
  parameter DWIDTH                                = 124,
  parameter RD_PORTS                              = 1,
  parameter WR_PORTS                              = 1,
  parameter CM_PORTS                              = 0,
  parameter BPHASE_RD                             = 0,
  parameter BPHASE_WR                             = 0,
  parameter BPHASE_CM                             = 0,
  parameter SEGMENTS                              = 0,
  parameter BITS_PER_SEGMENT                      = 0,
  parameter SDL_INITVAL                           = {1'b0},
  parameter ADDRESS_OFFSET                        = 0,
  parameter NO_CAM_LATENCY                        = 0,
  parameter NO_CAM_LSB                            = 0,
  parameter NUM_FLCP_FD                           = 3,
  parameter NUM_FLCP_RD                           = 3,
//  parameter BYPASS_CTECH                          = 0,
  parameter COL_REPAIR_WIDTH                      = 13,
  parameter ROW_REPAIR_WIDTH                      = 13,
  parameter NUM_FUSE_MISC                         = 20,
  parameter NUM_PWR_MGMT_MISC                     = 4,
  parameter BYPASS_RD_CLK_MUX                     = 1,//default 1
  parameter BYPASS_WR_CLK_MUX                     = 1,//default 1
  parameter BYPASS_CM_CLK_MUX                     = 1,//default 1
  parameter BYPASS_RST_B_SYNC                     = 1,//default 1
  parameter BYPASS_AFD_SYNC                       = 1,//default 1
  parameter CLOCK_METHODOLOGY                     = 1,//CTMESH == 1
  parameter RD_OUTPUT_MODE                        = 0,
  // ------------------------------
  // parameters for redundancy
  // either redundancy with physical elements or synthesis elements can be on at the same time
  // redundany with physical elements can be on only with matching array having redundancy elements
  // please contact sdg rf team or rtl primary contact for details
  // ------------------------------

  parameter NUM_COL_REPAIR                        = 1,
  parameter BYPASS_REPAIR_LATCHES                 = 0,
  parameter BYPASS_TRIM_LATCHES                   = 0,
  parameter NUM_ROW_REPAIR                        = 1,
  parameter REDUNDANCY_COL_CTECH                  = 0,
  parameter REDUNDANCY_ROW_CTECH                  = 0,
  parameter int OBS_XOR_SIZE                      = 3


)
(
  
//------------------------------------------------------------------------------------------------------------------------
// interfaces
//------------------------------------------------------------------------------------------------------------------------

  //------------------------------
  // functional read interfaces
  //------------------------------
  
  input   logic                           FUNC_RD_CLK_IN_P0,
  input   logic                           FUNC_RD_EN_IN_P0,
  output  logic   [DWIDTH-1:0]            DATA_OUT_P0,
  input   logic   [AWIDTH-1:0]            FUNC_RD_ADDR_IN_P0,



  //------------------------------
  // functional write interfaces
  //------------------------------

  input   logic                           FUNC_WR_CLK_IN_P0,
  input   logic                           FUNC_WR_EN_IN_P0,
  input   logic   [DWIDTH-1:0]            FUNC_WR_DATA_IN_P0,
  input   logic   [AWIDTH-1:0]            FUNC_WR_ADDR_IN_P0,



  //------------------------------
  // bist read interfaces
  //------------------------------
   
  input   logic                           BIST_RD_CLK_IN_P0,
  input   logic                           BIST_RD_EN_IN_P0,
  input   logic   [AWIDTH-1:0]            BIST_RD_ADDR_IN_P0,

  //------------------------------
  // bist write interfaces
  //------------------------------

  input   logic                           BIST_WR_CLK_IN_P0,
  input   logic                           BIST_WR_EN_IN_P0,
  input   logic   [DWIDTH-1:0]            BIST_WR_DATA_IN_P0,
  input   logic   [AWIDTH-1:0]            BIST_WR_ADDR_IN_P0,  


  
  //------------------------------
  // bist interfaces
  //------------------------------
  input   logic                           BIST_ENABLE,

  //------------------------------
  // rcb interfaces
  //------------------------------
  input   logic   [NUM_FLCP_FD-1:0]       flcp_fd,
  input   logic   [NUM_FLCP_RD-1:0]       flcp_rd,

  //------------------------------
  // dfx interfaces
  //------------------------------

  input   logic                           WRAPPER_RD_CLK_EN_P0,

  input   logic	                          WRAPPER_WR_CLK_EN_P0,

  input   logic                           IP_RESET_B,
  input   logic                           ARRAY_FREEZE,
  input   logic   [COL_REPAIR_WIDTH-1:0]  COL_REPAIR_IN,
  input   logic   [ROW_REPAIR_WIDTH-1:0]  ROW_REPAIR_IN,
  input   logic                           GLOBAL_RROW_EN_IN_RD_P0,
  input   logic                           OUTPUT_RESET_P0,
  input   logic                           GLOBAL_RROW_EN_IN_WR_P0,

  //------------------------------
  // scan interfaces
  //------------------------------
  input   logic                           FSCAN_CLKUNGATE,
  input   logic                           FSCAN_RAM_RDIS_B,
  input   logic                           FSCAN_RAM_WDIS_B,
  input   logic                           FSCAN_RAM_BYPSEL,
  input   logic                           FSCAN_RAM_INIT_EN,
  input   logic                           FSCAN_RAM_INIT_VAL,

  //------------------------------
  // fuse interfaces
  //------------------------------
  input   logic   [NUM_FUSE_MISC-1:0]     TRIM_FUSE_IN,
  input   logic                           ISOLATION_CONTROL_IN,
  input   logic                           SLEEP_FUSE_IN,

  //------------------------------
  // power management interfaces
  //------------------------------
  input   logic   [NUM_PWR_MGMT_MISC-1:0] PWR_MGMT_IN,
  output  logic   [NUM_PWR_MGMT_MISC-1:0] PWR_MGMT_OUT


);


  `ifndef INTEL_FAKE_MEM

// LV_pragma translate_off

  //------------------------------
  // array information
  //------------------------------
  localparam HB_BITS                = 128;  
  localparam HB_ENTRIES             = 256;  
  localparam HB_DWIDTH              = 128;  
  localparam HB_AWIDTH              = 8;  

  //------------------------------
  // redundancy information
  //------------------------------
  localparam RDN_ELEMENTS_COL       = 1;
  localparam RDN_ELEMENTS_ROW       = 0;

  localparam REDUNDANCY_PHY_COL_ON  = 1;
  localparam REDUNDANCY_PHY_ROW_ON  = 0;

  localparam SPARE_ENTRIES          = 0;
  localparam SPARE_ENTRIES_IO_HACK  = 0;

  localparam RDN_BITS               = (REDUNDANCY_PHY_COL_ON == 1) ? (BITS + (2*RDN_ELEMENTS_COL)) : (BITS);
  localparam RDN_ENTRIES            = (REDUNDANCY_PHY_ROW_ON == 1) ? (ENTRIES + RDN_ELEMENTS_ROW - SPARE_ENTRIES) : (ENTRIES);
  localparam RDN_DWIDTH             = (REDUNDANCY_PHY_COL_ON == 1) ? (BITS + (2*RDN_ELEMENTS_COL)) : (BITS);
  localparam RDN_AWIDTH             = (REDUNDANCY_PHY_ROW_ON == 1) ? $clog2(ENTRIES + RDN_ELEMENTS_ROW - SPARE_ENTRIES) : $clog2(ENTRIES);

  localparam DWIDTH_DELTA           = HB_DWIDTH - RDN_DWIDTH;
  localparam ADDR_RDN_COL           = RDN_BITS - 1;
  //localparam AWIDTH_DELTA           = HB_AWIDTH - RDN_AWIDTH;
  localparam AWIDTH_DELTA           = HB_AWIDTH - AWIDTH;
  localparam ADDR_RDN_ROW           = RDN_ENTRIES - 1;

  localparam EXTRA_BITS             = HB_BITS - RDN_BITS;
  localparam EXTRA_ENTRIES          = HB_ENTRIES - RDN_ENTRIES;

  //------------------------------
  // dfx_misc_rf_in redundancy fuse information
  //------------------------------
  localparam COL_REPAIR_IN_CREN    = 0;
  localparam COL_REPAIR_IN_CRMIN   = 1;
  localparam COL_REPAIR_IN_CRMAX   = $clog2(BITS)+2-1;
  localparam ROW_REPAIR_IN_RREN    = 1;
  localparam ROW_REPAIR_IN_RRMIN   = 2;
  localparam ROW_REPAIR_IN_RRMAX   = $clog2(ENTRIES-SPARE_ENTRIES)+2-1;
  localparam int OBS_FLOP_NUM_WR   = ((BITS+AWIDTH)/OBS_XOR_SIZE)+(((BITS+AWIDTH)%OBS_XOR_SIZE)>0);
  localparam int OBS_FLOP_NUM_RD   = (AWIDTH/OBS_XOR_SIZE)+((AWIDTH%OBS_XOR_SIZE)>0);
  //------------------------------
  // nets for combining nets with lintra dangling violation in various modes
  //------------------------------
  wire                          lintra_dangling_mswt_mode;
  wire                          lintra_dangling_bypass_bist_en_sync;

  
  wire                          FUNC_RD_CLK_BYPOBS_GATED_P0;
  wire                          lintra_dangling_bypass_rd_clk_mux_P0;

  wire                          FUNC_WR_CLK_BYPOBS_GATED_P0;
  wire                          lintra_dangling_bypass_wr_clk_mux_P0;


  wire   [OBS_FLOP_NUM_WR-1:0]  mem_bypass_obs_P0;
  wire   [BITS-1:0]             mem_bypass_obs_repli_P0;

//  if (RD_OUTPUT_MODE == 0)
//  begin: read_output_mode

  //------------------------------
  // declarations
  //------------------------------
  
  //------------------------------
  // nets to clock sync mux
  //------------------------------

  wire afd_sync_wr_clk_phase_a_p0;
  wire afd_sync_wr_clk_phase_b_p0;
  wire bist_en_wr_phase_a_p0;
  wire bist_en_wr_phase_b_p0;
  wire lcb_fr_wr_clk_to_afd_sync_P0;

  wire bist_en_rd_phase_a_p0;
  wire bist_en_rd_phase_b_p0;
  wire rst_b_sync_rd_clk_phase_a_P0;
  wire rst_b_sync_rd_clk_phase_b_P0;
  wire lcb_fr_rd_clk_to_rst_b_sync_P0;



  //------------------------------
  // nets to func/bist mux
  //------------------------------

  wire                          FUNC_RD_EN_IN_P0_toMUX                ;
  wire                          BIST_RD_EN_IN_P0_toMUX                ;
  wire [AWIDTH-1:0]             FUNC_RD_ADDR_IN_P0_toMUX              ;
  wire [AWIDTH-1:0]             BIST_RD_ADDR_IN_P0_toMUX              ;

  wire                          FUNC_WR_EN_IN_P0_toMUX                ;
  wire                          BIST_WR_EN_IN_P0_toMUX                ;
  wire [AWIDTH-1:0]             FUNC_WR_ADDR_IN_P0_toMUX              ;
  wire [AWIDTH-1:0]             BIST_WR_ADDR_IN_P0_toMUX              ;
  wire [DWIDTH-1:0]             FUNC_WR_DATA_IN_P0_toMUX              ;
  wire [DWIDTH-1:0]             BIST_WR_DATA_IN_P0_toMUX              ;

  //------------------------------
  // nets to/from memory
  //------------------------------

  wire                          RD_CLK_IN_P0_toMEM            ;
  wire                          RD_EN_IN_P0_toMEM             ;
  wire  [AWIDTH-1:0]            RD_ADDR_IN_P0_toRRL           ;
  logic [HB_AWIDTH-1:0]         RD_ADDR_IN_P0_toMEM           ;
  wire  [HB_DWIDTH-1:0]         DATA_OUT_P0_fromMEM           ;
  wire  [DWIDTH-1:0]            DATA_OUT_P0_fromCRL           ;
  wire  [BITS-1:0]              DATA_OUTmx_P0                 ;
  reg   [DWIDTH-1:0]            DATA_OUT_P0_to_outmux         ;

  wire                          WR_CLK_IN_P0_toMEM            ;
  wire                          WR_EN_IN_P0_toMEM             ;
  wire  [AWIDTH-1:0]            WR_ADDR_IN_P0_toRRL           ;
  logic [HB_AWIDTH-1:0]         WR_ADDR_IN_P0_toMEM           ;
  wire  [DWIDTH-1:0]            WR_DATA_IN_P0_toCRL           ;
  wire  [HB_DWIDTH-1:0]         WR_DATA_IN_P0_toMEM           ;
  wire                          no_global_rrow_en_in_wr_P0    ;
 
  wire                          sdl_init_fromCBL_P0           ;
  wire                          sdl_init_toMEM_array_P0       ;
  wire                          sdl_initp0_toMEM              ;
  wire                          no_global_rrow_en_in_rd_P0    ;

  logic [COL_REPAIR_WIDTH-1:0]  col_repair_in_l_no_scan       ;
  logic [NUM_FUSE_MISC-1:0]     trim_fuse_in_l_no_scan        ;
  wire  [NUM_PWR_MGMT_MISC-1:0] pwr_mgmt_in_l_no_scan         ;
  wire  [NUM_PWR_MGMT_MISC-1:0] pwr_mgmt_out_l_no_scan        ;
  logic                         no_sleep_fuse_in              ;
  logic		                    no_isolation_control	      ;

  wire [COL_REPAIR_WIDTH-1:0]   col_repair_in_l_no_scan_toMEM ;
  wire [NUM_FUSE_MISC-1:0]      trim_fuse_in_l_no_scan_toMEM  ;
  wire [NUM_PWR_MGMT_MISC-1:0]  pwr_mgmt_in_l_no_scan_toMEM   ;


 
  //SOFT ROW REPAIR nets
  reg   [DWIDTH-1:0]            row_red_0_array_no_scan;  // redundant row
  logic                         row_repair_en0;
  logic [AWIDTH-1:0]            row_repair_addr0;
  wire                          row_red_0_wr_match_p0;
  wire                          row_red_0_wen_laoutp0;
  reg                           row_red_0_gwclkp0;
  

  wire                          row_red_wr_clk_p0; 
  
  wire                          row_red_0_rd_match_p0; 
  reg                           row_red_0_rd_match_ff_p0_no_scan;
  reg                           sdl_init_row_repair_0_reset_p0_no_scan;
  reg   [DWIDTH-1:0]            sdl_init_rr0_out_p0_no_scan;
  

  wire                          row_red_rd_clk_p0;
  logic                         sdl_init_regrr_p0; 
  wire                          row_red_ren_laoutp0;
  reg                           row_red_grclkp0;
    

  //------------------------------
  // logics
  //------------------------------
  //------------------------------
  //(CLOCK_METHODOLGY == 1) 
  //------------------------------
  //    if (BYPASS_CTECH == 0)
  //    begin: ctech
  //    if (CLOCK_METHODOLOGY == 1)begin:CTMESH_clock_macro
  generate

  wire rcb_rd_clk_en_p0;
  wire RCB_RD_EnableP0;
  wire rcb_rd_clk_p0;
  wire lcb_fr_rd_clk_P0;
  wire lcb_obs_rd_clk_P0;
  wire bist_en_rd_phase_a_toMux_p0  ;
  wire bist_en_rd_phase_b_toMux_p0  ;
  wire bist_en_rd_fromMux_phase_a_p0;
  wire bist_en_rd_fromMux_phase_b_p0;

  wire rst_b_sync_rd_clk_to_phase_a_P0 ;
  wire rst_b_sync_rd_clk_to_phase_b_P0 ;
  wire rst_b_sync_rd_clk_from_phase_b_P0;

  wire rcb_wr_clk_en_p0;
  wire RCB_WR_EnableP0;
  wire rcb_wr_clk_p0;  
  wire lcb_fr_wr_clk_P0;
  wire lcb_obs_wr_clk_P0;
  wire bist_en_wr_phase_a_toMux_p0;  
  wire bist_en_wr_phase_b_toMux_p0;  
  wire bist_en_wr_fromMux_phase_a_p0; 
  wire bist_en_wr_fromMux_phase_b_p0; 

  wire afd_sync_wr_clk_to_phase_a_p0;
  wire afd_sync_wr_clk_to_phase_b_p0;
  wire afd_sync_wr_clk_from_phase_b_p0;

  
  assign RCB_RD_EnableP0 = WRAPPER_RD_CLK_EN_P0 | FSCAN_CLKUNGATE;
  assign rcb_rd_clk_en_p0  = RCB_RD_EnableP0;

  assign RCB_WR_EnableP0 = WRAPPER_WR_CLK_EN_P0 | FSCAN_CLKUNGATE;
  assign rcb_wr_clk_en_p0  = RCB_WR_EnableP0;


  //--------------------------
  //READ RCB/LCB freerunning and observation
  //-------------------------- 

  arf124b256e1r1w0cbbehcaa4acw_clk_and instance_rcb_rd_p0 (.en(rcb_rd_clk_en_p0), .clk(FUNC_RD_CLK_IN_P0), .clkout(rcb_rd_clk_p0));
  arf124b256e1r1w0cbbehcaa4acw_clk_and instance_lcb_obs_rd_p0 (.clk(rcb_rd_clk_p0), .en(FSCAN_CLKUNGATE), .clkout(lcb_obs_rd_clk_P0));
  assign FUNC_RD_CLK_BYPOBS_GATED_P0 = lcb_obs_rd_clk_P0;//read obs gated clock

  if ((BYPASS_RST_B_SYNC == 0) || (BPHASE_RD == 1)) begin:lcb_fr_rd_clk

    arf124b256e1r1w0cbbehcaa4acw_clk_and instance_lcb_fr_rd_p0 (.en(1'b1), .clk(rcb_rd_clk_p0), .clkout(lcb_fr_rd_clk_P0));
    assign lcb_fr_rd_clk_to_rst_b_sync_P0 = lcb_fr_rd_clk_P0;// freerunning clock to ip_reset_b sync
  end:lcb_fr_rd_clk
    
  //-------------------------
  //WRITE RCB/LCB freeruning and observation
  //-------------------------

  arf124b256e1r1w0cbbehcaa4acw_clk_and instance_rcb_wr_p0 (.en(rcb_wr_clk_en_p0), .clk(FUNC_WR_CLK_IN_P0), .clkout(rcb_wr_clk_p0));
  arf124b256e1r1w0cbbehcaa4acw_clk_and instance_lcb_obs_wr_p0 (.clk(rcb_wr_clk_p0), .en(FSCAN_CLKUNGATE), .clkout(lcb_obs_wr_clk_P0));   
  assign FUNC_WR_CLK_BYPOBS_GATED_P0 = lcb_obs_wr_clk_P0;//write obs clock

  if ((BYPASS_AFD_SYNC == 0) || (BPHASE_WR == 1)) begin:lcb_fr_wr_clk

    arf124b256e1r1w0cbbehcaa4acw_clk_and instance_lcb_fr_wr_p0 (.en(1'b1), .clk(rcb_wr_clk_p0), .clkout(lcb_fr_wr_clk_P0));
    assign lcb_fr_wr_clk_to_afd_sync_P0 = lcb_fr_wr_clk_P0; // freerunning clk to afd sync

  end:lcb_fr_wr_clk




  //-----------------------------------
  // BISTENABLE logic
  //-----------------------------------

  //assign bist_en_phase_a = BIST_ENABLE;

  //---------------
  // BIST WR Latch
  //---------------
  if (BPHASE_WR == 1) begin:b_phase_write
    arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_bist_en_wr_p0 (.o(bist_en_wr_phase_b_toMux_p0), .d(BIST_ENABLE), .clkb(lcb_fr_wr_clk_to_afd_sync_P0));
    arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_bist_en_sync_wr_clk_p0 ( .d1(FSCAN_RAM_INIT_VAL), .d2(bist_en_wr_phase_b_toMux_p0), .s(FSCAN_RAM_INIT_EN), .o(bist_en_wr_fromMux_phase_b_p0) );
    assign bist_en_wr_phase_b_p0 = bist_en_wr_fromMux_phase_b_p0;
  end:b_phase_write

  if (BPHASE_WR == 0) begin:a_phase_write
    arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_bist_en_sync_wr_clk_p0 ( .d1(FSCAN_RAM_INIT_VAL), .d2(BIST_ENABLE), .s(FSCAN_RAM_INIT_EN), .o(bist_en_wr_fromMux_phase_a_p0));
    assign bist_en_wr_phase_a_p0 = bist_en_wr_fromMux_phase_a_p0;
  end:a_phase_write

  //---------------
  // BIST RD Latch
  //---------------
  if (BPHASE_RD == 1) begin:b_phase_read
    arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_bist_en_rd_p0 (.o(bist_en_rd_phase_b_toMux_p0), .d(BIST_ENABLE), .clkb(lcb_fr_rd_clk_to_rst_b_sync_P0));
    arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_bist_en_sync_rd_clk_p0 ( .d1(FSCAN_RAM_INIT_VAL), .d2(bist_en_rd_phase_b_toMux_p0), .s(FSCAN_RAM_INIT_EN), .o(bist_en_rd_fromMux_phase_b_p0) );
    assign bist_en_rd_phase_b_p0 = bist_en_rd_fromMux_phase_b_p0;
  end:b_phase_read

  if (BPHASE_RD == 0) begin:a_phase_read
    arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_bist_en_sync_rd_clk_p0 ( .d1(FSCAN_RAM_INIT_VAL), .d2(BIST_ENABLE), .s(FSCAN_RAM_INIT_EN), .o(bist_en_rd_fromMux_phase_a_p0));
    assign bist_en_rd_phase_a_p0 = bist_en_rd_fromMux_phase_a_p0;
  end:a_phase_read

       
       
  //------------------------------
  // ctech ARRAY FREEZE synchronizer
  //------------------------------
  if (BYPASS_AFD_SYNC == 0 ) begin: ctech_afd_sync
    if (BPHASE_WR == 1) begin:ip_afd_b_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_sync instance_ctech_afd_wr_clk_p0 ( .clk(lcb_fr_wr_clk_to_afd_sync_P0), .d(ARRAY_FREEZE), .o(afd_sync_wr_clk_to_phase_b_p0));
      arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_afd_sync_wr_clk_p0 (.o(afd_sync_wr_clk_from_phase_b_p0), .d(afd_sync_wr_clk_to_phase_b_p0), .clkb(lcb_fr_wr_clk_to_afd_sync_P0));                                        
      assign afd_sync_wr_clk_phase_b_p0 = afd_sync_wr_clk_from_phase_b_p0;
    end:ip_afd_b_latch
    
    if (BPHASE_WR == 0) begin:ip_afd_to_a_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_sync instance_ctech_afd_wr_clk_p0 ( .clk(lcb_fr_wr_clk_to_afd_sync_P0), .d(ARRAY_FREEZE), .o(afd_sync_wr_clk_to_phase_a_p0));
      assign afd_sync_wr_clk_phase_a_p0 = afd_sync_wr_clk_to_phase_a_p0;
    end:ip_afd_to_a_latch
  end: ctech_afd_sync  
   
  //------------------------------
  // bypass ARRAY FREEZE synchronizer
  //------------------------------
  if (BYPASS_AFD_SYNC == 1) begin: ctech_bypass_afd_sync
    if (BPHASE_WR == 1) begin:ip_afd_b_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_afd_sync_wr_clk_p0 (.o(afd_sync_wr_clk_from_phase_b_p0), .d(ARRAY_FREEZE), .clkb(lcb_fr_wr_clk_to_afd_sync_P0));
      assign afd_sync_wr_clk_phase_b_p0 = afd_sync_wr_clk_from_phase_b_p0;
    end:ip_afd_b_latch
    if (BPHASE_WR == 0) begin:if_byp_afd_b_latch
      assign afd_sync_wr_clk_phase_a_p0 = ARRAY_FREEZE;
    end:if_byp_afd_b_latch 
  end: ctech_bypass_afd_sync
      
  //------------------------------
  // ctech IP_RESET_B synchronizer
  //------------------------------
  if (BYPASS_RST_B_SYNC == 0) begin: ctech_rst_b_sync
    if (BPHASE_RD == 1) begin:ip_rst_b_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_sync instance_ctech_rst_b_rd_clk_p0 ( .clk(lcb_fr_rd_clk_to_rst_b_sync_P0), .d(IP_RESET_B), .o(rst_b_sync_rd_clk_to_phase_b_P0));
      arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_rst_b_sync_rd_clk_p0 (.o(rst_b_sync_rd_clk_from_phase_b_P0), .d(rst_b_sync_rd_clk_to_phase_b_P0), .clkb(lcb_fr_rd_clk_to_rst_b_sync_P0));
      assign rst_b_sync_rd_clk_phase_b_P0 = rst_b_sync_rd_clk_from_phase_b_P0;
    end:ip_rst_b_latch
        
    if (BPHASE_RD == 0) begin:ip_rst_to_a_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_sync instance_ctech_rst_b_rd_clk_p0 ( .clk(lcb_fr_rd_clk_to_rst_b_sync_P0), .d(IP_RESET_B), .o(rst_b_sync_rd_clk_to_phase_a_P0) );
      assign rst_b_sync_rd_clk_phase_a_P0 = rst_b_sync_rd_clk_to_phase_a_P0;
    end:ip_rst_to_a_latch
  end: ctech_rst_b_sync
          
  //------------------------------
  // bypass IP_RESET_B synchronizer
  //------------------------------
  if (BYPASS_RST_B_SYNC == 1) begin: ctech_bypass_rst_b_sync
    if (BPHASE_RD == 1) begin:ip_byp_rst_b_latch
      arf124b256e1r1w0cbbehcaa4acw_ctech_latch_p instance_ctech_latch_p_rst_b_sync_rd_clk_p0 (.o(rst_b_sync_rd_clk_from_phase_b_P0), .d(IP_RESET_B), .clkb(lcb_fr_rd_clk_to_rst_b_sync_P0));
      assign rst_b_sync_rd_clk_phase_b_P0 = rst_b_sync_rd_clk_from_phase_b_P0;
    end:ip_byp_rst_b_latch

    if (BPHASE_RD == 0) begin:ip_byp_rst_to_a_latch
      assign rst_b_sync_rd_clk_phase_a_P0 = IP_RESET_B;
    end:ip_byp_rst_to_a_latch
  end:ctech_bypass_rst_b_sync

  //------------------------------
  // ctech read clock synchronizer mux
  //------------------------------
  if (BYPASS_RD_CLK_MUX == 0) begin:bypass_rd_clk_mux_off 
    arf124b256e1r1w0cbbehcaa4acw_ctech_clk_mux instance_ctech_rd_clk_mux_p0 ( .clk2(FUNC_RD_CLK_IN_P0), .clk1(BIST_RD_CLK_IN_P0), .s(bist_en_rd_phase_b_p0), .clkout(RD_CLK_IN_P0_toMEM));
  end:bypass_rd_clk_mux_off 

  //------------------------------
  // ctech bypass read clock synchronizer mux
  //------------------------------
  if (BYPASS_RD_CLK_MUX == 1) begin:bypass_rd_clk_mux_on
    assign RD_CLK_IN_P0_toMEM = FUNC_RD_CLK_IN_P0;
    assign lintra_dangling_bypass_rd_clk_mux_P0 = BIST_RD_CLK_IN_P0;
  end:bypass_rd_clk_mux_on  

  //------------------------------
  // ctech write clock synchronizer mux
  //------------------------------
  if (BYPASS_WR_CLK_MUX == 0) begin:bypass_wr_clk_mux_off 
    arf124b256e1r1w0cbbehcaa4acw_ctech_clk_mux instance_ctech_wr_clk_mux_p0 ( .clk2(FUNC_WR_CLK_IN_P0), .clk1(BIST_WR_CLK_IN_P0), .s(bist_en_wr_phase_a_p0), .clkout(WR_CLK_IN_P0_toMEM) );
  end:bypass_wr_clk_mux_off 

  //------------------------------
  // ctech bypass write clock synchronizer mux
  //------------------------------
  if (BYPASS_WR_CLK_MUX == 1) begin:bypass_wr_clk_mux_on
    assign WR_CLK_IN_P0_toMEM = FUNC_WR_CLK_IN_P0;
    assign lintra_dangling_bypass_wr_clk_mux_P0 = BIST_WR_CLK_IN_P0;
  end:bypass_wr_clk_mux_on    

  

  

  //------------------------------
  // logics fscan read disable before mux for read interfaces
  //------------------------------
  assign FUNC_RD_EN_IN_P0_toMUX = FUNC_RD_EN_IN_P0;
  assign BIST_RD_EN_IN_P0_toMUX = BIST_RD_EN_IN_P0;

  //------------------------------
  // logics fscan write disable before mux for write interfaces
  //------------------------------
  assign FUNC_WR_EN_IN_P0_toMUX = FUNC_WR_EN_IN_P0;
  assign BIST_WR_EN_IN_P0_toMUX  = BIST_WR_EN_IN_P0;

  

  //------------------------------
  //logics FUNC/BIST ADDR and DATA
  //------------------------------
  assign FUNC_RD_ADDR_IN_P0_toMUX = FUNC_RD_ADDR_IN_P0;
  assign BIST_RD_ADDR_IN_P0_toMUX = BIST_RD_ADDR_IN_P0;
  assign BIST_WR_ADDR_IN_P0_toMUX = BIST_WR_ADDR_IN_P0;
  assign FUNC_WR_ADDR_IN_P0_toMUX = FUNC_WR_ADDR_IN_P0;
  assign FUNC_WR_DATA_IN_P0_toMUX = FUNC_WR_DATA_IN_P0;
  assign BIST_WR_DATA_IN_P0_toMUX = BIST_WR_DATA_IN_P0;
 
  //------------------------------
  // logics to assert sdl_init
  //------------------------------ 
  assign sdl_init_fromCBL_P0 = (~( FSCAN_RAM_INIT_EN | rst_b_sync_rd_clk_phase_a_P0 )) | FSCAN_RAM_BYPSEL  | OUTPUT_RESET_P0;
  assign sdl_init_toMEM_array_P0 =  sdl_init_fromCBL_P0;   
  assign sdl_initp0_toMEM = sdl_init_toMEM_array_P0;

  //------------------------------
  // logics mux for read interfaces
  //------------------------------ 
  assign RD_EN_IN_P0_toMEM   = ( bist_en_rd_phase_a_p0 ? BIST_RD_EN_IN_P0_toMUX : FUNC_RD_EN_IN_P0_toMUX) & FSCAN_RAM_RDIS_B ;
  assign RD_ADDR_IN_P0_toRRL = bist_en_rd_phase_a_p0 ?  BIST_RD_ADDR_IN_P0_toMUX : FUNC_RD_ADDR_IN_P0_toMUX;



  //------------------------------
  //logics mux for DATA OUT
  //------------------------------   

  if (RD_OUTPUT_MODE==0) begin : rd_data_mux  
   
    genvar j;
    for (j=0; j<BITS; j++) begin : bypass_replica                        
       assign mem_bypass_obs_repli_P0[j] = mem_bypass_obs_P0[j%OBS_FLOP_NUM_WR];
    end : bypass_replica

    `ifdef INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
    assign DATA_OUTmx_P0 = FSCAN_RAM_BYPSEL ? mem_bypass_obs_repli_P0 :  DATA_OUT_P0_to_outmux;
    assign DATA_OUT_P0 = DATA_OUTmx_P0;

    `else // INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
    assign DATA_OUTmx_P0 = FSCAN_RAM_BYPSEL ? mem_bypass_obs_repli_P0 :  DATA_OUT_P0_to_outmux;
    arf124b256e1r1w0cbbehcaa4acw_ctech_buf ctech_buf_from_mux_P0[BITS-1:0] (.a(DATA_OUTmx_P0), .o(DATA_OUT_P0));

    `endif // INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES

  end : rd_data_mux      
  else begin : no_rd_data_mux

    `ifdef INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
    assign DATA_OUTmx_P0 =  DATA_OUT_P0_to_outmux;
    assign DATA_OUT_P0 = DATA_OUTmx_P0;

    `else  // INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
    assign DATA_OUTmx_P0 =  DATA_OUT_P0_to_outmux;
    arf124b256e1r1w0cbbehcaa4acw_ctech_buf ctech_buf_P0[BITS-1:0] (.a(DATA_OUTmx_P0), .o(DATA_OUT_P0));

    `endif // INTC_MEM_ARF124B256E1R1W0CBBEHCAA4ACW_DISABLE_CTECH_SCAN_FEATURES
  end : no_rd_data_mux

  //------------------------------
  // logics mux for write interfaces
  //------------------------------ 
  assign WR_EN_IN_P0_toMEM   = ( bist_en_wr_phase_a_p0 ? BIST_WR_EN_IN_P0_toMUX : FUNC_WR_EN_IN_P0_toMUX ) & (~afd_sync_wr_clk_phase_a_p0 & FSCAN_RAM_WDIS_B);
  assign WR_ADDR_IN_P0_toRRL = bist_en_wr_phase_a_p0 ? BIST_WR_ADDR_IN_P0_toMUX : FUNC_WR_ADDR_IN_P0_toMUX;
  
  assign WR_DATA_IN_P0_toCRL = bist_en_wr_phase_a_p0 ? BIST_WR_DATA_IN_P0_toMUX : FUNC_WR_DATA_IN_P0_toMUX; 

  


  //------------------------------
  // logics for col_repair_in
  //------------------------------
  if (BYPASS_REPAIR_LATCHES == 0) begin:Repair_latches_on
    always_latch begin: latch_no_scan_COL_REPAIR_IN
      if (~FSCAN_RAM_INIT_EN) begin
        col_repair_in_l_no_scan <= COL_REPAIR_IN; 
        row_repair_en0 <= ROW_REPAIR_IN[0] & (~|ROW_REPAIR_IN[ROW_REPAIR_WIDTH-1:(AWIDTH+1)]);
        row_repair_addr0 <= ROW_REPAIR_IN[AWIDTH:1]; 
      end
    end: latch_no_scan_COL_REPAIR_IN 
    assign col_repair_in_l_no_scan_toMEM = col_repair_in_l_no_scan;
  end:Repair_latches_on
  else if (BYPASS_REPAIR_LATCHES == 1) begin : no_col_repair_fuse_latch
    assign col_repair_in_l_no_scan = COL_REPAIR_IN;
    assign col_repair_in_l_no_scan_toMEM = col_repair_in_l_no_scan; 
    assign row_repair_en0 = ROW_REPAIR_IN[0] & (~|ROW_REPAIR_IN[ROW_REPAIR_WIDTH-1:(AWIDTH+1)]);
    assign row_repair_addr0 = ROW_REPAIR_IN[AWIDTH:1]; 
  end 

  //------------------------------
  // logics for fuse miscellaneous
  //------------------------------
  if (BYPASS_TRIM_LATCHES == 0) begin:Trim_latches_on
    always_latch begin: latch_no_scan_TRIM_FUSE_IN
      if (~FSCAN_RAM_INIT_EN) begin
        trim_fuse_in_l_no_scan <= TRIM_FUSE_IN;
      end
    end: latch_no_scan_TRIM_FUSE_IN
  end:Trim_latches_on
  else if (BYPASS_TRIM_LATCHES == 1) begin : no_trim_fuse_latch
    assign trim_fuse_in_l_no_scan = TRIM_FUSE_IN;
  end

  //------------------------------
  // logics for power management miscellaneous
  //------------------------------
  assign pwr_mgmt_in_l_no_scan = PWR_MGMT_IN;
  //assign PWR_MGMT_OUT[NUM_PWR_MGMT_MISC-1:0] = {(NUM_PWR_MGMT_MISC-0){1'b0}}; 
  //if power gating is not requested pwr mgmt out is assigned from pwr mgmt in
  assign pwr_mgmt_out_l_no_scan = pwr_mgmt_in_l_no_scan;

  assign PWR_MGMT_OUT = pwr_mgmt_out_l_no_scan;

  assign  no_sleep_fuse_in           = SLEEP_FUSE_IN   ;
  assign  no_isolation_control       = ISOLATION_CONTROL_IN	        ;

  //------------------------------
  // logics for column redundancy
  //------------------------------
   
  if ((NUM_COL_REPAIR == 1) && ((REDUNDANCY_PHY_COL_ON == 1))) begin: logics_col_redundancy_on 
  //------------------------------
  // ctech logics for column redundancy
  //------------------------------
  if (REDUNDANCY_COL_CTECH) begin: logics_col_redundancy_ctech
   
    wire [DWIDTH-1:0] ctech_mux_2to1_din_d1_p0;
    wire [DWIDTH-1:0] ctech_mux_2to1_din_d2_p0;
    wire [DWIDTH-1:0] ctech_mux_2to1_din_s_p0;
    wire [DWIDTH-1:0] ctech_mux_2to1_dout_d1_p0;
    wire [DWIDTH-1:0] ctech_mux_2to1_dout_d2_p0;
    wire [DWIDTH-1:0] ctech_mux_2to1_dout_s_p0;
  
    for (genvar i = 0; (i < (DWIDTH/2)); i++) begin: logics_col_redundancy_on_rd_for_loop
	  
      assign ctech_mux_2to1_dout_d1_p0[2*i+0] = DATA_OUT_P0_fromMEM[2*i+0+2];
      assign ctech_mux_2to1_dout_d2_p0[2*i+0] = DATA_OUT_P0_fromMEM[2*i+0];
      assign ctech_mux_2to1_dout_s_p0[2*i+0]  = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i+0) >= col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN])));
      
      assign ctech_mux_2to1_dout_d1_p0[2*i+1] = DATA_OUT_P0_fromMEM[2*i+1+2];
      assign ctech_mux_2to1_dout_d2_p0[2*i+1] = DATA_OUT_P0_fromMEM[2*i+1];
      assign ctech_mux_2to1_dout_s_p0[2*i+1]  = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i+1) >= col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN])));
       
      arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_dout_p0 (
        .o(DATA_OUT_P0_fromCRL[2*i+0]),
        .d1(ctech_mux_2to1_dout_d1_p0[2*i+0]),
        .d2(ctech_mux_2to1_dout_d2_p0[2*i+0]), 
        .s(ctech_mux_2to1_dout_s_p0[2*i+0]));
      
      arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_dout2_p0 (
        .o(DATA_OUT_P0_fromCRL[2*i+1]),
        .d1(ctech_mux_2to1_dout_d1_p0[2*i+1]),
        .d2(ctech_mux_2to1_dout_d2_p0[2*i+1]), 
        .s(ctech_mux_2to1_dout_s_p0[2*i+1]));
    end: logics_col_redundancy_on_rd_for_loop

	
    assign WR_DATA_IN_P0_toMEM[0] = WR_DATA_IN_P0_toCRL[0];
    assign WR_DATA_IN_P0_toMEM[1] = WR_DATA_IN_P0_toCRL[1];
      
    for (genvar i = 2; (i <= (DWIDTH/2)); i++) begin: logics_col_redundancy_on_wr_for_loop
      assign ctech_mux_2to1_din_d1_p0[2*i-2] = WR_DATA_IN_P0_toCRL[2*i-4];
      assign ctech_mux_2to1_din_d2_p0[2*i-2] = WR_DATA_IN_P0_toCRL[2*i-2];
      assign ctech_mux_2to1_din_s_p0[2*i-2]  = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i-2) > col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN])));
      
      assign ctech_mux_2to1_din_d1_p0[2*i-2+1] = WR_DATA_IN_P0_toCRL[2*i-4+1];
      assign ctech_mux_2to1_din_d2_p0[2*i-2+1] = WR_DATA_IN_P0_toCRL[2*i-2+1];
      assign ctech_mux_2to1_din_s_p0[2*i-2+1]  = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i-2+1) > col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN]))); 

      arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_din_p0 (
        .o(WR_DATA_IN_P0_toMEM[2*i-2]),
        .d1(ctech_mux_2to1_din_d1_p0[2*i-2]),
        .d2(ctech_mux_2to1_din_d2_p0[2*i-2]), 
        .s(ctech_mux_2to1_din_s_p0[2*i-2]));
      
      arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_din2_p0 (
        .o(WR_DATA_IN_P0_toMEM[2*i-2+1]),
        .d1(ctech_mux_2to1_din_d1_p0[2*i-2+1]),
        .d2(ctech_mux_2to1_din_d2_p0[2*i-2+1]), 
        .s(ctech_mux_2to1_din_s_p0[2*i-2+1])); 

    
    end: logics_col_redundancy_on_wr_for_loop  

   
	assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1-1-1] = WR_DATA_IN_P0_toCRL[DWIDTH-1-1];
	assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1-1]   = WR_DATA_IN_P0_toCRL[DWIDTH-1]; 
    assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1]     = WR_DATA_IN_P0_toCRL[DWIDTH-1-1];
    assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1]       = WR_DATA_IN_P0_toCRL[DWIDTH-1];
  end: logics_col_redundancy_ctech

  //------------------------------
  // non ctech logics for column redundancy
  //------------------------------
  else begin: logics_col_redundancy_non_ctech
   
    for (genvar i = 0; (i < (DWIDTH/2)); i++) begin: logics_col_redundancy_on_rd_for_loop
	
      assign DATA_OUT_P0_fromCRL[2*i+0] = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i+0) >= col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN]))) ? DATA_OUT_P0_fromMEM[2*i+0+2] : DATA_OUT_P0_fromMEM[2*i+0];
      assign DATA_OUT_P0_fromCRL[2*i+1] = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i+1) >= col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN]))) ? DATA_OUT_P0_fromMEM[2*i+1+2] : DATA_OUT_P0_fromMEM[2*i+1];
    end: logics_col_redundancy_on_rd_for_loop

    
    assign WR_DATA_IN_P0_toMEM[0] = WR_DATA_IN_P0_toCRL[0];
    assign WR_DATA_IN_P0_toMEM[1] = WR_DATA_IN_P0_toCRL[1];

    for (genvar i = 2; (i <= (DWIDTH/2)); i++) begin: logics_col_redundancy_on_wr_for_loop
      assign WR_DATA_IN_P0_toMEM[2*i-2] = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i-2) > col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN]))) ? WR_DATA_IN_P0_toCRL[2*i-4] : WR_DATA_IN_P0_toCRL[2*i-2];
      assign WR_DATA_IN_P0_toMEM[2*i-2+1] = ((col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CREN] && ((2*i-2+1) > col_repair_in_l_no_scan_toMEM[COL_REPAIR_IN_CRMAX:COL_REPAIR_IN_CRMIN]))) ? WR_DATA_IN_P0_toCRL[2*i-4+1] : WR_DATA_IN_P0_toCRL[2*i-2+1];
    end: logics_col_redundancy_on_wr_for_loop      

   
	assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1-1-1] = WR_DATA_IN_P0_toCRL[DWIDTH-1-1];
	assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1-1]   = WR_DATA_IN_P0_toCRL[DWIDTH-1]; 
    assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1-1]     = WR_DATA_IN_P0_toCRL[DWIDTH-1-1];
    assign WR_DATA_IN_P0_toMEM[HB_DWIDTH-1]       = WR_DATA_IN_P0_toCRL[DWIDTH-1];
  end: logics_col_redundancy_non_ctech
  end: logics_col_redundancy_on
  else
  begin: logics_col_redundancy_off
     
    assign DATA_OUT_P0_fromCRL = DATA_OUT_P0_fromMEM[DWIDTH-1:0];
    
    assign WR_DATA_IN_P0_toMEM = {{DWIDTH_DELTA{WR_DATA_IN_P0_toCRL[HB_DWIDTH-EXTRA_BITS-1-1-1]}},{(2*RDN_ELEMENTS_COL){WR_DATA_IN_P0_toCRL[HB_DWIDTH-EXTRA_BITS-1-1-1]}},WR_DATA_IN_P0_toCRL};
   
  end: logics_col_redundancy_off 

  //------------------------------
  // logics for row redundancy
  //------------------------------
 
   
  if (NUM_ROW_REPAIR == 1) begin: logics_row_redundancy_on
    if (BPHASE_RD == 1) begin:rd_b_phase_rr
      arf124b256e1r1w0cbbehcaa4acw_ctech_clk_inv rd_clk_inv_p0 (.clk(RD_CLK_IN_P0_toMEM), .clkout(row_red_rd_clk_p0));
    end:rd_b_phase_rr

    if (BPHASE_RD == 0) begin:rd_a_phase_rr
      assign row_red_rd_clk_p0 = RD_CLK_IN_P0_toMEM;
    end:rd_a_phase_rr

    if (BPHASE_WR == 1) begin:wr_b_phase_rr
      arf124b256e1r1w0cbbehcaa4acw_ctech_clk_inv wr_clk_inv_p0 (.clk(WR_CLK_IN_P0_toMEM), .clkout(row_red_wr_clk_p0));
    end:wr_b_phase_rr

    if (BPHASE_WR == 0) begin:wr_a_phase_rr
      assign row_red_wr_clk_p0 = WR_CLK_IN_P0_toMEM;
    end:wr_a_phase_rr

    
    always_ff @(posedge  row_red_rd_clk_p0) sdl_init_regrr_p0 <= sdl_init_fromCBL_P0;
    assign sdl_init_row_repair_0_reset_p0_no_scan = ~row_repair_en0 | sdl_init_regrr_p0;

    assign RD_ADDR_IN_P0_toMEM = {{AWIDTH_DELTA{1'b0}},RD_ADDR_IN_P0_toRRL};

    
    assign WR_ADDR_IN_P0_toMEM = {{AWIDTH_DELTA{1'b0}},WR_ADDR_IN_P0_toRRL};

    
    assign row_red_0_wen_laoutp0 = WR_EN_IN_P0_toMEM & row_repair_en0 & row_red_0_wr_match_p0;
    assign row_red_ren_laoutp0 =  RD_EN_IN_P0_toMEM;
    
    
    arf124b256e1r1w0cbbehcaa4acw_clk_and instance_ctech_clk_and_row_red_0_gwclkp0 (.clk(row_red_wr_clk_p0), .en(row_red_0_wen_laoutp0), .clkout(row_red_0_gwclkp0));
    
    arf124b256e1r1w0cbbehcaa4acw_clk_and instance_ctech_clk_and_row_red_grclkp0 (.clk(row_red_rd_clk_p0), .en(row_red_ren_laoutp0), .clkout(row_red_grclkp0));

   
    
    assign row_red_0_wr_match_p0 = GLOBAL_RROW_EN_IN_WR_P0 | (row_repair_en0 & (WR_ADDR_IN_P0_toMEM==row_repair_addr0));
    
    assign row_red_0_rd_match_p0 = GLOBAL_RROW_EN_IN_RD_P0 | (row_repair_en0 & (RD_ADDR_IN_P0_toMEM==row_repair_addr0));   
    always_ff @(posedge row_red_0_gwclkp0) begin                                  
       row_red_0_array_no_scan <= row_red_0_wr_match_p0 ? WR_DATA_IN_P0_toCRL : row_red_0_array_no_scan;
    end  

    
      
    always_ff @(posedge row_red_grclkp0, posedge sdl_init_row_repair_0_reset_p0_no_scan) begin        
      if (sdl_init_row_repair_0_reset_p0_no_scan) begin
        sdl_init_rr0_out_p0_no_scan <= {DWIDTH{1'b0}};
        row_red_0_rd_match_ff_p0_no_scan <= 1'b0;
      end else begin
        sdl_init_rr0_out_p0_no_scan <= row_red_0_rd_match_p0 ? row_red_0_array_no_scan : sdl_init_rr0_out_p0_no_scan;
        row_red_0_rd_match_ff_p0_no_scan <= row_red_0_rd_match_p0;
      end
    end
	  
     
    
    for (genvar i=0; (i<DWIDTH); i++) begin : data_out_0_row_r_on
      arf124b256e1r1w0cbbehcaa4acw_ctech_mux_2to1 instance_ctech_mux_2to1_data_out_p0_to_mux (.d1(sdl_init_rr0_out_p0_no_scan[i]), .d2(DATA_OUT_P0_fromCRL[i]), .s(row_red_0_rd_match_ff_p0_no_scan), .o(DATA_OUT_P0_to_outmux[i]));
    end : data_out_0_row_r_on       	  	
    
     
  end: logics_row_redundancy_on
  if ((NUM_ROW_REPAIR == 0) && (REDUNDANCY_PHY_ROW_ON == 0)) begin: logics_row_redundancy_off
    assign DATA_OUT_P0_to_outmux = DATA_OUT_P0_fromCRL; 
    assign RD_ADDR_IN_P0_toMEM = {{AWIDTH_DELTA{1'b0}},RD_ADDR_IN_P0_toRRL};
    assign  no_global_rrow_en_in_rd_P0 = GLOBAL_RROW_EN_IN_RD_P0;
  
    assign WR_ADDR_IN_P0_toMEM = {{AWIDTH_DELTA{1'b0}},WR_ADDR_IN_P0_toRRL};
    assign  no_global_rrow_en_in_wr_P0 = GLOBAL_RROW_EN_IN_WR_P0;
  
  end: logics_row_redundancy_off

 

  //------------------------------------------------
  // instantiation arf124b256e1r1w0cbbehcaa4acw
  //------------------------------------------------
  arf124b256e1r1w0cbbehcaa4acw array (

    //------------------------------
    // read interfaces
    //------------------------------
     .ckrdp0           ( RD_CLK_IN_P0_toMEM    )
    ,.rdenp0           ( RD_EN_IN_P0_toMEM     )
    ,.rdaddrp0         ( RD_ADDR_IN_P0_toMEM   )
    ,.rddatap0         ( DATA_OUT_P0_fromMEM   )
    ,.sdl_initp0       ( sdl_initp0_toMEM      )

    //------------------------------
    // write interfaces
    //------------------------------
    ,.ckwrp0           ( WR_CLK_IN_P0_toMEM    )
    ,.wrenp0           ( WR_EN_IN_P0_toMEM     )
    ,.wraddrp0         ( WR_ADDR_IN_P0_toMEM   )
    ,.wrdatap0         ( WR_DATA_IN_P0_toMEM   )

  

    //------------------------------
    // rcb interfaces
    //------------------------------
    ,.rdaddrp0_fd      ( flcp_fd[0] )
    ,.rdaddrp0_rd      ( flcp_rd[0] )
    ,.wraddrp0_fd      ( flcp_fd[1] )
    ,.wraddrp0_rd      ( flcp_rd[1] )
    ,.wrdatap0_fd      ( flcp_fd[2] )
    ,.wrdatap0_rd      ( flcp_rd[2] )
  );
 
  endgenerate

  //------------------------------------------------------------------------------------------------------------------------
  // swt observe flops
  //------------------------------------------------------------------------------------------------------------------------

    
  //------------------------------
  // swt observe flops for read interfaces
  //------------------------------ 
  
  arf124b256e1r1w0cbbehcaa4acw_swt_obs_ff_phase_a # (
    .OBS_PIN_NUM (AWIDTH),
    .OBS_XOR_SIZE (OBS_XOR_SIZE),
    .OBS_FLOP_NUM(OBS_FLOP_NUM_RD))
  instance_swt_obs_ff_phase_a_rd_p0 (
    .clock  ( {FUNC_RD_CLK_BYPOBS_GATED_P0} ),
    .in     ( {RD_ADDR_IN_P0_toRRL} ),
    .out    ( ));

  //------------------------------
  // swt observe flops for write interfaces
  //------------------------------ 
  
  arf124b256e1r1w0cbbehcaa4acw_swt_obs_ff_phase_a # (
    .OBS_PIN_NUM (BITS+AWIDTH),
    .OBS_XOR_SIZE (OBS_XOR_SIZE),
    .OBS_FLOP_NUM(OBS_FLOP_NUM_WR))
  instance_swt_obs_ff_phase_a_wr_p0 (
    .clock  ( {FUNC_WR_CLK_BYPOBS_GATED_P0} ),
    .in     ( {WR_DATA_IN_P0_toCRL, WR_ADDR_IN_P0_toRRL} ),
    .out    (mem_bypass_obs_P0));
  




// LV_pragma translate_on
`else //INTEL_FAKE_MEM

  (* memory *) reg [BITS-1:0] mem_array [ENTRIES-1:0] /* synthesis syn_ramstyle = "block_ram" */;

  assign PWR_MGMT_OUT = PWR_MGMT_IN;
  wire [DWIDTH-1:0]                        DATA_OUT_P0;
  //Read and Write with not
  reg [DWIDTH-1:0]                        DATA_OUT_P0_n;
  wire [DWIDTH-1:0]                        FUNC_WR_DATA_IN_P0_n;
  assign DATA_OUT_P0 = ~DATA_OUT_P0_n;
  assign FUNC_WR_DATA_IN_P0_n = ~FUNC_WR_DATA_IN_P0;
  always @(posedge FUNC_WR_CLK_IN_P0) begin
    if (FUNC_WR_EN_IN_P0) begin
      mem_array[FUNC_WR_ADDR_IN_P0] <= FUNC_WR_DATA_IN_P0_n;
    end
  end
  
  always @(posedge FUNC_RD_CLK_IN_P0) begin
    if (FUNC_RD_EN_IN_P0) begin
      DATA_OUT_P0_n <= mem_array[FUNC_RD_ADDR_IN_P0];
    end
  end
  `endif //INTEL_FAKE_MEM
endmodule // end module arf124b256e1r1w0cbbehcaa4acw_dfx_wrapper
`endif // endif ifndef ARF124B256E1R1W0CBBEHCAA4ACW_DFX_WRAPPER_SV 
