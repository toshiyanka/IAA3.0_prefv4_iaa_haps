VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf096b192e1r1w0cbbeheaa4acw
  CLASS BLOCK ;
  FOREIGN arf096b192e1r1w0cbbeheaa4acw ;
  ORIGIN 0 0 ;
  SIZE 34.2 BY 41.28 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 21.48 10.028 22.68 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 19.56 10.028 20.76 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 21.48 11.616 22.68 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 21.48 11.916 22.68 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 21.48 12.172 22.68 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 21.48 12.428 22.68 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 21.48 12.728 22.68 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 21.48 12.988 22.68 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 21.48 13.156 22.68 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 21.48 13.416 22.68 ;
    END
  END rdaddrp0[7]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 21.48 10.628 22.68 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 21.48 10.928 22.68 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 21.48 11.188 22.68 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 21.48 11.356 22.68 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 19.56 11.916 20.76 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 19.56 12.172 20.76 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 19.56 12.428 20.76 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 19.56 12.728 20.76 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 19.56 12.988 20.76 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 19.56 13.156 20.76 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 19.56 13.416 20.76 ;
    END
  END wraddrp0[6]
  PIN wraddrp0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 19.56 13.716 20.76 ;
    END
  END wraddrp0[7]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.584 19.56 10.628 20.76 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 19.56 10.928 20.76 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 9.984 0.24 10.028 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 3.84 13.072 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 3.84 13.156 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 4.56 13.628 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 4.56 13.716 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 5.28 14.056 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 5.28 14.228 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 6 14.616 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 6 10.116 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 6.72 10.928 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 6.72 11.016 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 0.24 10.116 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 7.44 11.528 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 7.44 11.616 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 8.16 12.088 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 8.16 12.172 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 8.88 12.516 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 8.88 12.728 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 9.6 13.072 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 9.6 13.156 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 10.32 13.628 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 10.32 13.716 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 0.96 11.016 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 11.04 14.056 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 11.04 14.228 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 11.76 14.616 12.96 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 11.76 10.116 12.96 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.884 12.48 10.928 13.68 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.972 12.48 11.016 13.68 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 13.2 11.528 14.4 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 13.2 11.616 14.4 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 13.92 12.088 15.12 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 13.92 12.172 15.12 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 0.96 11.188 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 14.64 12.516 15.84 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 14.64 12.728 15.84 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 15.36 13.072 16.56 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 15.36 13.156 16.56 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 16.08 13.628 17.28 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 16.08 13.716 17.28 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 16.8 14.056 18 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 16.8 14.228 18 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 17.52 14.616 18.72 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 17.52 10.116 18.72 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 1.68 11.528 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 23.28 10.288 24.48 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 23.28 10.372 24.48 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 24 11.188 25.2 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 24 11.272 25.2 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 24.72 11.616 25.92 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 24.72 11.828 25.92 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 25.44 12.172 26.64 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 25.44 12.256 26.64 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 26.16 12.728 27.36 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 26.16 12.816 27.36 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 1.68 11.616 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 26.88 13.156 28.08 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 26.88 13.328 28.08 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 27.6 13.716 28.8 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 27.6 13.888 28.8 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 28.32 14.228 29.52 ;
    END
  END wrdatap0[64]
  PIN wrdatap0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 28.32 14.316 29.52 ;
    END
  END wrdatap0[65]
  PIN wrdatap0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 29.04 10.116 30.24 ;
    END
  END wrdatap0[66]
  PIN wrdatap0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 29.04 10.288 30.24 ;
    END
  END wrdatap0[67]
  PIN wrdatap0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 29.76 11.188 30.96 ;
    END
  END wrdatap0[68]
  PIN wrdatap0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 29.76 11.272 30.96 ;
    END
  END wrdatap0[69]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 2.4 12.088 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 30.48 11.616 31.68 ;
    END
  END wrdatap0[70]
  PIN wrdatap0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 30.48 11.828 31.68 ;
    END
  END wrdatap0[71]
  PIN wrdatap0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 31.2 12.172 32.4 ;
    END
  END wrdatap0[72]
  PIN wrdatap0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 31.2 12.256 32.4 ;
    END
  END wrdatap0[73]
  PIN wrdatap0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 31.92 12.728 33.12 ;
    END
  END wrdatap0[74]
  PIN wrdatap0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 31.92 12.816 33.12 ;
    END
  END wrdatap0[75]
  PIN wrdatap0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 32.64 13.156 33.84 ;
    END
  END wrdatap0[76]
  PIN wrdatap0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 32.64 13.328 33.84 ;
    END
  END wrdatap0[77]
  PIN wrdatap0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 33.36 13.716 34.56 ;
    END
  END wrdatap0[78]
  PIN wrdatap0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 33.36 13.888 34.56 ;
    END
  END wrdatap0[79]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 2.4 12.172 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 34.08 14.228 35.28 ;
    END
  END wrdatap0[80]
  PIN wrdatap0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 34.08 14.316 35.28 ;
    END
  END wrdatap0[81]
  PIN wrdatap0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.072 34.8 10.116 36 ;
    END
  END wrdatap0[82]
  PIN wrdatap0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 34.8 10.288 36 ;
    END
  END wrdatap0[83]
  PIN wrdatap0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 35.52 11.188 36.72 ;
    END
  END wrdatap0[84]
  PIN wrdatap0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 35.52 11.272 36.72 ;
    END
  END wrdatap0[85]
  PIN wrdatap0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 36.24 11.616 37.44 ;
    END
  END wrdatap0[86]
  PIN wrdatap0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 36.24 11.828 37.44 ;
    END
  END wrdatap0[87]
  PIN wrdatap0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.128 36.96 12.172 38.16 ;
    END
  END wrdatap0[88]
  PIN wrdatap0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 36.96 12.256 38.16 ;
    END
  END wrdatap0[89]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 3.12 12.516 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 37.68 12.728 38.88 ;
    END
  END wrdatap0[90]
  PIN wrdatap0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 37.68 12.816 38.88 ;
    END
  END wrdatap0[91]
  PIN wrdatap0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.112 38.4 13.156 39.6 ;
    END
  END wrdatap0[92]
  PIN wrdatap0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 38.4 13.328 39.6 ;
    END
  END wrdatap0[93]
  PIN wrdatap0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.672 39.12 13.716 40.32 ;
    END
  END wrdatap0[94]
  PIN wrdatap0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 39.12 13.888 40.32 ;
    END
  END wrdatap0[95]
  PIN wrdatap0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.184 39.84 14.228 41.04 ;
    END
  END wrdatap0[96]
  PIN wrdatap0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 39.84 14.316 41.04 ;
    END
  END wrdatap0[97]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.684 3.12 12.728 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 19.56 11.356 20.76 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.572 19.56 11.616 20.76 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 19.56 11.188 20.76 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 0.24 10.288 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 3.84 13.328 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 3.84 13.416 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 4.56 13.888 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 4.56 13.972 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 5.28 14.316 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 5.28 14.528 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 6 10.288 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 6 10.372 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 6.72 11.188 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 6.72 11.272 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 0.24 10.372 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 7.44 11.828 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 7.44 11.916 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 8.16 12.256 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 8.16 12.428 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 8.88 12.816 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 8.88 12.988 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 9.6 13.328 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 9.6 13.416 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 10.32 13.888 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 10.32 13.972 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 0.96 11.272 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 11.04 14.316 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 11.04 14.528 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 11.76 10.288 12.96 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 11.76 10.372 12.96 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.144 12.48 11.188 13.68 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.228 12.48 11.272 13.68 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 13.2 11.828 14.4 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 13.2 11.916 14.4 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 13.92 12.256 15.12 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 13.92 12.428 15.12 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 0.96 11.356 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 14.64 12.816 15.84 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 14.64 12.988 15.84 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.284 15.36 13.328 16.56 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 15.36 13.416 16.56 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.844 16.08 13.888 17.28 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 16.08 13.972 17.28 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.272 16.8 14.316 18 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 16.8 14.528 18 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.244 17.52 10.288 18.72 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 17.52 10.372 18.72 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.784 1.68 11.828 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 23.28 10.456 24.48 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.672 23.28 10.716 24.48 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 24 11.356 25.2 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 24 11.528 25.2 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 24.72 11.916 25.92 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 24.72 12.088 25.92 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 25.44 12.428 26.64 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 25.44 12.516 26.64 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 26.16 12.988 27.36 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 26.16 13.072 27.36 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 1.68 11.916 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 26.88 13.416 28.08 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 26.88 13.628 28.08 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 27.6 13.972 28.8 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 27.6 14.056 28.8 ;
    END
  END rddatap0[63]
  PIN rddatap0[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 28.32 14.528 29.52 ;
    END
  END rddatap0[64]
  PIN rddatap0[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 28.32 14.616 29.52 ;
    END
  END rddatap0[65]
  PIN rddatap0[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 29.04 10.372 30.24 ;
    END
  END rddatap0[66]
  PIN rddatap0[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 29.04 10.456 30.24 ;
    END
  END rddatap0[67]
  PIN rddatap0[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 29.76 11.356 30.96 ;
    END
  END rddatap0[68]
  PIN rddatap0[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 29.76 11.528 30.96 ;
    END
  END rddatap0[69]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.212 2.4 12.256 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 30.48 11.916 31.68 ;
    END
  END rddatap0[70]
  PIN rddatap0[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 30.48 12.088 31.68 ;
    END
  END rddatap0[71]
  PIN rddatap0[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 31.2 12.428 32.4 ;
    END
  END rddatap0[72]
  PIN rddatap0[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 31.2 12.516 32.4 ;
    END
  END rddatap0[73]
  PIN rddatap0[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 31.92 12.988 33.12 ;
    END
  END rddatap0[74]
  PIN rddatap0[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 31.92 13.072 33.12 ;
    END
  END rddatap0[75]
  PIN rddatap0[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 32.64 13.416 33.84 ;
    END
  END rddatap0[76]
  PIN rddatap0[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 32.64 13.628 33.84 ;
    END
  END rddatap0[77]
  PIN rddatap0[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 33.36 13.972 34.56 ;
    END
  END rddatap0[78]
  PIN rddatap0[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 33.36 14.056 34.56 ;
    END
  END rddatap0[79]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 2.4 12.428 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 34.08 14.528 35.28 ;
    END
  END rddatap0[80]
  PIN rddatap0[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 34.08 14.616 35.28 ;
    END
  END rddatap0[81]
  PIN rddatap0[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.328 34.8 10.372 36 ;
    END
  END rddatap0[82]
  PIN rddatap0[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 10.412 34.8 10.456 36 ;
    END
  END rddatap0[83]
  PIN rddatap0[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.312 35.52 11.356 36.72 ;
    END
  END rddatap0[84]
  PIN rddatap0[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.484 35.52 11.528 36.72 ;
    END
  END rddatap0[85]
  PIN rddatap0[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.872 36.24 11.916 37.44 ;
    END
  END rddatap0[86]
  PIN rddatap0[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.044 36.24 12.088 37.44 ;
    END
  END rddatap0[87]
  PIN rddatap0[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.384 36.96 12.428 38.16 ;
    END
  END rddatap0[88]
  PIN rddatap0[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.472 36.96 12.516 38.16 ;
    END
  END rddatap0[89]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.772 3.12 12.816 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 37.68 12.988 38.88 ;
    END
  END rddatap0[90]
  PIN rddatap0[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.028 37.68 13.072 38.88 ;
    END
  END rddatap0[91]
  PIN rddatap0[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.372 38.4 13.416 39.6 ;
    END
  END rddatap0[92]
  PIN rddatap0[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.584 38.4 13.628 39.6 ;
    END
  END rddatap0[93]
  PIN rddatap0[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 13.928 39.12 13.972 40.32 ;
    END
  END rddatap0[94]
  PIN rddatap0[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.012 39.12 14.056 40.32 ;
    END
  END rddatap0[95]
  PIN rddatap0[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.484 39.84 14.528 41.04 ;
    END
  END rddatap0[96]
  PIN rddatap0[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 14.572 39.84 14.616 41.04 ;
    END
  END rddatap0[97]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 12.944 3.12 12.988 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 41.22 ;
        RECT 2.662 0.06 2.738 41.22 ;
        RECT 4.462 0.06 4.538 41.22 ;
        RECT 6.262 0.06 6.338 41.22 ;
        RECT 8.062 0.06 8.138 41.22 ;
        RECT 9.862 0.06 9.938 41.22 ;
        RECT 11.662 0.06 11.738 41.22 ;
        RECT 13.462 0.06 13.538 41.22 ;
        RECT 15.262 0.06 15.338 41.22 ;
        RECT 17.062 0.06 17.138 41.22 ;
        RECT 18.862 0.06 18.938 41.22 ;
        RECT 20.662 0.06 20.738 41.22 ;
        RECT 22.462 0.06 22.538 41.22 ;
        RECT 24.262 0.06 24.338 41.22 ;
        RECT 26.062 0.06 26.138 41.22 ;
        RECT 27.862 0.06 27.938 41.22 ;
        RECT 29.662 0.06 29.738 41.22 ;
        RECT 31.462 0.06 31.538 41.22 ;
        RECT 33.262 0.06 33.338 41.22 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 41.22 ;
        RECT 3.562 0.06 3.638 41.22 ;
        RECT 5.362 0.06 5.438 41.22 ;
        RECT 7.162 0.06 7.238 41.22 ;
        RECT 8.962 0.06 9.038 41.22 ;
        RECT 10.762 0.06 10.838 41.22 ;
        RECT 12.562 0.06 12.638 41.22 ;
        RECT 14.362 0.06 14.438 41.22 ;
        RECT 16.162 0.06 16.238 41.22 ;
        RECT 17.962 0.06 18.038 41.22 ;
        RECT 19.762 0.06 19.838 41.22 ;
        RECT 21.562 0.06 21.638 41.22 ;
        RECT 23.362 0.06 23.438 41.22 ;
        RECT 25.162 0.06 25.238 41.22 ;
        RECT 26.962 0.06 27.038 41.22 ;
        RECT 28.762 0.06 28.838 41.22 ;
        RECT 30.562 0.06 30.638 41.22 ;
        RECT 32.362 0.06 32.438 41.22 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 34.216 41.294 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 34.22 41.3 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 34.2705 41.318 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 34.235 41.35 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 34.27 41.318 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 34.259 41.37 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 34.29 41.342 ;
    LAYER m7 SPACING 0 ;
      RECT 33.338 41.34 34.24 41.4 ;
      RECT 33.338 -0.06 34.292 41.34 ;
      RECT 33.338 -0.12 34.24 -0.06 ;
      RECT 32.438 -0.12 33.262 41.4 ;
      RECT 31.538 -0.12 32.362 41.4 ;
      RECT 30.638 -0.12 31.462 41.4 ;
      RECT 29.738 -0.12 30.562 41.4 ;
      RECT 28.838 -0.12 29.662 41.4 ;
      RECT 27.938 -0.12 28.762 41.4 ;
      RECT 27.038 -0.12 27.862 41.4 ;
      RECT 26.138 -0.12 26.962 41.4 ;
      RECT 25.238 -0.12 26.062 41.4 ;
      RECT 24.338 -0.12 25.162 41.4 ;
      RECT 23.438 -0.12 24.262 41.4 ;
      RECT 22.538 -0.12 23.362 41.4 ;
      RECT 21.638 -0.12 22.462 41.4 ;
      RECT 20.738 -0.12 21.562 41.4 ;
      RECT 19.838 -0.12 20.662 41.4 ;
      RECT 18.938 -0.12 19.762 41.4 ;
      RECT 18.038 -0.12 18.862 41.4 ;
      RECT 17.138 -0.12 17.962 41.4 ;
      RECT 16.238 -0.12 17.062 41.4 ;
      RECT 15.338 -0.12 16.162 41.4 ;
      RECT 14.438 41.04 15.262 41.4 ;
      RECT 14.438 39.84 14.484 41.04 ;
      RECT 14.528 39.84 14.572 41.04 ;
      RECT 14.616 39.84 15.262 41.04 ;
      RECT 14.438 35.28 15.262 39.84 ;
      RECT 14.438 34.08 14.484 35.28 ;
      RECT 14.528 34.08 14.572 35.28 ;
      RECT 14.616 34.08 15.262 35.28 ;
      RECT 14.438 29.52 15.262 34.08 ;
      RECT 14.438 28.32 14.484 29.52 ;
      RECT 14.528 28.32 14.572 29.52 ;
      RECT 14.616 28.32 15.262 29.52 ;
      RECT 14.438 18.72 15.262 28.32 ;
      RECT 14.438 18 14.572 18.72 ;
      RECT 14.616 17.52 15.262 18.72 ;
      RECT 14.528 17.52 14.572 18 ;
      RECT 14.438 16.8 14.484 18 ;
      RECT 14.528 16.8 15.262 17.52 ;
      RECT 14.438 12.96 15.262 16.8 ;
      RECT 14.438 12.24 14.572 12.96 ;
      RECT 14.616 11.76 15.262 12.96 ;
      RECT 14.528 11.76 14.572 12.24 ;
      RECT 14.438 11.04 14.484 12.24 ;
      RECT 14.528 11.04 15.262 11.76 ;
      RECT 14.438 7.2 15.262 11.04 ;
      RECT 14.438 6.48 14.572 7.2 ;
      RECT 14.616 6 15.262 7.2 ;
      RECT 14.528 6 14.572 6.48 ;
      RECT 14.438 5.28 14.484 6.48 ;
      RECT 14.528 5.28 15.262 6 ;
      RECT 14.438 -0.12 15.262 5.28 ;
      RECT 13.538 41.04 14.362 41.4 ;
      RECT 13.538 40.32 14.184 41.04 ;
      RECT 14.228 39.84 14.272 41.04 ;
      RECT 14.316 39.84 14.362 41.04 ;
      RECT 14.056 39.84 14.184 40.32 ;
      RECT 13.538 39.6 13.672 40.32 ;
      RECT 13.716 39.12 13.844 40.32 ;
      RECT 13.888 39.12 13.928 40.32 ;
      RECT 13.972 39.12 14.012 40.32 ;
      RECT 14.056 39.12 14.362 39.84 ;
      RECT 13.628 39.12 13.672 39.6 ;
      RECT 13.538 38.4 13.584 39.6 ;
      RECT 13.628 38.4 14.362 39.12 ;
      RECT 13.538 35.28 14.362 38.4 ;
      RECT 13.538 34.56 14.184 35.28 ;
      RECT 14.228 34.08 14.272 35.28 ;
      RECT 14.316 34.08 14.362 35.28 ;
      RECT 14.056 34.08 14.184 34.56 ;
      RECT 13.538 33.84 13.672 34.56 ;
      RECT 13.716 33.36 13.844 34.56 ;
      RECT 13.888 33.36 13.928 34.56 ;
      RECT 13.972 33.36 14.012 34.56 ;
      RECT 14.056 33.36 14.362 34.08 ;
      RECT 13.628 33.36 13.672 33.84 ;
      RECT 13.538 32.64 13.584 33.84 ;
      RECT 13.628 32.64 14.362 33.36 ;
      RECT 13.538 29.52 14.362 32.64 ;
      RECT 13.538 28.8 14.184 29.52 ;
      RECT 14.228 28.32 14.272 29.52 ;
      RECT 14.316 28.32 14.362 29.52 ;
      RECT 14.056 28.32 14.184 28.8 ;
      RECT 13.538 28.08 13.672 28.8 ;
      RECT 13.716 27.6 13.844 28.8 ;
      RECT 13.888 27.6 13.928 28.8 ;
      RECT 13.972 27.6 14.012 28.8 ;
      RECT 14.056 27.6 14.362 28.32 ;
      RECT 13.628 27.6 13.672 28.08 ;
      RECT 13.538 26.88 13.584 28.08 ;
      RECT 13.628 26.88 14.362 27.6 ;
      RECT 13.538 20.76 14.362 26.88 ;
      RECT 13.538 19.56 13.672 20.76 ;
      RECT 13.716 19.56 14.362 20.76 ;
      RECT 13.538 18 14.362 19.56 ;
      RECT 13.538 17.28 14.012 18 ;
      RECT 14.056 16.8 14.184 18 ;
      RECT 14.228 16.8 14.272 18 ;
      RECT 14.316 16.8 14.362 18 ;
      RECT 13.972 16.8 14.012 17.28 ;
      RECT 13.538 16.08 13.584 17.28 ;
      RECT 13.628 16.08 13.672 17.28 ;
      RECT 13.716 16.08 13.844 17.28 ;
      RECT 13.888 16.08 13.928 17.28 ;
      RECT 13.972 16.08 14.362 16.8 ;
      RECT 13.538 12.24 14.362 16.08 ;
      RECT 13.538 11.52 14.012 12.24 ;
      RECT 14.056 11.04 14.184 12.24 ;
      RECT 14.228 11.04 14.272 12.24 ;
      RECT 14.316 11.04 14.362 12.24 ;
      RECT 13.972 11.04 14.012 11.52 ;
      RECT 13.538 10.32 13.584 11.52 ;
      RECT 13.628 10.32 13.672 11.52 ;
      RECT 13.716 10.32 13.844 11.52 ;
      RECT 13.888 10.32 13.928 11.52 ;
      RECT 13.972 10.32 14.362 11.04 ;
      RECT 13.538 6.48 14.362 10.32 ;
      RECT 13.538 5.76 14.012 6.48 ;
      RECT 14.056 5.28 14.184 6.48 ;
      RECT 14.228 5.28 14.272 6.48 ;
      RECT 14.316 5.28 14.362 6.48 ;
      RECT 13.972 5.28 14.012 5.76 ;
      RECT 13.538 4.56 13.584 5.76 ;
      RECT 13.628 4.56 13.672 5.76 ;
      RECT 13.716 4.56 13.844 5.76 ;
      RECT 13.888 4.56 13.928 5.76 ;
      RECT 13.972 4.56 14.362 5.28 ;
      RECT 13.538 -0.12 14.362 4.56 ;
      RECT 12.638 39.6 13.462 41.4 ;
      RECT 12.638 38.88 13.112 39.6 ;
      RECT 13.156 38.4 13.284 39.6 ;
      RECT 13.328 38.4 13.372 39.6 ;
      RECT 13.416 38.4 13.462 39.6 ;
      RECT 13.072 38.4 13.112 38.88 ;
      RECT 12.638 37.68 12.684 38.88 ;
      RECT 12.728 37.68 12.772 38.88 ;
      RECT 12.816 37.68 12.944 38.88 ;
      RECT 12.988 37.68 13.028 38.88 ;
      RECT 13.072 37.68 13.462 38.4 ;
      RECT 12.638 33.84 13.462 37.68 ;
      RECT 12.638 33.12 13.112 33.84 ;
      RECT 13.156 32.64 13.284 33.84 ;
      RECT 13.328 32.64 13.372 33.84 ;
      RECT 13.416 32.64 13.462 33.84 ;
      RECT 13.072 32.64 13.112 33.12 ;
      RECT 12.638 31.92 12.684 33.12 ;
      RECT 12.728 31.92 12.772 33.12 ;
      RECT 12.816 31.92 12.944 33.12 ;
      RECT 12.988 31.92 13.028 33.12 ;
      RECT 13.072 31.92 13.462 32.64 ;
      RECT 12.638 28.08 13.462 31.92 ;
      RECT 12.638 27.36 13.112 28.08 ;
      RECT 13.156 26.88 13.284 28.08 ;
      RECT 13.328 26.88 13.372 28.08 ;
      RECT 13.416 26.88 13.462 28.08 ;
      RECT 13.072 26.88 13.112 27.36 ;
      RECT 12.638 26.16 12.684 27.36 ;
      RECT 12.728 26.16 12.772 27.36 ;
      RECT 12.816 26.16 12.944 27.36 ;
      RECT 12.988 26.16 13.028 27.36 ;
      RECT 13.072 26.16 13.462 26.88 ;
      RECT 12.638 22.68 13.462 26.16 ;
      RECT 12.638 21.48 12.684 22.68 ;
      RECT 12.728 21.48 12.944 22.68 ;
      RECT 12.988 21.48 13.112 22.68 ;
      RECT 13.156 21.48 13.372 22.68 ;
      RECT 13.416 21.48 13.462 22.68 ;
      RECT 12.638 20.76 13.462 21.48 ;
      RECT 12.638 19.56 12.684 20.76 ;
      RECT 12.728 19.56 12.944 20.76 ;
      RECT 12.988 19.56 13.112 20.76 ;
      RECT 13.156 19.56 13.372 20.76 ;
      RECT 13.416 19.56 13.462 20.76 ;
      RECT 12.638 16.56 13.462 19.56 ;
      RECT 12.638 15.84 13.028 16.56 ;
      RECT 13.072 15.36 13.112 16.56 ;
      RECT 13.156 15.36 13.284 16.56 ;
      RECT 13.328 15.36 13.372 16.56 ;
      RECT 13.416 15.36 13.462 16.56 ;
      RECT 12.988 15.36 13.028 15.84 ;
      RECT 12.638 14.64 12.684 15.84 ;
      RECT 12.728 14.64 12.772 15.84 ;
      RECT 12.816 14.64 12.944 15.84 ;
      RECT 12.988 14.64 13.462 15.36 ;
      RECT 12.638 10.8 13.462 14.64 ;
      RECT 12.638 10.08 13.028 10.8 ;
      RECT 13.072 9.6 13.112 10.8 ;
      RECT 13.156 9.6 13.284 10.8 ;
      RECT 13.328 9.6 13.372 10.8 ;
      RECT 13.416 9.6 13.462 10.8 ;
      RECT 12.988 9.6 13.028 10.08 ;
      RECT 12.638 8.88 12.684 10.08 ;
      RECT 12.728 8.88 12.772 10.08 ;
      RECT 12.816 8.88 12.944 10.08 ;
      RECT 12.988 8.88 13.462 9.6 ;
      RECT 12.638 5.04 13.462 8.88 ;
      RECT 12.638 4.32 13.028 5.04 ;
      RECT 13.072 3.84 13.112 5.04 ;
      RECT 13.156 3.84 13.284 5.04 ;
      RECT 13.328 3.84 13.372 5.04 ;
      RECT 13.416 3.84 13.462 5.04 ;
      RECT 12.988 3.84 13.028 4.32 ;
      RECT 12.638 3.12 12.684 4.32 ;
      RECT 12.728 3.12 12.772 4.32 ;
      RECT 12.816 3.12 12.944 4.32 ;
      RECT 12.988 3.12 13.462 3.84 ;
      RECT 12.638 -0.12 13.462 3.12 ;
      RECT 11.738 38.16 12.562 41.4 ;
      RECT 11.738 37.44 12.128 38.16 ;
      RECT 12.172 36.96 12.212 38.16 ;
      RECT 12.256 36.96 12.384 38.16 ;
      RECT 12.428 36.96 12.472 38.16 ;
      RECT 12.516 36.96 12.562 38.16 ;
      RECT 12.088 36.96 12.128 37.44 ;
      RECT 11.738 36.24 11.784 37.44 ;
      RECT 11.828 36.24 11.872 37.44 ;
      RECT 11.916 36.24 12.044 37.44 ;
      RECT 12.088 36.24 12.562 36.96 ;
      RECT 11.738 32.4 12.562 36.24 ;
      RECT 11.738 31.68 12.128 32.4 ;
      RECT 12.172 31.2 12.212 32.4 ;
      RECT 12.256 31.2 12.384 32.4 ;
      RECT 12.428 31.2 12.472 32.4 ;
      RECT 12.516 31.2 12.562 32.4 ;
      RECT 12.088 31.2 12.128 31.68 ;
      RECT 11.738 30.48 11.784 31.68 ;
      RECT 11.828 30.48 11.872 31.68 ;
      RECT 11.916 30.48 12.044 31.68 ;
      RECT 12.088 30.48 12.562 31.2 ;
      RECT 11.738 26.64 12.562 30.48 ;
      RECT 11.738 25.92 12.128 26.64 ;
      RECT 12.172 25.44 12.212 26.64 ;
      RECT 12.256 25.44 12.384 26.64 ;
      RECT 12.428 25.44 12.472 26.64 ;
      RECT 12.516 25.44 12.562 26.64 ;
      RECT 12.088 25.44 12.128 25.92 ;
      RECT 11.738 24.72 11.784 25.92 ;
      RECT 11.828 24.72 11.872 25.92 ;
      RECT 11.916 24.72 12.044 25.92 ;
      RECT 12.088 24.72 12.562 25.44 ;
      RECT 11.738 22.68 12.562 24.72 ;
      RECT 11.738 21.48 11.872 22.68 ;
      RECT 11.916 21.48 12.128 22.68 ;
      RECT 12.172 21.48 12.384 22.68 ;
      RECT 12.428 21.48 12.562 22.68 ;
      RECT 11.738 20.76 12.562 21.48 ;
      RECT 11.738 19.56 11.872 20.76 ;
      RECT 11.916 19.56 12.128 20.76 ;
      RECT 12.172 19.56 12.384 20.76 ;
      RECT 12.428 19.56 12.562 20.76 ;
      RECT 11.738 15.84 12.562 19.56 ;
      RECT 11.738 15.12 12.472 15.84 ;
      RECT 12.516 14.64 12.562 15.84 ;
      RECT 12.428 14.64 12.472 15.12 ;
      RECT 11.738 14.4 12.044 15.12 ;
      RECT 12.088 13.92 12.128 15.12 ;
      RECT 12.172 13.92 12.212 15.12 ;
      RECT 12.256 13.92 12.384 15.12 ;
      RECT 12.428 13.92 12.562 14.64 ;
      RECT 11.916 13.92 12.044 14.4 ;
      RECT 11.738 13.2 11.784 14.4 ;
      RECT 11.828 13.2 11.872 14.4 ;
      RECT 11.916 13.2 12.562 13.92 ;
      RECT 11.738 10.08 12.562 13.2 ;
      RECT 11.738 9.36 12.472 10.08 ;
      RECT 12.516 8.88 12.562 10.08 ;
      RECT 12.428 8.88 12.472 9.36 ;
      RECT 11.738 8.64 12.044 9.36 ;
      RECT 12.088 8.16 12.128 9.36 ;
      RECT 12.172 8.16 12.212 9.36 ;
      RECT 12.256 8.16 12.384 9.36 ;
      RECT 12.428 8.16 12.562 8.88 ;
      RECT 11.916 8.16 12.044 8.64 ;
      RECT 11.738 7.44 11.784 8.64 ;
      RECT 11.828 7.44 11.872 8.64 ;
      RECT 11.916 7.44 12.562 8.16 ;
      RECT 11.738 4.32 12.562 7.44 ;
      RECT 11.738 3.6 12.472 4.32 ;
      RECT 12.516 3.12 12.562 4.32 ;
      RECT 12.428 3.12 12.472 3.6 ;
      RECT 11.738 2.88 12.044 3.6 ;
      RECT 12.088 2.4 12.128 3.6 ;
      RECT 12.172 2.4 12.212 3.6 ;
      RECT 12.256 2.4 12.384 3.6 ;
      RECT 12.428 2.4 12.562 3.12 ;
      RECT 11.916 2.4 12.044 2.88 ;
      RECT 11.738 1.68 11.784 2.88 ;
      RECT 11.828 1.68 11.872 2.88 ;
      RECT 11.916 1.68 12.562 2.4 ;
      RECT 11.738 -0.12 12.562 1.68 ;
      RECT 10.838 37.44 11.662 41.4 ;
      RECT 10.838 36.72 11.572 37.44 ;
      RECT 11.616 36.24 11.662 37.44 ;
      RECT 11.528 36.24 11.572 36.72 ;
      RECT 10.838 35.52 11.144 36.72 ;
      RECT 11.188 35.52 11.228 36.72 ;
      RECT 11.272 35.52 11.312 36.72 ;
      RECT 11.356 35.52 11.484 36.72 ;
      RECT 11.528 35.52 11.662 36.24 ;
      RECT 10.838 31.68 11.662 35.52 ;
      RECT 10.838 30.96 11.572 31.68 ;
      RECT 11.616 30.48 11.662 31.68 ;
      RECT 11.528 30.48 11.572 30.96 ;
      RECT 10.838 29.76 11.144 30.96 ;
      RECT 11.188 29.76 11.228 30.96 ;
      RECT 11.272 29.76 11.312 30.96 ;
      RECT 11.356 29.76 11.484 30.96 ;
      RECT 11.528 29.76 11.662 30.48 ;
      RECT 10.838 25.92 11.662 29.76 ;
      RECT 10.838 25.2 11.572 25.92 ;
      RECT 11.616 24.72 11.662 25.92 ;
      RECT 11.528 24.72 11.572 25.2 ;
      RECT 10.838 24 11.144 25.2 ;
      RECT 11.188 24 11.228 25.2 ;
      RECT 11.272 24 11.312 25.2 ;
      RECT 11.356 24 11.484 25.2 ;
      RECT 11.528 24 11.662 24.72 ;
      RECT 10.838 22.68 11.662 24 ;
      RECT 10.838 21.48 10.884 22.68 ;
      RECT 10.928 21.48 11.144 22.68 ;
      RECT 11.188 21.48 11.312 22.68 ;
      RECT 11.356 21.48 11.572 22.68 ;
      RECT 11.616 21.48 11.662 22.68 ;
      RECT 10.838 20.76 11.662 21.48 ;
      RECT 10.838 19.56 10.884 20.76 ;
      RECT 10.928 19.56 11.144 20.76 ;
      RECT 11.188 19.56 11.312 20.76 ;
      RECT 11.356 19.56 11.572 20.76 ;
      RECT 11.616 19.56 11.662 20.76 ;
      RECT 10.838 14.4 11.662 19.56 ;
      RECT 10.838 13.68 11.484 14.4 ;
      RECT 11.528 13.2 11.572 14.4 ;
      RECT 11.616 13.2 11.662 14.4 ;
      RECT 11.272 13.2 11.484 13.68 ;
      RECT 10.838 12.48 10.884 13.68 ;
      RECT 10.928 12.48 10.972 13.68 ;
      RECT 11.016 12.48 11.144 13.68 ;
      RECT 11.188 12.48 11.228 13.68 ;
      RECT 11.272 12.48 11.662 13.2 ;
      RECT 10.838 8.64 11.662 12.48 ;
      RECT 10.838 7.92 11.484 8.64 ;
      RECT 11.528 7.44 11.572 8.64 ;
      RECT 11.616 7.44 11.662 8.64 ;
      RECT 11.272 7.44 11.484 7.92 ;
      RECT 10.838 6.72 10.884 7.92 ;
      RECT 10.928 6.72 10.972 7.92 ;
      RECT 11.016 6.72 11.144 7.92 ;
      RECT 11.188 6.72 11.228 7.92 ;
      RECT 11.272 6.72 11.662 7.44 ;
      RECT 10.838 2.88 11.662 6.72 ;
      RECT 10.838 2.16 11.484 2.88 ;
      RECT 11.528 1.68 11.572 2.88 ;
      RECT 11.616 1.68 11.662 2.88 ;
      RECT 11.356 1.68 11.484 2.16 ;
      RECT 10.838 0.96 10.972 2.16 ;
      RECT 11.016 0.96 11.144 2.16 ;
      RECT 11.188 0.96 11.228 2.16 ;
      RECT 11.272 0.96 11.312 2.16 ;
      RECT 11.356 0.96 11.662 1.68 ;
      RECT 10.838 -0.12 11.662 0.96 ;
      RECT 9.938 36 10.762 41.4 ;
      RECT 9.938 34.8 10.072 36 ;
      RECT 10.116 34.8 10.244 36 ;
      RECT 10.288 34.8 10.328 36 ;
      RECT 10.372 34.8 10.412 36 ;
      RECT 10.456 34.8 10.762 36 ;
      RECT 9.938 30.24 10.762 34.8 ;
      RECT 9.938 29.04 10.072 30.24 ;
      RECT 10.116 29.04 10.244 30.24 ;
      RECT 10.288 29.04 10.328 30.24 ;
      RECT 10.372 29.04 10.412 30.24 ;
      RECT 10.456 29.04 10.762 30.24 ;
      RECT 9.938 24.48 10.762 29.04 ;
      RECT 9.938 23.28 10.244 24.48 ;
      RECT 10.288 23.28 10.328 24.48 ;
      RECT 10.372 23.28 10.412 24.48 ;
      RECT 10.456 23.28 10.672 24.48 ;
      RECT 10.716 23.28 10.762 24.48 ;
      RECT 9.938 22.68 10.762 23.28 ;
      RECT 9.938 21.48 9.984 22.68 ;
      RECT 10.028 21.48 10.584 22.68 ;
      RECT 10.628 21.48 10.762 22.68 ;
      RECT 9.938 20.76 10.762 21.48 ;
      RECT 9.938 19.56 9.984 20.76 ;
      RECT 10.028 19.56 10.584 20.76 ;
      RECT 10.628 19.56 10.762 20.76 ;
      RECT 9.938 18.72 10.762 19.56 ;
      RECT 9.938 17.52 10.072 18.72 ;
      RECT 10.116 17.52 10.244 18.72 ;
      RECT 10.288 17.52 10.328 18.72 ;
      RECT 10.372 17.52 10.762 18.72 ;
      RECT 9.938 12.96 10.762 17.52 ;
      RECT 9.938 11.76 10.072 12.96 ;
      RECT 10.116 11.76 10.244 12.96 ;
      RECT 10.288 11.76 10.328 12.96 ;
      RECT 10.372 11.76 10.762 12.96 ;
      RECT 9.938 7.2 10.762 11.76 ;
      RECT 9.938 6 10.072 7.2 ;
      RECT 10.116 6 10.244 7.2 ;
      RECT 10.288 6 10.328 7.2 ;
      RECT 10.372 6 10.762 7.2 ;
      RECT 9.938 1.44 10.762 6 ;
      RECT 9.938 0.24 9.984 1.44 ;
      RECT 10.028 0.24 10.072 1.44 ;
      RECT 10.116 0.24 10.244 1.44 ;
      RECT 10.288 0.24 10.328 1.44 ;
      RECT 10.372 0.24 10.762 1.44 ;
      RECT 9.938 -0.12 10.762 0.24 ;
      RECT 9.038 -0.12 9.862 41.4 ;
      RECT 8.138 -0.12 8.962 41.4 ;
      RECT 7.238 -0.12 8.062 41.4 ;
      RECT 6.338 -0.12 7.162 41.4 ;
      RECT 5.438 -0.12 6.262 41.4 ;
      RECT 4.538 -0.12 5.362 41.4 ;
      RECT 3.638 -0.12 4.462 41.4 ;
      RECT 2.738 -0.12 3.562 41.4 ;
      RECT 1.838 -0.12 2.662 41.4 ;
      RECT 0.938 -0.12 1.762 41.4 ;
      RECT -0.04 41.34 0.862 41.4 ;
      RECT -0.092 -0.06 0.862 41.34 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 33.458 0 34.12 41.28 ;
      RECT 32.558 0 33.142 41.28 ;
      RECT 31.658 0 32.242 41.28 ;
      RECT 30.758 0 31.342 41.28 ;
      RECT 29.858 0 30.442 41.28 ;
      RECT 28.958 0 29.542 41.28 ;
      RECT 28.058 0 28.642 41.28 ;
      RECT 27.158 0 27.742 41.28 ;
      RECT 26.258 0 26.842 41.28 ;
      RECT 25.358 0 25.942 41.28 ;
      RECT 24.458 0 25.042 41.28 ;
      RECT 23.558 0 24.142 41.28 ;
      RECT 22.658 0 23.242 41.28 ;
      RECT 21.758 0 22.342 41.28 ;
      RECT 20.858 0 21.442 41.28 ;
      RECT 19.958 0 20.542 41.28 ;
      RECT 19.058 0 19.642 41.28 ;
      RECT 18.158 0 18.742 41.28 ;
      RECT 17.258 0 17.842 41.28 ;
      RECT 16.358 0 16.942 41.28 ;
      RECT 15.458 0 16.042 41.28 ;
      RECT 14.558 41.16 15.142 41.28 ;
      RECT 14.736 39.72 15.142 41.16 ;
      RECT 14.558 35.4 15.142 39.72 ;
      RECT 14.736 33.96 15.142 35.4 ;
      RECT 14.558 29.64 15.142 33.96 ;
      RECT 14.736 28.2 15.142 29.64 ;
      RECT 14.558 18.84 15.142 28.2 ;
      RECT 14.736 17.4 15.142 18.84 ;
      RECT 14.648 16.68 15.142 17.4 ;
      RECT 14.558 13.08 15.142 16.68 ;
      RECT 14.736 11.64 15.142 13.08 ;
      RECT 14.648 10.92 15.142 11.64 ;
      RECT 14.558 7.32 15.142 10.92 ;
      RECT 14.736 5.88 15.142 7.32 ;
      RECT 14.648 5.16 15.142 5.88 ;
      RECT 14.558 0 15.142 5.16 ;
      RECT 13.658 41.16 14.242 41.28 ;
      RECT 13.658 40.44 14.064 41.16 ;
      RECT 12.758 39.72 13.342 41.28 ;
      RECT 12.758 39 12.992 39.72 ;
      RECT 11.858 38.28 12.442 41.28 ;
      RECT 11.858 37.56 12.008 38.28 ;
      RECT 10.958 37.56 11.542 41.28 ;
      RECT 10.958 36.84 11.452 37.56 ;
      RECT 10.958 35.4 11.024 36.84 ;
      RECT 10.958 31.8 11.542 35.4 ;
      RECT 10.958 31.08 11.452 31.8 ;
      RECT 10.958 29.64 11.024 31.08 ;
      RECT 10.958 26.04 11.542 29.64 ;
      RECT 10.958 25.32 11.452 26.04 ;
      RECT 10.958 23.88 11.024 25.32 ;
      RECT 10.958 22.8 11.542 23.88 ;
      RECT 10.058 36.12 10.642 41.28 ;
      RECT 10.576 34.68 10.642 36.12 ;
      RECT 10.058 30.36 10.642 34.68 ;
      RECT 10.576 28.92 10.642 30.36 ;
      RECT 10.058 24.6 10.642 28.92 ;
      RECT 10.058 23.16 10.124 24.6 ;
      RECT 10.058 22.8 10.642 23.16 ;
      RECT 10.148 21.36 10.464 22.8 ;
      RECT 10.058 20.88 10.642 21.36 ;
      RECT 10.148 19.44 10.464 20.88 ;
      RECT 10.058 18.84 10.642 19.44 ;
      RECT 10.492 17.4 10.642 18.84 ;
      RECT 10.058 13.08 10.642 17.4 ;
      RECT 10.492 11.64 10.642 13.08 ;
      RECT 10.058 7.32 10.642 11.64 ;
      RECT 10.492 5.88 10.642 7.32 ;
      RECT 10.058 1.56 10.642 5.88 ;
      RECT 10.492 0.12 10.642 1.56 ;
      RECT 10.058 0 10.642 0.12 ;
      RECT 9.158 0 9.742 41.28 ;
      RECT 8.258 0 8.842 41.28 ;
      RECT 7.358 0 7.942 41.28 ;
      RECT 6.458 0 7.042 41.28 ;
      RECT 5.558 0 6.142 41.28 ;
      RECT 4.658 0 5.242 41.28 ;
      RECT 3.758 0 4.342 41.28 ;
      RECT 2.858 0 3.442 41.28 ;
      RECT 1.958 0 2.542 41.28 ;
      RECT 1.058 0 1.642 41.28 ;
      RECT 0.08 0 0.742 41.28 ;
      RECT 14.176 39 14.242 39.72 ;
      RECT 13.748 38.28 14.242 39 ;
      RECT 13.658 35.4 14.242 38.28 ;
      RECT 13.658 34.68 14.064 35.4 ;
      RECT 13.192 37.56 13.342 38.28 ;
      RECT 12.758 33.96 13.342 37.56 ;
      RECT 12.758 33.24 12.992 33.96 ;
      RECT 12.208 36.12 12.442 36.84 ;
      RECT 11.858 32.52 12.442 36.12 ;
      RECT 11.858 31.8 12.008 32.52 ;
      RECT 14.176 33.24 14.242 33.96 ;
      RECT 13.748 32.52 14.242 33.24 ;
      RECT 13.658 29.64 14.242 32.52 ;
      RECT 13.658 28.92 14.064 29.64 ;
      RECT 13.192 31.8 13.342 32.52 ;
      RECT 12.758 28.2 13.342 31.8 ;
      RECT 12.758 27.48 12.992 28.2 ;
      RECT 12.208 30.36 12.442 31.08 ;
      RECT 11.858 26.76 12.442 30.36 ;
      RECT 11.858 26.04 12.008 26.76 ;
      RECT 14.176 27.48 14.242 28.2 ;
      RECT 13.748 26.76 14.242 27.48 ;
      RECT 13.658 20.88 14.242 26.76 ;
      RECT 13.836 19.44 14.242 20.88 ;
      RECT 13.658 18.12 14.242 19.44 ;
      RECT 13.658 17.4 13.892 18.12 ;
      RECT 13.192 26.04 13.342 26.76 ;
      RECT 12.758 22.8 13.342 26.04 ;
      RECT 12.208 24.6 12.442 25.32 ;
      RECT 11.858 22.8 12.442 24.6 ;
      RECT 12.758 20.88 13.342 21.36 ;
      RECT 11.858 20.88 12.442 21.36 ;
      RECT 10.958 20.88 11.542 21.36 ;
      RECT 12.758 16.68 13.342 19.44 ;
      RECT 12.758 15.96 12.908 16.68 ;
      RECT 11.858 15.96 12.442 19.44 ;
      RECT 11.858 15.24 12.352 15.96 ;
      RECT 11.858 14.52 11.924 15.24 ;
      RECT 10.958 14.52 11.542 19.44 ;
      RECT 10.958 13.8 11.364 14.52 ;
      RECT 14.092 15.96 14.242 16.68 ;
      RECT 13.658 12.36 14.242 15.96 ;
      RECT 13.658 11.64 13.892 12.36 ;
      RECT 13.108 14.52 13.342 15.24 ;
      RECT 12.758 10.92 13.342 14.52 ;
      RECT 12.758 10.2 12.908 10.92 ;
      RECT 12.036 13.08 12.442 13.8 ;
      RECT 11.858 10.2 12.442 13.08 ;
      RECT 11.858 9.48 12.352 10.2 ;
      RECT 11.858 8.76 11.924 9.48 ;
      RECT 11.392 12.36 11.542 13.08 ;
      RECT 10.958 8.76 11.542 12.36 ;
      RECT 10.958 8.04 11.364 8.76 ;
      RECT 14.092 10.2 14.242 10.92 ;
      RECT 13.658 6.6 14.242 10.2 ;
      RECT 13.658 5.88 13.892 6.6 ;
      RECT 13.108 8.76 13.342 9.48 ;
      RECT 12.758 5.16 13.342 8.76 ;
      RECT 12.758 4.44 12.908 5.16 ;
      RECT 12.036 7.32 12.442 8.04 ;
      RECT 11.858 4.44 12.442 7.32 ;
      RECT 11.858 3.72 12.352 4.44 ;
      RECT 11.858 3 11.924 3.72 ;
      RECT 11.392 6.6 11.542 7.32 ;
      RECT 10.958 3 11.542 6.6 ;
      RECT 10.958 2.28 11.364 3 ;
      RECT 14.092 4.44 14.242 5.16 ;
      RECT 13.658 0 14.242 4.44 ;
      RECT 13.108 3 13.342 3.72 ;
      RECT 12.758 0 13.342 3 ;
      RECT 12.036 1.56 12.442 2.28 ;
      RECT 11.858 0 12.442 1.56 ;
      RECT 11.476 0.84 11.542 1.56 ;
      RECT 10.958 0 11.542 0.84 ;
    LAYER m0 ;
      RECT 0 0.002 34.2 41.278 ;
    LAYER m1 ;
      RECT 0 0 34.2 41.28 ;
    LAYER m2 ;
      RECT 0 0.015 34.2 41.265 ;
    LAYER m3 ;
      RECT 0.015 0 34.185 41.28 ;
    LAYER m4 ;
      RECT 0 0.02 34.2 41.26 ;
    LAYER m5 ;
      RECT 0.012 0 34.188 41.28 ;
    LAYER m6 ;
      RECT 0 0.012 34.2 41.268 ;
  END
  PROPERTY hpml_layer "7" ;
  PROPERTY heml_layer "7" ;
END arf096b192e1r1w0cbbeheaa4acw

END LIBRARY
