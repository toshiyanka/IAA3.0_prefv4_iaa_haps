module ctech_lib_inv (
   input logic a,
   output logic o1
);
   d04inn00ln0c5 ctech_lib_dcszo (.a(a), .o1(o1));
endmodule
