module ctech_lib_clk_firewall_ls_and (o, a, en);
   input logic a,en;
   output logic o;
   d04sca00ld0b0 ctech_lib_dcszo (.a(a),.o(o),.en(en));
endmodule
