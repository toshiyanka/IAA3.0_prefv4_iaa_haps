//-----------------------------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2015 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to the source code
// ("Material") are owned by Intel Corporation or its suppliers or licensors. Title to the Material
// remains with Intel Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its suppliers and licensors.
// The Material is protected by worldwide copyright and trade secret laws and treaty provisions.
// No part of the Material may be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual property right is
// granted to or conferred upon you by disclosure or delivery of the Materials, either expressly, by
// implication, inducement, estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//-----------------------------------------------------------------------------------------------------
//-- Test
//-----------------------------------------------------------------------------------------------------
`ifndef hqm_iosf_prim_mem_wr_badparity_seq__SV
`define hqm_iosf_prim_mem_wr_badparity_seq__SV

import IosfPkg::*;

//-------------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------------
class hqm_iosf_prim_mem_wr_badparity_seq extends IosfSendTxnSeq;

  `ovm_sequence_utils(hqm_iosf_prim_mem_wr_badparity_seq,IosfAgtSeqr)

  rand logic [63:0]     iosf_addr;
  rand Iosf::data_t     iosf_data[];
  rand logic [7:0]      iosf_sai;
  static logic [7:0]    iosf_tag = 0;


   rand bit m_driveBadCmdParity; ; // toggles cmd parity signal
   rand bit m_driveBadDataParity; //  toggles data[0] when set
   rand int unsigned m_driveBadDataParityCycle;// bad parity data cycle
   rand int unsigned m_driveBadDataParityPct; // more than one cycle


  constraint deflt { soft iosf_sai == 8'h03; }

  extern                function        new(string name = "hqm_iosf_prim_mem_wr_badparity_seq");
  extern virtual        task            body();

endclass : hqm_iosf_prim_mem_wr_badparity_seq

function hqm_iosf_prim_mem_wr_badparity_seq::new(string name = "hqm_iosf_prim_mem_wr_badparity_seq");
  super.new(name);
endfunction

//------------------
//-- body
//------------------
task hqm_iosf_prim_mem_wr_badparity_seq::body();
  IosfTxn               iosfTxn;
  Iosf::data_t          data_i[];

  iosfTxn = new("iosfTxn");

  data_i = iosf_data;

  iosfTxn.set_sequencer (get_sequencer());
  iosfTxn.cmd               = (iosf_addr[63:32] == 32'h0) ? Iosf::MWr32 : Iosf::MWr64;
  iosfTxn.reqChId           = 0;
  iosfTxn.trafficClass      = 0;
  iosfTxn.reqID             = 0;
  iosfTxn.reqType           = Iosf::getReqTypeFromCmd (iosfTxn.cmd);
  iosfTxn.procHint          = 0;
  iosfTxn.length            = data_i.size();
  iosfTxn.address           = iosf_addr;
  iosfTxn.byteEnWithData    = 0;
  iosfTxn.data              = data_i;
  iosfTxn.first_byte_en     = 4'hf;
  iosfTxn.last_byte_en      = (data_i.size() > 1) ? 4'hf : 4'h0;
  iosfTxn.reqLocked         = 0;  
  iosfTxn.compareType       = Iosf::CMP_EQ;
  iosfTxn.compareCompletion = 0;
  iosfTxn.waitForCompletion = 0;
  iosfTxn.pollingMode       = 0;
  iosfTxn.tag               = iosf_tag;
  iosfTxn.expectRsp         = 0;
  iosfTxn.driveBadCmdParity = m_driveBadCmdParity;
  iosfTxn.driveBadDataParity = m_driveBadDataParity;
  iosfTxn.driveBadDataParityCycle = m_driveBadDataParityCycle;
  iosfTxn.driveBadDataParityPct   = m_driveBadDataParityPct;
  iosfTxn.reqGap            =  0;
  iosfTxn.chain             =  1'b0;
  iosfTxn.sai               =  iosf_sai;

  iosf_tag++;

  `ovm_send (iosfTxn)

  ovm_report_info(get_full_name(), $psprintf("MWr64 Address=0x%x SAI=0x%02x Data=0x%08x",iosf_addr,iosf_sai,data_i[0]), OVM_LOW);

endtask : body  

`endif
