.DFX_NUM_OF_FEATURES_TO_SECURE         (DFXSECURE_DFX_NUM_OF_FEATURES_TO_SECURE),
.DFX_SECURE_WIDTH                      (DFXSECURE_DFX_SECURE_WIDTH),
.DFX_USE_SB_OVR                        (DFXSECURE_DFX_USE_SB_OVR),
.DFX_VISA_BLACK                        (DFXSECURE_DFX_VISA_BLACK),
.DFX_VISA_GREEN                        (DFXSECURE_DFX_VISA_GREEN),
.DFX_VISA_ORANGE                       (DFXSECURE_DFX_VISA_ORANGE),
.DFX_VISA_RED                          (DFXSECURE_DFX_VISA_RED),
.DFX_EARLYBOOT_FEATURE_ENABLE          (DFXSECURE_DFX_EARLYBOOT_FEATURE_ENABLE),
.DFX_SECURE_POLICY_MATRIX              (DFXSECURE_DFX_SECURE_POLICY_MATRIX)
