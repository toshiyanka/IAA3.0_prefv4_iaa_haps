VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf054b128e1r1w0cbbehraa4acw
  CLASS BLOCK ;
  FOREIGN arf054b128e1r1w0cbbehraa4acw ;
  ORIGIN 0 0 ;
  SIZE 23.4 BY 24.96 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 2.52 0.472 3.72 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 0.6 0.472 1.8 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 2.52 2.272 3.72 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 2.52 2.616 3.72 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 2.52 2.916 3.72 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.52 3.428 3.72 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 2.52 3.728 3.72 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 2.52 4.072 3.72 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 2.52 0.728 3.72 ;
    END
  END rdaddrp0[6]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 2.52 0.816 3.72 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 2.52 1.116 3.72 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 2.52 1.628 3.72 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 2.52 1.928 3.72 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 0.6 2.616 1.8 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.6 2.916 1.8 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.6 3.428 1.8 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.6 3.728 1.8 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 0.6 4.072 1.8 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 0.6 0.728 1.8 ;
    END
  END wraddrp0[5]
  PIN wraddrp0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 0.6 1.028 1.8 ;
    END
  END wraddrp0[6]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 0.6 0.816 1.8 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 0.6 1.116 1.8 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 4.08 2.528 5.28 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 7.68 2.272 8.88 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 7.68 2.616 8.88 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 8.4 2.528 9.6 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 8.4 2.828 9.6 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 9.12 2.272 10.32 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 9.12 2.616 10.32 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 9.84 2.528 11.04 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 9.84 2.828 11.04 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 10.56 2.272 11.76 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 10.56 2.616 11.76 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 4.08 2.828 5.28 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 11.28 2.528 12.48 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 11.28 2.828 12.48 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 12 2.272 13.2 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 12 2.616 13.2 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 12.72 2.528 13.92 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12.72 2.828 13.92 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 13.44 2.272 14.64 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 13.44 2.616 14.64 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 14.16 2.528 15.36 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 14.16 2.828 15.36 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 4.8 2.272 6 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 14.88 2.272 16.08 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 14.88 2.616 16.08 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 15.6 2.528 16.8 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 15.6 2.828 16.8 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 16.32 2.272 17.52 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 16.32 2.616 17.52 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 17.04 2.528 18.24 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 17.04 2.828 18.24 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 17.76 2.272 18.96 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 17.76 2.616 18.96 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 4.8 2.616 6 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 18.48 2.528 19.68 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 18.48 2.828 19.68 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 19.2 2.272 20.4 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.2 2.616 20.4 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 19.92 2.528 21.12 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 19.92 2.828 21.12 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 20.64 2.272 21.84 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 20.64 2.616 21.84 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 21.36 2.528 22.56 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 21.36 2.828 22.56 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 5.52 2.528 6.72 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 22.08 2.272 23.28 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 22.08 2.616 23.28 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 22.8 2.528 24 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 22.8 2.828 24 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 23.52 2.272 24.72 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 23.52 2.616 24.72 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.52 2.828 6.72 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 6.24 2.272 7.44 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 6.24 2.616 7.44 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6.96 2.528 8.16 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 6.96 2.828 8.16 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.6 1.928 1.8 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.6 2.272 1.8 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 0.6 1.628 1.8 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 4.08 4.328 5.28 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 7.68 4.072 8.88 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 7.68 3.428 8.88 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 8.4 4.328 9.6 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.4 3.516 9.6 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 9.12 4.072 10.32 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9.12 3.428 10.32 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.84 4.328 11.04 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 9.84 3.516 11.04 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 10.56 4.072 11.76 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 10.56 3.428 11.76 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 4.08 3.516 5.28 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 11.28 4.328 12.48 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.28 3.516 12.48 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 12 4.072 13.2 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 12 3.428 13.2 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 12.72 4.328 13.92 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.72 3.516 13.92 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 13.44 4.072 14.64 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 13.44 3.428 14.64 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 14.16 4.328 15.36 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 14.16 3.516 15.36 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 4.8 4.072 6 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 14.88 4.072 16.08 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 14.88 3.428 16.08 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 15.6 4.328 16.8 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 15.6 3.516 16.8 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 16.32 4.072 17.52 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.32 3.428 17.52 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 17.04 4.328 18.24 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 17.04 3.516 18.24 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 17.76 4.072 18.96 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 17.76 3.428 18.96 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.8 3.428 6 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 18.48 4.328 19.68 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 18.48 3.516 19.68 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 19.2 4.072 20.4 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 19.2 3.428 20.4 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 19.92 4.328 21.12 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 19.92 3.516 21.12 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 20.64 4.072 21.84 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.64 3.428 21.84 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 21.36 4.328 22.56 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 21.36 3.516 22.56 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 5.52 4.328 6.72 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 22.08 4.072 23.28 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 22.08 3.428 23.28 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 22.8 4.328 24 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 22.8 3.516 24 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 23.52 4.072 24.72 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 23.52 3.428 24.72 ;
    END
  END rddatap0[55]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.52 3.516 6.72 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.24 4.072 7.44 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6.24 3.428 7.44 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6.96 4.328 8.16 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 6.96 3.516 8.16 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 24.9 ;
        RECT 2.662 0.06 2.738 24.9 ;
        RECT 4.462 0.06 4.538 24.9 ;
        RECT 6.262 0.06 6.338 24.9 ;
        RECT 8.062 0.06 8.138 24.9 ;
        RECT 9.862 0.06 9.938 24.9 ;
        RECT 11.662 0.06 11.738 24.9 ;
        RECT 13.462 0.06 13.538 24.9 ;
        RECT 15.262 0.06 15.338 24.9 ;
        RECT 17.062 0.06 17.138 24.9 ;
        RECT 18.862 0.06 18.938 24.9 ;
        RECT 20.662 0.06 20.738 24.9 ;
        RECT 22.462 0.06 22.538 24.9 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 24.9 ;
        RECT 3.562 0.06 3.638 24.9 ;
        RECT 5.362 0.06 5.438 24.9 ;
        RECT 7.162 0.06 7.238 24.9 ;
        RECT 8.962 0.06 9.038 24.9 ;
        RECT 10.762 0.06 10.838 24.9 ;
        RECT 12.562 0.06 12.638 24.9 ;
        RECT 14.362 0.06 14.438 24.9 ;
        RECT 16.162 0.06 16.238 24.9 ;
        RECT 17.962 0.06 18.038 24.9 ;
        RECT 19.762 0.06 19.838 24.9 ;
        RECT 21.562 0.06 21.638 24.9 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 23.416 24.974 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 23.42 24.98 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 23.4705 24.998 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 23.435 25.03 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 23.47 24.998 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 23.459 25.05 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 23.49 25.022 ;
    LAYER m7 SPACING 0 ;
      RECT 22.538 25.02 23.44 25.08 ;
      RECT 22.538 -0.06 23.492 25.02 ;
      RECT 22.538 -0.12 23.44 -0.06 ;
      RECT 21.638 -0.12 22.462 25.08 ;
      RECT 20.738 -0.12 21.562 25.08 ;
      RECT 19.838 -0.12 20.662 25.08 ;
      RECT 18.938 -0.12 19.762 25.08 ;
      RECT 18.038 -0.12 18.862 25.08 ;
      RECT 17.138 -0.12 17.962 25.08 ;
      RECT 16.238 -0.12 17.062 25.08 ;
      RECT 15.338 -0.12 16.162 25.08 ;
      RECT 14.438 -0.12 15.262 25.08 ;
      RECT 13.538 -0.12 14.362 25.08 ;
      RECT 12.638 -0.12 13.462 25.08 ;
      RECT 11.738 -0.12 12.562 25.08 ;
      RECT 10.838 -0.12 11.662 25.08 ;
      RECT 9.938 -0.12 10.762 25.08 ;
      RECT 9.038 -0.12 9.862 25.08 ;
      RECT 8.138 -0.12 8.962 25.08 ;
      RECT 7.238 -0.12 8.062 25.08 ;
      RECT 6.338 -0.12 7.162 25.08 ;
      RECT 5.438 -0.12 6.262 25.08 ;
      RECT 4.538 -0.12 5.362 25.08 ;
      RECT 3.638 24.72 4.462 25.08 ;
      RECT 4.072 24 4.462 24.72 ;
      RECT 3.638 23.52 4.028 24.72 ;
      RECT 4.072 23.52 4.284 24 ;
      RECT 3.638 23.28 4.284 23.52 ;
      RECT 4.328 22.8 4.462 24 ;
      RECT 4.072 22.8 4.284 23.28 ;
      RECT 4.072 22.56 4.462 22.8 ;
      RECT 3.638 22.08 4.028 23.28 ;
      RECT 4.072 22.08 4.284 22.56 ;
      RECT 3.638 21.84 4.284 22.08 ;
      RECT 4.328 21.36 4.462 22.56 ;
      RECT 4.072 21.36 4.284 21.84 ;
      RECT 4.072 21.12 4.462 21.36 ;
      RECT 3.638 20.64 4.028 21.84 ;
      RECT 4.072 20.64 4.284 21.12 ;
      RECT 3.638 20.4 4.284 20.64 ;
      RECT 4.328 19.92 4.462 21.12 ;
      RECT 4.072 19.92 4.284 20.4 ;
      RECT 4.072 19.68 4.462 19.92 ;
      RECT 3.638 19.2 4.028 20.4 ;
      RECT 4.072 19.2 4.284 19.68 ;
      RECT 3.638 18.96 4.284 19.2 ;
      RECT 4.328 18.48 4.462 19.68 ;
      RECT 4.072 18.48 4.284 18.96 ;
      RECT 4.072 18.24 4.462 18.48 ;
      RECT 3.638 17.76 4.028 18.96 ;
      RECT 4.072 17.76 4.284 18.24 ;
      RECT 3.638 17.52 4.284 17.76 ;
      RECT 4.328 17.04 4.462 18.24 ;
      RECT 4.072 17.04 4.284 17.52 ;
      RECT 4.072 16.8 4.462 17.04 ;
      RECT 3.638 16.32 4.028 17.52 ;
      RECT 4.072 16.32 4.284 16.8 ;
      RECT 3.638 16.08 4.284 16.32 ;
      RECT 4.328 15.6 4.462 16.8 ;
      RECT 4.072 15.6 4.284 16.08 ;
      RECT 4.072 15.36 4.462 15.6 ;
      RECT 3.638 14.88 4.028 16.08 ;
      RECT 4.072 14.88 4.284 15.36 ;
      RECT 3.638 14.64 4.284 14.88 ;
      RECT 4.328 14.16 4.462 15.36 ;
      RECT 4.072 14.16 4.284 14.64 ;
      RECT 4.072 13.92 4.462 14.16 ;
      RECT 3.638 13.44 4.028 14.64 ;
      RECT 4.072 13.44 4.284 13.92 ;
      RECT 3.638 13.2 4.284 13.44 ;
      RECT 4.328 12.72 4.462 13.92 ;
      RECT 4.072 12.72 4.284 13.2 ;
      RECT 4.072 12.48 4.462 12.72 ;
      RECT 3.638 12 4.028 13.2 ;
      RECT 4.072 12 4.284 12.48 ;
      RECT 3.638 11.76 4.284 12 ;
      RECT 4.328 11.28 4.462 12.48 ;
      RECT 4.072 11.28 4.284 11.76 ;
      RECT 4.072 11.04 4.462 11.28 ;
      RECT 3.638 10.56 4.028 11.76 ;
      RECT 4.072 10.56 4.284 11.04 ;
      RECT 3.638 10.32 4.284 10.56 ;
      RECT 4.328 9.84 4.462 11.04 ;
      RECT 4.072 9.84 4.284 10.32 ;
      RECT 4.072 9.6 4.462 9.84 ;
      RECT 3.638 9.12 4.028 10.32 ;
      RECT 4.072 9.12 4.284 9.6 ;
      RECT 3.638 8.88 4.284 9.12 ;
      RECT 4.328 8.4 4.462 9.6 ;
      RECT 4.072 8.4 4.284 8.88 ;
      RECT 4.072 8.16 4.462 8.4 ;
      RECT 3.638 7.68 4.028 8.88 ;
      RECT 4.072 7.68 4.284 8.16 ;
      RECT 3.638 7.44 4.284 7.68 ;
      RECT 4.328 6.96 4.462 8.16 ;
      RECT 4.072 6.96 4.284 7.44 ;
      RECT 4.072 6.72 4.462 6.96 ;
      RECT 3.638 6.24 4.028 7.44 ;
      RECT 4.072 6.24 4.284 6.72 ;
      RECT 3.638 6 4.284 6.24 ;
      RECT 4.328 5.52 4.462 6.72 ;
      RECT 4.072 5.52 4.284 6 ;
      RECT 4.072 5.28 4.462 5.52 ;
      RECT 3.638 4.8 4.028 6 ;
      RECT 4.072 4.8 4.284 5.28 ;
      RECT 4.328 4.08 4.462 5.28 ;
      RECT 3.638 4.08 4.284 4.8 ;
      RECT 3.638 3.72 4.462 4.08 ;
      RECT 3.638 2.52 3.684 3.72 ;
      RECT 3.728 2.52 4.028 3.72 ;
      RECT 4.072 2.52 4.462 3.72 ;
      RECT 3.638 1.8 4.462 2.52 ;
      RECT 3.638 0.6 3.684 1.8 ;
      RECT 3.728 0.6 4.028 1.8 ;
      RECT 4.072 0.6 4.462 1.8 ;
      RECT 3.638 -0.12 4.462 0.6 ;
      RECT 2.738 24.72 3.562 25.08 ;
      RECT 2.738 24 3.384 24.72 ;
      RECT 3.428 24 3.562 24.72 ;
      RECT 2.828 23.52 3.384 24 ;
      RECT 3.428 23.52 3.472 24 ;
      RECT 2.828 23.28 3.472 23.52 ;
      RECT 2.738 22.8 2.784 24 ;
      RECT 3.516 22.8 3.562 24 ;
      RECT 2.828 22.8 3.384 23.28 ;
      RECT 3.428 22.8 3.472 23.28 ;
      RECT 2.738 22.56 3.384 22.8 ;
      RECT 3.428 22.56 3.562 22.8 ;
      RECT 2.828 22.08 3.384 22.56 ;
      RECT 3.428 22.08 3.472 22.56 ;
      RECT 2.828 21.84 3.472 22.08 ;
      RECT 2.738 21.36 2.784 22.56 ;
      RECT 3.516 21.36 3.562 22.56 ;
      RECT 2.828 21.36 3.384 21.84 ;
      RECT 3.428 21.36 3.472 21.84 ;
      RECT 2.738 21.12 3.384 21.36 ;
      RECT 3.428 21.12 3.562 21.36 ;
      RECT 2.828 20.64 3.384 21.12 ;
      RECT 3.428 20.64 3.472 21.12 ;
      RECT 2.828 20.4 3.472 20.64 ;
      RECT 2.738 19.92 2.784 21.12 ;
      RECT 3.516 19.92 3.562 21.12 ;
      RECT 2.828 19.92 3.384 20.4 ;
      RECT 3.428 19.92 3.472 20.4 ;
      RECT 2.738 19.68 3.384 19.92 ;
      RECT 3.428 19.68 3.562 19.92 ;
      RECT 2.828 19.2 3.384 19.68 ;
      RECT 3.428 19.2 3.472 19.68 ;
      RECT 2.828 18.96 3.472 19.2 ;
      RECT 2.738 18.48 2.784 19.68 ;
      RECT 3.516 18.48 3.562 19.68 ;
      RECT 2.828 18.48 3.384 18.96 ;
      RECT 3.428 18.48 3.472 18.96 ;
      RECT 2.738 18.24 3.384 18.48 ;
      RECT 3.428 18.24 3.562 18.48 ;
      RECT 2.828 17.76 3.384 18.24 ;
      RECT 3.428 17.76 3.472 18.24 ;
      RECT 2.828 17.52 3.472 17.76 ;
      RECT 2.738 17.04 2.784 18.24 ;
      RECT 3.516 17.04 3.562 18.24 ;
      RECT 2.828 17.04 3.384 17.52 ;
      RECT 3.428 17.04 3.472 17.52 ;
      RECT 2.738 16.8 3.384 17.04 ;
      RECT 3.428 16.8 3.562 17.04 ;
      RECT 2.828 16.32 3.384 16.8 ;
      RECT 3.428 16.32 3.472 16.8 ;
      RECT 2.828 16.08 3.472 16.32 ;
      RECT 2.738 15.6 2.784 16.8 ;
      RECT 3.516 15.6 3.562 16.8 ;
      RECT 2.828 15.6 3.384 16.08 ;
      RECT 3.428 15.6 3.472 16.08 ;
      RECT 2.738 15.36 3.384 15.6 ;
      RECT 3.428 15.36 3.562 15.6 ;
      RECT 2.828 14.88 3.384 15.36 ;
      RECT 3.428 14.88 3.472 15.36 ;
      RECT 2.828 14.64 3.472 14.88 ;
      RECT 2.738 14.16 2.784 15.36 ;
      RECT 3.516 14.16 3.562 15.36 ;
      RECT 2.828 14.16 3.384 14.64 ;
      RECT 3.428 14.16 3.472 14.64 ;
      RECT 2.738 13.92 3.384 14.16 ;
      RECT 3.428 13.92 3.562 14.16 ;
      RECT 2.828 13.44 3.384 13.92 ;
      RECT 3.428 13.44 3.472 13.92 ;
      RECT 2.828 13.2 3.472 13.44 ;
      RECT 2.738 12.72 2.784 13.92 ;
      RECT 3.516 12.72 3.562 13.92 ;
      RECT 2.828 12.72 3.384 13.2 ;
      RECT 3.428 12.72 3.472 13.2 ;
      RECT 2.738 12.48 3.384 12.72 ;
      RECT 3.428 12.48 3.562 12.72 ;
      RECT 2.828 12 3.384 12.48 ;
      RECT 3.428 12 3.472 12.48 ;
      RECT 2.828 11.76 3.472 12 ;
      RECT 2.738 11.28 2.784 12.48 ;
      RECT 3.516 11.28 3.562 12.48 ;
      RECT 2.828 11.28 3.384 11.76 ;
      RECT 3.428 11.28 3.472 11.76 ;
      RECT 2.738 11.04 3.384 11.28 ;
      RECT 3.428 11.04 3.562 11.28 ;
      RECT 2.828 10.56 3.384 11.04 ;
      RECT 3.428 10.56 3.472 11.04 ;
      RECT 2.828 10.32 3.472 10.56 ;
      RECT 2.738 9.84 2.784 11.04 ;
      RECT 3.516 9.84 3.562 11.04 ;
      RECT 2.828 9.84 3.384 10.32 ;
      RECT 3.428 9.84 3.472 10.32 ;
      RECT 2.738 9.6 3.384 9.84 ;
      RECT 3.428 9.6 3.562 9.84 ;
      RECT 2.828 9.12 3.384 9.6 ;
      RECT 3.428 9.12 3.472 9.6 ;
      RECT 2.828 8.88 3.472 9.12 ;
      RECT 2.738 8.4 2.784 9.6 ;
      RECT 3.516 8.4 3.562 9.6 ;
      RECT 2.828 8.4 3.384 8.88 ;
      RECT 3.428 8.4 3.472 8.88 ;
      RECT 2.738 8.16 3.384 8.4 ;
      RECT 3.428 8.16 3.562 8.4 ;
      RECT 2.828 7.68 3.384 8.16 ;
      RECT 3.428 7.68 3.472 8.16 ;
      RECT 2.828 7.44 3.472 7.68 ;
      RECT 2.738 6.96 2.784 8.16 ;
      RECT 3.516 6.96 3.562 8.16 ;
      RECT 2.828 6.96 3.384 7.44 ;
      RECT 3.428 6.96 3.472 7.44 ;
      RECT 2.738 6.72 3.384 6.96 ;
      RECT 3.428 6.72 3.562 6.96 ;
      RECT 2.828 6.24 3.384 6.72 ;
      RECT 3.428 6.24 3.472 6.72 ;
      RECT 2.828 6 3.472 6.24 ;
      RECT 2.738 5.52 2.784 6.72 ;
      RECT 3.516 5.52 3.562 6.72 ;
      RECT 2.828 5.52 3.384 6 ;
      RECT 3.428 5.52 3.472 6 ;
      RECT 2.738 5.28 3.384 5.52 ;
      RECT 3.428 5.28 3.562 5.52 ;
      RECT 2.828 4.8 3.384 5.28 ;
      RECT 3.428 4.8 3.472 5.28 ;
      RECT 2.738 4.08 2.784 5.28 ;
      RECT 3.516 4.08 3.562 5.28 ;
      RECT 2.828 4.08 3.472 4.8 ;
      RECT 2.738 3.72 3.562 4.08 ;
      RECT 2.738 2.52 2.872 3.72 ;
      RECT 2.916 2.52 3.384 3.72 ;
      RECT 3.428 2.52 3.562 3.72 ;
      RECT 2.738 1.8 3.562 2.52 ;
      RECT 2.738 0.6 2.872 1.8 ;
      RECT 2.916 0.6 3.384 1.8 ;
      RECT 3.428 0.6 3.562 1.8 ;
      RECT 2.738 -0.12 3.562 0.6 ;
      RECT 1.838 24.72 2.662 25.08 ;
      RECT 2.272 24 2.572 24.72 ;
      RECT 1.838 23.52 2.228 24.72 ;
      RECT 2.616 23.52 2.662 24.72 ;
      RECT 2.272 23.52 2.484 24 ;
      RECT 2.528 23.52 2.572 24 ;
      RECT 1.838 23.28 2.484 23.52 ;
      RECT 2.528 23.28 2.662 23.52 ;
      RECT 2.272 22.8 2.484 23.28 ;
      RECT 2.528 22.8 2.572 23.28 ;
      RECT 2.272 22.56 2.572 22.8 ;
      RECT 1.838 22.08 2.228 23.28 ;
      RECT 2.616 22.08 2.662 23.28 ;
      RECT 2.272 22.08 2.484 22.56 ;
      RECT 2.528 22.08 2.572 22.56 ;
      RECT 1.838 21.84 2.484 22.08 ;
      RECT 2.528 21.84 2.662 22.08 ;
      RECT 2.272 21.36 2.484 21.84 ;
      RECT 2.528 21.36 2.572 21.84 ;
      RECT 2.272 21.12 2.572 21.36 ;
      RECT 1.838 20.64 2.228 21.84 ;
      RECT 2.616 20.64 2.662 21.84 ;
      RECT 2.272 20.64 2.484 21.12 ;
      RECT 2.528 20.64 2.572 21.12 ;
      RECT 1.838 20.4 2.484 20.64 ;
      RECT 2.528 20.4 2.662 20.64 ;
      RECT 2.272 19.92 2.484 20.4 ;
      RECT 2.528 19.92 2.572 20.4 ;
      RECT 2.272 19.68 2.572 19.92 ;
      RECT 1.838 19.2 2.228 20.4 ;
      RECT 2.616 19.2 2.662 20.4 ;
      RECT 2.272 19.2 2.484 19.68 ;
      RECT 2.528 19.2 2.572 19.68 ;
      RECT 1.838 18.96 2.484 19.2 ;
      RECT 2.528 18.96 2.662 19.2 ;
      RECT 2.272 18.48 2.484 18.96 ;
      RECT 2.528 18.48 2.572 18.96 ;
      RECT 2.272 18.24 2.572 18.48 ;
      RECT 1.838 17.76 2.228 18.96 ;
      RECT 2.616 17.76 2.662 18.96 ;
      RECT 2.272 17.76 2.484 18.24 ;
      RECT 2.528 17.76 2.572 18.24 ;
      RECT 1.838 17.52 2.484 17.76 ;
      RECT 2.528 17.52 2.662 17.76 ;
      RECT 2.272 17.04 2.484 17.52 ;
      RECT 2.528 17.04 2.572 17.52 ;
      RECT 2.272 16.8 2.572 17.04 ;
      RECT 1.838 16.32 2.228 17.52 ;
      RECT 2.616 16.32 2.662 17.52 ;
      RECT 2.272 16.32 2.484 16.8 ;
      RECT 2.528 16.32 2.572 16.8 ;
      RECT 1.838 16.08 2.484 16.32 ;
      RECT 2.528 16.08 2.662 16.32 ;
      RECT 2.272 15.6 2.484 16.08 ;
      RECT 2.528 15.6 2.572 16.08 ;
      RECT 2.272 15.36 2.572 15.6 ;
      RECT 1.838 14.88 2.228 16.08 ;
      RECT 2.616 14.88 2.662 16.08 ;
      RECT 2.272 14.88 2.484 15.36 ;
      RECT 2.528 14.88 2.572 15.36 ;
      RECT 1.838 14.64 2.484 14.88 ;
      RECT 2.528 14.64 2.662 14.88 ;
      RECT 2.272 14.16 2.484 14.64 ;
      RECT 2.528 14.16 2.572 14.64 ;
      RECT 2.272 13.92 2.572 14.16 ;
      RECT 1.838 13.44 2.228 14.64 ;
      RECT 2.616 13.44 2.662 14.64 ;
      RECT 2.272 13.44 2.484 13.92 ;
      RECT 2.528 13.44 2.572 13.92 ;
      RECT 1.838 13.2 2.484 13.44 ;
      RECT 2.528 13.2 2.662 13.44 ;
      RECT 2.272 12.72 2.484 13.2 ;
      RECT 2.528 12.72 2.572 13.2 ;
      RECT 2.272 12.48 2.572 12.72 ;
      RECT 1.838 12 2.228 13.2 ;
      RECT 2.616 12 2.662 13.2 ;
      RECT 2.272 12 2.484 12.48 ;
      RECT 2.528 12 2.572 12.48 ;
      RECT 1.838 11.76 2.484 12 ;
      RECT 2.528 11.76 2.662 12 ;
      RECT 2.272 11.28 2.484 11.76 ;
      RECT 2.528 11.28 2.572 11.76 ;
      RECT 2.272 11.04 2.572 11.28 ;
      RECT 1.838 10.56 2.228 11.76 ;
      RECT 2.616 10.56 2.662 11.76 ;
      RECT 2.272 10.56 2.484 11.04 ;
      RECT 2.528 10.56 2.572 11.04 ;
      RECT 1.838 10.32 2.484 10.56 ;
      RECT 2.528 10.32 2.662 10.56 ;
      RECT 2.272 9.84 2.484 10.32 ;
      RECT 2.528 9.84 2.572 10.32 ;
      RECT 2.272 9.6 2.572 9.84 ;
      RECT 1.838 9.12 2.228 10.32 ;
      RECT 2.616 9.12 2.662 10.32 ;
      RECT 2.272 9.12 2.484 9.6 ;
      RECT 2.528 9.12 2.572 9.6 ;
      RECT 1.838 8.88 2.484 9.12 ;
      RECT 2.528 8.88 2.662 9.12 ;
      RECT 2.272 8.4 2.484 8.88 ;
      RECT 2.528 8.4 2.572 8.88 ;
      RECT 2.272 8.16 2.572 8.4 ;
      RECT 1.838 7.68 2.228 8.88 ;
      RECT 2.616 7.68 2.662 8.88 ;
      RECT 2.272 7.68 2.484 8.16 ;
      RECT 2.528 7.68 2.572 8.16 ;
      RECT 1.838 7.44 2.484 7.68 ;
      RECT 2.528 7.44 2.662 7.68 ;
      RECT 2.272 6.96 2.484 7.44 ;
      RECT 2.528 6.96 2.572 7.44 ;
      RECT 2.272 6.72 2.572 6.96 ;
      RECT 1.838 6.24 2.228 7.44 ;
      RECT 2.616 6.24 2.662 7.44 ;
      RECT 2.272 6.24 2.484 6.72 ;
      RECT 2.528 6.24 2.572 6.72 ;
      RECT 1.838 6 2.484 6.24 ;
      RECT 2.528 6 2.662 6.24 ;
      RECT 2.272 5.52 2.484 6 ;
      RECT 2.528 5.52 2.572 6 ;
      RECT 2.272 5.28 2.572 5.52 ;
      RECT 1.838 4.8 2.228 6 ;
      RECT 2.616 4.8 2.662 6 ;
      RECT 2.272 4.8 2.484 5.28 ;
      RECT 2.528 4.8 2.572 5.28 ;
      RECT 1.838 4.08 2.484 4.8 ;
      RECT 2.528 4.08 2.662 4.8 ;
      RECT 1.838 3.72 2.662 4.08 ;
      RECT 1.838 2.52 1.884 3.72 ;
      RECT 1.928 2.52 2.228 3.72 ;
      RECT 2.272 2.52 2.572 3.72 ;
      RECT 2.616 2.52 2.662 3.72 ;
      RECT 1.838 1.8 2.662 2.52 ;
      RECT 1.838 0.6 1.884 1.8 ;
      RECT 1.928 0.6 2.228 1.8 ;
      RECT 2.272 0.6 2.572 1.8 ;
      RECT 2.616 0.6 2.662 1.8 ;
      RECT 1.838 -0.12 2.662 0.6 ;
      RECT 0.938 3.72 1.762 25.08 ;
      RECT 0.938 2.52 1.072 3.72 ;
      RECT 1.116 2.52 1.584 3.72 ;
      RECT 1.628 2.52 1.762 3.72 ;
      RECT 0.938 1.8 1.762 2.52 ;
      RECT 0.938 0.6 0.984 1.8 ;
      RECT 1.028 0.6 1.072 1.8 ;
      RECT 1.116 0.6 1.584 1.8 ;
      RECT 1.628 0.6 1.762 1.8 ;
      RECT 0.938 -0.12 1.762 0.6 ;
      RECT -0.04 25.02 0.862 25.08 ;
      RECT -0.092 3.72 0.862 25.02 ;
      RECT -0.092 2.52 0.428 3.72 ;
      RECT 0.472 2.52 0.684 3.72 ;
      RECT 0.728 2.52 0.772 3.72 ;
      RECT 0.816 2.52 0.862 3.72 ;
      RECT -0.092 1.8 0.862 2.52 ;
      RECT -0.092 0.6 0.428 1.8 ;
      RECT 0.472 0.6 0.684 1.8 ;
      RECT 0.728 0.6 0.772 1.8 ;
      RECT 0.816 0.6 0.862 1.8 ;
      RECT -0.092 -0.06 0.862 0.6 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 22.658 0 23.32 24.96 ;
      RECT 21.758 0 22.342 24.96 ;
      RECT 20.858 0 21.442 24.96 ;
      RECT 19.958 0 20.542 24.96 ;
      RECT 19.058 0 19.642 24.96 ;
      RECT 18.158 0 18.742 24.96 ;
      RECT 17.258 0 17.842 24.96 ;
      RECT 16.358 0 16.942 24.96 ;
      RECT 15.458 0 16.042 24.96 ;
      RECT 14.558 0 15.142 24.96 ;
      RECT 13.658 0 14.242 24.96 ;
      RECT 12.758 0 13.342 24.96 ;
      RECT 11.858 0 12.442 24.96 ;
      RECT 10.958 0 11.542 24.96 ;
      RECT 10.058 0 10.642 24.96 ;
      RECT 9.158 0 9.742 24.96 ;
      RECT 8.258 0 8.842 24.96 ;
      RECT 7.358 0 7.942 24.96 ;
      RECT 6.458 0 7.042 24.96 ;
      RECT 5.558 0 6.142 24.96 ;
      RECT 4.658 0 5.242 24.96 ;
      RECT 3.758 24.84 4.342 24.96 ;
      RECT 4.192 24.12 4.342 24.84 ;
      RECT 3.758 4.68 3.908 24.84 ;
      RECT 3.758 3.96 4.164 4.68 ;
      RECT 3.758 3.84 4.342 3.96 ;
      RECT 3.848 2.4 3.908 3.84 ;
      RECT 4.192 2.4 4.342 3.84 ;
      RECT 3.758 1.92 4.342 2.4 ;
      RECT 3.848 0.48 3.908 1.92 ;
      RECT 4.192 0.48 4.342 1.92 ;
      RECT 3.758 0 4.342 0.48 ;
      RECT 2.858 24.84 3.442 24.96 ;
      RECT 2.858 24.12 3.264 24.84 ;
      RECT 2.948 4.68 3.264 24.12 ;
      RECT 2.948 3.96 3.352 4.68 ;
      RECT 2.858 3.84 3.442 3.96 ;
      RECT 3.036 2.4 3.264 3.84 ;
      RECT 2.858 1.92 3.442 2.4 ;
      RECT 3.036 0.48 3.264 1.92 ;
      RECT 2.858 0 3.442 0.48 ;
      RECT 1.958 24.84 2.542 24.96 ;
      RECT 2.392 24.12 2.452 24.84 ;
      RECT 1.958 4.68 2.108 24.84 ;
      RECT 1.958 3.96 2.364 4.68 ;
      RECT 1.958 3.84 2.542 3.96 ;
      RECT 2.048 2.4 2.108 3.84 ;
      RECT 2.392 2.4 2.452 3.84 ;
      RECT 1.958 1.92 2.542 2.4 ;
      RECT 2.048 0.48 2.108 1.92 ;
      RECT 2.392 0.48 2.452 1.92 ;
      RECT 1.958 0 2.542 0.48 ;
      RECT 1.058 3.84 1.642 24.96 ;
      RECT 1.236 2.4 1.464 3.84 ;
      RECT 1.058 1.92 1.642 2.4 ;
      RECT 1.236 0.48 1.464 1.92 ;
      RECT 1.058 0 1.642 0.48 ;
      RECT 0.08 3.84 0.742 24.96 ;
      RECT 0.08 2.4 0.308 3.84 ;
      RECT 0.08 1.92 0.742 2.4 ;
      RECT 0.08 0.48 0.308 1.92 ;
      RECT 0.08 0 0.742 0.48 ;
    LAYER m0 ;
      RECT 0 0.002 23.4 24.958 ;
    LAYER m1 ;
      RECT 0 0 23.4 24.96 ;
    LAYER m2 ;
      RECT 0 0.015 23.4 24.945 ;
    LAYER m3 ;
      RECT 0.015 0 23.385 24.96 ;
    LAYER m4 ;
      RECT 0 0.02 23.4 24.94 ;
    LAYER m5 ;
      RECT 0.012 0 23.388 24.96 ;
    LAYER m6 ;
      RECT 0 0.012 23.4 24.948 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf054b128e1r1w0cbbehraa4acw

END LIBRARY
