parameter TARGETREG=1;
parameter DEASSERT_CLK_SIGS=0;
parameter ASYNCEQDEPTH=22;
parameter NPQUEUEDEPTH=10;
parameter RELATIVE_PLACEMENT_EN=0;
parameter MAXNPMSTR=0;
parameter SB_PARITY_REQUIRED=0;
parameter TX_EXT_HEADER_SUPPORT=1;
parameter MATCHED_INTERNAL_WIDTH=0;
parameter IOSFSB_EP_SPEC_REV=11;
parameter SIDE_USYNC_DELAY=1;
parameter DUMMY_CLKBUF=0;
parameter DO_SERR_MASTER=0;
parameter LATCHQUEUES=0;
parameter EXPECTED_COMPLETIONS_COUNTER=0;
parameter NUM_REPEATER=0;
parameter VARIABLE_CLAIM_DELAY=0;
parameter GLOBAL_EP=0;
parameter VALONLYMODEL=0;
parameter USYNC_ENABLE=0;
parameter NUMBER_OF_BITS_PER_LANE=8;
parameter RX_EXT_HEADER_SUPPORT=1;
parameter UNIQUE_EXT_HEADERS=1;
parameter SBE_VISA_ID_PARAM=11;
parameter NUM_CLAIM_REPEATER=0;
parameter NUMBER_OF_VISAMUX_MODULES=1;
parameter MAXPCTRGT=0;
parameter MAXTRGTDATA=63;
parameter AGENT_USYNC_DELAY=1;
parameter ASYNCENDPT=0;
parameter MAXPLDBIT=31;
parameter PIPEINPS=0;
parameter RX_EXT_HEADER_IDS=44;
parameter RSWIDTH=0;
parameter SAIWIDTH=8;
parameter MAXMSTRDATA=63;
parameter PCQUEUEDEPTH=16;
parameter ASYNCIQDEPTH=26;
parameter SKIP_ACTIVEREQ=1;
parameter DISABLE_COMPLETION_FENCING=0;
parameter ISM_COMPLETION_FENCING=0;
parameter FAB_CLK_PERIOD=4478;
parameter MAXMSTRADDR=47;
parameter MASTERREG=1;
parameter IOSFSB_FBRC_SPEC_REV=11;
parameter CLKREQDEFAULT=1;
parameter FBRC_EXT_HEADER_SUPPORT=1;
parameter PIPEISMS=0;
parameter MAXNPTRGT=0;
parameter NUM_RX_EXT_HEADERS=0+1;
parameter AGT_CLK_PERIOD=7263;
parameter AGT_EXT_HEADER_SUPPORT=1;
parameter BULKRDWR=0;
parameter NUMBER_OF_OUTPUT_LANES=1;
parameter MAXPCMSTR=0;
parameter NUM_TX_EXT_HEADERS=0+1;
parameter CUP2PUT1CYC=0;
parameter MAXTRGTADDR=15;
parameter GLOBAL_EP_IS_STRAP=0;
parameter BULK_PERF=0;

