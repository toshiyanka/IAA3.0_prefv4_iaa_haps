// File output was printed on: Thursday, March 21, 2013 4:21:02 PM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
//             TAP                SlvIDcode       IDcode      IR_Width  Node  Sec_connections  Hybrid_en  Dfx_Security  Hierarchy_Level  PositionOfTap  IsVendorTap    VendorIdOpcode 
Create_TAP_LUT (IPLEVEL_STAP,  32'h0400_0001,  32'h1234_5679, 'd8,     'd0,       'd0,         'd0,       GREEN,           1,               0,             1,             'h0C);
