// CCTypes begin

	typedef class CCAgent;
	typedef class CCAgentSequencer;
	//typedef class CCAgentMonitor;
	typedef class CCAgentDriver;
	//typedef class CCAgentPrinter;
	typedef class CCAgentSeqItem;
	//typedef class CCAgentResponseVSequencer;
	typedef class CCAgentResponder;
	typedef class CCAgentSIPResponder;

	//typedef class CCAgentBaseResponseVSeq;
	typedef class CCAgentResponseSeqItem;
	typedef class CCAgentArbiter;
	typedef class CCAgentSIPFSM;
	typedef class CCAgentFabricFSM;

//	typedef class CCAgentFETFSM;
//	typedef class CCAgentFETState;


