//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//
//  -- Intel Proprietary
//  -- Copyright (C) 2015 Intel Corporation
//  -- All Rights Reserved
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2009-2020 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code (Material) are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//
//
//  Collateral Description:
//  IOSF - Sideband Channel IP
//
//  Source organization:
//  SEG / SIP / IOSF IP Engineering
//
//  Support Information:
//  WEB: http://moss.amr.ith.intel.com/sites/SoftIP/Shared%20Documents/Forms/AllItems.aspx
//  HSD: https://vthsd.fm.intel.com/hsd/seg_softip/default.aspx
//
//  Revision:
//  2020WW22_PICr33
//
//  Module <sTAP> :  < put your functional description here in plain text >
//
//------------------------------------------------------------------------------

//----------------------------------------------------------------------
// Intel Proprietary -- Copyright 2009 Intel -- All rights reserved
//----------------------------------------------------------------------
// NOTE: Log history is at end of file.
//----------------------------------------------------------------------
//
//    FILENAME    : stap_irdecoder.sv
//    DESIGNER    : Sunjiv Sachan
//    PROJECT     : sTAP
//    
//    
//    PURPOSE     : sTAP IR Decoder Logic
//    DESCRIPTION :
//       This module generated decoder enable signals. This is generated by
//       comparing instruction address with address defined by parameter.
//----------------------------------------------------------------------
//    LOCAL PARAMETERS:
//
//    HIGH
//       This is 1 bit one value
//
//    LOW
//       This is 1 bit zero value
//
//    ONE
//       This is number 1 to and is declared just to avoid lint warnings
//
//    TWO
//       This is number 2 to and is declared just to avoid lint warnings
//
//    IRDECODER_STAP_ADDRESS_OF_USERCODE
//       This is address of optional USERCODE register.
//----------------------------------------------------------------------
module stap_irdecoder
   #(
   parameter IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION       = 8,
   parameter IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS      = 0,
   parameter IRDECODER_STAP_INSTRUCTION_FOR_DATA_REGISTERS = 0,
   parameter IRDECODER_STAP_ADDRESS_OF_CLAMP               = 0,
   parameter IRDECODER_STAP_MINIMUM_SIZEOF_INSTRUCTION     = 0,
   parameter IRDECODER_STAP_ENABLE_BSCAN                   = 0
   )
   (
   input  logic                                                    powergoodrst_trst_b, //kbbhagwa cdc fix
   input  logic [(IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  stap_irreg_ireg,

   input  logic [(IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION - 1):0]  stap_irreg_ireg_nxt,//kbbhagwa cdc fix 
   input  logic                                                    ftap_tck, //kbbhagwa cdc fix
   output logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] stap_irdecoder_drselect,
   output logic                                                    stap_and_all_bits_irreg,
   output logic                                                    stap_or_all_bits_irreg
   );

   // *********************************************************************
   // Local parameters
   // *********************************************************************
   localparam DRREG_STAP_POSITION_OF_SLVIDCODE   = (IRDECODER_STAP_ENABLE_BSCAN == 1) ? 5 : 2; //kbbhagwa cdc fix
   localparam HIGH                               = 1'b1;
   localparam LOW                                = 1'b0;
   localparam ONE                                = 1;
   localparam TWO                                = 2;
   //localparam IRDECODER_STAP_POSITION_OF_IDCODE  = 3;
   localparam IRDECODER_STAP_POSITION_OF_HIGHZ   = 3;
   localparam IRDECODER_STAP_POSITION_OF_EXTEST  = 4;
   //localparam IRDECODER_STAP_POSITION_OF_RESIRA  = 6;
   //localparam IRDECODER_STAP_POSITION_OF_RESIRB  = 7;
   //localparam IRDECODER_STAP_ADDRESS_OF_USERCODE = (IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION == 8) ? 8'h05 :
   //   {{(IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION -
   //      IRDECODER_STAP_MINIMUM_SIZEOF_INSTRUCTION + 4){LOW}}, 4'h5};

   // *********************************************************************
   // Internal signals
   // *********************************************************************
   logic                                                    and_all_bits_irreg_nxt; //kbbhagwa cdc fix
   logic                                                    or_all_bits_irreg_nxt; //kbbhagwa cdc fix
   //logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] drselect_reset_value;
   //

   logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] irdecoder_drselect_nxt;
   logic [(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - 1):0] decoder_drselect;
   //kbbhagwa cdc fix

   logic                                                    decode_clamp;
   //logic                                                    decode_usercode;

   // *********************************************************************
   // Generate construct is used to generate number of decoded output lines
   // which is equal to IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS
   // *********************************************************************
   generate
      for (genvar i = 0; i < IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS; i = i + 1)
      begin
         stap_decoder #(
                        .DECODER_INSTRUCTION_TO_DECODE
                           (IRDECODER_STAP_INSTRUCTION_FOR_DATA_REGISTERS[
                              (((i * IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION) +
                                IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION) - 1):
                              (i * IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION)]),
                        .DECODER_STAP_SIZE_OF_EACH_INSTRUCTION
                           (IRDECODER_STAP_SIZE_OF_EACH_INSTRUCTION)
                       )
         i_stap_decoder (
//                         .stap_irreg_ireg  (stap_irreg_ireg),
                         .stap_irreg_ireg  (stap_irreg_ireg_nxt), //kbbhagwa cdc fix
                         .decoder_drselect (decoder_drselect[i])
                        );
      end
   endgenerate

always_ff @(negedge ftap_tck or negedge powergoodrst_trst_b)
  if ( ~ powergoodrst_trst_b )
      for ( integer i = 0; i <= (IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS -1 ); i++ ) 
      begin
         if ( i == DRREG_STAP_POSITION_OF_SLVIDCODE )
             stap_irdecoder_drselect[DRREG_STAP_POSITION_OF_SLVIDCODE] <= 1'b1;
         else
             stap_irdecoder_drselect[i] <= 1'b0;
      end
  else 
        stap_irdecoder_drselect <= irdecoder_drselect_nxt;
//kbbhagwa cdc fix

   // *********************************************************************
   // Decoding of some of the Instructions
   // *********************************************************************
   assign stap_and_all_bits_irreg = &(stap_irreg_ireg);
   assign stap_or_all_bits_irreg  = |(stap_irreg_ireg);

   assign and_all_bits_irreg_nxt = &(stap_irreg_ireg_nxt);
   assign or_all_bits_irreg_nxt  = |(stap_irreg_ireg_nxt);

   generate
      if (IRDECODER_STAP_ENABLE_BSCAN == 1)
      begin
         assign decode_clamp =
// (stap_irreg_ireg == IRDECODER_STAP_ADDRESS_OF_CLAMP)    ? HIGH : LOW;
// kbbhagwa cdc fix
            (stap_irreg_ireg_nxt == IRDECODER_STAP_ADDRESS_OF_CLAMP)    ? HIGH : LOW;
         //assign decode_usercode =
         //   (stap_irreg_ireg == IRDECODER_STAP_ADDRESS_OF_USERCODE) ? HIGH : LOW;
         // *********************************************************************
         // Default value of decoder select points to BYPASS register
         // *********************************************************************
// kbbhagwa cdc fix assign stap_irdecoder_drselect =
         assign irdecoder_drselect_nxt =
            (and_all_bits_irreg_nxt == HIGH)                                       ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            (or_all_bits_irreg_nxt == LOW )                                        ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - TWO){LOW}}, HIGH, LOW} :
            (decode_clamp == HIGH)                                                  ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
         //   (decode_usercode == HIGH)                                               ?
         //      {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            (decoder_drselect == {IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS{LOW}})   ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            //(decoder_drselect[IRDECODER_STAP_POSITION_OF_IDCODE] == HIGH)           ?
               //{{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            (decoder_drselect[IRDECODER_STAP_POSITION_OF_HIGHZ]  == HIGH)           ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            //(decoder_drselect[IRDECODER_STAP_POSITION_OF_RESIRA] == HIGH)           ?
               //{{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            //(decoder_drselect[IRDECODER_STAP_POSITION_OF_RESIRB] == HIGH)           ?
               //{{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            decoder_drselect;
      end
      else
      begin
         assign irdecoder_drselect_nxt =
            (and_all_bits_irreg_nxt == HIGH)                                       ?
//kbbhagwa cdc fix  (stap_and_all_bits_irreg == HIGH)                                       ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            (or_all_bits_irreg_nxt == LOW )                                        ?
//            (stap_or_all_bits_irreg == LOW )                                        ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - TWO){LOW}}, HIGH, LOW} :
            (decoder_drselect == {IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS{LOW}})   ?
               {{(IRDECODER_STAP_NUMBER_OF_TOTAL_REGISTERS - ONE){LOW}}, HIGH}      :
            decoder_drselect;
      end
   endgenerate

endmodule
