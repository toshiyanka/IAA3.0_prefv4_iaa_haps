//-----------------------------------------------------------------
// Intel Proprietary -- Copyright 2013 Intel -- All rights reserved 
//-----------------------------------------------------------------
// Author       : rahul Ramaswami
// Date Created : 06-2014
//-----------------------------------------------------------------
// Description:
// DNV topology picker
//------------------------------------------------------------------
// Define & register this picker with shr_tb


`picker_class_begin(socket_picker, base_socket_picker)


`picker_class_end
