//------------------------------------------------------------------------------------------------------------------------
//
//  INTEL CONFIDENTIAL
//
//  Copyright 2023 Intel Corporation All Rights Reserved.
//
//  The source code contained or described herein and all documents related
//  to the source code ("Material") are owned by Intel Corporation or its
//  suppliers or licensors. Title to the Material remains with Intel
//  Corporation or its suppliers and licensors. The Material contains trade
//  secrets and proprietary and confidential information of Intel or its
//  suppliers and licensors. The Material is protected by worldwide copyright
//  and trade secret laws and treaty provisions. No part of the Material may
//  be used, copied, reproduced, modified, published, uploaded, posted,
//  transmitted, distributed, or disclosed in any way without Intel's prior
//  express written permission.
//
//  No license under any patent, copyright, trade secret or other intellectual
//  property right is granted to or conferred upon you by disclosure or
//  delivery of the Materials, either expressly, by implication, inducement,
//  estoppel or otherwise. Any license under such intellectual property rights
//  must be express and approved by Intel in writing.
//

//------------------------------------------------------------------------------------------------------------------------
// Intel Proprietary        Intel Confidential        Intel Proprietary        Intel Confidential        Intel Proprietary
//------------------------------------------------------------------------------------------------------------------------
// Generated by                  : cudoming
// Generated on                  : April 19, 2023
//------------------------------------------------------------------------------------------------------------------------
// General Information:
// ------------------------------
// 2r2w0c standard array for SDG server designs.
// Behavioral modeling of a parameterized register file core with no DFX features.
// RTL is written in SystemVerilog.
//------------------------------------------------------------------------------------------------------------------------
// Detail Information:
// ------------------------------
// Addresses        : RD/WR addresses are encoded.
//                    Input addresses will be valid at the array in 1 phases after being driven.
//                    Address latency of 1 is corresponding to a B-latch.
// Enables          : RD/WR enables are used to condition the clock and wordlines.
//                  : Input enables will be valid at the array in 1 phases after being driven.
//                    Enable latency of 1 is corresponding to a B-latch.
// Write Data       : Write data will be valid at the array 2 phases after being driven.
//                    Write data latency of 2 is corresponding to a rising-edge flop. 
// Read Data        : Read data will be valid at the output of a SDL 1 phase after being read.
//                    Read data latency of 1 is corresponding to a B-latch.
// Address Offset   : 
//------------------------------------------------------------------------------------------------------------------------

//------------------------------------------------------------------------------------------------------------------------
// Other Information:
// ------------------------------
// SDG RFIP RTL Release Path:
// /p/hdk/rtl/ip_releases/shdk74/array_macro_module
//
//------------------------------------------------------------------------------------------------------------------------


/// Parent Module    : arf156b040e2r2w0cbbehbaa4acw_dfx_wrapper
/// Child Module     : array_generic_rwx_std

`ifndef ARF156B040E2R2W0CBBEHBAA4ACW_SV
`define ARF156B040E2R2W0CBBEHBAA4ACW_SV

//------------------------------------------------------------------------------------------------------------------------
// module arf156b040e2r2w0cbbehbaa4acw
//------------------------------------------------------------------------------------------------------------------------
module arf156b040e2r2w0cbbehbaa4acw #(

//------------------------------------------------------------------------------------------------------------------------
// local parameters
//------------------------------------------------------------------------------------------------------------------------
  localparam MODULE                 = "arf156b040e2r2w0cbbehbaa4acw",
  localparam BITS                   = 160,
  localparam ENTRIES                = 40,
  localparam DWIDTH                 = 160,
  localparam AWIDTH                 = 6,
  localparam RD_PORTS               = 2,
  localparam WR_PORTS               = 2,
  localparam CM_PORTS               = 0,
  localparam BPHASE_RD              = 0,
  localparam BPHASE_WR              = 0,
  localparam BPHASE_CM              = 0,
  localparam SEGMENTS               = 0,
  localparam BITS_PER_SEGMENT       = 0,
  localparam SDL_INITVAL            = {1'b0,1'b0},
  localparam ADDRESS_OFFSET         = 0,
  localparam NO_CAM_LATENCY         = 0,
  localparam NO_CAM_LSB             = 0
)
(

//------------------------------------------------------------------------------------------------------------------------
// interfaces
//------------------------------------------------------------------------------------------------------------------------

  //------------------------------
  // read interfaces
  //------------------------------
  input   wire                            ckrdp0,
  input   wire                            rdenp0,
  input   wire    [AWIDTH-1:0]            rdaddrp0,
  output  wire    [DWIDTH-1:0]            rddatap0,
  input   wire                            sdl_initp0,
  input   wire                            ckrdp1,
  input   wire                            rdenp1,
  input   wire    [AWIDTH-1:0]            rdaddrp1,
  output  wire    [DWIDTH-1:0]            rddatap1,
  input   wire                            sdl_initp1,

  //------------------------------
  // write interfaces
  //------------------------------
  input   wire                            ckwrp0,
  input   wire                            wrenp0,
  input   wire    [AWIDTH-1:0]            wraddrp0,
  input   wire    [DWIDTH-1:0]            wrdatap0,
  input   wire                            ckwrp1,
  input   wire                            wrenp1,
  input   wire    [AWIDTH-1:0]            wraddrp1,
  input   wire    [DWIDTH-1:0]            wrdatap1,



  //------------------------------
  // rcb interfaces
  //------------------------------
  input   wire                            rdaddrp0_fd,
  input   wire                            rdaddrp0_rd,
  input   wire                            rdaddrp1_fd,
  input   wire                            rdaddrp1_rd,
  input   wire                            wraddrp0_fd,
  input   wire                            wraddrp0_rd,
  input   wire                            wrdatap0_fd,
  input   wire                            wrdatap0_rd,
  input   wire                            wraddrp1_fd,
  input   wire                            wraddrp1_rd,
  input   wire                            wrdatap1_fd,
  input   wire                            wrdatap1_rd

);



//------------------------------------------------------------------------------------------------------------------------
// instantiation array_generic_rwx_std
//------------------------------------------------------------------------------------------------------------------------
arf156b040e2r2w0cbbehbaa4acw_array_generic_rwx_std #
(

  .MODULE                     (MODULE),
  .BITS                       (BITS),
  .ENTRIES                    (ENTRIES),
  .AWIDTH                     (AWIDTH),
  .DWIDTH                     (DWIDTH),
  .RD_PORTS                   (RD_PORTS),
  .WR_PORTS                   (WR_PORTS),
  .CM_PORTS                   (CM_PORTS),
  .BPHASE_RD                  (BPHASE_RD),
  .BPHASE_WR                  (BPHASE_WR),
  .BPHASE_CM                  (BPHASE_CM),
  .SEGMENTS                   (SEGMENTS),
  .BITS_PER_SEGMENT           (BITS_PER_SEGMENT),
  .SDL_INITVAL                (SDL_INITVAL),
  .ADDRESS_OFFSET             (ADDRESS_OFFSET),
  .NO_CAM_LATENCY             (NO_CAM_LATENCY),
  .NO_CAM_LSB                 (NO_CAM_LSB)

)
array_generic
(

  //------------------------------
  // read interfaces
  //------------------------------
  .ckrd             ( {>>{ ckrdp0, ckrdp1  }} ),
  .rden             ( {>>{ rdenp0, rdenp1 }} ),
  .rdaddr           ( {>>{ rdaddrp0, rdaddrp1 }} ),
  .rddata           ( {>>{ rddatap0, rddatap1 }} ),
  .sdl_init         ( {>>{ sdl_initp0, sdl_initp1 }} ),

  //------------------------------
  // write interfaces
  //------------------------------
  .ckwr             ( {>>{ ckwrp0, ckwrp1 }} ),
  .wren             ( {>>{ wrenp0, wrenp1 }} ),
  .wraddr           ( {>>{ wraddrp0, wraddrp1 }} ),
  .wrdata           ( {>>{ wrdatap0, wrdatap1 }} ),



  //------------------------------
  // rcb interfaces
  //------------------------------
  .rdaddr_fd        ( {>>{ rdaddrp0_fd, rdaddrp1_fd }} ),
  .rdaddr_rd        ( {>>{ rdaddrp0_rd, rdaddrp1_rd }} ),
  .wraddr_fd        ( {>>{ wraddrp0_fd, wraddrp1_fd }} ),
  .wraddr_rd        ( {>>{ wraddrp0_rd, wraddrp1_rd }} ),
  .wrdata_fd        ( {>>{ wrdatap0_fd, wrdatap1_fd }} ),
  .wrdata_rd        ( {>>{ wrdatap0_rd, wrdatap1_rd }} )


);

`ifdef INTC_MEM_GLS

  //err variables
  logic errSDL_INITP0, errSDL_INITP1;
  logic errsdl_initp0, errsdl_initp1;
  logic errRDENP0, errRDENP1;
  logic errrdenp0, errrdenp1;
  logic errRDADDRP0, errRDADDRP1;
  logic errrdaddrp0, errrdaddrp1;
  
  logic errWRENP0, errWRENP1;
  logic errwrenp0, errwrenp1;
  logic errWRADDRP0, errWRADDRP1;
  logic errwraddrp0, errwraddrp1;
  logic errWRDATAP0, errWRDATAP1;
  logic errwrdatap0, errwrdatap1;


  always @(errSDL_INITP0) errsdl_initp0 = 1'b1;
  always @(errRDENP0) errrdenp0 = 1'b1;
  always @(errRDADDRP0) errrdaddrp0 = 1'b1;

  always @(errSDL_INITP1) errsdl_initp1 = 1'b1;
  always @(errRDENP1) errrdenp1 = 1'b1;
  always @(errRDADDRP1) errrdaddrp1 = 1'b1;

  always @(errWRENP0) errwrenp0 = 1'b1;
  always @(errWRADDRP0) errwraddrp0 = 1'b1;
  always @(errWRDATAP0) errwrdatap0 = 1'b1;

  always @(errWRENP1) errwrenp1 = 1'b1;
  always @(errWRADDRP1) errwraddrp1 = 1'b1;
  always @(errWRDATAP1) errwrdatap1 = 1'b1;

  always @(negedge ckrdp0) begin
    errsdl_initp0 = 1'b0;
    errrdenp0 = 1'b0;
    errrdaddrp0 = 1'b0;
  end

  always @(negedge ckrdp1) begin
    errsdl_initp1 = 1'b0;
    errrdenp1 = 1'b0;
    errrdaddrp1 = 1'b0;
  end

  always @(negedge ckwrp0) begin
    errwrenp0 = 1'b0;
    errwraddrp0 = 1'b0;
    errwrdatap0 = 1'b0;
  end

  always @(negedge ckwrp1) begin
    errwrenp1 = 1'b0;
    errwraddrp1 = 1'b0;
    errwrdatap1 = 1'b0;
  end


specify
  specparam trddatap0_r = 0.00:0.00:0.00;
  specparam trddatap0_f = 0.00:0.00:0.00;

  specparam trddatap1_r = 0.00:0.00:0.00;
  specparam trddatap1_f = 0.00:0.00:0.00;

  specparam tsdl_initp0_sr = 0.00:0.00:0.00;
  specparam tsdl_initp0_sf = 0.00:0.00:0.00;
  specparam tsdl_initp0_hr = 0.00:0.00:0.00;
  specparam tsdl_initp0_hf = 0.00:0.00:0.00;

  specparam tsdl_initp1_sr = 0.00:0.00:0.00;
  specparam tsdl_initp1_sf = 0.00:0.00:0.00;
  specparam tsdl_initp1_hr = 0.00:0.00:0.00;
  specparam tsdl_initp1_hf = 0.00:0.00:0.00;

  specparam trdenp0_sr = 0.00:0.00:0.00;
  specparam trdenp0_sf = 0.00:0.00:0.00;
  specparam trdenp0_hr = 0.00:0.00:0.00;
  specparam trdenp0_hf = 0.00:0.00:0.00;

  specparam trdenp1_sr = 0.00:0.00:0.00;
  specparam trdenp1_sf = 0.00:0.00:0.00;
  specparam trdenp1_hr = 0.00:0.00:0.00;
  specparam trdenp1_hf = 0.00:0.00:0.00;

  specparam trdaddrp0_sr = 0.00:0.00:0.00;
  specparam trdaddrp0_sf = 0.00:0.00:0.00;
  specparam trdaddrp0_hr = 0.00:0.00:0.00;
  specparam trdaddrp0_hf = 0.00:0.00:0.00;

  specparam trdaddrp1_sr = 0.00:0.00:0.00;
  specparam trdaddrp1_sf = 0.00:0.00:0.00;
  specparam trdaddrp1_hr = 0.00:0.00:0.00;
  specparam trdaddrp1_hf = 0.00:0.00:0.00;

  specparam twrenp0_sr = 0.00:0.00:0.00;
  specparam twrenp0_sf = 0.00:0.00:0.00;
  specparam twrenp0_hr = 0.00:0.00:0.00;
  specparam twrenp0_hf = 0.00:0.00:0.00;

  specparam twrenp1_sr = 0.00:0.00:0.00;
  specparam twrenp1_sf = 0.00:0.00:0.00;
  specparam twrenp1_hr = 0.00:0.00:0.00;
  specparam twrenp1_hf = 0.00:0.00:0.00;

  specparam twraddrp0_sr = 0.00:0.00:0.00;
  specparam twraddrp0_sf = 0.00:0.00:0.00;
  specparam twraddrp0_hr = 0.00:0.00:0.00;
  specparam twraddrp0_hf = 0.00:0.00:0.00;
  specparam twraddrp1_sr = 0.00:0.00:0.00;
  specparam twraddrp1_sf = 0.00:0.00:0.00;
  specparam twraddrp1_hr = 0.00:0.00:0.00;
  specparam twraddrp1_hf = 0.00:0.00:0.00;
  
  specparam twrdatap0_sr = 0.00:0.00:0.00;
  specparam twrdatap0_sf = 0.00:0.00:0.00;
  specparam twrdatap0_hr = 0.00:0.00:0.00;
  specparam twrdatap0_hf = 0.00:0.00:0.00;  
  specparam twrdatap1_sr = 0.00:0.00:0.00;
  specparam twrdatap1_sf = 0.00:0.00:0.00;
  specparam twrdatap1_hr = 0.00:0.00:0.00;
  specparam twrdatap1_hf = 0.00:0.00:0.00;

  //sdl_init
  $setuphold(posedge ckrdp0, posedge sdl_initp0, tsdl_initp0_sr, tsdl_initp0_hr, errSDL_INITP0);
  $setuphold(posedge ckrdp0, negedge sdl_initp0, tsdl_initp0_sf, tsdl_initp0_hf, errSDL_INITP0);

  $setuphold(posedge ckrdp1, posedge sdl_initp1, tsdl_initp1_sr, tsdl_initp1_hr, errSDL_INITP1);
  $setuphold(posedge ckrdp1, negedge sdl_initp1, tsdl_initp1_sf, tsdl_initp1_hf, errSDL_INITP1);


  //rden
  $setuphold(posedge ckrdp0, posedge rdenp0, trdenp0_sr, trdenp0_hr, errRDENP0);
  $setuphold(posedge ckrdp0, negedge rdenp0, trdenp0_sf, trdenp0_hf, errRDENP0);

  $setuphold(posedge ckrdp1, posedge rdenp1, trdenp1_sr, trdenp1_hr, errRDENP1);
  $setuphold(posedge ckrdp1, negedge rdenp1, trdenp1_sf, trdenp1_hf, errRDENP1);

  
  //rdaddr
  $setuphold(posedge ckrdp0, posedge rdaddrp0[5], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[5], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[4], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[4], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[3], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[3], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[2], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[2], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[1], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[1], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);
  $setuphold(posedge ckrdp0, posedge rdaddrp0[0], trdaddrp0_sr, trdaddrp0_hr, errRDADDRP0);
  $setuphold(posedge ckrdp0, negedge rdaddrp0[0], trdaddrp0_sf, trdaddrp0_hf, errRDADDRP0);

  $setuphold(posedge ckrdp1, posedge rdaddrp1[5], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[5], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[4], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[4], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[3], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[3], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[2], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[2], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[1], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[1], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);
  $setuphold(posedge ckrdp1, posedge rdaddrp1[0], trdaddrp1_sr, trdaddrp1_hr, errRDADDRP1);
  $setuphold(posedge ckrdp1, negedge rdaddrp1[0], trdaddrp1_sf, trdaddrp1_hf, errRDADDRP1);


  //wren
  $setuphold(posedge ckwrp0, posedge wrenp0, twrenp0_sr, twrenp0_hr, errWRENP0);
  $setuphold(posedge ckwrp0, negedge wrenp0, twrenp0_sf, twrenp0_hf, errWRENP0);

  $setuphold(posedge ckwrp1, posedge wrenp1, twrenp1_sr, twrenp1_hr, errWRENP1);
  $setuphold(posedge ckwrp1, negedge wrenp1, twrenp1_sf, twrenp1_hf, errWRENP1);

 
  //wraddr
  $setuphold(posedge ckwrp0, posedge wraddrp0[5], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[5], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[4], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[4], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[3], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[3], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[2], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[2], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[1], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[1], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);
  $setuphold(posedge ckwrp0, posedge wraddrp0[0], twraddrp0_sr, twraddrp0_hr, errWRADDRP0);
  $setuphold(posedge ckwrp0, negedge wraddrp0[0], twraddrp0_sf, twraddrp0_hf, errWRADDRP0);

  $setuphold(posedge ckwrp1, posedge wraddrp1[5], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[5], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[4], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[4], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[3], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[3], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[2], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[2], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[1], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[1], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);
  $setuphold(posedge ckwrp1, posedge wraddrp1[0], twraddrp1_sr, twraddrp1_hr, errWRADDRP1);
  $setuphold(posedge ckwrp1, negedge wraddrp1[0], twraddrp1_sf, twraddrp1_hf, errWRADDRP1);

  
  //wrdata
  $setuphold(posedge ckwrp0, posedge wrdatap0[159], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[159], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[158], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[158], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[157], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[157], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[156], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[156], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[155], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[155], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[154], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[154], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[153], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[153], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[152], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[152], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[151], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[151], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[150], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[150], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[149], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[149], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[148], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[148], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[147], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[147], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[146], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[146], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[145], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[145], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[144], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[144], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[143], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[143], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[142], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[142], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[141], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[141], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[140], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[140], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[139], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[139], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[138], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[138], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[137], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[137], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[136], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[136], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[135], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[135], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[134], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[134], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[133], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[133], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[132], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[132], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[131], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[131], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[130], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[130], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[129], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[129], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[128], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[128], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[127], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[127], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[126], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[126], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[125], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[125], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[124], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[124], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[123], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[123], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[122], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[122], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[121], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[121], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[120], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[120], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[119], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[119], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[118], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[118], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[117], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[117], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[116], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[116], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[115], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[115], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[114], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[114], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[113], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[113], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[112], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[112], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[111], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[111], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[110], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[110], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[109], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[109], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[108], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[108], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[107], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[107], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[106], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[106], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[105], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[105], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[104], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[104], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[103], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[103], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[102], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[102], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[101], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[101], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[100], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[100], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[99], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[99], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[98], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[98], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[97], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[97], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[96], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[96], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[95], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[95], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[94], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[94], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[93], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[93], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[92], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[92], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[91], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[91], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[90], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[90], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[89], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[89], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[88], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[88], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[87], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[87], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[86], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[86], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[85], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[85], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[84], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[84], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[83], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[83], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[82], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[82], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[81], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[81], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[80], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[80], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[79], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[79], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[78], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[78], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[77], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[77], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[76], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[76], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[75], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[75], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[74], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[74], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[73], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[73], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[72], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[72], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[71], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[71], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[70], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[70], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[69], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[69], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[68], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[68], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[67], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[67], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[66], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[66], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[65], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[65], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[64], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[64], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[63], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[63], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[62], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[62], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[61], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[61], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[60], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[60], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[59], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[59], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[58], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[58], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[57], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[57], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[56], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[56], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[55], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[55], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[54], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[54], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[53], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[53], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[52], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[52], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[51], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[51], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[50], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[50], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[49], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[49], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[48], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[48], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[47], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[47], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[46], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[46], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[45], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[45], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[44], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[44], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[43], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[43], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[42], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[42], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[41], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[41], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[40], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[40], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[39], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[39], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[38], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[38], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[37], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[37], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[36], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[36], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[35], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[35], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[34], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[34], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[33], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[33], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[32], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[32], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[31], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[31], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[30], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[30], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[29], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[29], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[28], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[28], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[27], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[27], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[26], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[26], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[25], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[25], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[24], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[24], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[23], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[23], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[22], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[22], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[21], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[21], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[20], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[20], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[19], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[19], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[18], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[18], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[17], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[17], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[16], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[16], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[15], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[15], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[14], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[14], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[13], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[13], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[12], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[12], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[11], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[11], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[10], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[10], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[9], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[9], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[8], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[8], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[7], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[7], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[6], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[6], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[5], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[5], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[4], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[4], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[3], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[3], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[2], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[2], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[1], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[1], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);
  $setuphold(posedge ckwrp0, posedge wrdatap0[0], twrdatap0_sr, twrdatap0_hr, errWRDATAP0);
  $setuphold(posedge ckwrp0, negedge wrdatap0[0], twrdatap0_sf, twrdatap0_hf, errWRDATAP0);

  $setuphold(posedge ckwrp1, posedge wrdatap1[159], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[159], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[158], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[158], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[157], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[157], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[156], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[156], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[155], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[155], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[154], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[154], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[153], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[153], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[152], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[152], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[151], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[151], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[150], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[150], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[149], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[149], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[148], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[148], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[147], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[147], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[146], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[146], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[145], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[145], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[144], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[144], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[143], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[143], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[142], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[142], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[141], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[141], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[140], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[140], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[139], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[139], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[138], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[138], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[137], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[137], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[136], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[136], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[135], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[135], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[134], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[134], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[133], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[133], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[132], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[132], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[131], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[131], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[130], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[130], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[129], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[129], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[128], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[128], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[127], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[127], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[126], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[126], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[125], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[125], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[124], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[124], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[123], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[123], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[122], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[122], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[121], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[121], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[120], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[120], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[119], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[119], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[118], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[118], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[117], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[117], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[116], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[116], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[115], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[115], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[114], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[114], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[113], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[113], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[112], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[112], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[111], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[111], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[110], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[110], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[109], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[109], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[108], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[108], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[107], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[107], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[106], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[106], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[105], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[105], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[104], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[104], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[103], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[103], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[102], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[102], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[101], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[101], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[100], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[100], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[99], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[99], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[98], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[98], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[97], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[97], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[96], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[96], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[95], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[95], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[94], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[94], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[93], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[93], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[92], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[92], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[91], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[91], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[90], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[90], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[89], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[89], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[88], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[88], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[87], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[87], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[86], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[86], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[85], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[85], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[84], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[84], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[83], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[83], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[82], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[82], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[81], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[81], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[80], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[80], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[79], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[79], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[78], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[78], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[77], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[77], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[76], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[76], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[75], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[75], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[74], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[74], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[73], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[73], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[72], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[72], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[71], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[71], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[70], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[70], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[69], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[69], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[68], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[68], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[67], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[67], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[66], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[66], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[65], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[65], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[64], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[64], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[63], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[63], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[62], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[62], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[61], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[61], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[60], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[60], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[59], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[59], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[58], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[58], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[57], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[57], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[56], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[56], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[55], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[55], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[54], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[54], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[53], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[53], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[52], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[52], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[51], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[51], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[50], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[50], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[49], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[49], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[48], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[48], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[47], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[47], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[46], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[46], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[45], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[45], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[44], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[44], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[43], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[43], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[42], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[42], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[41], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[41], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[40], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[40], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[39], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[39], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[38], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[38], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[37], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[37], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[36], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[36], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[35], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[35], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[34], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[34], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[33], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[33], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[32], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[32], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[31], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[31], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[30], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[30], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[29], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[29], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[28], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[28], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[27], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[27], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[26], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[26], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[25], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[25], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[24], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[24], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[23], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[23], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[22], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[22], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[21], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[21], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[20], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[20], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[19], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[19], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[18], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[18], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[17], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[17], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[16], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[16], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[15], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[15], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[14], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[14], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[13], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[13], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[12], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[12], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[11], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[11], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[10], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[10], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[9], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[9], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[8], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[8], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[7], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[7], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[6], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[6], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[5], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[5], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[4], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[4], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[3], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[3], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[2], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[2], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[1], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[1], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);
  $setuphold(posedge ckwrp1, posedge wrdatap1[0], twrdatap1_sr, twrdatap1_hr, errWRDATAP1);
  $setuphold(posedge ckwrp1, negedge wrdatap1[0], twrdatap1_sf, twrdatap1_hf, errWRDATAP1);


  //q 
  (posedge ckrdp0 => rddatap0[159]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[158]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[157]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[156]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[155]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[154]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[153]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[152]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[151]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[150]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[149]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[148]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[147]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[146]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[145]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[144]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[143]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[142]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[141]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[140]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[139]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[138]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[137]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[136]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[135]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[134]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[133]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[132]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[131]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[130]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[129]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[128]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[127]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[126]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[125]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[124]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[123]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[122]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[121]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[120]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[119]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[118]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[117]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[116]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[115]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[114]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[113]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[112]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[111]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[110]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[109]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[108]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[107]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[106]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[105]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[104]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[103]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[102]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[101]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[100]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[99]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[98]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[97]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[96]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[95]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[94]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[93]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[92]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[91]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[90]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[89]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[88]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[87]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[86]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[85]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[84]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[83]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[82]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[81]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[80]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[79]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[78]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[77]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[76]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[75]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[74]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[73]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[72]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[71]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[70]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[69]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[68]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[67]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[66]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[65]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[64]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[63]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[62]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[61]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[60]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[59]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[58]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[57]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[56]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[55]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[54]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[53]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[52]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[51]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[50]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[49]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[48]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[47]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[46]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[45]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[44]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[43]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[42]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[41]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[40]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[39]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[38]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[37]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[36]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[35]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[34]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[33]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[32]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[31]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[30]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[29]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[28]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[27]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[26]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[25]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[24]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[23]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[22]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[21]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[20]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[19]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[18]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[17]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[16]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[15]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[14]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[13]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[12]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[11]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[10]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[9]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[8]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[7]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[6]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[5]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[4]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[3]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[2]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[1]) = (trddatap0_r, trddatap0_f); 
  (posedge ckrdp0 => rddatap0[0]) = (trddatap0_r, trddatap0_f);
 
  (posedge ckrdp1 => rddatap1[159]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[158]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[157]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[156]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[155]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[154]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[153]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[152]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[151]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[150]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[149]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[148]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[147]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[146]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[145]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[144]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[143]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[142]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[141]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[140]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[139]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[138]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[137]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[136]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[135]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[134]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[133]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[132]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[131]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[130]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[129]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[128]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[127]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[126]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[125]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[124]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[123]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[122]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[121]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[120]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[119]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[118]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[117]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[116]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[115]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[114]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[113]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[112]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[111]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[110]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[109]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[108]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[107]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[106]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[105]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[104]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[103]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[102]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[101]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[100]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[99]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[98]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[97]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[96]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[95]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[94]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[93]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[92]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[91]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[90]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[89]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[88]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[87]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[86]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[85]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[84]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[83]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[82]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[81]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[80]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[79]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[78]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[77]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[76]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[75]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[74]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[73]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[72]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[71]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[70]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[69]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[68]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[67]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[66]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[65]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[64]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[63]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[62]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[61]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[60]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[59]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[58]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[57]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[56]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[55]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[54]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[53]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[52]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[51]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[50]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[49]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[48]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[47]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[46]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[45]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[44]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[43]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[42]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[41]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[40]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[39]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[38]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[37]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[36]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[35]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[34]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[33]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[32]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[31]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[30]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[29]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[28]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[27]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[26]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[25]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[24]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[23]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[22]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[21]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[20]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[19]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[18]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[17]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[16]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[15]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[14]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[13]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[12]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[11]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[10]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[9]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[8]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[7]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[6]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[5]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[4]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[3]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[2]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[1]) = (trddatap1_r, trddatap1_f); 
  (posedge ckrdp1 => rddatap1[0]) = (trddatap1_r, trddatap1_f);

endspecify

`endif



endmodule // end module arf156b040e2r2w0cbbehbaa4acw
`endif // endif ifndef ARF156B040E2R2W0CBBEHBAA4ACW_SV
