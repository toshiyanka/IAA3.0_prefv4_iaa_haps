VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf028b032e2r2w0cbbehraa4acw
  CLASS BLOCK ;
  FOREIGN arf028b032e2r2w0cbbehraa4acw ;
  ORIGIN 0 0 ;
  SIZE 18 BY 20.16 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 3.24 0.388 4.44 ;
    END
  END ckrdp0
  PIN ckrdp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 3.24 2.916 4.44 ;
    END
  END ckrdp1
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.344 0.84 0.388 2.04 ;
    END
  END ckwrp0
  PIN ckwrp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 0.84 3.172 2.04 ;
    END
  END ckwrp1
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 3.24 1.628 4.44 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 3.24 1.928 4.44 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 3.24 2.188 4.44 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 3.24 2.356 4.44 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.24 2.616 4.44 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 3.24 0.556 4.44 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 3.24 0.816 4.44 ;
    END
  END rdaddrp0_rd
  PIN rdaddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 3.24 4.156 4.44 ;
    END
  END rdaddrp1[0]
  PIN rdaddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 3.24 4.416 4.44 ;
    END
  END rdaddrp1[1]
  PIN rdaddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 3.24 4.716 4.44 ;
    END
  END rdaddrp1[2]
  PIN rdaddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 3.24 4.972 4.44 ;
    END
  END rdaddrp1[3]
  PIN rdaddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 3.24 5.228 4.44 ;
    END
  END rdaddrp1[4]
  PIN rdaddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 3.24 3.172 4.44 ;
    END
  END rdaddrp1_fd
  PIN rdaddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 3.24 3.428 4.44 ;
    END
  END rdaddrp1_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 3.24 1.116 4.44 ;
    END
  END rdenp0
  PIN rdenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.24 3.728 4.44 ;
    END
  END rdenp1
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 3.24 1.372 4.44 ;
    END
  END sdl_initp0
  PIN sdl_initp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 3.24 3.988 4.44 ;
    END
  END sdl_initp1
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.84 1.928 2.04 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.144 0.84 2.188 2.04 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.312 0.84 2.356 2.04 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 0.84 2.616 2.04 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.84 2.916 2.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.512 0.84 0.556 2.04 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 0.84 0.816 2.04 ;
    END
  END wraddrp0_rd
  PIN wraddrp1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 0.84 4.716 2.04 ;
    END
  END wraddrp1[0]
  PIN wraddrp1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 0.84 4.972 2.04 ;
    END
  END wraddrp1[1]
  PIN wraddrp1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.184 0.84 5.228 2.04 ;
    END
  END wraddrp1[2]
  PIN wraddrp1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 0.84 5.528 2.04 ;
    END
  END wraddrp1[3]
  PIN wraddrp1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 0.84 5.788 2.04 ;
    END
  END wraddrp1[4]
  PIN wraddrp1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.84 3.428 2.04 ;
    END
  END wraddrp1_fd
  PIN wraddrp1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.84 3.728 2.04 ;
    END
  END wraddrp1_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 5.16 3.256 6.36 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 9.96 4.888 11.16 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 9.96 4.972 11.16 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 10.92 4.156 12.12 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 10.92 4.328 12.12 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 11.88 3.728 13.08 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 11.88 3.816 13.08 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 12.84 3.428 14.04 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 12.84 3.516 14.04 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 13.8 4.972 15 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 13.8 3.172 15 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.16 3.516 6.36 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 14.76 4.416 15.96 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 14.76 4.628 15.96 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 15.72 3.728 16.92 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 15.72 3.816 16.92 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 16.68 3.428 17.88 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.68 3.516 17.88 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 17.64 4.972 18.84 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 17.64 3.172 18.84 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 18.6 4.416 19.8 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 18.6 4.628 19.8 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 6.12 4.716 7.32 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 6.12 4.888 7.32 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 7.08 3.988 8.28 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 7.08 4.072 8.28 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.04 3.516 9.24 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 8.04 3.728 9.24 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 9 3.256 10.2 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9 3.428 10.2 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 0.84 1.372 2.04 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 0.84 1.628 2.04 ;
    END
  END wrdatap0_rd
  PIN wrdatap1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 5.16 3.816 6.36 ;
    END
  END wrdatap1[0]
  PIN wrdatap1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 9.96 3.172 11.16 ;
    END
  END wrdatap1[10]
  PIN wrdatap1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 9.96 3.516 11.16 ;
    END
  END wrdatap1[11]
  PIN wrdatap1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 10.92 4.416 12.12 ;
    END
  END wrdatap1[12]
  PIN wrdatap1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.584 10.92 4.628 12.12 ;
    END
  END wrdatap1[13]
  PIN wrdatap1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 11.88 3.988 13.08 ;
    END
  END wrdatap1[14]
  PIN wrdatap1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 11.88 4.072 13.08 ;
    END
  END wrdatap1[15]
  PIN wrdatap1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 12.84 4.156 14.04 ;
    END
  END wrdatap1[16]
  PIN wrdatap1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 12.84 4.328 14.04 ;
    END
  END wrdatap1[17]
  PIN wrdatap1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 13.8 3.256 15 ;
    END
  END wrdatap1[18]
  PIN wrdatap1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 13.8 3.728 15 ;
    END
  END wrdatap1[19]
  PIN wrdatap1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 5.16 4.072 6.36 ;
    END
  END wrdatap1[1]
  PIN wrdatap1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 14.76 4.716 15.96 ;
    END
  END wrdatap1[20]
  PIN wrdatap1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 14.76 4.888 15.96 ;
    END
  END wrdatap1[21]
  PIN wrdatap1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 15.72 3.988 16.92 ;
    END
  END wrdatap1[22]
  PIN wrdatap1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 15.72 4.072 16.92 ;
    END
  END wrdatap1[23]
  PIN wrdatap1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 16.68 4.156 17.88 ;
    END
  END wrdatap1[24]
  PIN wrdatap1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 16.68 4.328 17.88 ;
    END
  END wrdatap1[25]
  PIN wrdatap1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.212 17.64 3.256 18.84 ;
    END
  END wrdatap1[26]
  PIN wrdatap1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 17.64 3.728 18.84 ;
    END
  END wrdatap1[27]
  PIN wrdatap1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.672 18.6 4.716 19.8 ;
    END
  END wrdatap1[28]
  PIN wrdatap1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.844 18.6 4.888 19.8 ;
    END
  END wrdatap1[29]
  PIN wrdatap1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.928 6.12 4.972 7.32 ;
    END
  END wrdatap1[2]
  PIN wrdatap1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 6.12 3.172 7.32 ;
    END
  END wrdatap1[3]
  PIN wrdatap1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 7.08 4.156 8.28 ;
    END
  END wrdatap1[4]
  PIN wrdatap1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 7.08 4.328 8.28 ;
    END
  END wrdatap1[5]
  PIN wrdatap1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 8.04 3.816 9.24 ;
    END
  END wrdatap1[6]
  PIN wrdatap1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 8.04 4.416 9.24 ;
    END
  END wrdatap1[7]
  PIN wrdatap1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 9 3.988 10.2 ;
    END
  END wrdatap1[8]
  PIN wrdatap1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 9 4.072 10.2 ;
    END
  END wrdatap1[9]
  PIN wrdatap1_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.112 0.84 4.156 2.04 ;
    END
  END wrdatap1_fd
  PIN wrdatap1_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.372 0.84 4.416 2.04 ;
    END
  END wrdatap1_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 0.84 1.116 2.04 ;
    END
  END wrenp0
  PIN wrenp1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.944 0.84 3.988 2.04 ;
    END
  END wrenp1
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 5.16 5.956 6.36 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 9.96 5.616 11.16 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 9.96 5.788 11.16 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 10.92 5.316 12.12 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 10.92 5.528 12.12 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 11.88 6.856 13.08 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 11.88 7.028 13.08 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 12.84 6.428 14.04 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 12.84 6.516 14.04 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 13.8 5.788 15 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 13.8 5.872 15 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 5.16 6.128 6.36 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 14.76 5.316 15.96 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 14.76 5.528 15.96 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 15.72 6.856 16.92 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 15.72 7.028 16.92 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 16.68 6.428 17.88 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 16.68 6.516 17.88 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 17.64 5.788 18.84 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 17.64 5.872 18.84 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 18.6 5.316 19.8 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 18.6 5.528 19.8 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 6.12 5.528 7.32 ;
    END
  END rddatap0[2]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 6.12 5.616 7.32 ;
    END
  END rddatap0[3]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.984 7.08 7.028 8.28 ;
    END
  END rddatap0[4]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.272 7.08 5.316 8.28 ;
    END
  END rddatap0[5]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 8.04 6.688 9.24 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 8.04 6.772 9.24 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 9 6.128 10.2 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 9 6.216 10.2 ;
    END
  END rddatap0[9]
  PIN rddatap1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 5.16 6.216 6.36 ;
    END
  END rddatap1[0]
  PIN rddatap1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 9.96 5.872 11.16 ;
    END
  END rddatap1[10]
  PIN rddatap1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 9.96 5.956 11.16 ;
    END
  END rddatap1[11]
  PIN rddatap1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 10.92 6.128 12.12 ;
    END
  END rddatap1[12]
  PIN rddatap1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 10.92 6.216 12.12 ;
    END
  END rddatap1[13]
  PIN rddatap1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 11.88 5.616 13.08 ;
    END
  END rddatap1[14]
  PIN rddatap1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 11.88 5.788 13.08 ;
    END
  END rddatap1[15]
  PIN rddatap1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 12.84 6.688 14.04 ;
    END
  END rddatap1[16]
  PIN rddatap1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 12.84 6.772 14.04 ;
    END
  END rddatap1[17]
  PIN rddatap1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 13.8 5.956 15 ;
    END
  END rddatap1[18]
  PIN rddatap1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 13.8 6.128 15 ;
    END
  END rddatap1[19]
  PIN rddatap1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 5.16 6.428 6.36 ;
    END
  END rddatap1[1]
  PIN rddatap1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 14.76 5.616 15.96 ;
    END
  END rddatap1[20]
  PIN rddatap1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 14.76 6.216 15.96 ;
    END
  END rddatap1[21]
  PIN rddatap1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 15.72 5.788 16.92 ;
    END
  END rddatap1[22]
  PIN rddatap1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 15.72 5.872 16.92 ;
    END
  END rddatap1[23]
  PIN rddatap1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.644 16.68 6.688 17.88 ;
    END
  END rddatap1[24]
  PIN rddatap1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.728 16.68 6.772 17.88 ;
    END
  END rddatap1[25]
  PIN rddatap1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 17.64 5.956 18.84 ;
    END
  END rddatap1[26]
  PIN rddatap1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 17.64 6.128 18.84 ;
    END
  END rddatap1[27]
  PIN rddatap1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.572 18.6 5.616 19.8 ;
    END
  END rddatap1[28]
  PIN rddatap1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.172 18.6 6.216 19.8 ;
    END
  END rddatap1[29]
  PIN rddatap1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.744 6.12 5.788 7.32 ;
    END
  END rddatap1[2]
  PIN rddatap1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.828 6.12 5.872 7.32 ;
    END
  END rddatap1[3]
  PIN rddatap1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.912 7.08 5.956 8.28 ;
    END
  END rddatap1[4]
  PIN rddatap1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.084 7.08 6.128 8.28 ;
    END
  END rddatap1[5]
  PIN rddatap1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.812 8.04 6.856 9.24 ;
    END
  END rddatap1[6]
  PIN rddatap1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 5.484 8.04 5.528 9.24 ;
    END
  END rddatap1[7]
  PIN rddatap1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.384 9 6.428 10.2 ;
    END
  END rddatap1[8]
  PIN rddatap1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 6.472 9 6.516 10.2 ;
    END
  END rddatap1[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 20.1 ;
        RECT 2.662 0.06 2.738 20.1 ;
        RECT 4.462 0.06 4.538 20.1 ;
        RECT 6.262 0.06 6.338 20.1 ;
        RECT 8.062 0.06 8.138 20.1 ;
        RECT 9.862 0.06 9.938 20.1 ;
        RECT 11.662 0.06 11.738 20.1 ;
        RECT 13.462 0.06 13.538 20.1 ;
        RECT 15.262 0.06 15.338 20.1 ;
        RECT 17.062 0.06 17.138 20.1 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 20.1 ;
        RECT 3.562 0.06 3.638 20.1 ;
        RECT 5.362 0.06 5.438 20.1 ;
        RECT 7.162 0.06 7.238 20.1 ;
        RECT 8.962 0.06 9.038 20.1 ;
        RECT 10.762 0.06 10.838 20.1 ;
        RECT 12.562 0.06 12.638 20.1 ;
        RECT 14.362 0.06 14.438 20.1 ;
        RECT 16.162 0.06 16.238 20.1 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 18.016 20.174 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 18.02 20.18 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 18.0705 20.198 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 18.035 20.23 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 18.07 20.198 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 18.059 20.25 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 18.09 20.222 ;
    LAYER m7 SPACING 0 ;
      RECT 17.138 20.22 18.04 20.28 ;
      RECT 17.138 -0.06 18.092 20.22 ;
      RECT 17.138 -0.12 18.04 -0.06 ;
      RECT 16.238 -0.12 17.062 20.28 ;
      RECT 15.338 -0.12 16.162 20.28 ;
      RECT 14.438 -0.12 15.262 20.28 ;
      RECT 13.538 -0.12 14.362 20.28 ;
      RECT 12.638 -0.12 13.462 20.28 ;
      RECT 11.738 -0.12 12.562 20.28 ;
      RECT 10.838 -0.12 11.662 20.28 ;
      RECT 9.938 -0.12 10.762 20.28 ;
      RECT 9.038 -0.12 9.862 20.28 ;
      RECT 8.138 -0.12 8.962 20.28 ;
      RECT 7.238 -0.12 8.062 20.28 ;
      RECT 6.338 17.88 7.162 20.28 ;
      RECT 6.772 16.92 7.162 17.88 ;
      RECT 6.338 16.68 6.384 17.88 ;
      RECT 6.428 16.68 6.472 17.88 ;
      RECT 6.516 16.68 6.644 17.88 ;
      RECT 6.688 16.68 6.728 17.88 ;
      RECT 6.772 16.68 6.812 16.92 ;
      RECT 6.856 15.72 6.984 16.92 ;
      RECT 7.028 15.72 7.162 16.92 ;
      RECT 6.338 15.72 6.812 16.68 ;
      RECT 6.338 14.04 7.162 15.72 ;
      RECT 6.772 13.08 7.162 14.04 ;
      RECT 6.338 12.84 6.384 14.04 ;
      RECT 6.428 12.84 6.472 14.04 ;
      RECT 6.516 12.84 6.644 14.04 ;
      RECT 6.688 12.84 6.728 14.04 ;
      RECT 6.772 12.84 6.812 13.08 ;
      RECT 6.856 11.88 6.984 13.08 ;
      RECT 7.028 11.88 7.162 13.08 ;
      RECT 6.338 11.88 6.812 12.84 ;
      RECT 6.338 10.2 7.162 11.88 ;
      RECT 6.516 9.24 7.162 10.2 ;
      RECT 6.338 9 6.384 10.2 ;
      RECT 6.428 9 6.472 10.2 ;
      RECT 6.516 9 6.644 9.24 ;
      RECT 6.856 8.28 7.162 9.24 ;
      RECT 6.688 8.04 6.728 9.24 ;
      RECT 6.772 8.04 6.812 9.24 ;
      RECT 6.338 8.04 6.644 9 ;
      RECT 6.856 8.04 6.984 8.28 ;
      RECT 7.028 7.08 7.162 8.28 ;
      RECT 6.338 7.08 6.984 8.04 ;
      RECT 6.338 6.36 7.162 7.08 ;
      RECT 6.338 5.16 6.384 6.36 ;
      RECT 6.428 5.16 7.162 6.36 ;
      RECT 6.338 -0.12 7.162 5.16 ;
      RECT 5.438 19.8 6.262 20.28 ;
      RECT 5.616 18.84 6.172 19.8 ;
      RECT 5.438 18.6 5.484 19.8 ;
      RECT 5.528 18.6 5.572 19.8 ;
      RECT 6.216 18.6 6.262 19.8 ;
      RECT 5.616 18.6 5.744 18.84 ;
      RECT 6.128 18.6 6.172 18.84 ;
      RECT 5.788 17.64 5.828 18.84 ;
      RECT 5.872 17.64 5.912 18.84 ;
      RECT 5.956 17.64 6.084 18.84 ;
      RECT 5.438 17.64 5.744 18.6 ;
      RECT 6.128 17.64 6.262 18.6 ;
      RECT 5.438 16.92 6.262 17.64 ;
      RECT 5.438 15.96 5.744 16.92 ;
      RECT 5.872 15.96 6.262 16.92 ;
      RECT 5.788 15.72 5.828 16.92 ;
      RECT 5.616 15.72 5.744 15.96 ;
      RECT 5.872 15.72 6.172 15.96 ;
      RECT 5.616 15 6.172 15.72 ;
      RECT 5.438 14.76 5.484 15.96 ;
      RECT 5.528 14.76 5.572 15.96 ;
      RECT 6.216 14.76 6.262 15.96 ;
      RECT 5.616 14.76 5.744 15 ;
      RECT 6.128 14.76 6.172 15 ;
      RECT 5.788 13.8 5.828 15 ;
      RECT 5.872 13.8 5.912 15 ;
      RECT 5.956 13.8 6.084 15 ;
      RECT 5.438 13.8 5.744 14.76 ;
      RECT 6.128 13.8 6.262 14.76 ;
      RECT 5.438 13.08 6.262 13.8 ;
      RECT 5.438 12.12 5.572 13.08 ;
      RECT 5.788 12.12 6.262 13.08 ;
      RECT 5.616 11.88 5.744 13.08 ;
      RECT 5.528 11.88 5.572 12.12 ;
      RECT 5.788 11.88 6.084 12.12 ;
      RECT 5.528 11.16 6.084 11.88 ;
      RECT 5.438 10.92 5.484 12.12 ;
      RECT 6.128 10.92 6.172 12.12 ;
      RECT 6.216 10.92 6.262 12.12 ;
      RECT 5.528 10.92 5.572 11.16 ;
      RECT 5.956 10.92 6.084 11.16 ;
      RECT 5.956 10.2 6.262 10.92 ;
      RECT 5.616 9.96 5.744 11.16 ;
      RECT 5.788 9.96 5.828 11.16 ;
      RECT 5.872 9.96 5.912 11.16 ;
      RECT 5.438 9.96 5.572 10.92 ;
      RECT 5.956 9.96 6.084 10.2 ;
      RECT 5.438 9.24 6.084 9.96 ;
      RECT 6.128 9 6.172 10.2 ;
      RECT 6.216 9 6.262 10.2 ;
      RECT 5.528 9 6.084 9.24 ;
      RECT 5.528 8.28 6.262 9 ;
      RECT 5.438 8.04 5.484 9.24 ;
      RECT 5.528 8.04 5.912 8.28 ;
      RECT 5.438 7.32 5.912 8.04 ;
      RECT 5.956 7.08 6.084 8.28 ;
      RECT 6.128 7.08 6.262 8.28 ;
      RECT 5.872 7.08 5.912 7.32 ;
      RECT 5.872 6.36 6.262 7.08 ;
      RECT 5.438 6.12 5.484 7.32 ;
      RECT 5.528 6.12 5.572 7.32 ;
      RECT 5.616 6.12 5.744 7.32 ;
      RECT 5.788 6.12 5.828 7.32 ;
      RECT 5.872 6.12 5.912 6.36 ;
      RECT 5.956 5.16 6.084 6.36 ;
      RECT 6.128 5.16 6.172 6.36 ;
      RECT 6.216 5.16 6.262 6.36 ;
      RECT 5.438 5.16 5.912 6.12 ;
      RECT 5.438 2.04 6.262 5.16 ;
      RECT 5.438 0.84 5.484 2.04 ;
      RECT 5.528 0.84 5.744 2.04 ;
      RECT 5.788 0.84 6.262 2.04 ;
      RECT 5.438 -0.12 6.262 0.84 ;
      RECT 4.538 19.8 5.362 20.28 ;
      RECT 4.888 18.84 5.272 19.8 ;
      RECT 4.538 18.6 4.584 19.8 ;
      RECT 4.628 18.6 4.672 19.8 ;
      RECT 4.716 18.6 4.844 19.8 ;
      RECT 5.316 18.6 5.362 19.8 ;
      RECT 4.888 18.6 4.928 18.84 ;
      RECT 4.972 18.6 5.272 18.84 ;
      RECT 4.538 17.64 4.928 18.6 ;
      RECT 4.972 17.64 5.362 18.6 ;
      RECT 4.538 15.96 5.362 17.64 ;
      RECT 4.888 15 5.272 15.96 ;
      RECT 4.538 14.76 4.584 15.96 ;
      RECT 4.628 14.76 4.672 15.96 ;
      RECT 4.716 14.76 4.844 15.96 ;
      RECT 5.316 14.76 5.362 15.96 ;
      RECT 4.888 14.76 4.928 15 ;
      RECT 4.972 14.76 5.272 15 ;
      RECT 4.538 13.8 4.928 14.76 ;
      RECT 4.972 13.8 5.362 14.76 ;
      RECT 4.538 12.12 5.362 13.8 ;
      RECT 4.628 11.16 5.272 12.12 ;
      RECT 4.538 10.92 4.584 12.12 ;
      RECT 5.316 10.92 5.362 12.12 ;
      RECT 4.628 10.92 4.844 11.16 ;
      RECT 4.972 10.92 5.272 11.16 ;
      RECT 4.888 9.96 4.928 11.16 ;
      RECT 4.538 9.96 4.844 10.92 ;
      RECT 4.972 9.96 5.362 10.92 ;
      RECT 4.538 8.28 5.362 9.96 ;
      RECT 4.538 7.32 5.272 8.28 ;
      RECT 5.316 7.08 5.362 8.28 ;
      RECT 4.972 7.08 5.272 7.32 ;
      RECT 4.538 6.12 4.672 7.32 ;
      RECT 4.716 6.12 4.844 7.32 ;
      RECT 4.888 6.12 4.928 7.32 ;
      RECT 4.972 6.12 5.362 7.08 ;
      RECT 4.538 4.44 5.362 6.12 ;
      RECT 4.538 3.24 4.672 4.44 ;
      RECT 4.716 3.24 4.928 4.44 ;
      RECT 4.972 3.24 5.184 4.44 ;
      RECT 5.228 3.24 5.362 4.44 ;
      RECT 4.538 2.04 5.362 3.24 ;
      RECT 4.538 0.84 4.672 2.04 ;
      RECT 4.716 0.84 4.928 2.04 ;
      RECT 4.972 0.84 5.184 2.04 ;
      RECT 5.228 0.84 5.362 2.04 ;
      RECT 4.538 -0.12 5.362 0.84 ;
      RECT 3.638 19.8 4.462 20.28 ;
      RECT 3.638 18.84 4.372 19.8 ;
      RECT 4.416 18.6 4.462 19.8 ;
      RECT 3.728 18.6 4.372 18.84 ;
      RECT 3.728 17.88 4.462 18.6 ;
      RECT 3.638 17.64 3.684 18.84 ;
      RECT 3.728 17.64 4.112 17.88 ;
      RECT 3.638 16.92 4.112 17.64 ;
      RECT 4.156 16.68 4.284 17.88 ;
      RECT 4.328 16.68 4.462 17.88 ;
      RECT 4.072 16.68 4.112 16.92 ;
      RECT 4.072 15.96 4.462 16.68 ;
      RECT 3.638 15.72 3.684 16.92 ;
      RECT 3.728 15.72 3.772 16.92 ;
      RECT 3.816 15.72 3.944 16.92 ;
      RECT 3.988 15.72 4.028 16.92 ;
      RECT 4.072 15.72 4.372 15.96 ;
      RECT 3.638 15 4.372 15.72 ;
      RECT 4.416 14.76 4.462 15.96 ;
      RECT 3.728 14.76 4.372 15 ;
      RECT 3.728 14.04 4.462 14.76 ;
      RECT 3.638 13.8 3.684 15 ;
      RECT 3.728 13.8 4.112 14.04 ;
      RECT 3.638 13.08 4.112 13.8 ;
      RECT 4.156 12.84 4.284 14.04 ;
      RECT 4.328 12.84 4.462 14.04 ;
      RECT 4.072 12.84 4.112 13.08 ;
      RECT 4.072 12.12 4.462 12.84 ;
      RECT 3.638 11.88 3.684 13.08 ;
      RECT 3.728 11.88 3.772 13.08 ;
      RECT 3.816 11.88 3.944 13.08 ;
      RECT 3.988 11.88 4.028 13.08 ;
      RECT 4.072 11.88 4.112 12.12 ;
      RECT 4.156 10.92 4.284 12.12 ;
      RECT 4.328 10.92 4.372 12.12 ;
      RECT 4.416 10.92 4.462 12.12 ;
      RECT 3.638 10.92 4.112 11.88 ;
      RECT 3.638 10.2 4.462 10.92 ;
      RECT 3.638 9.24 3.944 10.2 ;
      RECT 4.072 9.24 4.462 10.2 ;
      RECT 3.988 9 4.028 10.2 ;
      RECT 3.816 9 3.944 9.24 ;
      RECT 4.072 9 4.372 9.24 ;
      RECT 3.816 8.28 4.372 9 ;
      RECT 3.638 8.04 3.684 9.24 ;
      RECT 3.728 8.04 3.772 9.24 ;
      RECT 4.416 8.04 4.462 9.24 ;
      RECT 3.816 8.04 3.944 8.28 ;
      RECT 4.328 8.04 4.372 8.28 ;
      RECT 3.988 7.08 4.028 8.28 ;
      RECT 4.072 7.08 4.112 8.28 ;
      RECT 4.156 7.08 4.284 8.28 ;
      RECT 3.638 7.08 3.944 8.04 ;
      RECT 4.328 7.08 4.462 8.04 ;
      RECT 3.638 6.36 4.462 7.08 ;
      RECT 3.638 5.16 3.772 6.36 ;
      RECT 3.816 5.16 4.028 6.36 ;
      RECT 4.072 5.16 4.462 6.36 ;
      RECT 3.638 4.44 4.462 5.16 ;
      RECT 3.638 3.24 3.684 4.44 ;
      RECT 3.728 3.24 3.944 4.44 ;
      RECT 3.988 3.24 4.112 4.44 ;
      RECT 4.156 3.24 4.372 4.44 ;
      RECT 4.416 3.24 4.462 4.44 ;
      RECT 3.638 2.04 4.462 3.24 ;
      RECT 3.638 0.84 3.684 2.04 ;
      RECT 3.728 0.84 3.944 2.04 ;
      RECT 3.988 0.84 4.112 2.04 ;
      RECT 4.156 0.84 4.372 2.04 ;
      RECT 4.416 0.84 4.462 2.04 ;
      RECT 3.638 -0.12 4.462 0.84 ;
      RECT 2.738 18.84 3.562 20.28 ;
      RECT 3.256 17.88 3.562 18.84 ;
      RECT 2.738 17.64 3.128 18.84 ;
      RECT 3.172 17.64 3.212 18.84 ;
      RECT 3.256 17.64 3.384 17.88 ;
      RECT 3.428 16.68 3.472 17.88 ;
      RECT 3.516 16.68 3.562 17.88 ;
      RECT 2.738 16.68 3.384 17.64 ;
      RECT 2.738 15 3.562 16.68 ;
      RECT 3.256 14.04 3.562 15 ;
      RECT 2.738 13.8 3.128 15 ;
      RECT 3.172 13.8 3.212 15 ;
      RECT 3.256 13.8 3.384 14.04 ;
      RECT 3.428 12.84 3.472 14.04 ;
      RECT 3.516 12.84 3.562 14.04 ;
      RECT 2.738 12.84 3.384 13.8 ;
      RECT 2.738 11.16 3.562 12.84 ;
      RECT 3.172 10.2 3.472 11.16 ;
      RECT 2.738 9.96 3.128 11.16 ;
      RECT 3.516 9.96 3.562 11.16 ;
      RECT 3.172 9.96 3.212 10.2 ;
      RECT 3.428 9.96 3.472 10.2 ;
      RECT 3.428 9.24 3.562 9.96 ;
      RECT 3.256 9 3.384 10.2 ;
      RECT 2.738 9 3.212 9.96 ;
      RECT 3.428 9 3.472 9.24 ;
      RECT 3.516 8.04 3.562 9.24 ;
      RECT 2.738 8.04 3.472 9 ;
      RECT 2.738 7.32 3.562 8.04 ;
      RECT 3.172 6.36 3.562 7.32 ;
      RECT 2.738 6.12 3.128 7.32 ;
      RECT 3.172 6.12 3.212 6.36 ;
      RECT 3.256 5.16 3.472 6.36 ;
      RECT 3.516 5.16 3.562 6.36 ;
      RECT 2.738 5.16 3.212 6.12 ;
      RECT 2.738 4.44 3.562 5.16 ;
      RECT 2.738 3.24 2.872 4.44 ;
      RECT 2.916 3.24 3.128 4.44 ;
      RECT 3.172 3.24 3.384 4.44 ;
      RECT 3.428 3.24 3.562 4.44 ;
      RECT 2.738 2.04 3.562 3.24 ;
      RECT 2.738 0.84 2.872 2.04 ;
      RECT 2.916 0.84 3.128 2.04 ;
      RECT 3.172 0.84 3.384 2.04 ;
      RECT 3.428 0.84 3.562 2.04 ;
      RECT 2.738 -0.12 3.562 0.84 ;
      RECT 1.838 4.44 2.662 20.28 ;
      RECT 1.838 3.24 1.884 4.44 ;
      RECT 1.928 3.24 2.144 4.44 ;
      RECT 2.188 3.24 2.312 4.44 ;
      RECT 2.356 3.24 2.572 4.44 ;
      RECT 2.616 3.24 2.662 4.44 ;
      RECT 1.838 2.04 2.662 3.24 ;
      RECT 1.838 0.84 1.884 2.04 ;
      RECT 1.928 0.84 2.144 2.04 ;
      RECT 2.188 0.84 2.312 2.04 ;
      RECT 2.356 0.84 2.572 2.04 ;
      RECT 2.616 0.84 2.662 2.04 ;
      RECT 1.838 -0.12 2.662 0.84 ;
      RECT 0.938 4.44 1.762 20.28 ;
      RECT 0.938 3.24 1.072 4.44 ;
      RECT 1.116 3.24 1.328 4.44 ;
      RECT 1.372 3.24 1.584 4.44 ;
      RECT 1.628 3.24 1.762 4.44 ;
      RECT 0.938 2.04 1.762 3.24 ;
      RECT 0.938 0.84 1.072 2.04 ;
      RECT 1.116 0.84 1.328 2.04 ;
      RECT 1.372 0.84 1.584 2.04 ;
      RECT 1.628 0.84 1.762 2.04 ;
      RECT 0.938 -0.12 1.762 0.84 ;
      RECT -0.04 20.22 0.862 20.28 ;
      RECT -0.092 4.44 0.862 20.22 ;
      RECT -0.092 3.24 0.344 4.44 ;
      RECT 0.388 3.24 0.512 4.44 ;
      RECT 0.556 3.24 0.772 4.44 ;
      RECT 0.816 3.24 0.862 4.44 ;
      RECT -0.092 2.04 0.862 3.24 ;
      RECT -0.092 0.84 0.344 2.04 ;
      RECT 0.388 0.84 0.512 2.04 ;
      RECT 0.556 0.84 0.772 2.04 ;
      RECT 0.816 0.84 0.862 2.04 ;
      RECT -0.092 -0.06 0.862 0.84 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 17.258 0 17.92 20.16 ;
      RECT 16.358 0 16.942 20.16 ;
      RECT 15.458 0 16.042 20.16 ;
      RECT 14.558 0 15.142 20.16 ;
      RECT 13.658 0 14.242 20.16 ;
      RECT 12.758 0 13.342 20.16 ;
      RECT 11.858 0 12.442 20.16 ;
      RECT 10.958 0 11.542 20.16 ;
      RECT 10.058 0 10.642 20.16 ;
      RECT 9.158 0 9.742 20.16 ;
      RECT 8.258 0 8.842 20.16 ;
      RECT 7.358 0 7.942 20.16 ;
      RECT 6.458 18 7.042 20.16 ;
      RECT 6.892 17.04 7.042 18 ;
      RECT 5.558 19.92 6.142 20.16 ;
      RECT 5.736 18.96 6.052 19.92 ;
      RECT 4.658 19.92 5.242 20.16 ;
      RECT 5.008 18.96 5.152 19.92 ;
      RECT 5.092 18.48 5.152 18.96 ;
      RECT 4.658 17.52 4.808 18.48 ;
      RECT 5.092 17.52 5.242 18.48 ;
      RECT 4.658 16.08 5.242 17.52 ;
      RECT 5.008 15.12 5.152 16.08 ;
      RECT 5.092 14.64 5.152 15.12 ;
      RECT 4.658 13.68 4.808 14.64 ;
      RECT 5.092 13.68 5.242 14.64 ;
      RECT 4.658 12.24 5.242 13.68 ;
      RECT 4.748 11.28 5.152 12.24 ;
      RECT 5.092 10.8 5.152 11.28 ;
      RECT 4.658 9.84 4.724 10.8 ;
      RECT 5.092 9.84 5.242 10.8 ;
      RECT 4.658 8.4 5.242 9.84 ;
      RECT 4.658 7.44 5.152 8.4 ;
      RECT 5.092 6.96 5.152 7.44 ;
      RECT 5.092 6 5.242 6.96 ;
      RECT 4.658 4.56 5.242 6 ;
      RECT 3.758 19.92 4.342 20.16 ;
      RECT 3.758 18.96 4.252 19.92 ;
      RECT 3.848 18.48 4.252 18.96 ;
      RECT 3.848 18 4.342 18.48 ;
      RECT 3.848 17.52 3.992 18 ;
      RECT 3.758 17.04 3.992 17.52 ;
      RECT 2.858 18.96 3.442 20.16 ;
      RECT 3.376 18 3.442 18.96 ;
      RECT 2.858 17.52 3.008 18.96 ;
      RECT 2.858 16.56 3.264 17.52 ;
      RECT 2.858 15.12 3.442 16.56 ;
      RECT 3.376 14.16 3.442 15.12 ;
      RECT 2.858 13.68 3.008 15.12 ;
      RECT 2.858 12.72 3.264 13.68 ;
      RECT 2.858 11.28 3.442 12.72 ;
      RECT 3.292 10.32 3.352 11.28 ;
      RECT 2.858 9.84 3.008 11.28 ;
      RECT 2.858 8.88 3.092 9.84 ;
      RECT 2.858 7.92 3.352 8.88 ;
      RECT 2.858 7.44 3.442 7.92 ;
      RECT 3.292 6.48 3.442 7.44 ;
      RECT 2.858 6 3.008 7.44 ;
      RECT 2.858 5.04 3.092 6 ;
      RECT 2.858 4.56 3.442 5.04 ;
      RECT 1.958 4.56 2.542 20.16 ;
      RECT 1.058 4.56 1.642 20.16 ;
      RECT 0.08 4.56 0.742 20.16 ;
      RECT 0.08 3.12 0.224 4.56 ;
      RECT 0.08 2.16 0.742 3.12 ;
      RECT 0.08 0.72 0.224 2.16 ;
      RECT 0.08 0 0.742 0.72 ;
      RECT 5.558 17.52 5.624 18.48 ;
      RECT 5.558 17.04 6.142 17.52 ;
      RECT 5.558 16.08 5.624 17.04 ;
      RECT 5.992 16.08 6.142 17.04 ;
      RECT 5.992 15.6 6.052 16.08 ;
      RECT 5.736 15.12 6.052 15.6 ;
      RECT 6.458 15.6 6.692 16.56 ;
      RECT 6.458 14.16 7.042 15.6 ;
      RECT 6.892 13.2 7.042 14.16 ;
      RECT 4.192 16.08 4.342 16.56 ;
      RECT 4.192 15.6 4.252 16.08 ;
      RECT 3.758 15.12 4.252 15.6 ;
      RECT 3.848 14.64 4.252 15.12 ;
      RECT 3.848 14.16 4.342 14.64 ;
      RECT 3.848 13.68 3.992 14.16 ;
      RECT 3.758 13.2 3.992 13.68 ;
      RECT 5.558 13.68 5.624 14.64 ;
      RECT 5.558 13.2 6.142 13.68 ;
      RECT 5.908 12.24 6.142 13.2 ;
      RECT 5.908 11.76 5.964 12.24 ;
      RECT 5.648 11.28 5.964 11.76 ;
      RECT 6.458 11.76 6.692 12.72 ;
      RECT 6.458 10.32 7.042 11.76 ;
      RECT 6.636 9.36 7.042 10.32 ;
      RECT 6.976 8.4 7.042 9.36 ;
      RECT 4.192 12.24 4.342 12.72 ;
      RECT 3.758 10.8 3.992 11.76 ;
      RECT 3.758 10.32 4.342 10.8 ;
      RECT 3.758 9.36 3.824 10.32 ;
      RECT 4.192 9.36 4.342 10.32 ;
      RECT 4.192 8.88 4.252 9.36 ;
      RECT 3.936 8.4 4.252 8.88 ;
      RECT 6.076 10.32 6.142 10.8 ;
      RECT 5.558 9.36 5.964 9.84 ;
      RECT 5.648 8.88 5.964 9.36 ;
      RECT 5.648 8.4 6.142 8.88 ;
      RECT 5.648 7.92 5.792 8.4 ;
      RECT 5.558 7.44 5.792 7.92 ;
      RECT 6.458 7.92 6.524 8.88 ;
      RECT 6.458 6.96 6.864 7.92 ;
      RECT 6.458 6.48 7.042 6.96 ;
      RECT 6.548 5.04 7.042 6.48 ;
      RECT 6.458 0 7.042 5.04 ;
      RECT 3.758 6.96 3.824 7.92 ;
      RECT 3.758 6.48 4.342 6.96 ;
      RECT 4.192 5.04 4.342 6.48 ;
      RECT 3.758 4.56 4.342 5.04 ;
      RECT 5.992 6.48 6.142 6.96 ;
      RECT 5.558 5.04 5.792 6 ;
      RECT 5.558 2.16 6.142 5.04 ;
      RECT 5.908 0.72 6.142 2.16 ;
      RECT 5.558 0 6.142 0.72 ;
      RECT 4.658 2.16 5.242 3.12 ;
      RECT 3.758 2.16 4.342 3.12 ;
      RECT 2.858 2.16 3.442 3.12 ;
      RECT 1.958 2.16 2.542 3.12 ;
      RECT 1.058 2.16 1.642 3.12 ;
      RECT 4.658 0 5.242 0.72 ;
      RECT 3.758 0 4.342 0.72 ;
      RECT 2.858 0 3.442 0.72 ;
      RECT 1.958 0 2.542 0.72 ;
      RECT 1.058 0 1.642 0.72 ;
    LAYER m0 ;
      RECT 0 0.002 18 20.158 ;
    LAYER m1 ;
      RECT 0 0 18 20.16 ;
    LAYER m2 ;
      RECT 0 0.015 18 20.145 ;
    LAYER m3 ;
      RECT 0.015 0 17.985 20.16 ;
    LAYER m4 ;
      RECT 0 0.02 18 20.14 ;
    LAYER m5 ;
      RECT 0.012 0 17.988 20.16 ;
    LAYER m6 ;
      RECT 0 0.012 18 20.148 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf028b032e2r2w0cbbehraa4acw

END LIBRARY
