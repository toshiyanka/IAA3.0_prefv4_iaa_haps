module ctech_lib_or2 (
   input logic a,
   input logic b,
   output logic o
);
   d04orn02ln0b0 ctech_lib_dcszo (.a(a), .b(b), .o(o));
endmodule
