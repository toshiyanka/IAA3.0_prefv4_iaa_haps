//               TAP              SlvIDcode   IR_Width  Node  Sec_connections  Hybrid_en  Dfx_Security  Hierarchy_Level  PositionOfTap
Create_TAP_LUT (IPLEVEL_STAP,  32'h1234_5679,   'h8,     'd0,       'd0,         'd0,       GREEN,           1,               0);
