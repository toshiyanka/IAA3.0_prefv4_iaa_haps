module dfxsecure_plugin_waiver_ctrl;
endmodule
