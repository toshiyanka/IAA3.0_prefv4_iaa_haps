`include "ep_base_chk_sig.svh"

   
`include "ep_reg_chk_sig.svh"

   
`include "ep_assumptions.svh"
