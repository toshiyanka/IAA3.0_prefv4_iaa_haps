VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

PROPERTYDEFINITIONS
  MACRO hpml_layer STRING ;
  MACRO heml_layer STRING ;
END PROPERTYDEFINITIONS

MACRO arf062b064e1r1w0cbbehsaa4acw
  CLASS BLOCK ;
  FOREIGN arf062b064e1r1w0cbbehsaa4acw ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 28.8 ;
  PIN ckrdp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 14.76 4.072 15.96 ;
    END
  END ckrdp0
  PIN ckwrp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 12.84 1.116 14.04 ;
    END
  END ckwrp0
  PIN rdaddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.984 14.76 1.028 15.96 ;
    END
  END rdaddrp0[0]
  PIN rdaddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.072 14.76 1.116 15.96 ;
    END
  END rdaddrp0[1]
  PIN rdaddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 14.76 1.372 15.96 ;
    END
  END rdaddrp0[2]
  PIN rdaddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 14.76 1.628 15.96 ;
    END
  END rdaddrp0[3]
  PIN rdaddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 14.76 1.716 15.96 ;
    END
  END rdaddrp0[4]
  PIN rdaddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 14.76 2.016 15.96 ;
    END
  END rdaddrp0[5]
  PIN rdaddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 14.76 4.328 15.96 ;
    END
  END rdaddrp0_fd
  PIN rdaddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.428 14.76 0.472 15.96 ;
    END
  END rdaddrp0_rd
  PIN rdenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.684 14.76 0.728 15.96 ;
    END
  END rdenp0
  PIN sdl_initp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 0.772 14.76 0.816 15.96 ;
    END
  END sdl_initp0
  PIN wraddrp0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 12.84 2.616 14.04 ;
    END
  END wraddrp0[0]
  PIN wraddrp0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 12.84 2.828 14.04 ;
    END
  END wraddrp0[1]
  PIN wraddrp0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 12.84 2.916 14.04 ;
    END
  END wraddrp0[2]
  PIN wraddrp0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 12.84 3.172 14.04 ;
    END
  END wraddrp0[3]
  PIN wraddrp0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 12.84 3.428 14.04 ;
    END
  END wraddrp0[4]
  PIN wraddrp0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 12.84 3.816 14.04 ;
    END
  END wraddrp0[5]
  PIN wraddrp0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.328 12.84 1.372 14.04 ;
    END
  END wraddrp0_fd
  PIN wraddrp0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.584 12.84 1.628 14.04 ;
    END
  END wraddrp0_rd
  PIN wrdatap0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 0.24 1.928 1.44 ;
    END
  END wrdatap0[0]
  PIN wrdatap0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 3.84 1.928 5.04 ;
    END
  END wrdatap0[10]
  PIN wrdatap0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 3.84 2.272 5.04 ;
    END
  END wrdatap0[11]
  PIN wrdatap0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 4.56 2.916 5.76 ;
    END
  END wrdatap0[12]
  PIN wrdatap0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 4.56 2.016 5.76 ;
    END
  END wrdatap0[13]
  PIN wrdatap0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 5.28 2.616 6.48 ;
    END
  END wrdatap0[14]
  PIN wrdatap0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 5.28 2.828 6.48 ;
    END
  END wrdatap0[15]
  PIN wrdatap0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 6 2.272 7.2 ;
    END
  END wrdatap0[16]
  PIN wrdatap0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 6 2.528 7.2 ;
    END
  END wrdatap0[17]
  PIN wrdatap0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 6.72 2.016 7.92 ;
    END
  END wrdatap0[18]
  PIN wrdatap0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 6.72 2.616 7.92 ;
    END
  END wrdatap0[19]
  PIN wrdatap0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 0.24 2.016 1.44 ;
    END
  END wrdatap0[1]
  PIN wrdatap0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 7.44 1.928 8.64 ;
    END
  END wrdatap0[20]
  PIN wrdatap0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 7.44 2.272 8.64 ;
    END
  END wrdatap0[21]
  PIN wrdatap0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 8.16 2.916 9.36 ;
    END
  END wrdatap0[22]
  PIN wrdatap0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 8.16 2.016 9.36 ;
    END
  END wrdatap0[23]
  PIN wrdatap0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 8.88 2.616 10.08 ;
    END
  END wrdatap0[24]
  PIN wrdatap0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 8.88 2.828 10.08 ;
    END
  END wrdatap0[25]
  PIN wrdatap0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 9.6 2.272 10.8 ;
    END
  END wrdatap0[26]
  PIN wrdatap0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 9.6 2.528 10.8 ;
    END
  END wrdatap0[27]
  PIN wrdatap0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 10.32 2.016 11.52 ;
    END
  END wrdatap0[28]
  PIN wrdatap0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 10.32 2.616 11.52 ;
    END
  END wrdatap0[29]
  PIN wrdatap0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 0.96 2.916 2.16 ;
    END
  END wrdatap0[2]
  PIN wrdatap0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 11.04 1.928 12.24 ;
    END
  END wrdatap0[30]
  PIN wrdatap0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 11.04 2.272 12.24 ;
    END
  END wrdatap0[31]
  PIN wrdatap0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 16.56 1.928 17.76 ;
    END
  END wrdatap0[32]
  PIN wrdatap0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 16.56 2.272 17.76 ;
    END
  END wrdatap0[33]
  PIN wrdatap0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 17.28 2.916 18.48 ;
    END
  END wrdatap0[34]
  PIN wrdatap0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 17.28 2.016 18.48 ;
    END
  END wrdatap0[35]
  PIN wrdatap0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 18 2.616 19.2 ;
    END
  END wrdatap0[36]
  PIN wrdatap0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 18 2.828 19.2 ;
    END
  END wrdatap0[37]
  PIN wrdatap0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 18.72 2.272 19.92 ;
    END
  END wrdatap0[38]
  PIN wrdatap0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 18.72 2.528 19.92 ;
    END
  END wrdatap0[39]
  PIN wrdatap0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 0.96 2.272 2.16 ;
    END
  END wrdatap0[3]
  PIN wrdatap0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 19.44 2.016 20.64 ;
    END
  END wrdatap0[40]
  PIN wrdatap0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 19.44 2.616 20.64 ;
    END
  END wrdatap0[41]
  PIN wrdatap0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 20.16 1.928 21.36 ;
    END
  END wrdatap0[42]
  PIN wrdatap0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 20.16 2.272 21.36 ;
    END
  END wrdatap0[43]
  PIN wrdatap0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 20.88 2.916 22.08 ;
    END
  END wrdatap0[44]
  PIN wrdatap0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 20.88 2.016 22.08 ;
    END
  END wrdatap0[45]
  PIN wrdatap0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 21.6 2.616 22.8 ;
    END
  END wrdatap0[46]
  PIN wrdatap0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 21.6 2.828 22.8 ;
    END
  END wrdatap0[47]
  PIN wrdatap0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 22.32 2.272 23.52 ;
    END
  END wrdatap0[48]
  PIN wrdatap0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 22.32 2.528 23.52 ;
    END
  END wrdatap0[49]
  PIN wrdatap0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 1.68 2.616 2.88 ;
    END
  END wrdatap0[4]
  PIN wrdatap0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 23.04 2.016 24.24 ;
    END
  END wrdatap0[50]
  PIN wrdatap0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 23.04 2.616 24.24 ;
    END
  END wrdatap0[51]
  PIN wrdatap0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 23.76 1.928 24.96 ;
    END
  END wrdatap0[52]
  PIN wrdatap0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 23.76 2.272 24.96 ;
    END
  END wrdatap0[53]
  PIN wrdatap0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.872 24.48 2.916 25.68 ;
    END
  END wrdatap0[54]
  PIN wrdatap0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 24.48 2.016 25.68 ;
    END
  END wrdatap0[55]
  PIN wrdatap0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 25.2 2.616 26.4 ;
    END
  END wrdatap0[56]
  PIN wrdatap0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 25.2 2.828 26.4 ;
    END
  END wrdatap0[57]
  PIN wrdatap0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 25.92 2.272 27.12 ;
    END
  END wrdatap0[58]
  PIN wrdatap0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 25.92 2.528 27.12 ;
    END
  END wrdatap0[59]
  PIN wrdatap0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.784 1.68 2.828 2.88 ;
    END
  END wrdatap0[5]
  PIN wrdatap0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 26.64 2.016 27.84 ;
    END
  END wrdatap0[60]
  PIN wrdatap0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 26.64 2.616 27.84 ;
    END
  END wrdatap0[61]
  PIN wrdatap0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.884 27.36 1.928 28.56 ;
    END
  END wrdatap0[62]
  PIN wrdatap0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 27.36 2.272 28.56 ;
    END
  END wrdatap0[63]
  PIN wrdatap0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.228 2.4 2.272 3.6 ;
    END
  END wrdatap0[6]
  PIN wrdatap0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 2.4 2.528 3.6 ;
    END
  END wrdatap0[7]
  PIN wrdatap0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 3.12 2.016 4.32 ;
    END
  END wrdatap0[8]
  PIN wrdatap0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.572 3.12 2.616 4.32 ;
    END
  END wrdatap0[9]
  PIN wrdatap0_fd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.972 12.84 2.016 14.04 ;
    END
  END wrdatap0_fd
  PIN wrdatap0_rd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 2.484 12.84 2.528 14.04 ;
    END
  END wrdatap0_rd
  PIN wrenp0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 1.672 12.84 1.716 14.04 ;
    END
  END wrenp0
  PIN rddatap0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 0.24 3.516 1.44 ;
    END
  END rddatap0[0]
  PIN rddatap0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 3.84 3.516 5.04 ;
    END
  END rddatap0[10]
  PIN rddatap0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 3.84 3.728 5.04 ;
    END
  END rddatap0[11]
  PIN rddatap0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 4.56 3.428 5.76 ;
    END
  END rddatap0[12]
  PIN rddatap0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 4.56 3.816 5.76 ;
    END
  END rddatap0[13]
  PIN rddatap0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 5.28 3.172 6.48 ;
    END
  END rddatap0[14]
  PIN rddatap0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 5.28 3.516 6.48 ;
    END
  END rddatap0[15]
  PIN rddatap0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 6 4.328 7.2 ;
    END
  END rddatap0[16]
  PIN rddatap0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 6 3.428 7.2 ;
    END
  END rddatap0[17]
  PIN rddatap0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 6.72 3.816 7.92 ;
    END
  END rddatap0[18]
  PIN rddatap0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 6.72 4.072 7.92 ;
    END
  END rddatap0[19]
  PIN rddatap0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 0.24 3.728 1.44 ;
    END
  END rddatap0[1]
  PIN rddatap0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 7.44 3.516 8.64 ;
    END
  END rddatap0[20]
  PIN rddatap0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 7.44 3.728 8.64 ;
    END
  END rddatap0[21]
  PIN rddatap0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 8.16 3.428 9.36 ;
    END
  END rddatap0[22]
  PIN rddatap0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 8.16 3.816 9.36 ;
    END
  END rddatap0[23]
  PIN rddatap0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 8.88 3.172 10.08 ;
    END
  END rddatap0[24]
  PIN rddatap0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 8.88 3.516 10.08 ;
    END
  END rddatap0[25]
  PIN rddatap0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 9.6 4.328 10.8 ;
    END
  END rddatap0[26]
  PIN rddatap0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 9.6 3.428 10.8 ;
    END
  END rddatap0[27]
  PIN rddatap0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 10.32 3.816 11.52 ;
    END
  END rddatap0[28]
  PIN rddatap0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 10.32 4.072 11.52 ;
    END
  END rddatap0[29]
  PIN rddatap0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 0.96 3.428 2.16 ;
    END
  END rddatap0[2]
  PIN rddatap0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 11.04 3.516 12.24 ;
    END
  END rddatap0[30]
  PIN rddatap0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 11.04 3.728 12.24 ;
    END
  END rddatap0[31]
  PIN rddatap0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 16.56 3.516 17.76 ;
    END
  END rddatap0[32]
  PIN rddatap0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 16.56 3.728 17.76 ;
    END
  END rddatap0[33]
  PIN rddatap0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 17.28 3.428 18.48 ;
    END
  END rddatap0[34]
  PIN rddatap0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 17.28 3.816 18.48 ;
    END
  END rddatap0[35]
  PIN rddatap0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 18 3.172 19.2 ;
    END
  END rddatap0[36]
  PIN rddatap0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 18 3.516 19.2 ;
    END
  END rddatap0[37]
  PIN rddatap0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 18.72 4.328 19.92 ;
    END
  END rddatap0[38]
  PIN rddatap0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 18.72 3.428 19.92 ;
    END
  END rddatap0[39]
  PIN rddatap0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 0.96 3.816 2.16 ;
    END
  END rddatap0[3]
  PIN rddatap0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 19.44 3.816 20.64 ;
    END
  END rddatap0[40]
  PIN rddatap0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 19.44 4.072 20.64 ;
    END
  END rddatap0[41]
  PIN rddatap0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 20.16 3.516 21.36 ;
    END
  END rddatap0[42]
  PIN rddatap0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 20.16 3.728 21.36 ;
    END
  END rddatap0[43]
  PIN rddatap0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 20.88 3.428 22.08 ;
    END
  END rddatap0[44]
  PIN rddatap0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 20.88 3.816 22.08 ;
    END
  END rddatap0[45]
  PIN rddatap0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 21.6 3.172 22.8 ;
    END
  END rddatap0[46]
  PIN rddatap0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 21.6 3.516 22.8 ;
    END
  END rddatap0[47]
  PIN rddatap0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 22.32 4.328 23.52 ;
    END
  END rddatap0[48]
  PIN rddatap0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 22.32 3.428 23.52 ;
    END
  END rddatap0[49]
  PIN rddatap0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 1.68 3.172 2.88 ;
    END
  END rddatap0[4]
  PIN rddatap0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 23.04 3.816 24.24 ;
    END
  END rddatap0[50]
  PIN rddatap0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 23.04 4.072 24.24 ;
    END
  END rddatap0[51]
  PIN rddatap0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 23.76 3.516 24.96 ;
    END
  END rddatap0[52]
  PIN rddatap0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 23.76 3.728 24.96 ;
    END
  END rddatap0[53]
  PIN rddatap0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 24.48 3.428 25.68 ;
    END
  END rddatap0[54]
  PIN rddatap0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 24.48 3.816 25.68 ;
    END
  END rddatap0[55]
  PIN rddatap0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.128 25.2 3.172 26.4 ;
    END
  END rddatap0[56]
  PIN rddatap0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 25.2 3.516 26.4 ;
    END
  END rddatap0[57]
  PIN rddatap0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 25.92 4.328 27.12 ;
    END
  END rddatap0[58]
  PIN rddatap0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 25.92 3.428 27.12 ;
    END
  END rddatap0[59]
  PIN rddatap0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 1.68 3.516 2.88 ;
    END
  END rddatap0[5]
  PIN rddatap0[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 26.64 3.816 27.84 ;
    END
  END rddatap0[60]
  PIN rddatap0[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 26.64 4.072 27.84 ;
    END
  END rddatap0[61]
  PIN rddatap0[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.472 27.36 3.516 28.56 ;
    END
  END rddatap0[62]
  PIN rddatap0[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.684 27.36 3.728 28.56 ;
    END
  END rddatap0[63]
  PIN rddatap0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.284 2.4 4.328 3.6 ;
    END
  END rddatap0[6]
  PIN rddatap0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.384 2.4 3.428 3.6 ;
    END
  END rddatap0[7]
  PIN rddatap0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 3.772 3.12 3.816 4.32 ;
    END
  END rddatap0[8]
  PIN rddatap0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.028 3.12 4.072 4.32 ;
    END
  END rddatap0[9]
  PIN vcc
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 0.862 0.06 0.938 28.74 ;
        RECT 2.662 0.06 2.738 28.74 ;
        RECT 4.462 0.06 4.538 28.74 ;
        RECT 6.262 0.06 6.338 28.74 ;
        RECT 8.062 0.06 8.138 28.74 ;
        RECT 9.862 0.06 9.938 28.74 ;
        RECT 11.662 0.06 11.738 28.74 ;
        RECT 13.462 0.06 13.538 28.74 ;
    END
  END vcc
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.762 0.06 1.838 28.74 ;
        RECT 3.562 0.06 3.638 28.74 ;
        RECT 5.362 0.06 5.438 28.74 ;
        RECT 7.162 0.06 7.238 28.74 ;
        RECT 8.962 0.06 9.038 28.74 ;
        RECT 10.762 0.06 10.838 28.74 ;
        RECT 12.562 0.06 12.638 28.74 ;
    END
  END vss
  OBS
    LAYER m0 SPACING 0 ;
      RECT -0.016 -0.014 14.416 28.814 ;
    LAYER m1 SPACING 0 ;
      RECT -0.02 -0.02 14.42 28.82 ;
    LAYER m2 SPACING 0 ;
      RECT -0.0705 -0.038 14.4705 28.838 ;
    LAYER m3 SPACING 0 ;
      RECT -0.035 -0.07 14.435 28.87 ;
    LAYER m4 SPACING 0 ;
      RECT -0.07 -0.038 14.47 28.838 ;
    LAYER m5 SPACING 0 ;
      RECT -0.059 -0.09 14.459 28.89 ;
    LAYER m6 SPACING 0 ;
      RECT -0.09 -0.062 14.49 28.862 ;
    LAYER m7 SPACING 0 ;
      RECT 13.538 28.86 14.44 28.92 ;
      RECT 13.538 -0.06 14.492 28.86 ;
      RECT 13.538 -0.12 14.44 -0.06 ;
      RECT 12.638 -0.12 13.462 28.92 ;
      RECT 11.738 -0.12 12.562 28.92 ;
      RECT 10.838 -0.12 11.662 28.92 ;
      RECT 9.938 -0.12 10.762 28.92 ;
      RECT 9.038 -0.12 9.862 28.92 ;
      RECT 8.138 -0.12 8.962 28.92 ;
      RECT 7.238 -0.12 8.062 28.92 ;
      RECT 6.338 -0.12 7.162 28.92 ;
      RECT 5.438 -0.12 6.262 28.92 ;
      RECT 4.538 -0.12 5.362 28.92 ;
      RECT 3.638 28.56 4.462 28.92 ;
      RECT 3.728 27.84 4.462 28.56 ;
      RECT 3.638 27.36 3.684 28.56 ;
      RECT 3.728 27.36 3.772 27.84 ;
      RECT 4.072 27.12 4.462 27.84 ;
      RECT 3.816 26.64 4.028 27.84 ;
      RECT 3.638 26.64 3.772 27.36 ;
      RECT 4.072 26.64 4.284 27.12 ;
      RECT 4.328 25.92 4.462 27.12 ;
      RECT 3.638 25.92 4.284 26.64 ;
      RECT 3.638 25.68 4.462 25.92 ;
      RECT 3.638 24.96 3.772 25.68 ;
      RECT 3.816 24.48 4.462 25.68 ;
      RECT 3.728 24.48 3.772 24.96 ;
      RECT 3.728 24.24 4.462 24.48 ;
      RECT 3.638 23.76 3.684 24.96 ;
      RECT 3.728 23.76 3.772 24.24 ;
      RECT 4.072 23.52 4.462 24.24 ;
      RECT 3.816 23.04 4.028 24.24 ;
      RECT 3.638 23.04 3.772 23.76 ;
      RECT 4.072 23.04 4.284 23.52 ;
      RECT 4.328 22.32 4.462 23.52 ;
      RECT 3.638 22.32 4.284 23.04 ;
      RECT 3.638 22.08 4.462 22.32 ;
      RECT 3.638 21.36 3.772 22.08 ;
      RECT 3.816 20.88 4.462 22.08 ;
      RECT 3.728 20.88 3.772 21.36 ;
      RECT 3.728 20.64 4.462 20.88 ;
      RECT 3.638 20.16 3.684 21.36 ;
      RECT 3.728 20.16 3.772 20.64 ;
      RECT 4.072 19.92 4.462 20.64 ;
      RECT 3.816 19.44 4.028 20.64 ;
      RECT 3.638 19.44 3.772 20.16 ;
      RECT 4.072 19.44 4.284 19.92 ;
      RECT 4.328 18.72 4.462 19.92 ;
      RECT 3.638 18.72 4.284 19.44 ;
      RECT 3.638 18.48 4.462 18.72 ;
      RECT 3.638 17.76 3.772 18.48 ;
      RECT 3.816 17.28 4.462 18.48 ;
      RECT 3.728 17.28 3.772 17.76 ;
      RECT 3.638 16.56 3.684 17.76 ;
      RECT 3.728 16.56 4.462 17.28 ;
      RECT 3.638 15.96 4.462 16.56 ;
      RECT 3.638 14.76 4.028 15.96 ;
      RECT 4.072 14.76 4.284 15.96 ;
      RECT 4.328 14.76 4.462 15.96 ;
      RECT 3.638 14.04 4.462 14.76 ;
      RECT 3.638 12.84 3.772 14.04 ;
      RECT 3.816 12.84 4.462 14.04 ;
      RECT 3.638 12.24 4.462 12.84 ;
      RECT 3.728 11.52 4.462 12.24 ;
      RECT 3.638 11.04 3.684 12.24 ;
      RECT 3.728 11.04 3.772 11.52 ;
      RECT 4.072 10.8 4.462 11.52 ;
      RECT 3.816 10.32 4.028 11.52 ;
      RECT 3.638 10.32 3.772 11.04 ;
      RECT 4.072 10.32 4.284 10.8 ;
      RECT 4.328 9.6 4.462 10.8 ;
      RECT 3.638 9.6 4.284 10.32 ;
      RECT 3.638 9.36 4.462 9.6 ;
      RECT 3.638 8.64 3.772 9.36 ;
      RECT 3.816 8.16 4.462 9.36 ;
      RECT 3.728 8.16 3.772 8.64 ;
      RECT 3.728 7.92 4.462 8.16 ;
      RECT 3.638 7.44 3.684 8.64 ;
      RECT 3.728 7.44 3.772 7.92 ;
      RECT 4.072 7.2 4.462 7.92 ;
      RECT 3.816 6.72 4.028 7.92 ;
      RECT 3.638 6.72 3.772 7.44 ;
      RECT 4.072 6.72 4.284 7.2 ;
      RECT 4.328 6 4.462 7.2 ;
      RECT 3.638 6 4.284 6.72 ;
      RECT 3.638 5.76 4.462 6 ;
      RECT 3.638 5.04 3.772 5.76 ;
      RECT 3.816 4.56 4.462 5.76 ;
      RECT 3.728 4.56 3.772 5.04 ;
      RECT 3.728 4.32 4.462 4.56 ;
      RECT 3.638 3.84 3.684 5.04 ;
      RECT 3.728 3.84 3.772 4.32 ;
      RECT 4.072 3.6 4.462 4.32 ;
      RECT 3.816 3.12 4.028 4.32 ;
      RECT 3.638 3.12 3.772 3.84 ;
      RECT 4.072 3.12 4.284 3.6 ;
      RECT 4.328 2.4 4.462 3.6 ;
      RECT 3.638 2.4 4.284 3.12 ;
      RECT 3.638 2.16 4.462 2.4 ;
      RECT 3.638 1.44 3.772 2.16 ;
      RECT 3.816 0.96 4.462 2.16 ;
      RECT 3.728 0.96 3.772 1.44 ;
      RECT 3.638 0.24 3.684 1.44 ;
      RECT 3.728 0.24 4.462 0.96 ;
      RECT 3.638 -0.12 4.462 0.24 ;
      RECT 2.738 28.56 3.562 28.92 ;
      RECT 2.738 27.36 3.472 28.56 ;
      RECT 3.516 27.36 3.562 28.56 ;
      RECT 2.738 27.12 3.562 27.36 ;
      RECT 2.738 26.4 3.384 27.12 ;
      RECT 3.428 26.4 3.562 27.12 ;
      RECT 3.172 25.92 3.384 26.4 ;
      RECT 3.428 25.92 3.472 26.4 ;
      RECT 2.828 25.68 3.128 26.4 ;
      RECT 3.172 25.68 3.472 25.92 ;
      RECT 2.738 25.2 2.784 26.4 ;
      RECT 3.516 25.2 3.562 26.4 ;
      RECT 2.828 25.2 2.872 25.68 ;
      RECT 2.916 25.2 3.128 25.68 ;
      RECT 3.172 25.2 3.384 25.68 ;
      RECT 3.428 25.2 3.472 25.68 ;
      RECT 3.428 24.96 3.562 25.2 ;
      RECT 2.738 24.48 2.872 25.2 ;
      RECT 2.916 24.48 3.384 25.2 ;
      RECT 3.428 24.48 3.472 24.96 ;
      RECT 3.516 23.76 3.562 24.96 ;
      RECT 2.738 23.76 3.472 24.48 ;
      RECT 2.738 23.52 3.562 23.76 ;
      RECT 2.738 22.8 3.384 23.52 ;
      RECT 3.428 22.8 3.562 23.52 ;
      RECT 3.172 22.32 3.384 22.8 ;
      RECT 3.428 22.32 3.472 22.8 ;
      RECT 2.828 22.08 3.128 22.8 ;
      RECT 3.172 22.08 3.472 22.32 ;
      RECT 2.738 21.6 2.784 22.8 ;
      RECT 3.516 21.6 3.562 22.8 ;
      RECT 2.828 21.6 2.872 22.08 ;
      RECT 2.916 21.6 3.128 22.08 ;
      RECT 3.172 21.6 3.384 22.08 ;
      RECT 3.428 21.6 3.472 22.08 ;
      RECT 3.428 21.36 3.562 21.6 ;
      RECT 2.738 20.88 2.872 21.6 ;
      RECT 2.916 20.88 3.384 21.6 ;
      RECT 3.428 20.88 3.472 21.36 ;
      RECT 3.516 20.16 3.562 21.36 ;
      RECT 2.738 20.16 3.472 20.88 ;
      RECT 2.738 19.92 3.562 20.16 ;
      RECT 2.738 19.2 3.384 19.92 ;
      RECT 3.428 19.2 3.562 19.92 ;
      RECT 3.172 18.72 3.384 19.2 ;
      RECT 3.428 18.72 3.472 19.2 ;
      RECT 2.828 18.48 3.128 19.2 ;
      RECT 3.172 18.48 3.472 18.72 ;
      RECT 2.738 18 2.784 19.2 ;
      RECT 3.516 18 3.562 19.2 ;
      RECT 2.828 18 2.872 18.48 ;
      RECT 2.916 18 3.128 18.48 ;
      RECT 3.172 18 3.384 18.48 ;
      RECT 3.428 18 3.472 18.48 ;
      RECT 3.428 17.76 3.562 18 ;
      RECT 2.738 17.28 2.872 18 ;
      RECT 2.916 17.28 3.384 18 ;
      RECT 3.428 17.28 3.472 17.76 ;
      RECT 3.516 16.56 3.562 17.76 ;
      RECT 2.738 16.56 3.472 17.28 ;
      RECT 2.738 14.04 3.562 16.56 ;
      RECT 2.738 12.84 2.784 14.04 ;
      RECT 2.828 12.84 2.872 14.04 ;
      RECT 2.916 12.84 3.128 14.04 ;
      RECT 3.172 12.84 3.384 14.04 ;
      RECT 3.428 12.84 3.562 14.04 ;
      RECT 2.738 12.24 3.562 12.84 ;
      RECT 2.738 11.04 3.472 12.24 ;
      RECT 3.516 11.04 3.562 12.24 ;
      RECT 2.738 10.8 3.562 11.04 ;
      RECT 2.738 10.08 3.384 10.8 ;
      RECT 3.428 10.08 3.562 10.8 ;
      RECT 3.172 9.6 3.384 10.08 ;
      RECT 3.428 9.6 3.472 10.08 ;
      RECT 2.828 9.36 3.128 10.08 ;
      RECT 3.172 9.36 3.472 9.6 ;
      RECT 2.738 8.88 2.784 10.08 ;
      RECT 3.516 8.88 3.562 10.08 ;
      RECT 2.828 8.88 2.872 9.36 ;
      RECT 2.916 8.88 3.128 9.36 ;
      RECT 3.172 8.88 3.384 9.36 ;
      RECT 3.428 8.88 3.472 9.36 ;
      RECT 3.428 8.64 3.562 8.88 ;
      RECT 2.738 8.16 2.872 8.88 ;
      RECT 2.916 8.16 3.384 8.88 ;
      RECT 3.428 8.16 3.472 8.64 ;
      RECT 3.516 7.44 3.562 8.64 ;
      RECT 2.738 7.44 3.472 8.16 ;
      RECT 2.738 7.2 3.562 7.44 ;
      RECT 2.738 6.48 3.384 7.2 ;
      RECT 3.428 6.48 3.562 7.2 ;
      RECT 3.172 6 3.384 6.48 ;
      RECT 3.428 6 3.472 6.48 ;
      RECT 2.828 5.76 3.128 6.48 ;
      RECT 3.172 5.76 3.472 6 ;
      RECT 2.738 5.28 2.784 6.48 ;
      RECT 3.516 5.28 3.562 6.48 ;
      RECT 2.828 5.28 2.872 5.76 ;
      RECT 2.916 5.28 3.128 5.76 ;
      RECT 3.172 5.28 3.384 5.76 ;
      RECT 3.428 5.28 3.472 5.76 ;
      RECT 3.428 5.04 3.562 5.28 ;
      RECT 2.738 4.56 2.872 5.28 ;
      RECT 2.916 4.56 3.384 5.28 ;
      RECT 3.428 4.56 3.472 5.04 ;
      RECT 3.516 3.84 3.562 5.04 ;
      RECT 2.738 3.84 3.472 4.56 ;
      RECT 2.738 3.6 3.562 3.84 ;
      RECT 2.738 2.88 3.384 3.6 ;
      RECT 3.428 2.88 3.562 3.6 ;
      RECT 3.172 2.4 3.384 2.88 ;
      RECT 3.428 2.4 3.472 2.88 ;
      RECT 2.828 2.16 3.128 2.88 ;
      RECT 3.172 2.16 3.472 2.4 ;
      RECT 2.738 1.68 2.784 2.88 ;
      RECT 3.516 1.68 3.562 2.88 ;
      RECT 2.828 1.68 2.872 2.16 ;
      RECT 2.916 1.68 3.128 2.16 ;
      RECT 3.172 1.68 3.384 2.16 ;
      RECT 3.428 1.68 3.472 2.16 ;
      RECT 3.428 1.44 3.562 1.68 ;
      RECT 2.738 0.96 2.872 1.68 ;
      RECT 2.916 0.96 3.384 1.68 ;
      RECT 3.428 0.96 3.472 1.44 ;
      RECT 3.516 0.24 3.562 1.44 ;
      RECT 2.738 0.24 3.472 0.96 ;
      RECT 2.738 -0.12 3.562 0.24 ;
      RECT 1.838 28.56 2.662 28.92 ;
      RECT 1.928 27.84 2.228 28.56 ;
      RECT 2.272 27.84 2.662 28.56 ;
      RECT 1.838 27.36 1.884 28.56 ;
      RECT 1.928 27.36 1.972 27.84 ;
      RECT 2.016 27.36 2.228 27.84 ;
      RECT 2.272 27.36 2.572 27.84 ;
      RECT 2.016 27.12 2.572 27.36 ;
      RECT 2.616 26.64 2.662 27.84 ;
      RECT 1.838 26.64 1.972 27.36 ;
      RECT 2.016 26.64 2.228 27.12 ;
      RECT 2.528 26.64 2.572 27.12 ;
      RECT 2.528 26.4 2.662 26.64 ;
      RECT 2.272 25.92 2.484 27.12 ;
      RECT 1.838 25.92 2.228 26.64 ;
      RECT 2.528 25.92 2.572 26.4 ;
      RECT 1.838 25.68 2.572 25.92 ;
      RECT 2.616 25.2 2.662 26.4 ;
      RECT 2.016 25.2 2.572 25.68 ;
      RECT 1.838 24.96 1.972 25.68 ;
      RECT 2.016 24.96 2.662 25.2 ;
      RECT 1.928 24.48 1.972 24.96 ;
      RECT 2.016 24.48 2.228 24.96 ;
      RECT 2.272 24.24 2.662 24.96 ;
      RECT 1.928 24.24 2.228 24.48 ;
      RECT 1.838 23.76 1.884 24.96 ;
      RECT 1.928 23.76 1.972 24.24 ;
      RECT 2.016 23.76 2.228 24.24 ;
      RECT 2.272 23.76 2.572 24.24 ;
      RECT 2.016 23.52 2.572 23.76 ;
      RECT 2.616 23.04 2.662 24.24 ;
      RECT 1.838 23.04 1.972 23.76 ;
      RECT 2.016 23.04 2.228 23.52 ;
      RECT 2.528 23.04 2.572 23.52 ;
      RECT 2.528 22.8 2.662 23.04 ;
      RECT 2.272 22.32 2.484 23.52 ;
      RECT 1.838 22.32 2.228 23.04 ;
      RECT 2.528 22.32 2.572 22.8 ;
      RECT 1.838 22.08 2.572 22.32 ;
      RECT 2.616 21.6 2.662 22.8 ;
      RECT 2.016 21.6 2.572 22.08 ;
      RECT 1.838 21.36 1.972 22.08 ;
      RECT 2.016 21.36 2.662 21.6 ;
      RECT 1.928 20.88 1.972 21.36 ;
      RECT 2.016 20.88 2.228 21.36 ;
      RECT 2.272 20.64 2.662 21.36 ;
      RECT 1.928 20.64 2.228 20.88 ;
      RECT 1.838 20.16 1.884 21.36 ;
      RECT 1.928 20.16 1.972 20.64 ;
      RECT 2.016 20.16 2.228 20.64 ;
      RECT 2.272 20.16 2.572 20.64 ;
      RECT 2.016 19.92 2.572 20.16 ;
      RECT 2.616 19.44 2.662 20.64 ;
      RECT 1.838 19.44 1.972 20.16 ;
      RECT 2.016 19.44 2.228 19.92 ;
      RECT 2.528 19.44 2.572 19.92 ;
      RECT 2.528 19.2 2.662 19.44 ;
      RECT 2.272 18.72 2.484 19.92 ;
      RECT 1.838 18.72 2.228 19.44 ;
      RECT 2.528 18.72 2.572 19.2 ;
      RECT 1.838 18.48 2.572 18.72 ;
      RECT 2.616 18 2.662 19.2 ;
      RECT 2.016 18 2.572 18.48 ;
      RECT 1.838 17.76 1.972 18.48 ;
      RECT 2.016 17.76 2.662 18 ;
      RECT 1.928 17.28 1.972 17.76 ;
      RECT 2.016 17.28 2.228 17.76 ;
      RECT 1.838 16.56 1.884 17.76 ;
      RECT 2.272 16.56 2.662 17.76 ;
      RECT 1.928 16.56 2.228 17.28 ;
      RECT 1.838 15.96 2.662 16.56 ;
      RECT 1.838 14.76 1.972 15.96 ;
      RECT 2.016 14.76 2.662 15.96 ;
      RECT 1.838 14.04 2.662 14.76 ;
      RECT 1.838 12.84 1.972 14.04 ;
      RECT 2.016 12.84 2.484 14.04 ;
      RECT 2.528 12.84 2.572 14.04 ;
      RECT 2.616 12.84 2.662 14.04 ;
      RECT 1.838 12.24 2.662 12.84 ;
      RECT 1.928 11.52 2.228 12.24 ;
      RECT 2.272 11.52 2.662 12.24 ;
      RECT 1.838 11.04 1.884 12.24 ;
      RECT 1.928 11.04 1.972 11.52 ;
      RECT 2.016 11.04 2.228 11.52 ;
      RECT 2.272 11.04 2.572 11.52 ;
      RECT 2.016 10.8 2.572 11.04 ;
      RECT 2.616 10.32 2.662 11.52 ;
      RECT 1.838 10.32 1.972 11.04 ;
      RECT 2.016 10.32 2.228 10.8 ;
      RECT 2.528 10.32 2.572 10.8 ;
      RECT 2.528 10.08 2.662 10.32 ;
      RECT 2.272 9.6 2.484 10.8 ;
      RECT 1.838 9.6 2.228 10.32 ;
      RECT 2.528 9.6 2.572 10.08 ;
      RECT 1.838 9.36 2.572 9.6 ;
      RECT 2.616 8.88 2.662 10.08 ;
      RECT 2.016 8.88 2.572 9.36 ;
      RECT 1.838 8.64 1.972 9.36 ;
      RECT 2.016 8.64 2.662 8.88 ;
      RECT 1.928 8.16 1.972 8.64 ;
      RECT 2.016 8.16 2.228 8.64 ;
      RECT 2.272 7.92 2.662 8.64 ;
      RECT 1.928 7.92 2.228 8.16 ;
      RECT 1.838 7.44 1.884 8.64 ;
      RECT 1.928 7.44 1.972 7.92 ;
      RECT 2.016 7.44 2.228 7.92 ;
      RECT 2.272 7.44 2.572 7.92 ;
      RECT 2.016 7.2 2.572 7.44 ;
      RECT 2.616 6.72 2.662 7.92 ;
      RECT 1.838 6.72 1.972 7.44 ;
      RECT 2.016 6.72 2.228 7.2 ;
      RECT 2.528 6.72 2.572 7.2 ;
      RECT 2.528 6.48 2.662 6.72 ;
      RECT 2.272 6 2.484 7.2 ;
      RECT 1.838 6 2.228 6.72 ;
      RECT 2.528 6 2.572 6.48 ;
      RECT 1.838 5.76 2.572 6 ;
      RECT 2.616 5.28 2.662 6.48 ;
      RECT 2.016 5.28 2.572 5.76 ;
      RECT 1.838 5.04 1.972 5.76 ;
      RECT 2.016 5.04 2.662 5.28 ;
      RECT 1.928 4.56 1.972 5.04 ;
      RECT 2.016 4.56 2.228 5.04 ;
      RECT 2.272 4.32 2.662 5.04 ;
      RECT 1.928 4.32 2.228 4.56 ;
      RECT 1.838 3.84 1.884 5.04 ;
      RECT 1.928 3.84 1.972 4.32 ;
      RECT 2.016 3.84 2.228 4.32 ;
      RECT 2.272 3.84 2.572 4.32 ;
      RECT 2.016 3.6 2.572 3.84 ;
      RECT 2.616 3.12 2.662 4.32 ;
      RECT 1.838 3.12 1.972 3.84 ;
      RECT 2.016 3.12 2.228 3.6 ;
      RECT 2.528 3.12 2.572 3.6 ;
      RECT 2.528 2.88 2.662 3.12 ;
      RECT 2.272 2.4 2.484 3.6 ;
      RECT 1.838 2.4 2.228 3.12 ;
      RECT 2.528 2.4 2.572 2.88 ;
      RECT 1.838 2.16 2.572 2.4 ;
      RECT 2.616 1.68 2.662 2.88 ;
      RECT 2.272 1.68 2.572 2.16 ;
      RECT 1.838 1.44 2.228 2.16 ;
      RECT 2.272 0.96 2.662 1.68 ;
      RECT 2.016 0.96 2.228 1.44 ;
      RECT 1.838 0.24 1.884 1.44 ;
      RECT 1.928 0.24 1.972 1.44 ;
      RECT 2.016 0.24 2.662 0.96 ;
      RECT 1.838 -0.12 2.662 0.24 ;
      RECT 0.938 15.96 1.762 28.92 ;
      RECT 0.938 14.76 0.984 15.96 ;
      RECT 1.028 14.76 1.072 15.96 ;
      RECT 1.116 14.76 1.328 15.96 ;
      RECT 1.372 14.76 1.584 15.96 ;
      RECT 1.628 14.76 1.672 15.96 ;
      RECT 1.716 14.76 1.762 15.96 ;
      RECT 0.938 14.04 1.762 14.76 ;
      RECT 0.938 12.84 1.072 14.04 ;
      RECT 1.116 12.84 1.328 14.04 ;
      RECT 1.372 12.84 1.584 14.04 ;
      RECT 1.628 12.84 1.672 14.04 ;
      RECT 1.716 12.84 1.762 14.04 ;
      RECT 0.938 -0.12 1.762 12.84 ;
      RECT -0.04 28.86 0.862 28.92 ;
      RECT -0.092 15.96 0.862 28.86 ;
      RECT -0.092 14.76 0.428 15.96 ;
      RECT 0.472 14.76 0.684 15.96 ;
      RECT 0.728 14.76 0.772 15.96 ;
      RECT 0.816 14.76 0.862 15.96 ;
      RECT -0.092 -0.06 0.862 14.76 ;
      RECT -0.04 -0.12 0.862 -0.06 ;
    LAYER m7 ;
      RECT 13.658 0 14.32 28.8 ;
      RECT 12.758 0 13.342 28.8 ;
      RECT 11.858 0 12.442 28.8 ;
      RECT 10.958 0 11.542 28.8 ;
      RECT 10.058 0 10.642 28.8 ;
      RECT 9.158 0 9.742 28.8 ;
      RECT 8.258 0 8.842 28.8 ;
      RECT 7.358 0 7.942 28.8 ;
      RECT 6.458 0 7.042 28.8 ;
      RECT 5.558 0 6.142 28.8 ;
      RECT 4.658 0 5.242 28.8 ;
      RECT 3.758 28.68 4.342 28.8 ;
      RECT 3.848 27.96 4.342 28.68 ;
      RECT 4.192 27.24 4.342 27.96 ;
      RECT 2.858 28.68 3.442 28.8 ;
      RECT 2.858 27.24 3.352 28.68 ;
      RECT 2.858 26.52 3.264 27.24 ;
      RECT 2.948 25.8 3.008 26.52 ;
      RECT 1.958 28.68 2.542 28.8 ;
      RECT 2.048 27.96 2.108 28.68 ;
      RECT 2.392 27.96 2.542 28.68 ;
      RECT 2.392 27.24 2.452 27.96 ;
      RECT 1.058 16.08 1.642 28.8 ;
      RECT 0.08 16.08 0.742 28.8 ;
      RECT 0.08 14.64 0.308 16.08 ;
      RECT 0.08 0 0.742 14.64 ;
      RECT 3.758 25.8 4.164 26.52 ;
      RECT 3.936 24.36 4.342 25.8 ;
      RECT 4.192 23.64 4.342 24.36 ;
      RECT 1.958 25.8 2.108 26.52 ;
      RECT 2.136 25.08 2.452 25.8 ;
      RECT 2.392 24.36 2.542 25.08 ;
      RECT 2.392 23.64 2.452 24.36 ;
      RECT 3.036 24.36 3.264 25.08 ;
      RECT 2.858 23.64 3.352 24.36 ;
      RECT 2.858 22.92 3.264 23.64 ;
      RECT 2.948 22.2 3.008 22.92 ;
      RECT 3.758 22.2 4.164 22.92 ;
      RECT 3.936 20.76 4.342 22.2 ;
      RECT 4.192 20.04 4.342 20.76 ;
      RECT 1.958 22.2 2.108 22.92 ;
      RECT 2.136 21.48 2.452 22.2 ;
      RECT 2.392 20.76 2.542 21.48 ;
      RECT 2.392 20.04 2.452 20.76 ;
      RECT 3.036 20.76 3.264 21.48 ;
      RECT 2.858 20.04 3.352 20.76 ;
      RECT 2.858 19.32 3.264 20.04 ;
      RECT 2.948 18.6 3.008 19.32 ;
      RECT 3.758 18.6 4.164 19.32 ;
      RECT 3.936 17.16 4.342 18.6 ;
      RECT 3.848 16.44 4.342 17.16 ;
      RECT 3.758 16.08 4.342 16.44 ;
      RECT 3.758 14.64 3.908 16.08 ;
      RECT 3.758 14.16 4.342 14.64 ;
      RECT 3.936 12.72 4.342 14.16 ;
      RECT 3.758 12.36 4.342 12.72 ;
      RECT 3.848 11.64 4.342 12.36 ;
      RECT 4.192 10.92 4.342 11.64 ;
      RECT 1.958 18.6 2.108 19.32 ;
      RECT 2.136 17.88 2.452 18.6 ;
      RECT 2.392 16.44 2.542 17.88 ;
      RECT 2.048 16.44 2.108 17.16 ;
      RECT 1.958 16.08 2.542 16.44 ;
      RECT 2.136 14.64 2.542 16.08 ;
      RECT 1.958 14.16 2.542 14.64 ;
      RECT 2.136 12.72 2.364 14.16 ;
      RECT 1.958 12.36 2.542 12.72 ;
      RECT 2.048 11.64 2.108 12.36 ;
      RECT 2.392 11.64 2.542 12.36 ;
      RECT 2.392 10.92 2.452 11.64 ;
      RECT 3.036 17.16 3.264 17.88 ;
      RECT 2.858 16.44 3.352 17.16 ;
      RECT 2.858 14.16 3.442 16.44 ;
      RECT 1.058 14.16 1.642 14.64 ;
      RECT 2.858 12.36 3.442 12.72 ;
      RECT 2.858 10.92 3.352 12.36 ;
      RECT 2.858 10.2 3.264 10.92 ;
      RECT 2.948 9.48 3.008 10.2 ;
      RECT 1.058 0 1.642 12.72 ;
      RECT 3.758 9.48 4.164 10.2 ;
      RECT 3.936 8.04 4.342 9.48 ;
      RECT 4.192 7.32 4.342 8.04 ;
      RECT 1.958 9.48 2.108 10.2 ;
      RECT 2.136 8.76 2.452 9.48 ;
      RECT 2.392 8.04 2.542 8.76 ;
      RECT 2.392 7.32 2.452 8.04 ;
      RECT 3.036 8.04 3.264 8.76 ;
      RECT 2.858 7.32 3.352 8.04 ;
      RECT 2.858 6.6 3.264 7.32 ;
      RECT 2.948 5.88 3.008 6.6 ;
      RECT 3.758 5.88 4.164 6.6 ;
      RECT 3.936 4.44 4.342 5.88 ;
      RECT 4.192 3.72 4.342 4.44 ;
      RECT 1.958 5.88 2.108 6.6 ;
      RECT 2.136 5.16 2.452 5.88 ;
      RECT 2.392 4.44 2.542 5.16 ;
      RECT 2.392 3.72 2.452 4.44 ;
      RECT 3.036 4.44 3.264 5.16 ;
      RECT 2.858 3.72 3.352 4.44 ;
      RECT 2.858 3 3.264 3.72 ;
      RECT 2.948 2.28 3.008 3 ;
      RECT 3.758 2.28 4.164 3 ;
      RECT 3.936 0.84 4.342 2.28 ;
      RECT 3.848 0.12 4.342 0.84 ;
      RECT 3.758 0 4.342 0.12 ;
      RECT 1.958 1.56 2.108 3 ;
      RECT 2.392 1.56 2.452 2.28 ;
      RECT 2.392 0.84 2.542 1.56 ;
      RECT 2.136 0.12 2.542 0.84 ;
      RECT 1.958 0 2.542 0.12 ;
      RECT 3.036 0.84 3.264 1.56 ;
      RECT 2.858 0.12 3.352 0.84 ;
      RECT 2.858 0 3.442 0.12 ;
    LAYER m0 ;
      RECT 0 0.002 14.4 28.798 ;
    LAYER m1 ;
      RECT 0 0 14.4 28.8 ;
    LAYER m2 ;
      RECT 0 0.015 14.4 28.785 ;
    LAYER m3 ;
      RECT 0.015 0 14.385 28.8 ;
    LAYER m4 ;
      RECT 0 0.02 14.4 28.78 ;
    LAYER m5 ;
      RECT 0.012 0 14.388 28.8 ;
    LAYER m6 ;
      RECT 0 0.012 14.4 28.788 ;
  END
  PROPERTY heml_layer "7" ;
  PROPERTY hpml_layer "7" ;
END arf062b064e1r1w0cbbehsaa4acw

END LIBRARY
