//-----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright (2013) (2013) Intel Corporation All Rights Reserved. 
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors. The
// Material is protected by worldwide copyright and trade secret laws and 
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or disclosed
// in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual 
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be 
// express and approved by Intel in writing.
//------------------------------------------------------------------------------
// File   : hcw_transaction.sv
// Author : Mike Betker
//
// Description :
//
// This class is derived form uvm_sequence_item and it represents the transaction 
// object being generated by sequence/sequencer and sent to the DUT through driver
//------------------------------------------------------------------------------
`ifndef HCW_TRANSACTION__SV
`define HCW_TRANSACTION__SV


`ifndef HQMCORE_DEBUG
 `define HCW_QID_WIDTH   8
`else
 `define HCW_QID_WIDTH   6
`endif

class hcw_transaction extends uvm_sequence_item;

 //------------------------- 
 //-- hcw transaction count
 //-------------------------
 static int     trans_count = 0;
 
 //------------------------- 
 //-- hcw info class
 //-------------------------
 hcw_transinfo  hcw_trinfo;

 
 //------------------------- 
 //-- hcw_fields
 //------------------------- 	 
 //-- controls
 rand bit	qe_valid;
 rand bit 	qe_orsp;
 rand bit	qe_uhl;
 rand bit	cq_pop;
 
 //-- atm/uno/ord/dir
 rand hcw_qtype qtype;
 
 
 //-- hcw_fields of ENQ hcw
 rand bit               dsi_error;
 rand bit               cq_int_rearm;
 rand logic [2:0]       msgtype;
 rand logic [3:0] 	cmp_id;
 rand bit               no_inflcnt_dec;
 rand logic [3:0] 	dbg;
 rand logic [1:0] 	wu;
 rand bit               meas; //--this is ts_flag field
 rand logic [15:0]   	lockid;
 rand logic [15:0]   	directinfo;
 rand logic [2:0]    	qpri;
 rand logic [hqm_pkg::DIR_QID_ARCH_WIDTH-1:0]    	qid;
 rand logic [15:0]   	idsi;

 rand logic [63:0]   	iptr; 
 
 //-- hcw_fields of SCH hcw
 rand logic [1:0]	qid_depth;
 rand logic             cq_gen;
 rand logic [hqm_pkg::DIR_PP_ARCH_WIDTH-1:0]	prod_port;  //-- this is ppid of enq   
 rand logic      	prod_isldb; //-- this is is_ldb of enq V2_TB
 
 
 //-- RSVD fields
 rand logic [15:0]       rsvd0;
 
           
                 
		
 //------------------------- 
 //-- hcw supporting fields
 //-------------------------  
 rand logic [7:0]       sai;                    // SAI value to be used when enqueuing/scheduling HCW
 rand bit         	is_error;               // bit from HCW
 rand bit         	is_ldb;                 // control PP for enqueue and field in scheduled HCW
 rand logic [7:0]    	rtn_credit_only;        // controls AXI user bit for hqm_core enqueue
 rand logic          	exp_rtn_credit_only;    // if set the scoreboard should verify that it detects the return credit only action for the HCW
 rand logic [(hqm_pkg::DIR_PP_ARCH_WIDTH-1):0]  ppid;                   // PP/CQ associated with enqueued/scheduled HCW
 rand logic [4:0]    	vasid;                  // VAS associated with enqueued/scheduled HCW
 rand logic [7:0]   	vfid;                   // dm_core testbench?
 rand logic [3:0]	frg_ldbnum;             // ?
 
 rand logic [7:0]   	pp_type_pp;             // {is_ldb, producer_port[6:0]}; lower 128 to represent dirpp{0:95}; upper 128 to represent ldbpp{0:63}
 rand logic [6:0]       pf_qid;

 rand bit               ingress_drop;           // identifies if the hcw will be dropped in hqm_system ingress logic (credit not returned to hqm_core)
 rand bit               exp_ingress_drop;       // identifies if it is expected that this HCW will be dropped in hqm_system ingress logic (credit not returned to hqm_core)
                                                //   - if set the scoreboard should verify that it has detected an HCW that should be dropped as a result of ingress checks
 rand bit               ingress_comp_nodrop;    // when ingress_drop=1 and ingress_comp_nodrop=1: this means ENQ is dropped, but completion is not
 rand bit               hcw_batch;              // Send HCWs in batch, if supported. Flush batched HCWs if 0.
 rand bit               is_vf;                  // identifies if the hcw is associated with a VF or PF
 rand bit               is_nm_pf;               // identifies if the hcw is going to be written through PF access window or PP address window
 rand bit [3:0]         vf_num;                 // VF number if HCW associated with a VF

 rand logic [7:0]       sch_cqid;               // Destination CQ of scheduled HCW
 rand logic [7:0]       sch_cq_occ_cq;          // unused?
 rand bit               sch_cq_occ;             // AXI user bit for scheduled HCW
 rand bit               sch_parity;             // AXI user bit for scheduled HCW
 rand bit               sch_error;              // AXI user bit for scheduled HCW
 rand bit               sch_qid_occ;            // unused?
 rand bit   [1:0]       sch_write_status;       // AXI user bit for scheduled HCW
 rand bit         	sch_is_ldb;             // Scheduled HCW is for a LDB CQ - AXI user bit for scheduled HCW
 rand logic [11:0]    	sch_addr;               // offset in CQ buffer 12-bit to support DIR4096

 bit			is_compled;
 bit			is_tokened;             // unused?
 bit                    is_sched;               //- when 1: it's HQM returned SCHED hcw_transaction (set when ATM HCW scheduled)
 bit			is_done;
 int                    ord_state; //-- 

 bit [1:0]          compare_type;  

 //------------------------- 
 //-- hcw embeded fields are passed to hcw_trinfo
 //-------------------------
 rand logic [63:0]	tbcnt; 

 rand logic [63:0]	tbcntsch;
 rand hcw_qtype         qtypesch;
 rand bit               isdir;  

      bit   [1:0]       enqattr;

 rand bit               is_ord;  //-- hqm_pp_cq_base_seq.sv cq_buffer_monitor() ::  read a SCHED HCW with qType=ORD => pend_comp_return.push(1); 
                                 //-- hqm_pp_cq_hqmproc_seq.sv                  ::  pop pend_comp_return, if it's 1  => is_ordered=1; and set is_ord=1 in generated ENQ HCW

 rand bit               reordenq_done;
 rand bit               reord;   //reord[1]=done(remove bit1); reord[0]=reordmark
 //-- old_version: rand logic [4:0]    	frg_cnt; //--09092016_newversionRTL supports upto 16K fragments, it reports intr when fragments > 16.
 rand logic [15:0]    	frg_cnt;
 rand logic [15:0]    	frg_num;
 rand logic [3:0]    	frg_ldbcnt;
 rand bit               frg_last;
 rand bit               frg_first;
 rand logic [15:0]	reordidx;
 rand bit               sch_frg_last;
 rand bit               sch_frg_first;
 rand logic [5:0]       ordqid;  //-- 
 rand logic [2:0]       ordpri;  //--
 rand logic [15:0]      ordlockid;  //-- 
 rand logic [63:0]      ordidx;  //-- track ordidx in the same ordqid      


 //-------------------------
 //-- performance mon
 //-------------------------
 time                   mea_start_time;
 int                    mea_latency_valid;

 //-------------------------
 //-- user field of Data mover ihcw interface write data channel
 //-------------------------
 rand logic [hqm_pkg::DIR_CQ_ARCH_WIDTH-1:0] 	cq;
 rand bit 					cq_parity;	
 rand logic [(8)-1:0] 		ecc_h;
 rand logic [(8)-1:0] 		ecc_l;

 //-------------------------
 //-- user field of Data mover thcw interface write data channel
 //-------------------------
 rand logic             vpp_vf_pf_parity;            // parity covers { is_pf, vf, vpp }
 rand logic             is_pf;                       // qid,vpp are physical
 rand logic [(4)-1:0]   vf;                          // virtual function
 rand logic [hqm_pkg::DIR_PP_ARCH_WIDTH-1:0]   vpp;  // virtual producer port (for tHCW enq)

 //-------------------------  
 //Constraints
 //-------------------------  
 
 constraint qtype_dir {
               //qtype == QDIR -> {lockid == 16'h0;} 
	       
       }

constraint c_vf {
                  soft is_vf == 1'b0;
                }

constraint c_hcw_batch {
                  soft hcw_batch == 1'b0;
                }

constraint c_ingress_drop {
                  soft ingress_drop == 1'b0;
                  soft exp_ingress_drop == 1'b0;
                  soft ingress_comp_nodrop == 1'b0;
                }

constraint c_exp_rtn_credit_only {
                  soft exp_rtn_credit_only == 1'b0;
                }

constraint c_is_nm_pf {
    soft is_nm_pf == 1'b0;
}
constraint c_frg {
    soft frg_first == 0;
    soft frg_last  == 0;
    soft frg_cnt   == 0;
}

 //-------------------------  
 //static constraint if any
 //-------------------------  
 //static constraint disable_type {xxx == 0;};
  
 

 //------------------------- 
 //-------------------------    
  `uvm_object_utils_begin(hcw_transaction)
     `uvm_field_int(sai,             UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ppid,            UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(vasid,           UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(is_error,        UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(is_ldb,          UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(is_vf,           UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(is_nm_pf,        UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(vf_num,          UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_cq_occ_cq,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_cq_occ,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_parity,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_error,       UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_qid_occ,     UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_write_status,  UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_is_ldb,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_addr,        UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(rtn_credit_only, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(exp_rtn_credit_only, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(hcw_batch,       UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ingress_drop,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(exp_ingress_drop,UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ingress_comp_nodrop,    UVM_ALL_ON | UVM_NOCOMPARE)

     `uvm_field_enum(hcw_qtype, qtype, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_enum(hcw_qtype, qtypesch, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qe_valid,  UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qe_orsp,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qe_uhl,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cq_pop,    UVM_ALL_ON | UVM_NOCOMPARE)
                    
     `uvm_field_int(dsi_error,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cq_int_rearm,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(dbg,       UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cmp_id,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(msgtype,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(directinfo,UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(lockid,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qpri,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qid,       UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(idsi,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(iptr,      UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(qid_depth, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cq_gen,    UVM_ALL_ON | UVM_NOCOMPARE)    
     `uvm_field_int(no_inflcnt_dec, UVM_ALL_ON | UVM_NOCOMPARE)                      
     `uvm_field_int(wu, UVM_ALL_ON | UVM_NOCOMPARE)                      
     `uvm_field_int(meas, UVM_ALL_ON | UVM_NOCOMPARE)                      
     `uvm_field_int(prod_port, UVM_ALL_ON | UVM_NOCOMPARE)                      
     `uvm_field_int(prod_isldb, UVM_ALL_ON | UVM_NOCOMPARE)                      

     `uvm_field_int(tbcnt,     UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(tbcntsch,UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(isdir,     UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(is_ord,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(enqattr,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(reord,     UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(reordenq_done,     UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(frg_cnt,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(frg_num,   UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(frg_ldbcnt,UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(frg_first, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(frg_last,  UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_frg_last,  UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(sch_frg_first, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ordpri,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ordqid,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ordlockid, UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ordidx,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(reordidx,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cq,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(cq_parity,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ecc_h,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(ecc_l,    UVM_ALL_ON | UVM_NOCOMPARE)
     `uvm_field_int(compare_type,    UVM_ALL_ON | UVM_NOCOMPARE)
  `uvm_object_utils_end
  
  
 
 //------------------------- 
 // Function: new 
 // Class constructor
 //------------------------- 
  function new (string name = "hcw_xaction_inst");
    super.new(name);
    
    hcw_trinfo          = new();
    compare_type        = 2'b0;
    is_vf               = 1'b0;
    is_nm_pf            = 1'b0;
    hcw_batch           = 1'b0;
    ingress_drop        = 1'b0;
    exp_ingress_drop    = 1'b0;
    ingress_comp_nodrop = 1'b0;
    exp_rtn_credit_only = 1'b0;

    set_transaction_id(trans_count);
    trans_count++;
  endfunction : new


 //------------------------- 
 // Function: post_randomize
 // SV function overload for randomizing this class
 //------------------------- 
 function void post_randomize();
   super.post_randomize();
 endfunction
   


 //------------------------- 
 //-- Note: by defualt, HQMCORE_DEBUG is not defined 
 //-- turn on HQMCORE_DEBUG if want to debug ORD, it will bring embedded fields to interface signals.
 //------------------------- 
 `ifndef HQMCORE_DEBUG
   `define HCW_ENQ_PACK_STRUCTURE_MACRO( ITEM ) \
               {``ITEM``.rsvd0[1:0],            \
                ``ITEM``.dsi_error,             \
                ``ITEM``.rsvd0[2],              \
                ``ITEM``.qe_valid,              \
                ``ITEM``.qe_orsp,               \
                ``ITEM``.qe_uhl,                \
                ``ITEM``.cq_pop,                \
                ``ITEM``.cmp_id[3:0],           \
                ``ITEM``.no_inflcnt_dec,        \
                ``ITEM``.wu[1:0],              \
                ``ITEM``.meas,                  \
                ``ITEM``.lockid[15:0],          \
                ``ITEM``.msgtype[2:0],          \
                ``ITEM``.qpri[2:0],             \
                ``ITEM``.qtype[1:0],            \
                ``ITEM``.qid[7:0],              \
                ``ITEM``.idsi[15:0],            \
                ``ITEM``.iptr[63:0]              \
                 }       

   
 `else
    //-- HQMCORE_DEBUG mode 
   `define HCW_ENQ_PACK_STRUCTURE_MACRO( ITEM ) \
               {``ITEM``.rsvd0[1:0],            \
                ``ITEM``.dsi_error,             \
                ``ITEM``.rsvd0[2],              \
                ``ITEM``.qe_valid,              \
                ``ITEM``.qe_orsp,               \
                ``ITEM``.qe_uhl,                \
                ``ITEM``.cq_pop,                \
                ``ITEM``.cmp_id[3:0],           \
                ``ITEM``.no_inflcnt_dec,        \
                ``ITEM``.wu[1:0],              \
                ``ITEM``.meas,                  \
                ``ITEM``.lockid[15:0],          \
                ``ITEM``.msgtype[2:0],          \
                ``ITEM``.qpri[2:0],             \
                ``ITEM``.qtype[1:0],            \
                ``ITEM``.rsvd0[4:3],            \
                ``ITEM``.qid[5:0],              \
                ``ITEM``.idsi[15:0],            \
                ``ITEM``.tbcnt[15:0],           \
                ``ITEM``.tbcntsch[15:0],        \
                ``ITEM``.qtypesch[1:0],         \
                ``ITEM``.isdir,                 \
                ``ITEM``.reord,                 \
                ``ITEM``.ingress_drop,          \
                ``ITEM``.frg_cnt[3:0],          \
                ``ITEM``.frg_last,              \
                ``ITEM``.ordqid[5:0],           \
                ``ITEM``.ordidx[15:0]           \
//                ``ITEM``.iptr[7:0]              \
                 }       
  
  
 `endif
 
 //-- 
 `ifndef HQMCORE_DEBUG
   `define HCW_SCH_PACK_STRUCTURE_MACRO( ITEM ) \
               {``ITEM``.rsvd0[1:0],            \
                ``ITEM``.is_error,              \
                ``ITEM``.rsvd0[3:2],            \
                ``ITEM``.qid_depth[1:0],        \
                ``ITEM``.cq_gen,                \
                ``ITEM``.cmp_id[3:0],           \
                ``ITEM``.dbg[0],                \
                ``ITEM``.wu[1:0],               \
                ``ITEM``.meas,                  \
                ``ITEM``.lockid[15:0],          \
                ``ITEM``.msgtype[2:0],          \
                ``ITEM``.qpri[2:0],             \
                ``ITEM``.qtype[1:0],            \
                ``ITEM``.qid[7:0],              \
                ``ITEM``.idsi[15:0],            \
                ``ITEM``.iptr[63:0]              \
                 }  
 `else
 
    //-- HQMCORE_DEBUG mode  
   `define HCW_SCH_PACK_STRUCTURE_MACRO( ITEM ) \
               {``ITEM``.rsvd0[1:0],            \
                ``ITEM``.is_error,              \
                ``ITEM``.rsvd0[3:2],            \
                ``ITEM``.qid_depth[1:0],        \
                ``ITEM``.cq_gen,                \
                ``ITEM``.cmp_id[3:0],           \
                ``ITEM``.dbg[0],                \
                ``ITEM``.wu[1:0],               \
                ``ITEM``.meas,                  \
                ``ITEM``.lockid[15:0],          \
                ``ITEM``.msgtype[2:0],          \
                ``ITEM``.qpri[2:0],             \
                ``ITEM``.qtype[1:0],            \
                ``ITEM``.rsvd0[5:4],            \
                ``ITEM``.qid[5:0],              \
                ``ITEM``.idsi[15:0],            \
                ``ITEM``.tbcnt[15:0],           \
                ``ITEM``.tbcntsch[15:0],        \
                ``ITEM``.qtypesch[1:0],         \
                ``ITEM``.isdir,                 \
                ``ITEM``.reord,                 \
                ``ITEM``.frg_cnt[4:0],          \
                ``ITEM``.frg_last,              \
                ``ITEM``.ordqid[5:0],           \
                ``ITEM``.ordidx[15:0]           \
//                ``ITEM``.iptr[7:0]              \
                 }  
 `endif

   
  //---------------------------------------------------------------------------- 
  //---------------------------------------------------------------------------- 
  //-- byte_size
  //----------------------------------------------------------------------------   
  virtual function int unsigned byte_size ( int kind = -1 ) ;
     return 16 ;
  endfunction : byte_size 

  
  //---------------------------------------------------------------------------- 
  //-- byte_pack (kind=0: ENQ hcw_xaction format; kind=1: SCH hcw_xaction format)
  //----------------------------------------------------------------------------  
  //virtual function int unsigned byte_pack ( ref logic[7:0] bytes[], input int kind = 0 ) ;
   virtual function logic[127:0] byte_pack ( input int kind = 0 ) ;
        logic [ 127:0 ] hcwdata ;
        int j ; 

	case (kind)
		'd0: begin
                       uvm_report_info(get_type_name(),$psprintf("hcw_xaction:byte_pack_pre: kind=%0d/tbcnt=%0d/tbcntsch=%0d, cmd=0x%0x/qtype=%0s/is_ldb=%0d/ppid=%0d/qid=0x%0x/lockid=0x%0x/iptr=0x%0x", kind, tbcnt, tbcntsch, {qe_valid,qe_orsp,qe_uhl,cq_pop}, qtype.name(), is_ldb, ppid, qid, lockid, iptr), UVM_MEDIUM); 
                       hcwdata = `HCW_ENQ_PACK_STRUCTURE_MACRO ( this ) ;
                     end 
		'd1: hcwdata = `HCW_SCH_PACK_STRUCTURE_MACRO ( this ) ; 
		default: hcwdata = `HCW_ENQ_PACK_STRUCTURE_MACRO ( this ) ;
	endcase
        			  
        uvm_report_info(get_type_name(),$psprintf("hcw_xaction:byte_pack kind=%0d/tbcnt=%0d/tbcntsch=%0d, hcwdata=0x%0x, cmd=0x%0x/qtype=%0s/is_ldb=%0d/ppid=%0d/qid=0x%0x/lockid=0x%0x/iptr=0x%0x", kind, tbcnt, tbcntsch, hcwdata, {qe_valid,qe_orsp,qe_uhl,cq_pop}, qtype.name(), is_ldb, ppid, qid, lockid, iptr), UVM_MEDIUM); 
        
        return hcwdata ;

    endfunction : byte_pack
 

  //---------------------------------------------------------------------------- 
  //-- byte_unpack (kind=0: ENQ hcw_xaction format; kind=1: SCH hcw_xaction format)
  //----------------------------------------------------------------------------  
    //virtual function int unsigned byte_unpack (const ref logic[7:0] bytes[],  input int kind = 0 ) ;
    virtual function byte_unpack (int kind = 0, logic[127:0] hcwdata ) ; 
        int j ;  
	
        // -- unpack
		case (kind)
           'd0: `HCW_ENQ_PACK_STRUCTURE_MACRO ( this ) =  hcwdata ; 
           'd1: `HCW_SCH_PACK_STRUCTURE_MACRO ( this ) =  hcwdata ; 			  
		   default: `HCW_ENQ_PACK_STRUCTURE_MACRO ( this ) =  hcwdata;
		endcase
	
        uvm_report_info(get_type_name(),$psprintf("hcw_xaction:byte_unpack kind=%0d/tbcnt=%0d/tbcntsch=%0d, hcwdata=0x%0x, qid=0x%0x/lockid=0x%0x/ordidx=%0d", kind, tbcnt, tbcntsch, hcwdata, qid, lockid, ordidx), UVM_MEDIUM); 


        //return bytes_tmp.size() ;
 
    endfunction : byte_unpack

    virtual function string sprint_hcw_enq();
      sprint_hcw_enq = $psprintf("rsvd0=0x%0x dsi_error=%01x qe_valid=%01x qe_orsp=%01x qe_uhl=%01x cq_pop=%01x cmp_id=0x%01x\n",
                                 rsvd0[4:0],
                                 dsi_error,
                                 qe_valid,
                                 qe_orsp,
                                 qe_uhl,
                                 cq_pop,
                                 cmp_id[3:0]
                                );

      sprint_hcw_enq = {sprint_hcw_enq,$psprintf("no_inflcnt_dec=%01x wu=%01x ts_flag=%0x lockid=0x%04x msgtype=%01x qpri=%01x qtype=%01x qid=0x%02x idsi=0x%04x iptr=0x%08x_%08x",
                                                 no_inflcnt_dec,
                                                 wu[1:0],
                                                 meas,
                                                 lockid[15:0],
                                                 msgtype[2:0],
                                                 qpri[2:0],
                                                 qtype[1:0],
                                                 qid[`HCW_QID_WIDTH-1:0],
                                                 idsi[15:0],
                                                 iptr[63:32],
                                                 iptr[31:0]
                                                )
                       };
    endfunction : sprint_hcw_enq

 
    virtual function string sprint_hcw_sch();
      sprint_hcw_sch = $psprintf("rsvd=%01x is_error=%01x rsvd=%01x qid_depth=%01x cq_gen=%01x cmp_id=%01x dbg=%01x meas=%01x \n",
                                 rsvd0[1:0],
                                 is_error,
                                 rsvd0[3:2],
                                 qid_depth,
                                 cq_gen,
                                 cmp_id[3:0],
                                 dbg[2:0],
                                 meas
                                );

      sprint_hcw_sch = {sprint_hcw_sch,$psprintf("is_ldb=%01x lockid=%0x msgtype=%01x qpri=%01x qtype=%01x qid=%02x idsi=%04x iptr=%08x_%08x",
                                                 is_ldb,
                                                 lockid[15:0],
                                                 msgtype[2:0],
                                                 qpri[2:0],
                                                 qtype[1:0],
                                                 qid,
                                                 idsi[15:0],
                                                 iptr[63:32],
                                                 iptr[31:0]
                                                )
                       };
    endfunction : sprint_hcw_sch

 
 
    virtual function string sprint_hcw_sch_rebuild();
      sprint_hcw_sch_rebuild = $psprintf("prod_isldb=%0d prod_prot=%0d cq=%0d qid=%0d pri=%0d lockid=0x%0x is_ord=%0d reord=%0d frg_cnt=%0d frg_first=%0d frg_last=%0d ordqid=%0d ordidx=%0d \n",
                                 prod_isldb,
                                 prod_port,
                                 ppid,
                                 qid,
                                 qpri,
                                 lockid,
                                 is_ord,
                                 reord,
                                 frg_cnt,
                                 frg_first,
                                 frg_last,
                                 ordqid,
                                 ordidx 
                                );
   endfunction : sprint_hcw_sch_rebuild
  //---------------------------------------------------------------------------- 

  //---------------------------------------------------------------------------- 
  //-- set_hcw_trinfo
  //----------------------------------------------------------------------------   
  virtual function set_hcw_trinfo (bit kind = 0) ;
      //hcw_trinfo = new();
      
      if( kind == 0 ) begin
         iptr                         = '0;
         iptr[63:48]                  = this.tbcnt[15:0]    ; //-- RTL uses 16-bit in seqnum tracing, keep this 16-bit  
      end 
      
      hcw_trinfo.info_msgtype         = this.msgtype;  
      hcw_trinfo.info_isdir   	      = this.isdir	    ;  
      hcw_trinfo.info_tbcnt	      = this.tbcnt	    ;  
      hcw_trinfo.info_qtypesch	      = this.qtypesch       ;  
      hcw_trinfo.info_tbcntsch	      = this.tbcntsch       ;    
      hcw_trinfo.info_lkid	      = this.lockid	    ;  
      hcw_trinfo.info_enqattr         = this.enqattr        ;	
      hcw_trinfo.info_reord	      = this.reord	    ;	
      hcw_trinfo.info_frg_cnt	      = this.frg_cnt        ; 
      hcw_trinfo.info_frg_ldbcnt      = this.frg_ldbcnt     ; 
      hcw_trinfo.info_frg_last	      = this.frg_last       ;  
      hcw_trinfo.info_ordpri	      = this.ordpri         ;  
      hcw_trinfo.info_ordqid	      = this.ordqid         ;  
      hcw_trinfo.info_ordlockid       = this.ordlockid      ;  
      hcw_trinfo.info_ordidx	      = this.ordidx         ;	
      hcw_trinfo.info_ppidx	      = this.ppid           ;	//--V2_TB
      hcw_trinfo.info_isldb	      = this.is_ldb         ;	//--V2_TB
      	 
        uvm_report_info(get_type_name(),$psprintf("hcw_xaction:set_hcw_trinfo info_tbcnt=%0d/info_ordqid=0x%0x/info_ordpri=%0d/info_ordidx=%0d/info_lockid=0x%0x/enqisldb=%0d/enqppid=%0d/iptr=0x%0x", 
                      hcw_trinfo.info_tbcnt, hcw_trinfo.info_ordqid,  hcw_trinfo.info_ordpri, hcw_trinfo.info_ordidx, hcw_trinfo.info_lkid, hcw_trinfo.info_isldb, hcw_trinfo.info_ppidx, iptr), UVM_DEBUG); 
	       
  endfunction : set_hcw_trinfo  


  //---------------------------------------------------------------------------- 
  //-- update_hcw_with_trinfo
  //----------------------------------------------------------------------------   
  virtual function update_hcw_with_trinfo (hcw_transinfo  hcw_trinfoupd) ; 
      
      this.msgtype     =    hcw_trinfoupd.info_msgtype	  ;  
      this.isdir       =    hcw_trinfoupd.info_isdir	  ;  
      this.tbcnt       =    hcw_trinfoupd.info_tbcnt	  ;  
      this.qtypesch    =    hcw_trinfoupd.info_qtypesch	  ;  
      this.tbcntsch    =    hcw_trinfoupd.info_tbcntsch	  ;    
      this.lockid      =    hcw_trinfoupd.info_lkid	  ;  
      this.enqattr     =    hcw_trinfoupd.info_enqattr	  ;   
      this.reord       =    hcw_trinfoupd.info_reord	  ;   
      this.frg_cnt     =    hcw_trinfoupd.info_frg_cnt	  ;  
      this.frg_ldbcnt  =    hcw_trinfoupd.info_frg_ldbcnt ;        
      this.frg_last    =    hcw_trinfoupd.info_frg_last   ;  
      this.ordqid      =    hcw_trinfoupd.info_ordqid	  ;  
      this.ordpri      =    hcw_trinfoupd.info_ordpri	  ;  
      this.ordlockid   =    hcw_trinfoupd.info_ordlockid  ;  
      this.ordidx      =    hcw_trinfoupd.info_ordidx	  ;  
      this.prod_port   =    hcw_trinfoupd.info_ppidx      ; //--V2_TB
      this.prod_isldb  =    hcw_trinfoupd.info_isldb      ; //--V2_TB
      
      this.hcw_trinfo.info_msgtype	   =    hcw_trinfoupd.info_msgtype    ; 
      this.hcw_trinfo.info_isdir	   =    hcw_trinfoupd.info_isdir      ; 
      this.hcw_trinfo.info_tbcnt	   =    hcw_trinfoupd.info_tbcnt      ; 
      this.hcw_trinfo.info_qtypesch	   =    hcw_trinfoupd.info_qtypesch   ; 
      this.hcw_trinfo.info_tbcntsch	   =    hcw_trinfoupd.info_tbcntsch   ; 
      this.hcw_trinfo.info_lkid 	   =    hcw_trinfoupd.info_lkid       ; 
      this.hcw_trinfo.info_enqattr         =    hcw_trinfoupd.info_enqattr    ; 
      this.hcw_trinfo.info_reord	   =    hcw_trinfoupd.info_reord      ; 
      this.hcw_trinfo.info_frg_cnt	   =    hcw_trinfoupd.info_frg_cnt    ; 
      this.hcw_trinfo.info_frg_ldbcnt      =    hcw_trinfoupd.info_frg_ldbcnt ;       
      this.hcw_trinfo.info_frg_last	   =    hcw_trinfoupd.info_frg_last   ; 
      this.hcw_trinfo.info_ordqid	   =    hcw_trinfoupd.info_ordqid     ; 
      this.hcw_trinfo.info_ordpri	   =    hcw_trinfoupd.info_ordpri     ; 
      this.hcw_trinfo.info_ordlockid       =    hcw_trinfoupd.info_ordlockid  ; 
      this.hcw_trinfo.info_ordidx	   =    hcw_trinfoupd.info_ordidx     ; 
      this.hcw_trinfo.info_ppidx           =    hcw_trinfoupd.info_ppidx      ; //--V2_TB
      this.hcw_trinfo.info_isldb           =    hcw_trinfoupd.info_isldb      ; //--V2_TB
      	 
        uvm_report_info(get_type_name(),$psprintf("hcw_xaction:update_hcw_with_trinfo iptr=0x%0x; info_tbcnt=%0d/info_ordqid=0x%0x/info_ordpri=%0d/info_ordidx=%0d/info_lockid=0x%0x; getting tbcnt=%0d/ordqid=0x%0x/ordpri=%0d/ordidx=0x%0x/lockid=0x%0x/enqis_ldb=%0d/enqprod_port=%0d", 
                      iptr, hcw_trinfoupd.info_tbcnt, hcw_trinfoupd.info_ordqid, hcw_trinfoupd.info_ordpri, hcw_trinfoupd.info_ordidx, hcw_trinfoupd.info_lkid, tbcnt, ordqid, ordpri, ordidx, lockid, prod_isldb, prod_port), UVM_DEBUG); 
	       
  endfunction : update_hcw_with_trinfo   
  

  //---------------------------------------------------------------------------- 
  //---------------------------------------------------------------------------- 
  //-- other supporting functions 
  //----------------------------------------------------------------------------   
  extern   virtual         function   void         do_copy(uvm_object rhs);
  extern   virtual         function   bit          do_compare(uvm_object rhs, uvm_comparer comparer);
                                
endclass : hcw_transaction


//----------------------------------------------------------------------------
//-- do_copy
//----------------------------------------------------------------------------
function void hcw_transaction::do_copy(uvm_object rhs);
    hcw_transaction rhs_;
    
    if (!$cast(rhs_, rhs)) begin
       uvm_report_error(get_full_name(), $psprintf("input is not a hcw_transaction"));
    end 

    super.do_copy(this);

    qe_valid = rhs_.qe_valid;
    qe_orsp  = rhs_.qe_orsp;
    qe_uhl   = rhs_.qe_uhl;
    cq_pop   = rhs_.cq_pop;
    qtype    = rhs_.qtype;
    qtypesch = rhs_.qtypesch;
    cmp_id   = rhs_.cmp_id;
    dbg      = rhs_.dbg;
    rsvd0    = rhs_.rsvd0;
    msgtype   = rhs_.msgtype;
    directinfo   = rhs_.directinfo;
    lockid   = rhs_.lockid;
    qpri     = rhs_.qpri;
    qid      = rhs_.qid;
    idsi     = rhs_.idsi;
    iptr     = rhs_.iptr;
    dsi_error    = rhs_.dsi_error;
    cq_int_rearm = rhs_.cq_int_rearm;
    
    is_error   = rhs_.is_error;
    is_ldb     = rhs_.is_ldb;
    is_vf      = rhs_.is_vf;
    is_nm_pf   = rhs_.is_nm_pf;
    vf_num     = rhs_.vf_num;
    sch_cq_occ_cq  = rhs_.sch_cq_occ_cq;
    sch_cq_occ     = rhs_.sch_cq_occ;
    sch_parity     = rhs_.sch_parity;
    sch_error      = rhs_.sch_error;
    sch_qid_occ    = rhs_.sch_qid_occ;
    sch_write_status = rhs_.sch_write_status;
    sch_is_ldb     = rhs_.sch_is_ldb;
    sch_addr       = rhs_.sch_addr;  
    rtn_credit_only       = rhs_.rtn_credit_only;
    exp_rtn_credit_only       = rhs_.exp_rtn_credit_only;
    hcw_batch      = rhs_.hcw_batch;
    ingress_drop   = rhs_.ingress_drop;
    exp_ingress_drop   = rhs_.exp_ingress_drop;
    ingress_comp_nodrop= rhs_.ingress_comp_nodrop;
    sai        = rhs_.sai;
    ppid       = rhs_.ppid;
    vasid      = rhs_.vasid;
    sch_cqid   = rhs_.sch_cqid;
    vfid       = rhs_.vfid;
    pp_type_pp = rhs_.pp_type_pp;
    pf_qid     = rhs_.pf_qid;
    frg_num    = rhs_.frg_num;
    frg_cnt    = rhs_.frg_cnt;     
    frg_ldbcnt = rhs_.frg_ldbcnt;     
    frg_first  = rhs_.frg_first;     
    frg_last   = rhs_.frg_last;     
    sch_frg_last   = rhs_.sch_frg_last;     
    sch_frg_first  = rhs_.sch_frg_first;     
    is_sched   = rhs_.is_sched;
    is_compled = rhs_.is_compled;
    is_tokened = rhs_.is_tokened;   
    is_done    = rhs_.is_done;
    ord_state  = rhs_.ord_state;
    tbcnt      = rhs_.tbcnt;                 
    tbcntsch   = rhs_.tbcntsch;                 
    isdir      = rhs_.isdir;                 
    is_ord     = rhs_.is_ord;                 
    enqattr    = rhs_.enqattr;                 
    reord      = rhs_.reord;                 
    reordenq_done = rhs_.reordenq_done;                 
    ordqid     = rhs_.ordqid;                 
    ordpri     = rhs_.ordpri;                 
    ordlockid  = rhs_.ordlockid;                 
    ordidx     = rhs_.ordidx;                 
    reordidx   = rhs_.reordidx;                 
    
    qid_depth = rhs_.qid_depth;
    cq_gen    = rhs_.cq_gen;
    wu        = rhs_.wu;
    meas      = rhs_.meas;
    no_inflcnt_dec      = rhs_.no_inflcnt_dec;
    prod_port = rhs_.prod_port;
    prod_isldb = rhs_.prod_isldb;
	cq		  = rhs_.cq;
	cq_parity = rhs_.cq_parity;
	ecc_h     = rhs_.ecc_h;
	ecc_l     = rhs_.ecc_l;
 
endfunction

  
 
//----------------------------------------------------------------------------
//-- do_compare
//----------------------------------------------------------------------------
function   bit    hcw_transaction::do_compare(uvm_object rhs, uvm_comparer comparer);

    hcw_transaction that;

    if (!$cast(that, rhs)) begin
      return 0;
    end 

    if(this.compare_type==2'b0) 
        return((super.do_compare(rhs, comparer) &&
            (this.qtype        == that.qtype) &&    
            (this.cmp_id       == that.cmp_id) &&    
            (this.dbg          == that.dbg) &&    
            (this.msgtype      == that.msgtype) &&    
            (this.lockid       == that.lockid) &&    
            (this.qpri         == that.qpri) &&    
            (this.qid          == that.qid) &&    
            (this.idsi         == that.idsi) &&    
            (this.tbcnt        == that.tbcnt) &&    
            (this.tbcntsch     == that.tbcntsch) &&    
            (this.qtypesch     == that.qtypesch) &&    
            (this.iptr         == that.iptr)  ));
     else if(this.compare_type == 2'b01)
        return((this.dsi_error  == that.dsi_error) &&    
            (this.cq_int_rearm  == that.cq_int_rearm) &&    
            (this.qe_valid      == that.qe_valid) &&    
            (this.qe_orsp       == that.qe_orsp) &&    
            (this.qe_uhl        == that.qe_uhl) &&    
            (this.cq_pop        == that.cq_pop) &&    
            (this.cmp_id        == that.cmp_id) &&    
            (this.dbg           == that.dbg) &&    
            (this.lockid        == that.lockid) &&    
            (this.idsi          == that.idsi) &&    
            (this.directinfo    == that.directinfo) &&  
            (this.iptr          == that.iptr));
     else if(this.compare_type  == 2'b10)
        return((this.dsi_error  == that.dsi_error) &&    
            (this.qe_valid      == that.qe_valid) &&    
            (this.qe_orsp       == that.qe_orsp) &&    
            (this.qe_uhl        == that.qe_uhl) &&    
            (this.cq_pop        == that.cq_pop) &&  
            (this.lockid[9:0]   == that.lockid[9:0]));    
     else 
        return((this.dsi_error  == that.dsi_error) &&    
            (this.cq_int_rearm  == that.cq_int_rearm) &&    
            (this.qe_valid      == that.qe_valid) &&    
            (this.qe_orsp       == that.qe_orsp) &&    
            (this.qe_uhl        == that.qe_uhl) &&    
            (this.cq_pop        == that.cq_pop) &&    
            (this.cmp_id        == that.cmp_id) &&    
            (this.dbg           == that.dbg) &&    
            (this.lockid        == that.lockid) &&    
            (this.idsi          == that.idsi) &&    
            (this.directinfo    == that.directinfo));
           
endfunction
	    
`endif
