//                  TapID,          Opcode,       DR_Width,       Dummy_Hi (int),      Dummy_lo (int),      IsTapLinkOp (bit) 
Create_Reg_Model (cltap,             14'h31,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'h32,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'h34,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'h36,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'h44,  8,      10,       0,      0);
Create_Reg_Model (cltap,             14'h48,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'hB1,  16,      10,       0,      0);
Create_Reg_Model (cltap,             14'hB2,  16,      10,       0,      0);
Create_Reg_Model (cltap,             14'hF3,  16,      10,       0,      0);
Create_Reg_Model (cltap,             14'hF4,  16,      10,       0,      0);
Create_Reg_Model (cltap,             14'h4A,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'hF5,  8,      10,       0,      0);
Create_Reg_Model (cltap,             14'hF1,  5,      10,       0,      0);
Create_Reg_Model (cltap,             14'hF0,  2,      10,       0,      0);
Create_Reg_Model (cltap,             14'h1E,  68,      10,       0,      0);
Create_Reg_Model (cltap,             14'h1D,  1,      10,       0,      0);
Create_Reg_Model (cltap,             14'h10,  1,      10,       0,      0);
Create_Reg_Model (cltap,             14'h07,  1,      10,       0,      0);
Create_Reg_Model (cltap,             14'h05,  1,      10,       0,      0);
Create_Reg_Model (cltap,             14'h12,  2,      10,       0,      0);
Create_Reg_Model (cltap,             14'h11,  2,      10,       0,      0);
Create_Reg_Model (cltap,             14'h02,  32,      10,       0,      0);
Create_Reg_Model (cltap,             14'h3fff,  1,      10,       0,      0);
Create_Reg_Model (dfx_aggregator,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (dfx_aggregator,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap0,             8'h31,    32,      10,       0,      0);
Create_Reg_Model (stap0,             8'h32,    32,      10,       0,      0);
Create_Reg_Model (stap0,             8'h34,    32,      10,       0,      0);
Create_Reg_Model (stap0,             8'h36,    32,      10,       0,      0);
Create_Reg_Model (stap0,             8'hB0,    16,      10,       0,      0);
Create_Reg_Model (stap0,             8'hB1,    16,      10,       0,      0);
Create_Reg_Model (stap0,             8'hB2,    16,      10,       0,      0);
Create_Reg_Model (stap0,             8'hB3,    16,      10,       0,      0);
Create_Reg_Model (stap0,             8'hB4,    16,      10,       0,      0);
Create_Reg_Model (stap0,             8'hD1,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hD2,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE0,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE1,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE2,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE6,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE7,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE8,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hEF,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hE9,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hEA,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'hEB,    8,      10,       0,      0);
Create_Reg_Model (stap0,             8'h13,    1,      10,       0,      0);
Create_Reg_Model (stap0,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap0,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap1,             8'h07,    1,      10,       0,      0);
Create_Reg_Model (stap1,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap1,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap3,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap3,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap4,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap4,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap5,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap5,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap6,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap6,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap7,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap7,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap8,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap8,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap_extr,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap_extr,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap_extr3,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap_extr3,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap_extr4,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap_extr4,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap_extr1,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap_extr1,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (stap_extr2,             8'hC,    32,      10,       0,      0);
Create_Reg_Model (stap_extr2,             8'hff,    1,      10,       0,      0);
Create_Reg_Model (cltap,            14'h70,   12,      10,     0,      1);
Create_Reg_Model (cltap,            14'h144,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h145,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h146,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h147,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h140,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h141,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h142,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h143,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h540,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h541,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h542,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h543,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h80,   4,      10,     0,      1);
Create_Reg_Model (cltap,            14'h148,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h149,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h14a,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h14b,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h84,   16,      10,     0,      1);
Create_Reg_Model (cltap,            14'h154,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h155,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h156,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h157,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h150,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h151,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h152,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h153,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h14C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h14d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h14e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h14f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h164,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h165,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h166,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h167,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h88,   4,      10,     0,      1);
Create_Reg_Model (cltap,            14'h158,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h159,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h15a,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h15b,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h71,   8,      10,     0,      1);
Create_Reg_Model (cltap,            14'h18C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h18d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h18e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h18f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h15C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h15d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h15e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h15f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h72,   8,      10,     0,      1);
Create_Reg_Model (cltap,            14'h38C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h38d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h38e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h38f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h35C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h35d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h35e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h35f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h73,   8,      10,     0,      1);
Create_Reg_Model (cltap,            14'h28C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h28d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h28e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h28f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h25C,    14,       10,      2,  1);
Create_Reg_Model (cltap,            14'h25d,    1,       10,      1,   1);
Create_Reg_Model (cltap,            14'h25e,   30,      10,       0,     1);
Create_Reg_Model (cltap,            14'h25f,   18,       10,     2,     1);
Create_Reg_Model (cltap,            14'h1A0,    14,        10,     1,     1);
Create_Reg_Model (cltap,            14'h1a1,    1,         10,     0,      1);
