// File output was printed on: Wednesday, March 20, 2013 9:00:22 AM
// Chassis TAP Tool version: 0.6.1.2
// ---------------------------------------------------- 
case (Node)
   'd0 : begin
            Tap_Info_Int.Next_Tap[0] = NOTAP;
        end
   'd1 : begin
            Tap_Info_Int.Next_Tap[0] = STAP0;
            Tap_Info_Int.Next_Tap[1] = STAP1;
            Tap_Info_Int.Next_Tap[2] = STAP20;
            Tap_Info_Int.Next_Tap[3] = STAP27;
            Tap_Info_Int.Next_Tap[4] = STAP28;
            Tap_Info_Int.Next_Tap[5] = STAP29;
        end
   'd2 : begin
            Tap_Info_Int.Next_Tap[0] = STAP2;
            Tap_Info_Int.Next_Tap[1] = STAP8;
        end
   'd3 : begin
            Tap_Info_Int.Next_Tap[0] = STAP3;
            Tap_Info_Int.Next_Tap[1] = STAP4;
            Tap_Info_Int.Next_Tap[2] = STAP7;
        end
   'd4 : begin
            Tap_Info_Int.Next_Tap[0] = STAP5;
            Tap_Info_Int.Next_Tap[1] = STAP6;
        end
   'd5 : begin
            Tap_Info_Int.Next_Tap[0] = STAP9;
            Tap_Info_Int.Next_Tap[1] = STAP10;
            Tap_Info_Int.Next_Tap[2] = STAP11;
            Tap_Info_Int.Next_Tap[3] = STAP12;
            Tap_Info_Int.Next_Tap[4] = STAP13;
        end
   'd6 : begin
            Tap_Info_Int.Next_Tap[0] = STAP14;
            Tap_Info_Int.Next_Tap[1] = STAP19;
        end
   'd7 : begin
            Tap_Info_Int.Next_Tap[0] = STAP15;
            Tap_Info_Int.Next_Tap[1] = STAP16;
            Tap_Info_Int.Next_Tap[2] = STAP17;
            Tap_Info_Int.Next_Tap[3] = STAP18;
        end
   'd8 : begin
            Tap_Info_Int.Next_Tap[0] = STAP21;
            Tap_Info_Int.Next_Tap[1] = STAP22;
            Tap_Info_Int.Next_Tap[2] = STAP23;
            Tap_Info_Int.Next_Tap[3] = STAP24;
        end
   'd9 : begin
            Tap_Info_Int.Next_Tap[0] = STAP25;
            Tap_Info_Int.Next_Tap[1] = STAP26;
        end
endcase


