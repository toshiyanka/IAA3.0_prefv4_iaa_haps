// File output was printed on: Thursday, March 21, 2013 4:21:02 PM
// Chassis TAP Tool version: 0.6.1.2
//----------------------------------------------------------------------
parameter NUMBER_OF_HIER  = 0;
parameter NUMBER_OF_STAPS = 0;
parameter NUMBER_OF_TERTIARY_PORTS = 0;
